Netlist to Test out the period "." separator for device model parameters
*
* this netlist is the "baseline" so it should not be run with any -hspice-ext options.
*
V1 1 0 0.5V
D1 1 2 DFOR
R1 2 0 10k
.MODEL DFOR D
+ IS = 2.355E-14 N = 1.112 BV = 1000 IBV = 0.001
+ RS = 0.137 CJO = 2.993E-10 VJ = 0.5033 M = 0.3144
+ FC = 0.5 EG = 1.11 XTI = 3 TT = 1.7E-07

.print DC V(1) V(2)  DFOR:IS  {DFOR:IS}
.dc V1 0.5V 0.5V 0.5V

.end
