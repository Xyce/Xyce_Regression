Simple RC circuit, with expressions on AC line
**********************************************************************
Isrc 1 0 AC 1 0 sin(0 1 1e+5 0 0)
R1 1 0 1e3
C1 1 0 2e-6

.param first=10
.param second=1
.param third=1e5

.AC DEC {first} {second} {third}

.print ac v(1)

.END
