*******************************************************
* Test that Xyce exits gracefully with a reasonable error
* message if the specified file, on a .LIB or .INC line,
* does not exist.
*
********************************************************

V1 1 0 SIN(0 1 1HZ)
R1 1 2 1
R2 2 0 2

.TRAN 0 1S
.PRINT TRAN V(2)

* Note: bogo.lib and bogo.lib1 files do not exist
.INC "bogo.lib"
.LIB "bogo1.lib" bogo

.END

