TL431 Circuit

*ALIAS  V(8)=VOUT
.PRINT TRAN  V(8)
* NOOP used to forego the operating point 
* This circuit does not perform as an oscillator if an operating point 
* calculation is done --- the transient solution simply has to start from
* an all-0 initial condition.
*
.TRAN 1U 1.5M 5U NOOP

R1 2 4 .978K
R2 2 1 2.65K
C1 1 11 4.7N 
*VC1 1 11 OP 0
R3 11 7 5.56K
R4 11 0 2.64K
R5 4 5 9.77K
V1 5 0 18
V2 6 0 10
C2 8 3 10U 
*VC2 8 3 OP 0
R6 8 0 10
R9 3 0 5M
R10 8 7 8.2
C5 6 0 .1U 
X8 6 4 8 AEI150
I1 8 0 PULSE 0 1 80U 1U 1U 500U 1M
X1 2 0 11 TL431

* Subcircuit and Model Definitions

.SUBCKT TL431 7 6 11
*             K A FDBK
.MODEL DCLAMP D (IS=13.5N RS=25M N=1.59 
+ CJO=45P VJ=.75 M=.302 TT=50.4N BV=34V IBV=1MA)
V1 1 6 2.495
R1 6 2 15.6
C1 2 6 .5U
R2 2 3 100
C2 3 4 .08U
R3 4 6 10
G2 6 8 3 6 1.73
D1 5 8 DCLAMP
D2 7 8 DCLAMP
V4 5 6 2
G1 6 2 1 11 0.11
.ENDS

.SUBCKT AEI150 3 1 60
.MODEL AEI150A NMOS(VTO=3.9 KP=8.932 RS=.015 RD=.015 LAMBDA=.003)
.MODEL DMAX D(CJO=7N VJ=.2 M=.669)
.MODEL DMIN D (CJO=7N)
C1 1 0 3.5N
C2 1 3 266P
D1 2 3 DMAX
D2 2 1 DMIN
RB 1 1 1
M1 3 1 6 6 AEI150A
LS 6 60 10N
.ENDS
.END


