Test of DC output for general external coupling code
* This version depends on the "general external" device to do the actual
* evaluation of the equations, and as such it MUST be run through the
* "GenCouplingSimulator" API with an appropriate "VectorComputeInterface"
* implementation.
* This is primarily intended to test the output handling

V1 1 0 DC 1
* 1K ohm Resistor implemented as external device
YGenExt R1 1 0 DPARAMS={NAME=R VALUE=1K}
.dc v1 0 5 .5
.print DC v(1) I(V1)
.end
