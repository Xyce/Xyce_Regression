* test of coupled inductor parameters on the .PRINT line, with .STEP
V1 1 0 SIN(0 1 1KHz)
R1 1 0 1
R2 2 0 1

* mutual inductor definition
L1 1 0 1e-3
L2 2 0 2mH
K1 L1 L2 0.75

.step L1:L list 1e-3 2e-3 3e-3

.TRAN 0 1ms 
.PRINT TRAN V(1) V(2) L1:L {L1:L}

.END 

