* RC ladder circuit

* Note that this netlist does not have the C1 device in it.
* This is because that capacitance is already included in the
* Y-parameter model used by YLIN_MOD1.

v1 1 0  sin  0 5 1e4
*C1 2 0 1e-2
Rgs 1 2 0.02
YLIN YLIN1 2 0 5 0 6 0 7 0 12 0 YLIN_MOD1
.MODEL YLIN_MOD1 LIN TSTONEFILE=ylin-5port-yparam.cir.y5p

.options hbint numfreq=10 tahb=0
.hb 1e4
.print hb v(1) v(2) v(5) v(6) v(7) v(12) i(v1)

.END
