* Test use of .OPTIONS OUTPUT ADD_STEPNUM_COL=TRUE
*
* See SON Bug 1209 for more details.
**************************************************

* Trivial high-pass filter

R2 c 0 1
R1 b c 1
C1 a b 1u
V1 a 0 DC 0V AC 1

.SENS OBJVARS=B PARAM=c1:c

* only output direct sensitivities
.options sensitivity direct=1 adjoint=0 stdoutput=1

.OPTIONS OUTPUT ADD_STEPNUM_COL=true

.print AC vr(b) vi(b) vp(b) vm(b) R1:R C1:C
.PRINT SENS vr(b) vi(b) vp(b) vm(b) R1:R R2:R C1:C
.PRINT SENS FORMAT=NOINDEX FILE=ac-sens-stepnum-col.cir.FD.SENS.noindex.prn
+ vr(b) vi(b) vp(b) vm(b) R1:R R2:R C1:C
.PRINT SENS FORMAT=GNUPLOT FILE=ac-sens-stepnum-col.cir.FD.SENS.gnuplot.prn
+ vr(b) vi(b) vp(b) vm(b) R1:R R2:R C1:C
.PRINT SENS FORMAT=SPLOT FILE=ac-sens-stepnum-col.cir.FD.SENS.splot.prn
+ vr(b) vi(b) vp(b) vm(b) R1:R R2:R C1:C
.ac dec 5 100Hz 1e6
.STEP C1 1u 5u 4u

.end
