Test of MOS3 initial conditions
* This test is a 42-inverter chain.  Without any ICs, the operating point
* fails to converge.
* This circuit, unlike the 50-inverter MOS1 chain, requires more help than
* just setting the state of the penultimate inverter.  Here, we need to set
* three inverters to their desired states using IC=.  This is done by having
* one subcircuit that represents an initial "output low" inverter, and 
* another initial "output high" inverter.
* The IC is applied only at the first newton step of the DCOP, and this
* nudge is enough to get convergence.

.subckt INVERTER IN OUT VDD GND
MN1 OUT IN GND GND CD4012_NMOS L=5u W=175u
MP1 OUT IN VDD VDD CD4012_PMOS L=5u W=270u
.ends

.subckt INVERTEROFF IN OUT VDD GND
MN1 OUT IN GND GND CD4012_NMOS L=5u W=175u IC=0,5
MP1 OUT IN VDD VDD CD4012_PMOS L=5u W=270u IC=-5,0
.ends

.subckt INVERTERON IN OUT VDD GND
MN1 OUT IN GND GND CD4012_NMOS L=5u W=175u IC=5,0
MP1 OUT IN VDD VDD CD4012_PMOS L=5u W=270u IC=0,-5
.ends

* A small load (R1, C1) is applied to the output node, VOUT. The input signal
* is at 5V for 1.5us and then at 0V for 1.5us. The voltage at VOUT is high (4.8V)
* when VIN1 is low and vice versa.
** Analysis setup **
*
.tran 20ns 30us
.print tran PRECISION=10 WIDTH=19 v(vout) v(in) v(1)

VDDdev 	VDD	0	5V
RIN	IN	1	1K
VIN1  1	0  5V PULSE (5V 0V 1.5us 5ns 5ns 1.5us 3.01us)
R1    VOUT  0  10K  
C2    VOUT  0  0.1p
XINV1 IN OUT2 VDD 0 INVERTER
XINV2 OUT2 OUT3 VDD 0 INVERTER
XINV3 OUT3 OUT4 VDD 0 INVERTER
XINV4 OUT4 OUT5 VDD 0 INVERTER
XINV5 OUT5 OUT6 VDD 0 INVERTER
XINV6 OUT6 OUT7 VDD 0 INVERTER
XINV7 OUT7 OUT8 VDD 0 INVERTER
XINV8 OUT8 OUT9 VDD 0 INVERTER
XINV9 OUT9 OUT10 VDD 0 INVERTER
XINV10 OUT10 OUT11 VDD 0 INVERTER
XINV11 OUT11 OUT12 VDD 0 INVERTER
XINV12 OUT12 OUT13 VDD 0 INVERTER
XINV13 OUT13 OUT14 VDD 0 INVERTER
XINV14 OUT14 OUT15 VDD 0 INVERTER
XINV15 OUT15 OUT16 VDD 0 INVERTER
XINV16 OUT16 OUT17 VDD 0 INVERTER
XINV17 OUT17 OUT18 VDD 0 INVERTER
XINV18 OUT18 OUT19 VDD 0 INVERTER
XINV19 OUT19 OUT20 VDD 0 INVERTER
XINV20 OUT20 OUT21 VDD 0 INVERTER
XINV21 OUT21 OUT22 VDD 0 INVERTER
XINV22 OUT22 OUT23 VDD 0 INVERTER
XINV23 OUT23 OUT24 VDD 0 INVERTER
XINV24 OUT24 OUT25 VDD 0 INVERTER
XINV25 OUT25 OUT26 VDD 0 INVERTER
XINV26 OUT26 OUT27 VDD 0 INVERTER
XINV27 OUT27 OUT28 VDD 0 INVERTER
XINV28 OUT28 OUT29 VDD 0 INVERTER
XINV29 OUT29 OUT30 VDD 0 INVERTER
XINV30 OUT30 OUT31 VDD 0 INVERTER
XINV31 OUT31 OUT32 VDD 0 INVERTER
XINV32 OUT32 OUT33 VDD 0 INVERTER
XINV33 OUT33 OUT34 VDD 0 INVERTER
*This inverter must have initial conditions just to get the 32-bit intel 
* build to converge
XINV34 OUT34 OUT35 VDD 0 INVERTERON
* These seven inverters need initial conditions to assure that the operating
* point converges.  All 7 are required on builds with the Intel 
* compiler, only the last 3 are required with GCC builds.
XINV35 OUT35 OUT36 VDD 0 INVERTEROFF
XINV36 OUT36 OUT37 VDD 0 INVERTERON
XINV37 OUT37 OUT38 VDD 0 INVERTEROFF
XINV38 OUT38 OUT39 VDD 0 INVERTERON
XINV39 OUT39 OUT40 VDD 0 INVERTEROFF
XINV40 OUT40 OUT41 VDD 0 INVERTERON
XINV41 OUT41 OUT42 VDD 0 INVERTEROFF
*
XINV42 OUT42 VOUT VDD 0 INVERTER
.MODEL cd4012_pmos PMOS (
+ LEVEL = 3  UO = 310  VTO = -1.6  TOX = 6E-08  NSUB = 5.701E+15
+ NSS = 0    VMAX = 5.374E+04   RS = 5.359   RD = 93.66   RSH = 0   IS = 1E-14
+ XJ = 7.9E-06   LD = 3E-08   DELTA = 0   THETA = 0.0278   ETA = 0.535   KAPPA = 0.643
+ KP = 1.711E-05 L=5u W=270u GAMMA=0.37 PHI=0.65 NFS=1E10
+ CBD=0.1P CBS=0.1P PB=0.81 CGSO=2P CGBO=4P CGDO=2P CJ=2E-4 MJ=0.5 CJSW=1E-9
+ MJSW=0.5 JS=1E-8 TPG=0 KF=1E-25 AF=1 FC=0.5 TNOM=27)
**************************
.MODEL cd4012_nmos NMOS (
+ LEVEL = 3 UO = 190   VTO = 1.679    TOX = 6E-08   NSUB = 8.601E+15
+ NSS = 0   RS = 13.21   RD = 11.59   RSH = 0   IS = 1E-14
+ VMAX = 4.206E+04 NFS=1E10  GAMMA=0.37 PHI=0.65 
+ XJ = 7.1E-06   LD = 8.6E-07   DELTA = 0   THETA = 0.0021   ETA = 0.057   KAPPA = 0.15
+ KP = 2.161E-05  L=5u W=175u
+ CBD=0.1P CBS=0.1P PB=0.81 CGSO=2P CGBO=4P CGDO=2P CJ=2E-4 MJ=0.5 CJSW=1E-9
+ MJSW=0.5 JS=1E-8 TPG=0 KF=1E-25 AF=1 FC=0.5 TNOM=27)
.END
