* test of coupled inductor parameters on the .PRINT line, when inside subcircuit
V1 1 0 SIN(0 1 1KHz)
R1 1 0 2
R2 2 0 2

X1 1 2 foo

.subckt foo a b
* mutual inductor definition
L1 a 0 1e-3
L2 b 0 2mH
K1 L1 L2 0.75
.ends

.TRAN 0 1ms 
.PRINT TRAN V(1) V(2) X1:L1:L {X1:L1:L} {2.0*X1:L1:L} {X1:L1:L**2} {(X1:L1:L)*R1:R}
.END 

