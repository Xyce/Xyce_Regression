Current-Contolled Switch Circuit Netlist
*
IS 0 1 DC 40mA
VMON 1 1A 0V
R1 1A 0 100
VMON1 2 3 0
R2 3 0 100
W1 1 2 VMON SW OFF
.MODEL SW ISWITCH (ION=10mA IOFF=0mA RON=1 ROFF=1E6)
.DC IS 0 40mA 1mA
.PRINT DC I(IS) I(VMON) I(VMON1)
.END


