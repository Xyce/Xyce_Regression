*Sample netlist for BSIM-MG 
*Drain current symmetry for nmos

*.options nonlin abstol=1e-6 reltol=1e-6 
.options device temp=25 


* --- Voltage Sources ---
vdrain drain 0 dc .1
esource source 0 drain 0 -1
vgate gate  0 pulse (0v 1v 0s 10n 10n 1u 5u) 
vbulk bulk 0 dc 0.0


* --- Transistor ---
M1 drain gate source bulk nmos1 TFIN=15n L=30n NFIN=10 NRS=1 NRD=1

.options nonlin-tran rhstol=1e-7
.tran 1n 5u

* The sources are all set up so that their branch currents have the opposite sign of the
* lead currents.
.print tran {-I(vdrain)-ID(M1)} {-I(vgate)-IG(M1)} {-I(ESOURCE)-IS(M1)} {-I(VBULK)-IE(M1)}

.measure tran maxmag1   max {abs(-I(vdrain)-ID(M1))} failvalue=1e-6
.measure tran totalrms1 rms {-I(vdrain)-ID(M1)} failvalue=1e-6  
.measure tran maxmag2   max {abs(-I(vgate)-IG(M1))} failvalue=1e-6
.measure tran totalrms2 rms {-I(vgate)-IG(M1)} failvalue=1e-6  
.measure tran maxmag3   max {abs(-I(ESOURCE)-IS(M1))} failvalue=1e-6
.measure tran totalrms3 rms {-I(ESOURCE)-IS(M1)} failvalue=1e-6 
.measure tran maxmag4   max {abs(-I(VBULK)-IE(M1))} failvalue=1e-6
.measure tran totalrms4 rms {-I(VBULK)-IE(M1)} failvalue=1e-6 

*comp {-I(vdrain)-ID(M1)} abstol=1.0e-6 zerotol=1.0e-7
*comp {-I(vgate)-IG(M1)} abstol=1.0e-6 zerotol=1.0e-7
*comp {-I(ESOURCE)-IS(M1)} abstol=1.0e-6 zerotol=1.0e-7
*comp {-I(VBULK)-IE(M1)} abstol=1.0e-6 zerotol=1.0e-7

******** BSIM-MG 105 Sample Modelcard for NMOS ********

** The BSIM-MG sample modelcard below was not extracted/obtained
** from/based on any real technologies. It should not be used for any
** other purposes except for benchmarking the implementation of BSIM-MG
** against BSIM Team's standard results

.model nmos1 nmos level=107
+ BULKMOD = 1
+ CAPMOD = 0
+ COREMOD = 0
+ CGEOMOD = 0
+ DEVTYPE = 1
+ GEOMOD = 0
+ GIDLMOD = 1
+ IGBMOD = 0
+ IGCMOD = 1
+ IIMOD = 0
+ NGATE  = 0
+ NQSMOD = 0
+ RDSMOD = 0
+ RGATEMOD = 0
+ RGEOMOD = 0
+ NSEG = 5
+ SDTERM = 0
+ SHMOD = 0
+ AGIDL = 1.00E-12
+ AGISL = 1.00E-12
+ AIGC = 0.014
+ AIGD = 0.0115
+ AIGS = 0.0115
+ AT  = 0.001
+ BG0SUB  = 1.17
+ BGIDL = 1.00E+07
+ BGISL = 1.00E+07
+ BIGC = 0.005
+ BIGD = 0.00332
+ BIGS = 0.00332
+ CDSC = 0.01
+ CDSCD = 0.01
+ CFD = 0.20E-10
+ CFS = 0.20E-10
+ CGBL  = 0
+ CGBO  = 0
+ CGDL  = 0
+ CGDO = 1e-10
+ CGSL  = 0
+ CGSO = 1e-10
+ CIGC = 0.25
+ CIGD = 0.35
+ CIGS = 0.35
+ CIT = 0
+ CKAPPAD  = 0.6
+ CKAPPAS  = 0.6
+ CTH0  = 0.000001243
+ DELTAVSAT  = 0.5
+ DELTAW  = 0
+ DELTAWCV  = 0
+ DLBIN  = 0
+ DLC  = 0
+ DLCIGD = 1.00E-09
+ DLCIGS = 1.00E-09
+ DROUT = 1
+ DSUB = 0.5
+ DVT0 = 0.05
+ DVT1 = 0.5
+ DVTSHIFT = 0
+ EASUB  = 4.05
+ EGIDL = 0.35
+ EGISL = 0.35
+ EOT  = 1.50E-09
+ EOTACC  = 1.0000001E-10
+ EOTBOX  = 1.40E-07
+ EPSROX  = 3.9
+ EPSRSP  = 3.9
+ EPSRSUB  = 11.9
+ ETA0  = 0.05
+ ETAMOB = 2
+ ETAQM  = 0.54
+ EU = 1.2
+ FPITCH  = 4.00E-08
+ HFIN  = 3.00E-08
+ IGT  = 2.5
+ K1RSCE = 0
+ KSATIV = 2
+ KT1 = 0
+ KT1L = 0
+ L  = 2.50E-08
+ LINT  = -2.00E-09
+ LPE0 = 0
+ LCDSCD = 5.00E-05
+ LCDSCDR = 5.00E-05
+ LRDSW = 0.2
+ LVSAT = 0
+ MEXP = 4
+ NBODY  = 1.00E+22
+ NC0SUB  = 2.86E+25
+ NI0SUB  = 1.10E+16
+ NIGC = 1
+ NSD  = 2.00E+26
+ PCLM = 0.05
+ PCLMCV = 0.013
+ PCLMG = 0
+ PCLMGCV = 0
+ PDIBL1 = 0
+ PDIBL2 = 0.002
+ PHIG  = 4.39
+ PHIN = 0.05
+ POXEDGE = 1.1
+ PQM  = 0.66
+ PRT  = 0
+ PRWG  = 0
+ PTWG  = 0
+ PTWGT  = 0.004
+ PVAG = 0
+ QM0  = 0.001
+ QMFACTOR  = 2.5
+ RDSW  = 200
+ RDSWMIN  = 0
+ RDWMIN  = 0
+ RSHD  = 0
+ RSHS  = 0
+ RSWMIN  = 0
+ RTH0  = 0.225
+ TBGASUB = 0.000473
+ TBGBSUB = 636
+ TFIN  = 1.40E-08
+ TGIDL  = -0.007
+ TMEXP  = 0
+ TNOM = 25
+ TOXP  = 2.10E-09
+ U0 = 0.025
+ UA = 0.55
+ UA1 = 0.001032
+ UCS = 1
+ UCSTE = -0.004775
+ UD = 0
+ UD1 = 0
+ UP = 0
+ UTE = -0.7
+ UTL = 0
+ VASAT = 0.2
+ VASATCV = 0.2
+ VSAT = 80000
+ WR  = 1
+ WTH0  = 2.60E-07
+ XL  = 0
.end
