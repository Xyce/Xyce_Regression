********************************************************
* The purpose of this test is to verify that Xyce 
* does not seg-fault if both of these things happen:
*
*  1) a model card has unrecognized parameters in it.
*
*  2) those unrecognized parameters are set via expressions.
*
* The exact circuit doesn't really matter.  This uses
* the Diode Clipper example from the Users Guide.
********************************************************
VCC 1 0 5V
VIN 3 0 SIN(0V 10V 1kHz)

.TRAN 2ns 2ms
.PRINT TRAN V(3) V(2) V(4)

D1 2 1 D1N3940
D2 0 2 D1N3940
R1 2 3 1K
R2 1 2 3.3K
R3 2 0 3.3K
R4 4 0 5.6K
C1 2 4 0.47u
*
* GENERIC FUNCTIONAL EQUIVALENT = 1N3940
* TYPE: DIODE
* SUBTYPE: RECTIFIER
.MODEL D1N3940 D(
+ IS = 4E-10
+ RS = .105
+ N = 1.48
+ TT = 8E-7
+ CJO = 1.95E-11
+ VJ = .4
+ M = .38
+ EG = 1.36
+ XTI = -8
+ KF = 0
+ AF = 1
+ FC = .9
+ BV = 600
+ IBV = 1E-4
+ BOGOPARAM={1+2} )

.END

