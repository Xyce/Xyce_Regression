Unit Test for DLTCH Digital Device

* Analysis Commands
.DC V4 0 3 3 
.DC V3 0 3 3 
.DC V2 0 3 3 
.DC V1 0 3 3

* Sources
V1 in_pre 0 3V
V2 in_clr 0 3V
V3 in_enable 0 3V
V4 in_data 0 3V

* Digital power and reference node
V5 dig_pn 0 3V 

* Output
.print DC v(in_pre) v(in_clr) v(in_enable) 
+ v(in_data) v(out_q) v(out_qbar)

* Set digital default parameters:
.param R1HI=5 R1LO=200 R0HI=200 R0LO=5 RIN=1000 R1=100
.param SW=5.e-9  CAPOUT=1.e-12  CAPIN=1.e-12
.param V_LO=0 V_HI=3

UDLTCH1 DLTCH dig_pn 0 in_pre in_clr in_enable in_data out_q out_qbar DMOD

R1 out_q 0 100K
R2 out_qbar 0 100K

.model DMOD DIG ( CLO=CAPOUT  CHI=CAPOUT
+ S0RLO=R0LO  S0RHI=R0HI  S0TSW=SW
+ S0VLO=-1  S0VHI=1.8
+ S1RLO=R1LO  S1RHI=R1HI  S1TSW=SW
+ S1VLO=1  S1VHI=3
+ RLOAD=RIN   CLOAD=CAPIN 
+ DELAY=20ns )

.end