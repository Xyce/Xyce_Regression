********************************************************
* Test that Xyce exits gracefully with a reasonable error
* message if the specified restart file is a directory
* rather than a file.
*
* The contents of this netlist doesn't really matter.
* The .OPTIONS RESTART line is reading from a directory, 
* rather than from a file.
*
*
*********************************************************
V1 1 0 SIN(0 1 1HZ)
R1 1 2 1
R2 2 0 2

.TRAN 0 1S
.PRINT TRAN V(2)

* attempting to read a restart file that is actually a directory
.OPTIONS RESTART FILE=. START_TIME=0

.END 
