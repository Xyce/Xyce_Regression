Test of series RLC circuit
* This version depends on the "general external" device to do the actual
* evaluation of the equations, and as such it MUST be run through the
* "GenCouplingSimulator" API with an appropriate "VectorComputeInterface"
* implementation.
*
* This tests three of the devices implemented by the test harness

V1 1 0 SIN (5v 5v 20MEG)  AC 1
* 1K ohm Resistor implemented as external device
YGenExt R1 1 1a DPARAMS={NAME=R VALUE=1K}
* RLC network implemented as external device
YGenExt rlc1 1a 0 DPARAMS={NAME=R,L,C VALUE=1K,1m,1p}

* Voltage-controlled current source implemented as external device
* NOTE:  Due to a limitation of the Xyce netlist parser, "optional"
* nodes are NOT processed correctly unless a model name is found on the
* instance line.  So it is necessary to specify one, even though
* there are no model parameters for this device.
YGenExt vccs1 2 0 1a 0  foobar DPARAMS={NAME=TRANSCONDUCTANCE VALUE=1}
R1 2 0 1

*Dummy model card just to get around Xyce parser limitation.
.model foobar genext
.ac dec 30 1 1e7
.print ac FILE=ACnoindex.prn FORMAT=NOINDEX v(1) v(1a) I(v1) V(2)
.print ac v(1) v(1a) I(v1) V(2)
.end
