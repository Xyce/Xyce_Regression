* Lead current test for E and H sources, and the
* voltage form of a B-source, for a .AC analysis

* RESISTOR DIVIDER
V1  1 0 DC 5.0 AC  1.0
R1  1 2 1
R2  2 0 1
*
* AMP AND LP FILTER
EAMP  3 0 2 0 1
RLP1  3 4 100
CLP1  4 0 1.59NF

H5 5 0 V1 1
R5 5 0 1

B6 6 0 V={V(4)}
R6 6 0 1

.OP
.AC DEC 5 100 100MEG
.PRINT AC V(4) I(V1) I(B6) I(EAMP) I(H5)

.END
