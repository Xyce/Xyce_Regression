RAW File Output test for Lumped Line
************************************************************
* This test has two purposes:
*   1) Verify that the variable types are correct. In 
*      this case, the Lumped Line contributes various
*      branch currents and voltages to the solution vector.  
*      The source code (N_DEV_TransLine.C) provides more details.
*
*   2) Verify that the data is actually correct for all of
*      the time-steps in the .RAW file output 
*
* The "gold" .RAW file output was generated by manually
* comparing that "gold" file with a .PRN file.  It was 
* generated for a limited set of fixed time-steps, so that
* a file comparison could be used to verify the test output's
* .RAW file against that "gold" .RAW file.
************************************************************
*                 v1 v2 td tr tf pw per
VsigGen 1 0 pulse(0.0 1.0 0.0 5ns 5ns 0.49e-6 1.0e-6)
RsigGen 1 1b 50

X_tl DUT  1b rlconeinch

.tran 0 1.0e-6
.options output initial_interval=5e-8
.options timeint method=gear 

* .PRINT statement is not actually used for .RAW output.
* It was included in the netslit so that the "gold" .RAW 
* file output could manually verified against a .PRN file
* during test development
.print tran V(1) V(1B) V(DUT) N(l:x_tl:x1:1_branch)
+ N(l:x_tl:x2:1_branch) N(l:x_tl:x3:1_branch)
+ I(VSIGGEN) N(x_tl:3) N(x_tl:4) N(x_tl:x1:3)
+ N(x_tl:x2:3) N(x_tl:x3:3)

* start of cable model
.param Rcable=1.0e-3; ohm/foot
.param Lcable=0.5u  ; H/foot
.param Ccable=60p   ; F/foot

.subckt rlclump I O 
L1 I 3  {Lcable*0.1/12.0}
C1 O 0  {Ccable*0.1/12.0}
R1 3 O  {Rcable*0.1/12.0}
.ends rlclump 

.subckt rlconeinch I O
x1 I 3 rlclump
x2 3 4 rlclump
x3 4 0 rlclump
.ends rlconeinch

.end