Regression test for simple uniform distribution propagation via regression PCE, .param version
*
.param testNorm={aunif(2k,1k)}
.param R1value={testNorm*2.0}

R2 1 0 6K
R1 1 2 {R1value}
v1 2 0 1000V

.dc v1 1000 1000 1

.print dc format=tecplot v(1)

.result {v(1)}
*
.SAMPLING useExpr=true

.options SAMPLES numsamples=10
+ regression_pce=true
+ order=5
+ outputs={v(1)}
+ sample_type=lhs
+ stdoutput=true
+ resample=true

.end
