*****************************************************
* Test FORMAT=GNUPLOT without .STEP.  This should 
* produce the same .FD.prn file as FORMAT=STD.
*
*****************************************************

* Trivial high-pass filter (V-C-R) circuit
R1 b 0 2
C1 a b 1u
V1 a 0 DC 0V AC 1

.print AC FORMAT=GNUPLOT R1:R C1:C vm(b) 
.ac dec 5 100Hz 1e6

.end

