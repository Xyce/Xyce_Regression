*** Test RAND in UDF
.GLOBAL_PARAM X=0
.FUNC MYFUNC(A) {RAND()+(0.0*A)}
.OP
.STEP X 0 2 1
.PRINT DC FORMAT=STD V(STEP) V(RAND)
VSTEP STEP 0 DC {X}
RSTEP STEP 0 1
VRAND RAND 0 DC {MYFUNC(1.0)}
RRAND RAND 0 1
.END

