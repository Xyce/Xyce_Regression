* test of coupled inductor parameters on the .PRINT line, with .STEP
V1 1 0 SIN(0 1 1KHz)
R1 1 0 2
R2 2 0 2

* mutual inductor definition
L1 1 0 100
L2 2 0 100
K1 L1 L2 1.00 nlcore

.model nlcore core level=2 c=0.001

.step L1:L list 100 200 300

.TRAN 0 1ms 
.PRINT TRAN V(1) V(2) L1:L {L1:L} {R1:R*L1:L}

.END 

