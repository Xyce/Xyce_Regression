* Xyce gold netlist 
.TRAN  0 1ms
.PRINT TRAN FORMAT=PROBE V(N04173) V(N03179)

R_R1  N04173 N03179  1k
R_R2  N03179  0 2K
V_V1  N04173 0 SIN(0 1 1KHz 0 0 0)

.END 
