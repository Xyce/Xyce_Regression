DC test of -r output format
*
* Trivial resistor circuit, just do a DC sweep and watch the output
*

R1 1 0 10
V1 1 0 DC 0V

.print DC v(1) I(v1)
.dc v1 0 10 .1
.step temp -10 10 10

.end
