 
.include copper.linear
.param a1=1e-5
R1  1 0 copper L=0.1 a={a1}
v1  1 0 5

 
.tran 0 1
.print tran R1:R R1:TEMP i(r1) r1:a
.end
