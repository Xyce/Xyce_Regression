RAW File Output test for Thermal Resistor, Inductor and Capacitor
************************************************************
* This test has two purposes:
*   1) Verify that the variable type (e.g., "current") and 
*      variable names are correct.  The inductor should 
*      contribute a branch current in each case.  The 
*      capacitor C2 should contribute a branch current since
*      it has an IC= instance parameter.
*
*   2) Verify that no contributions in the raw file header
*      appear from a current source (I device) or a level 2
*      thermal resistor.
*
*   3) Verify that the data is actually correct for all of
*      the time-steps in the .RAW file output 
*
* The "gold" .RAW file output was generated by manually
* comparing that "gold" file with a .PRN file.  It was 
* generated for a limited set of fixed time-steps, so that
* a file comparison could be used to verify the test output's
* .RAW file against that "gold" .RAW file.
************************************************************

* capacitor does not have an IC instance parameter
V1   1 0 SIN(0 2 10 0)
R1   1 2 1
C1   2 3 1u
L1   3 0 1m

* capacitor does have an IC instance parameter
V2   4 0 SIN(0 2 10 0)
R2   4 5 5
C2   5 6 1u IC=0.0
L2   6 0 1m

* circuit and subcircuit definition for I and thermal resistor test
I1  7 0 sin(0 2 10 0 ) 
R3  7 0 copper L=0.1 a=1e-5

* Thermal / resistivity properties for copper
* resistivity is in units of ohm*m
.model copper r ( level=2
+ resistivity=
+ {table(temp+273.15,
+      0,         0.5e-9,
+      100,        3e-9,
+      1000,       6.6e-8
+  )} 

* heat capacity is in units or J/K/m**3
* density (8.92e+3 kg/m**3) times table in J/K/kg
+ heatcapacity={8.92e+3*table(temp+273.15,
+      0,         1,
+      1000,      1500 
+  )} )

.options output initial_interval=5ms
.TRAN 0.5U 100ms

* .PRINT statement is not actually used for .RAW output.
* It was included in the netslit so that the "gold" .RAW 
* file output could manually verified against a .PRN file
* during test development
.PRINT TRAN v(1) v(2) v(3) v(4) v(5) v(6) v(7)
+ N(c2_branch) N(l1_branch) N(l2_branch) 
+ I(V1) I(V2) 

.END
