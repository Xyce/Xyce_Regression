A test of the TEAM memristor device

vsrc n1 0  sin( 0 1 1000 0 )

.options timeint reltol= 1e-4
*rload n1 n2 100

.model mrm1 memristor level=2 ron=50 roff=1000 koff=1.46e-18 kon=-4.68e-22 alphaoff=10 alphaon=10 wc=1.0e-12 ioff=115e-6 ion=-8.9e-6 xscaling=1.0e9 wt=4
ymemristor mr1 n1 n2 mrm1

rptg n2 0 50 

*COMP v(n1) abstol=1.0e-5 
*COMP v(n2) offset=1
*COMP i(rptg) abstol=0.002
*COMP n(ymemristor!mr1_x) abstol=0.01
*COMP n(ymemristor!mr1:r)  reltol=0.02

.print tran v(n1)  v(n2) i(rptg) n(ymemristor!mr1_x) n(ymemristor!mr1:r)
.tran 0 10e-3

.end

