* TRAN test of FORMAT=CSV output format

V1 1 0 SIN(0 1 1)
R1 1 2 1
R2 2 0 1

.OPTIONS OUTPUT SNAPSHOTS=true INITIAL_INTERVAL=0.01
.PRINT TRAN PRECISION=10 FORMAT= CSV V(1) V(2)
.TRAN 0 1

.END


