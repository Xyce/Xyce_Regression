Test of various types of solution variables in Bsrc expressions

R1 1 node 990
V1 1 0 1

B1 node 0 I={V(node)/10}
H2  2  0  V1  -200
E3  3  0  1  0   3
B4  4  0  V={V(node)*100}
R2  2  0  1
R3  3  0  1
R4  4  0  1

BSUM  SUM  0  V={1+5*I(H2)/v(1)-I(E3)/4-I(B4)/4}
RSUM  SUM  0  1

.DC V1 1 10 1
.PRINT DC V(1) V(2) V(3) V(node) I(H2) I(E3) I(B4) V(SUM) {1+5*I(H2)/v(1)-I(E3)/4-I(B4)/4}

.END
