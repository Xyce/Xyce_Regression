********************************************************
* Test that Xyce exits gracefully with a reasonable error
* message if the specified save file is a directory
* rather than a file.
*
* The contents of this netlist doesn't really matter.
* The .SAVE line is writing to a directory rather than
* to a file.
*
*
*********************************************************
V1 1 0 SIN(0 1 1HZ)
R1 1 2 1
R2 2 0 2

.TRAN 0 1S
.PRINT TRAN V(2)

* attempting to write the Save file to a directory
.SAVE TYPE=IC FILE=.

.END 
