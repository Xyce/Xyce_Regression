*******************************************************
* Test that parameters and global parameters work when
* the TEMP variable is a dependent parameter.  This uses
* the default temperature of 27C.
*
* See SON Bug 1203 for more details.
*******************************************************

.PARAM ptemp=37
.GLOBAL_PARAM DTEMP=10
.GLOBAL_PARAM GTEMP=37

* R1:R should be 2
V1 1 0 1
R1 1 0 1  TC=0.1 temp={ptemp}

* R2:R should be 3
V2 2 0 1
R2 2 0 1 TC=0.1 temp={GTEMP+DTEMP}

.DC V2 1 5 1
.PRINT DC V(2) I(R1) R1:TEMP I(R2) R2:TEMP

.END
