Testing .MEASURE lines that are mismatched with the Analysis Types
*********************************************************************
* This tests the error messages that should occur if an AC, NOISE or
* DC mode measure is requested for a netlist that is doing a
* .TRAN analysis. 
* 
* See SON Bug 889 for more details.
*
*
*********************************************************************
VS  1  0  SIN(0 1.0 1KHZ 0 0)
R1  1  0  100
.TRAN 0 1ms
.PRINT TRAN FORMAT=NOINDEX V(1) 

* Test what happens when a DC or AC measure is requested for a .TRAN netlist
.MEASURE DC dcmax max v(1)
.MEASURE AC acmax max v(1)
.MEASURE NOISE noisemax max v(1)

.END

