CHEBYSHEV HIGH-PASS FILTER
********************************************************************************
* Tier No.: 3
* Directory/Circuit Name:SANDLER9/sandler9.cir
* Description:  Chebyshev high-pass filter circuit netlist developed by Steve
*       Sandler to compare the validity of simulations using three different
*       circuit simulation tools. The results were compared to measured data.
* Input: V2
* Output: VDB(5) VP(5)
********************************************************************************
*
* MAIN CIRCUIT DEFINITION
*
R3 10 0 2.35K
X2 7 5 6 8 5 UA741T
C3 3 2 .1U
C4 2 7 .1U
R6 7 0 46.5K
R7 2 5 1.32K
V2 4 0 AC 1
V3 6 0 15
V4 0 8 15
X3 10 3 6 8 3 UA741T
C1 4 10 .1U
*
* ANALYSIS AND OPTIONS
*
.AC DEC 40 10HZ 10K
*ALIAS  V(5)=OUT
*.PRINT AC  VDB(5)  VP(5) 
.PRINT AC  V(5) 
*.OPTION ACCT
*
* SUBCIRCUIT DEFINITION
*
.SUBCKT UA741T    1 2 3 4 5
*
C1   11 12 4.664E-12
C2    6  7 20.00E-12
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
*BEGND 99  0 V={POLY(2) V(3) V(4) 0 .5 .5}
BEGND 99  0 V=.5*V(3)+.5*V(4)
*BFB    7 99 I={POLY(5) I(VB) I(VC) I(VE) I(VLP) I(VLN) 0 10.61E6 -10E6 10E6 10E6 -10E6}
BFB    7 99 I=10.61e6*I(VB)-10e6*I(VC)+10e6*I(VE)+10e6*I(VLP)-10e6*I(VLN)
GA 6  0 11 12 137.7E-6
GCM 0  6 10 99 2.574E-9
IEE  10  4 DC 10.16E-6
HLIM 90  0 VLIM 1K
Q1   11  2 13 QX
Q2   12  1 14 QX
R2    6  9 100.0E3
RC1   3 11 7.957E3
RC2   3 12 7.957E3
RE1  13 10 2.740E3
RE2  14 10 2.740E3
REE  10 99 19.69E6
RO1   8  5 150
RO2   7 99 150
RP    3  4 18.11E3
VB    9  0 DC 0
VC 3 53 DC 2.600
VE   54  4 DC 2.600
VLIM  7  8 DC 0
VLP  91  0 DC 25
VLN   0 92 DC 25
.MODEL DX D(IS=800.0E-18)
.MODEL QX NPN(IS=800.0E-18 BF=62.50)
.ENDS
.END

