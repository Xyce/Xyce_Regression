*David Vigliano
*Sandia National Labs
*9/23/2014

*This netlis creates a pair of voltages divider.  Both are driven by a pulse but one of them has rf on top of them.  This is done to test out the noise cancellation technique 

*This source creates the sources

vp vp 0 PULSE(0 5 1us 6ns 6ns 2.029us 3.666us)
vrf vinrf vp SIN(0 5 10Meg)
vin vin 0 PULSE(0 5 1us 6ns 6ns 2.029us 3.666us)

*This section adds in the voltage dividers
R1 vinrf voutrf 1k
R2 voutrf 0 1k
R3 vin vout 1k
R4 vout 0 1k

*This section defines the simulation type
.TRAN .1ns 4us 0s .1ns
*.TRAN .1ns 10ns 0s .1ns


*This section generates the output data
.OPTIONS OUTPUT INITIAL_INTERVAL = .1ns
.print TRAN v(vinrf) v(voutrf) v(vin) v(vout) 
