* This netlist is used to test the return codes from the
* Python initialize() method for the -norun case.
* Note: this test currently causes the Python interface
* to segfault.  See SON Bug 1065 for more details.

V1 1 0 SIN(0 1 1)
R1 1 0 1

.TRAN 0 1
.PRINT TRAN V(1)

.END

