Window Detector Circuit
********************************************************************************
* Tier No.: 3
* Directory/Circuit Name:SANDLER25/sandler25.cir
* Description:  The window detector circuit netlist was developed 
*       by Steve Sandler to compare the validity of simulations 
*       using 3 different circuit simulation tools.  The results 
*       were compared to measured data.
* Input: V_IN=V(2)
* Output: V(2), V(10)
********************************************************************************
*
* MAIN CIRCUIT DEFINITION
*
R1 7 3 100
R2 7 34 1K
R3 5 0 149.2K
R4 5 7 9.72K
R5 34 6 4.7K
R6 3 10 6.8K
R7 2 1 2.2K
R8 7 4 9.72K
D1 0 7 ZN4733
Q1 10 6 0 QN2222A
X4 4 1 3 0 34 0 LM111T
X5 1 5 3 0 34 0 LM111T
V1 3 0 10
V_IN 2 0 PULSE(2 5 2.25M 1U 1U 2.75M 3M)
*
* ANALYSIS AND OPTION STATEMENTS
*
.OPTIONS NONLIN-TRAN SEARCHMETHOD=0

.TRAN 1U 16M 6M 
.PRINT TRAN precision=12 V(2)  V(10)
*ALIAS  V(2)=IN V(10)=OUT2
*******************************************************
* MODEL DEFINITIONS
*******************************************************
.MODEL ZN4733 D (IS=.703F RS=.871 N=1 BV=5.059 IBV=49M
+ CJO=189P VJ=.75 M=.33 TT=50.1N)
* MOTOROLA 5.1 VOLT  1 WATT  ZENER DIODE  06-15-1993
.MODEL QN2222A NPN (IS=81.1F NF=1 BF=205 VAF=113 IKF=.5
+ ISE=10.6P NE=2 BR=4 NR=1 VAR=24 IKR=.225 RE=.343 RB=1.37
+ RC=.137 XTB=1.5 CJE=29.5P CJC=15.2P TF=397P TR=85N)
*   MOTOROLA 40 VOLT  .8 AMP  400 MHZ  SINPN  TRANSISTOR  04-11-1991
*******************************************************
* SUBCIRCUIT DEFINITIONS
*******************************************************
.SUBCKT LM111T    1 2 3 4 5 6
*
*F1    9  3 V1 1
BF1 9 3 I={I(V1)}
IEE   3  7 DC 100.0E-6
VI1  21  1 DC .45
VI2  22  2 DC .45
Q1    9 21  7 QIN
Q2    8 22  7 QIN
Q3    9  8  4 QMO
Q4    8  8  4 QMI
.MODEL QIN PNP(IS=800.0E-18 BF=666.7)
.MODEL QMI NPN(IS=800.0E-18 BF=1002)
.MODEL QMO NPN(IS=800.0E-18 BF=1000 CJC=1E-15 TR=102.5E-9)
E1   10  6  9  4  1
V1   10 11 DC 0
Q5    5 11  6 QOC
.MODEL QOC NPN(IS=800.0E-18 BF=103.5E3 CJC=1E-15 TF=11.60E-12 TR=48.19E-9)
DP    4  3 DX
RP    3  4 6.667E3
.MODEL DX  D(IS=800.0E-18)
*
.ENDS
**********************************************************
.END

