*******************************************************************************
* This netlist is equivalent to Step 3 for the AverageTest.cir netlist.
* It has VS1:VA=2 and VS3:V0=-0.5
*
*******************************************************************************
*
* a few sources of different types
VS1  1  0  SIN(0 2.0 100HZ 0 0)
VP   2  0  PULSE( 0 100 2ms 2ms 2ms 10ms 20ms )
VS3  3  0  SIN(-0.5 1.0 100HZ 0 0.5)
VS4  4  0  SIN(0.5 -1.0 100HZ 0 0.5)

R1  1  0  100
R2  2  0  100
R3  3  0  100
R4  4  0  100

.TRAN 0  0.5
.PRINT TRAN FORMAT=NOINDEX V(1) V(2) V(3) V(4)

.measure tran averageAll avg V(1) 
.measure tran averageTop AVG V(2)

* add TO-FROM modifiers
.measure tran sineHalfInterval Avg V(1) FROM=0 TO=0.25

* mix in TDs before and after FROM value.
.measure tran sineTDbetween avg V(1) FROM=0 TO=0.25 TD=0.1
.measure tran sineTDbefore avg V(1) FROM=0.15 TO=0.25 TD=0.1

* this test should return -1
.measure tran returnNegOne avg V(1) FROM=0.2e-3 TO=0.25e-3 TD=0.5e-3

* add tests for rise/fall/cross.  V3 and VS4 have a DC offset
* and are damped sinusoids
.measure tran avgv3fall2 avg v(3) fall=2
.measure tran avgv4rise1 avg v(4) rise=1
.measure tran avgv3cross2 avg v(3) cross=2

* test LAST for rise/fall/cross
.measure tran avg3falllast avg v(3) fall=last
.measure tran avg4riselast avg v(4) rise=last
.measure tran avg3crosslast avg v(3) cross=last
.measure tran avg4crosslast avg v(4) cross=last

* test RFC_LEVEL keyword
.measure tran avg1Rise1RFClevel50 avg V(1) RFC_LEVEL=0.5 RISE=1
.measure tran avg1Fall1RFClevel50 avg V(1) RFC_LEVEL=0.5 FALL=1
.measure tran avg1Cross1RFClevel50 avg V(1) RFC_LEVEL=0.5 CROSS=1 

*test Failed measures for rise/fall/cross
.measure tran avg3fallfail avg v(3) fall=250
.measure tran avg4risefail avg v(4) rise=250
.measure tran avgv3crossfail avg v(3) cross=250

.END

