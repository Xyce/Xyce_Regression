Xyce netlist for Diode clipper circuit with transient analysis statement
*
* Voltage Sources
V1 N04104 0 5V
V2 N04173 0 SIN(0V 10V 1kHz)
* Analysis Command
.TRAN 0 2ms
* Output
*.PRINT TRAN FORMAT=PROBE V(N04173) V(N03179) V(N03334) W(D_D1) V(N04104)
.PRINT TRAN FORMAT=PROBE V(N04173) V(N03179) V(N03334) V(N04104)
* Diodes
D_D1 N03179 N04104 D1N3940
D_D2 0 N03179 D1N3940
* Resistors
R1 N03179 N04173 1K
R2 N04104 N03179 3.3K
R3 N03179 0 3.3K
R4 N03334 0 5.6K
* Capacitor
C1 N03179 N03334 0.47u
*
* GENERIC FUNCTIONAL EQUIVALENT = 1N3940
* TYPE: DIODE
* SUBTYPE: RECTIFIER
.MODEL D1N3940 D(
+ IS = 4E-10
+ RS = .105
+ N = 1.48
+ TT = 8E-7
+ CJO = 1.95E-11
+ VJ = .4
+ M = .38
+ EG = 1.36
+ XTI = -8
+ KF = 0
+ AF = 1
+ FC = .9
+ BV = 600
+ IBV = 1E-4)
*
.END
