power test for level 2 diode 
* This is based on the Level2_Temp_Dep_Breakdown.cir test from the DIODE subdirectory
VIN 1 0 pulse ( 7.5 10 1m 1 1 3 6)
R1  1 2 1k
DZR1 0 2 DZR  

R2 1 3 1K
DZR2 3 0 DZR

.MODEL DZR D( level=2
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 1P
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 7.255;7.25 yields vout=5V @25C;6.9504;Vref determines Vout
+        IBV = .001
+ tbv1 = 0.00013
+ tbv2 = -5e-8
+        
+ )

.TRAN 0 1 0 100m
.options timeint method=trap
.options nonlin-tran rhstol=1.0e-7

.PRINT TRAN v(2) i(dzr1) {i(dzr1)*(v(0)-v(2))} w(dzr1) p(dzr1) 
+ v(3) i(dzr2) {i(dzr2)*(v(3)-v(0))} w(dzr2) p(dzr2) 

.END
