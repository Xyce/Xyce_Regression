* Transient sensitivity example, PWL source, finite difference version
.param cap=1u
.param res=1K
.param v0=0
.param v1=1
.param v2=-1
.param v3=-0.5
.param v4=0.25
.param v5=0.75
.param v6=0.0

c1 1 0 cap
c2 2 0 cap
R1 1 3 res
R2 1 2 res

Vin 3 0 PWL(
+ 0 {v0}
+ 1ms {v1}
+ 2ms {v2}
+ 3ms {v3}
+ 4ms {v4}
+ 5ms {v5}
+ 6ms {v6}  )

* Transient commands
.tran 0 10ms 
.options timeint reltol=1e-6 abstol=1e-6

.print tran v(2)

* Sensitivity commands
.print sens 
.SENS objfunc={V(2)} param=v0,v1,v2, v3,v4,v5,v6
.options SENSITIVITY direct=1 adjoint=0 forcefd=true
.end

