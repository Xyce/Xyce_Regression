********************************************************
* Netlist to test Noise output in STD format 
* with .STEP
*
********************************************************

* NOISE ANALYSIS: RESISTOR DIVIDER, AMP, AND LP FILTER
*
* RESISTOR DIVIDER
V1  1 0 DC 5.0 AC  1.0   
R1  1 2 100K
R2  2 0 100K
*
* AMP AND LP FILTER
EAMP  3 0 2 0 1
RLP1  3 4 100
CLP1  4 0 1.59NF

.STEP RLP1 1e3 1e4 9e3
.NOISE  V(4)  V1  DEC  5 100 100MEG 1
.PRINT NOISE V(4) VR(4) VI(4) INOISE ONOISE

.END
