* A gilbert cell mixer, taken from a schematic off a ham radio web page
* http://engphys.mcmaster.ca/~elmer101/swgilb.html
* The original was used in a PSPICE simulation.  I had to guess at the
* transistors used, so I just used a model for a 2n2222 out of the SPUDS
* database.
R5 1 2 100
X3 3 2 4 PDEBJT
X4 5 6 4 PDEBJT
X5 3 6 8 PDEBJT
X6 5 2 8 PDEBJT
R6 2 1 100
*the local oscillator
VLO 6 2 DC 0 SIN(0 .05V 4e6 0 0)
X1 4 10 11 PDEBJT
R1 11 12 10
R2 12 13 10
* input bias current
I1 12 0 DC 1.8mA
X2 8 15 13 PDEBJT
R4 15 16 1500
R3 16 10 1500
V1 16 0 DC 1.8V
*the input voltage to be mixed with the LO
V5 15 10 DC 0 sin(0 .05V 3e6 0 0)
R7 5 17 1500
R8 3 17 1500
V3 17 0 DC 8V
V2 1 0 DC 6V

*--------------------------------------------------------------------------------
.subckt PDEBJT col bas emi
ypde npnop3 col bas emi pdebjt    
+ C0=1.0e+17
+ tecplotlevel=0 
+ gnuplotlevel=0
*+ mobmodel=philips
*+ fielddep=true
+ l=9.0e-4 nx=80
* DOPING REGIONS:
+ region={name       =            reg1,  reg2
+         function   =            file, file
+         file       =       boron.dat, phos.dat
+         nmaxchop   =         1.5e+18, 3.3e+19
+         type       =           ptype,  ntype
+         species    =              BM,  PP }
*
* ELECTRODES:
+ node={name           = collector,      base,  emitter
+       bc             = dirichlet, dirichlet,  dirichlet
+       side           =     right,    middle,  left
+       area           =    1.0e-3,    1.0e-3,  1.0e-3
+       location       =    9.0e-4,    3.0e-4,  0.0 }
*
.MODEL pdebjt ZOD  level=1
*--------------------------------------------------------------------------------
.ends

.options nonlin continuation=gmin
.options device debuglevel=-1000
.options LINSOL type=klu
.options timeint reltol=1e-4

.TRAN 1ns 1us 
* v(6,2) should be the LO voltage, v(15,10) is the input
* output is viewed as difference between collector voltages of Q4/Q6 and Q3/Q5.
* Basically the output should be the product of LO and input voltage, but 
* not exactly.  A fourier transform will show extra frequency components.
* Spurious mixer products (harmonics) are inevitable, although minimized 
* by lower input amplitudes.  
.PRINT TRAN {v(6,2)+0.1} {v(15,10)+0.1} {v(5,3)+1.5}
*.save v(6,2) v(15,10) v(5,3)
*.PLOT TRAN v(5,3)
.four 1MEG v(5,3)
.end
