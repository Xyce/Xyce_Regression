* DC simulation for xyce
.options device temp=27 gmin=1e-15
.subckt mysub d_x g_x s_x b_x tnode_x
e_d d_v 0 d_x 0 1
v_d d_v d 0
f_d d_x 0 v_d   -1
e_g g_v 0 g_x 0 1
v_g g_v g 0
f_g g_x 0 v_g   -1
e_s s_v 0 s_x 0 1
v_s s_v s 0
f_s s_x 0 v_s   -1
e_b b_v 0 b_x 0 1
v_b b_v b 0
f_b b_x 0 v_b   -1
v_tnode tnode tnode_x 0
m1 d g s b tnode mymodel
+ W=10.0e-6
+ L=0.1e-6
+ ASOURCE=5e-12
+ ADRAIN=5e-12
+ PSOURCE=21e-6
+ PDRAIN=21e-6
+ SA=0.5e-6
+ SB=0.5e-6
+ SD=0.2e-6
+ NF=1
+ MULT=1
+ DELVTO=0
+ FACTUO=1
.model mymodel pmos level=10240 TYPE=-1
+ SWSCALE=1
+ VERSION=102.4
+ TMAX=1000
+ SWIGN=1
+ SWJUNASYM=1
+ QMC=1.000000000
+ TR=25.00000000
+ LVARO=0.000000000
+ LVARL=0.000000000
+ LVARW=0.000000000
+ LAP=0.000000000
+ WVARO=0.000000000
+ WVARL=0.000000000
+ WVARW=0.000000000
+ WOT=0.000000000
+ DLQ=-4.10000000E-09
+ DWQ=0.000000000
+ TOXEO=0.910000000E-09
+ TSIO=6.600000000E-09
+ XGEO=0.000000000
+ TBOXO=25.40000000E-09
+ NCHO=5.000000000E+17
+ NSUBO=-0.730000000E+18
+ CTO=30.67249414E-03
+ TOXPO=2.000000000E-09
+ NOVO=3.000000000E+20
+ NOVDO=1.000000000E+20
+ VFBO=-85.0000000E-03
+ VFBL=-36.27000000E-06
+ VFBLEXP=2.000000000
+ VFBL2=0.000000000
+ VFBLEXP2=2.000000000
+ VFBW=0.000000000
+ VFBLW=0.000000000
+ VFBBO=0.000000000
+ VFBLBO=0.000000000
+ STVFBO=38.30000000E-06
+ STVFBL=-11.37932375E-03
+ STVFBW=0.000000000
+ STVFBLW=0.000000000
+ CICFO=1.000000000
+ CICO=1.000000000
+ PSCEL=0.553385193
+ PSCELEXP=2.000000000
+ PSCEW=0.000000000
+ PSCEBO=165.5916660E-03
+ NSDDCO=2.530103064E+19
+ PSCEDLBO=2.091746736E-03
+ PNCEW=0.000000000
+ CFL=1.660000000
+ CFLEXP=2.200000000
+ CFW=0.000000000
+ CFBO=1.000000000
+ STCFL=0.000000000
+ CFDO=300.0000000E-03
+ CFDLL=15.00000000E-03
+ CFDLW=0.000000000
+ CFDLBO=1.300000000E-03
+ UO=33.87331005E-03
+ FBET1=-866.6296939E-03
+ FBET1W=0.000000000
+ LP1=10.00000000E-09
+ LP1W=0.000000000
+ FBET2=0.000000000
+ LP2=10.00000000E-09
+ BETW1=0.000000000
+ BETW2=0.000000000
+ WBET=10.00000000E-09
+ BETNBO=1.245000000
+ STBETO=1.500000000
+ STBETL=-6.512771960E-03
+ STBETW=0.000000000
+ STBETLW=0.000000000
+ CSO=1.995520150
+ CSL=105.9306025E-03
+ CSLEXP=1.000000000
+ CSW=0.000000000
+ CSLW=0.000000000
+ CSFIO=72.24225909E-03
+ CSBIO=0.000000000
+ STCSO=2.500000000
+ STCSL=0.000000000
+ STCSW=0.000000000
+ STCSLW=0.000000000
+ THECSO=1.228510856
+ STTHECSO=187.0000000E-03
+ CSTHRO=4.319569985
+ CSTHRBO=1.037523586
+ MUEO=3.107732193
+ STMUEO=1.389237021
+ THEMUO=1.670000000
+ STTHEMUO=-507.6786970E-03
+ XCORO=-15.40016781E-03
+ XCORL=205.0000000E-06
+ XCORLEXP=1.000000000
+ XCORW=0.000000000
+ XCORLW=0.000000000
+ XCORBO=1.000000000
+ STXCORO=0.000000000
+ FETAO=1.000000000
+ RSW1=146.0000000
+ RSW2=0.000000000
+ RSIGO=0.000000000
+ STRSO=-2.534816734E-03
+ RSGO=14.73876165E-03
+ THERSGO=910.5509649E-03
+ RSBO=1.600000000E-03
+ THESATO=35.08000000
+ THESATL=17.00000000
+ THESATLEXP=570.0000000E-03
+ THESATW=0.000000000
+ THESATLW=0.000000000
+ STTHESATO=-400.0000000E-03
+ STTHESATL=0.000000000
+ STTHESATW=0.000000000
+ STTHESATLW=0.000000000
+ THESATGO=444.0902099E-12
+ THESATBO=60.00000000E-03
+ AXO=8.000000000
+ AXL=45.79000000E-03
+ AXLEXP=1.000000000
+ AXL2=2.00000000E-03
+ AXLEXP2=1.700000000
+ ALPL1=7.074000000E-03
+ ALPLEXP=700.0000000E-03
+ ALPL2=0.000000000
+ ALPLEXP2=2.000000000
+ ALPW=0.000000000
+ ALP1L1=4.600000000E-06
+ ALP1LEXP=500.0000000E-03
+ ALP1L2=0.000000000
+ ALP1LEXP2=1.500000000
+ ALP1W=0.000000000
+ ALPBO=0.000000000
+ VPO=1.000000000E-03
+ VPGO=7.600000000E-03
+ GCOO=0.000000000
+ IGINVLW=180.0000000E+03
+ IGOVINVW=4.560668843E-03
+ IGOVINVDW=0.000000000
+ IGOVACCW=0.000000000
+ IGOVACCDW=0.000000000
+ STIGO=0.000000000
+ GC2CHO=1.100000000
+ GC3CHO=63.00000000E-03
+ GC2OVINVO=1.742285026
+ GC3OVINVO=-365.6683549E-03
+ GC2OVACCO=375.0000000E-03
+ GC3OVACCO=63.00000000E-03
+ GCDOVL=40.00000000E-03
+ GCVDOVO=-1.500000000
+ CHIBO=3.100000000
+ NIGINVO=47.00000000E-03
+ FNOVINVW=1.000000000E+04
+ FNOVINVDW=0.000000000
+ GCOVINVFNO=0.300000000
+ STIGFNO=0.000000000
+ AGIDLO=1.500000000E-10
+ AGIDLW=1.320000000E-09
+ AGIDLDW=7.2000000000E-10
+ BGIDLO=18.160000000
+ BGIDLDO=14.900000000
+ STBGIDLO=0.000000E+00
+ STBGIDLDO=0.000000E+00
+ CGIDLO=0.000000E+00
+ CGIDLDO=0.000000E+00
+ DGIDLO=8.00000000E-03
+ DGIDLL=12.00000000E-03
+ DGIDLDL=0.000000000
+ A1O=5.000000000
+ A1L=0.000000000
+ A1W=0.000000000
+ A2O=2.000000000
+ STA2O=0.000000000
+ A3O=1.000000000
+ A3L=0.000000000
+ A3W=0.000000000
+ CGBOVO=0.000000000
+ CGBOVL=4.000000000E-17
+ FIFW=0.300000000
+ NSDACO=5.000000000E+19
+ LOVO=0.520000000E-09
+ LOVDO=0.000000000
+ COVDLO=27.20000000E-03
+ COVDLW=0.000000000
+ COVDLBO=0.000000000
+ DVFBOVO=0.000000000
+ CFRO=0.000000000
+ CFRDO=0.000000000
+ CFRW=162.8000000E-18
+ CFRDW=0.000000000
+ CSDO=1.000000000
+ CSDBPO=0.000000000
+ RTHO=259.4000000E+03
+ RTHL=29.70000000
+ RTHW=5.800000000
+ RTHLW=11.80000000
+ STRTHO=0.000000000
+ CTHO=11.80000000E-15
+ LAMBTHO=148.0000000E-9
+ FTHO=0.755000000
+ FNTO=1.000000000
+ FNTEXCL=1.000000000
+ FNTEXCLEXP=2.000000000
+ NFAW=0.000000000
+ NFALW=8.000000000E+22
+ NFBLW=30.00000000E+06
+ NFCLW=0.000000000
+ NFEO=0.000000000
+ NFEBO=0.000000000
+ EFO=1.000000000
+ SAREF=1.000000000E-06
+ SBREF=1.000000000E-06
+ WLOD=0.000000000
+ KUO=2.000000000E-08
+ KVSAT=0.100000000
+ TKUO=0.000000000
+ LKUO=0.000000000
+ WKUO=0.000000000
+ PKUO=0.000000000
+ LLODKUO=0.000000000
+ WLODKUO=0.000000000
+ KVTHO=2.000000000E-09
+ LKVTHO=0.000000000
+ WKVTHO=0.000000000
+ PKVTHO=0.000000000
+ LLODVTH=0.000000000
+ WLODVTH=0.000000000
+ STETAO=0.000000000
+ LODETAO=1.000000000
+ STRLAMBDA=100.0000000E-09
+ STRALPHA=3.000000000
+ STRDVFBO=-0.100000000
+ STRWDVFBO=0.000000000
+ STRDCFL=0.100000000
+ STRRUO=-1.200000000
+ STRTRUO=0.000000000
+ STRRVSAT=0.100000000
+ SWIGATE=0
+ SWGIDL=0
+ SWSHE=0
+ SWSUBDEP=0
+ SWSTRESS=0
+ SWIMPACT=0
.ends
v_d d 0 -1.0
v_g g 0 1.01
v_s s 0 0
v_b b 0 0
i_tnode tnode 0 0
x1 d g s b tnode mysub
.dc v_g 1.0 -1.2 -0.01
.step v_d list -.05 -1.0
.print dc V(g) v(d) i(v_d) i(v_g)  i(v_s)
.end
