Simple RC circuit
*
* Eric Keiter, SNL
*
* Tests simultaneous sweeps of frequency, magnitude and phase, using a
* data table to specify frequency, magnitude and phase.

.global_param mag=1
.global_param phase=0.1

Isrc 1 0 AC {mag} {phase} 
R1 1 0 1e3
C1 1 0 2e-6


.data table
+ mag phase freq
+  1.0   0.1  1.0e0
+  2.0   0.2  1.0e1
+  3.0   0.3  1.0e2
+  4.0   0.4  1.0e3
+  5.0   0.5  1.0e4
+  6.0   0.6  1.0e5
.enddata


.print ac 
+ {Isrc:acmag}
+ {Isrc:acphase}
+ v(1)

.AC data=table

.END
