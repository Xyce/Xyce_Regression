test multiplier

Vin 1 0 1.0
Rin 1 2 1.0

.param Mval=2

Xtest1 2 3 testA
Xtest2 3 0 testA

.subckt testA A B 
Xtest A B testB  M={Mval/30}
.ends

.subckt testB A B PARAMS: M=30
R1 A B 0.5 M=30
.ends

.dc Mval list 50 60 70
.PRINT DC Mval V(1) V(2) V(3) I(Vin)  { Xtest1:Xtest:R1:R } { Xtest2:Xtest:R1:R }

