* D:\Data\Toyon\TL431_Infineon.asc
VREF 1 N002 2.495V
RE 1 REF 1Meg
C1 1 REF 1pF
RCMPLUS 1 N002 1G
RCMMINUS REF N002 1G
BG1 N002 4 I={IF(40*V(1,REF)<V(CATHODE),40*V(1,REF),V(CATHODE))}
Rd 4 N002 1k
Cd 4 N002 10nF
BG2 N002 5 I={IF(V(4)>0, 0.1*V(4), 0)}
R2 5 N002 0.1
Dinvaus N002 CATHODE Dein
D1 6 5 Daus
Raus 6 CATHODE 0.1
Rmasse N002 0 0.0001
V1 N001 0 SIN(5 5 1k) AC 1
R1 CATHODE REF 10k
R3 REF 0 10k
R4 CATHODE N001 1k
*.TRAN 1n 10m
*.PRINT TRAN  V(CATHODE) V(4) V(1,REF)
.ac dec 1000 100 10Meg
.PRINT AC V(CATHODE) V(4) V(1,REF)
.MODEL Dein D RS=3 N=7.3 IS=100000000p
* IS = 100uA !!!
.MODEL Daus D RS=0.0001 
*CJO=10PF
.end
