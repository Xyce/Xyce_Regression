* test circuit

V1 1 0 1
R1 1 2 50
YLIN YLIN1 2 3 YLIN_MOD1
YLIN YLIN2 3 4 YLIN_MOD2
YLIN YLIN3 4 5 YLIN_MOD3
YLIN YLIN4 5 6 YLIN_MOD4
YLIN YLIN5 6 0 YLIN_MOD5

.MODEL YLIN_MOD1 LIN TSTONEFILE=sparam.cir.s1p
.MODEL YLIN_MOD2 LIN TSTONEFILE=sparam.cir.ma.s1p
.MODEL YLIN_MOD3 LIN TSTONEFILE=sparam.cir.db.s1p
.MODEL YLIN_MOD4 LIN TSTONEFILE=yparams.ts2.cir.s2p
.MODEL YLIN_MOD5 LIN TSTONEFILE=sparams.ts2.cir.s3p


.DC V1 1 5 1
.PRINT DC V(1) V(2) V(3) V(4) V(5) V(6)

.END
