Test of source sweeps

*Analysis directives: 
.dc vin 1 8 .1
.print dc v(1) v(2)
.print homotopy v(1) v(2)

.options device debuglevel=-100
.options device timeint=-100

************************************
* **** Start Homotopy Setup ****
************************************
.options nonlin nlstrategy=0 searchmethod=0
+ maxstep=50 maxsearchstep=20 in_forcing=0 AZ_Tol=1.0e-6 memory=0
+ continuation=1

.options loca stepper=0 predictor=0 stepcontrol=0
+ conparam=vsrcscale
+ initialvalue=0.0 minvalue=-1.0 maxvalue=1.0
+ initialstepsize=0.2 minstepsize=1.0e-4 maxstepsize=0.2
+ aggressiveness=1.0
+ maxsteps=5000 maxnliters=200
**********************************
* **** End Homotopy Setup ****
**********************************

VIN 1 0 DC 8
R1 1 2 2K
c1 2 0 1uF 

.END
