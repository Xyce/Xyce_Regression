Power test for F-source (Current Controlled Current Source)
* Use a B-source as the controlling voltage source
B1   1 0 V={2.0*sin(2*pi*TIME) }
R1   1 2 1K
R2   0 2 100

* Test both linear and POLY formats
FLIN  3 0 B1 1
R3    3 4 1K
R4    0 4 100

FPOLY  5 0 POLY(1) B1 0 1
R5     5 6 1K
R6     0 6 100

.options timeint method=trap
.options nonlin-tran rhstol=1.0e-7
.TRAN 0 1.0
.PRINT TRAN FORMAT=noindex v(3) I(Flin) {I(Flin)*v(3)} p(Flin) W(Flin)
+ v(5) I(Fpoly) {I(Fpoly)*v(5)} p(Fpoly) W(Fpoly)

.END
