simple RC
*

*.tran 0 1.0e-3 0 1e-6
.hb 1e5
.print tran  v(1) v(2) 
*i(v4)

*.options mpdeint ic=2 auton2=true saveicdata=1  diff=0 wampde=1 phase=0 phasecoeff=0  T2=1e-5 oscout=1
.options hbint numfreq=21 saveicdata=1 
*.options timeint maxord=1 
*.options timeint reltol=1e-3
*.options timeint-mpde erroption=1
*.options timeint method=7 reltol=1e-3   DEBUGLEVEL=0 
*.options timeint erroption=1
.options linsol type=aztecoo AZ_precond=0 use_ifpack_precond=0
*.options nonlin maxstep=10
*.options device voltlim=0

v0 1 0 sin 0 1v 1e5 0 0
*v0 n0 0 sin 0 1v 1e5 0 0
*v1 n1 n0 sin 0 1v 2e5 0 0
*v2 n2 n1 sin 0 1v 3e5 0 0
*v3 n3 n2 sin 0 1v 4e5 0 0
*v4 1 n3 sin 0 1V 5e5 0 0
*v1 1 0 DC 3.7V
r1 1 2 1k
c1 2 0 2u

.end
