* Unit Test of Series Power Grid Branch Devices, in PQ Rectangular format

* vary the voltage at bus 1 to check if the answers match theory,
* given on pg.250-254 of Kundar. Ammeter is defined so that power
* flows from bus 1 into the branch between buses 1 and 2
V1R bus1R ammBus1P 1V
V1I bus1I ammBus1Q 0V
Vamm1P 0 ammBus1P 0V
Vamm1Q 0 ammBus1Q 0V

* initial conditions ("flat start") at bus 2
.NODESET V(bus2R)=1 V(bus2I)=0

* Have bus 3 be the slack bus. Ammeter is defined so that power 
* flows from branch between buses 2 and 3 into bus 3, so as to match
* equations in Kundar.
V3R bus3R ammBus3P 1V
V3I bus3I ammBus3Q 0V
Vamm3P ammBus3P 0 0V
Vamm3Q ammBus3Q 0 0V

* two series branches should give same answer as one branch with X=2
YPowerGridBranch pg12 bus1R bus2R bus1I bus2I AT=PQR R=0.0 X=1.0 B=0.0
YPowerGridBranch pg23 bus2R bus3R bus2I bus3I AT=PQR R=0.0 X=1.0 B=0.0

.DC V1I -0.5 1.0 0.5 V1R -0.5 1.0 0.5
.PRINT DC width=10 precision=6 V(bus1R) V(bus1I) 
+ I(Vamm1P) I(Vamm1Q) I(Vamm3P) I(Vamm3Q)
 
.end
