Test of Python+Tensorflow series RLC circuit
* This version depends on the "general external" device to do the actual
* evaluation of the equations, and as such it MUST be run through the
* "GenCouplingSimulator" API with an appropriate "VectorComputeInterface"
* implementation.
*
* This tests three of the devices implemented by the test harness

V1 1 0 SIN (5v 5v 20MEG)
* 1K ohm Resistor implemented as external device
YGenExt PY1 1 1a DPARAMS={NAME=R VALUE=1K}
+ SPARAMS={NAME=MODULENAME VALUE=./models/resistor.py}
* RLC network implemented as external device
YGenExt PY2 1a 0 DPARAMS={NAME=R,L,C VALUE=1K,1m,1p}
+ SPARAMS={NAME=MODULENAME VALUE=./models/rlc.py}

* Voltage-controlled current source implemented as external device
* NOTE:  Due to a limitation of the Xyce netlist parser, "optional"
* nodes are NOT processed correctly unless a model name is found on the
* instance line.  So it is necessary to specify one, even though
* there are no model parameters for this device.
YGenExt PY3 2 0 1a 0  foobar DPARAMS={NAME=TRANSCONDUCTANCE VALUE=1}
+ SPARAMS={NAME=MODULENAME VALUE=./models/tf_dnn_vccs.py}
R1 2 0 1

*Dummy model card just to get around Xyce parser limitation.
.model foobar genext
.tran 1n 4u
*COMP V(1) offset=.1
*COMP V(1a) offset=.1
*COMP I(v1) abstol=1.25e-6 offset=9e-5
*COMP V(2) offset=-.1
* Note:  Order is important here, because xyce_verify can't handle
* multiple .print tran lines and gets cornfused.
.print tran file=starvar.prn v(*) I(*)
.print tran PRECISION=16 v(1) v(1a) I(v1) V(2)
.end
