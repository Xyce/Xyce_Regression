*** simple solar cell eq. circuit 

*** circuit layout 
* solar cell grain model 
* voltage source 
Vdd n1 0 1 


*** model definition
.MODEL dm1 D (LEVEL=1 IS=8.9393e-09 N=1.682) 
.MODEL dm2 D (LEVEL=1 IS=1.0700e-06 N=1.660) 
.MODEL dm3 D (LEVEL=1 IS=2.3600e-08 N=1.820) 
.MODEL dm4 D (LEVEL=1 IS=5.0600e-15 N=1.940) 
.MODEL dm5 D (LEVEL=1 IS=2.8600e-06 N=1.650) 
.MODEL dm6 D (LEVEL=1 IS=1.6000e-04 N=1.270) 
.MODEL dm7 D (LEVEL=1 IS=1.5100e-08 N=1.770) 
.MODEL dm8 D (LEVEL=1 IS=2.7300e-16 N=1.950) 
.MODEL dm9 D (LEVEL=1 IS=1.0300e-16 N=1.650) 
.MODEL dm10 D (LEVEL=1 IS=2.0100e-08 N=1.270) 
.MODEL dm11 D (LEVEL=1 IS=2.5900e-06 N=1.770) 
.MODEL dm12 D (LEVEL=1 IS=1.5500e-11 N=1.950) 
.MODEL dm13 D (LEVEL=1 IS=0.0000e+00 N=2.000) 
.MODEL dm14 D (LEVEL=1 IS=0.0000e+00 N=2.000) 

*** diode definition
D2 n3 0 dm1 AREA=4.190e-07
D3 n4 0 dm1 AREA=3.064e-07
D4 n5 0 dm1 AREA=5.062e-07
D5 n6 0 dm1 AREA=2.541e-07
D6 n7 0 dm1 AREA=4.298e-07
D7 n8 0 dm1 AREA=8.625e-07
D8 n9 0 dm1 AREA=9.339e-07
D9 n10 0 dm1 AREA=5.878e-07
D10 n11 0 dm1 AREA=1.559e-06
D11 n12 0 dm1 AREA=1.225e-06
D12 n13 0 dm1 AREA=1.127e-06
D13 n14 0 dm1 AREA=6.810e-07
D14 n15 0 dm1 AREA=9.285e-07
D15 n16 0 dm1 AREA=1.314e-06
D16 n17 0 dm1 AREA=6.018e-07
D17 n18 0 dm1 AREA=1.235e-06
D18 n19 0 dm1 AREA=2.556e-07
D19 n20 0 dm1 AREA=4.861e-07
D20 n21 0 dm1 AREA=1.103e-06
D21 n22 0 dm1 AREA=5.660e-07
D22 n23 0 dm1 AREA=4.605e-07
D23 n24 0 dm1 AREA=6.236e-07
D24 n25 0 dm1 AREA=6.088e-07
D25 n26 0 dm1 AREA=1.298e-06
D26 n27 0 dm1 AREA=7.569e-07
D27 n28 0 dm1 AREA=3.530e-07
D28 n29 0 dm1 AREA=4.491e-07
D29 n30 0 dm1 AREA=6.631e-07
D30 n31 0 dm1 AREA=1.128e-06
D31 n32 0 dm1 AREA=8.167e-07
D32 n33 0 dm1 AREA=7.455e-07
D33 n34 0 dm1 AREA=7.323e-07
D34 n35 0 dm1 AREA=9.119e-07
D35 n36 0 dm1 AREA=4.246e-07
D36 n37 0 dm1 AREA=7.176e-07
D37 n38 0 dm1 AREA=1.426e-06
D38 n39 0 dm1 AREA=1.314e-06
D39 n40 0 dm1 AREA=1.214e-06
D40 n41 0 dm1 AREA=1.936e-06
D41 n42 0 dm1 AREA=6.377e-07
D42 n43 0 dm1 AREA=9.413e-07
D43 n44 0 dm1 AREA=7.136e-07
D44 n45 0 dm1 AREA=1.331e-06
D45 n46 0 dm1 AREA=7.655e-07
D46 n47 0 dm1 AREA=7.247e-07
D47 n48 0 dm1 AREA=2.307e-07
D48 n49 0 dm1 AREA=1.277e-06
D49 n50 0 dm1 AREA=2.119e-06
D50 n51 0 dm1 AREA=7.286e-07
D51 n52 0 dm1 AREA=4.096e-07
D52 n53 0 dm1 AREA=4.957e-07
D53 n54 0 dm1 AREA=6.202e-07
D54 n55 0 dm1 AREA=8.884e-07
D55 n56 0 dm1 AREA=1.846e-06
D56 n57 0 dm1 AREA=5.088e-07
D57 n58 0 dm1 AREA=1.370e-06
D58 n59 0 dm1 AREA=9.885e-07
D59 n60 0 dm1 AREA=7.307e-07
D60 n61 0 dm1 AREA=1.574e-06
D61 n62 0 dm1 AREA=4.701e-07
D62 n63 0 dm1 AREA=3.521e-07
D63 n64 0 dm1 AREA=1.134e-06
D64 n65 0 dm1 AREA=6.607e-07
D65 n66 0 dm1 AREA=6.719e-07
D66 n67 0 dm1 AREA=2.565e-06
D67 n68 0 dm1 AREA=3.700e-07
D68 n69 0 dm1 AREA=1.314e-06
D69 n70 0 dm1 AREA=1.633e-06
D70 n71 0 dm1 AREA=1.193e-06
D71 n72 0 dm1 AREA=8.711e-07
D72 n73 0 dm1 AREA=6.286e-07
D73 n74 0 dm1 AREA=3.611e-07
D74 n75 0 dm1 AREA=1.399e-06
D75 n76 0 dm1 AREA=1.387e-06
D76 n77 0 dm1 AREA=1.630e-06
D77 n78 0 dm1 AREA=6.776e-07
D78 n79 0 dm1 AREA=1.236e-06
D79 n80 0 dm1 AREA=6.540e-07
D80 n81 0 dm1 AREA=9.424e-07
D81 n82 0 dm1 AREA=1.068e-06
D82 n83 0 dm1 AREA=8.713e-07
D83 n84 0 dm1 AREA=1.235e-06
D84 n85 0 dm1 AREA=1.127e-06
D85 n86 0 dm1 AREA=9.646e-07
D86 n87 0 dm1 AREA=5.929e-07
D87 n88 0 dm1 AREA=8.341e-07
D88 n89 0 dm1 AREA=4.546e-07
D89 n90 0 dm1 AREA=1.055e-06
D90 n91 0 dm1 AREA=8.806e-07
D91 n92 0 dm1 AREA=7.549e-07
D92 n93 0 dm1 AREA=6.124e-07
D93 n94 0 dm1 AREA=1.046e-06
D94 n95 0 dm1 AREA=7.094e-07
D95 n96 0 dm1 AREA=7.010e-07
D96 n97 0 dm1 AREA=9.498e-07
D97 n98 0 dm1 AREA=6.611e-07
D98 n99 0 dm1 AREA=1.736e-06
D99 n100 0 dm1 AREA=1.062e-06
D100 n101 0 dm1 AREA=5.478e-07
D101 n102 0 dm1 AREA=1.304e-06
D102 n103 0 dm1 AREA=1.498e-06
D103 n104 0 dm1 AREA=9.375e-07
D104 n105 0 dm1 AREA=1.111e-06
D105 n106 0 dm1 AREA=6.419e-07
D106 n107 0 dm1 AREA=7.029e-07
D107 n108 0 dm1 AREA=1.010e-06
D108 n109 0 dm1 AREA=2.309e-06
D109 n110 0 dm1 AREA=1.723e-06
D110 n111 0 dm1 AREA=1.128e-06
D111 n112 0 dm1 AREA=8.483e-07
D112 n113 0 dm1 AREA=1.161e-06
D113 n114 0 dm1 AREA=9.833e-07
D114 n115 0 dm1 AREA=7.142e-07
D115 n116 0 dm1 AREA=1.951e-06
D116 n117 0 dm1 AREA=9.904e-07
D117 n118 0 dm1 AREA=1.572e-06
D118 n119 0 dm1 AREA=9.237e-07
D119 n120 0 dm1 AREA=9.627e-07
D120 n121 0 dm1 AREA=7.365e-07
D121 n122 0 dm1 AREA=1.908e-06
D122 n123 0 dm1 AREA=1.114e-06
D123 n124 0 dm1 AREA=5.429e-07
D124 n125 0 dm1 AREA=8.227e-07
D125 n126 0 dm1 AREA=5.163e-07
D126 n127 0 dm1 AREA=9.082e-07
D127 n128 0 dm1 AREA=1.799e-06
D128 n129 0 dm1 AREA=7.372e-07
D129 n130 0 dm1 AREA=1.142e-06
D130 n131 0 dm1 AREA=2.547e-07
D131 n132 0 dm1 AREA=2.459e-06
D132 n133 0 dm1 AREA=1.634e-06
D133 n134 0 dm1 AREA=6.828e-07
D134 n135 0 dm1 AREA=1.258e-06
D135 n136 0 dm1 AREA=9.633e-07
D136 n137 0 dm1 AREA=1.437e-06
D137 n138 0 dm1 AREA=9.349e-07
D138 n139 0 dm1 AREA=1.189e-06
D139 n140 0 dm1 AREA=6.119e-07
D140 n141 0 dm1 AREA=6.820e-07
D141 n142 0 dm1 AREA=3.288e-07
D142 n143 0 dm1 AREA=7.578e-07
D143 n144 0 dm1 AREA=1.446e-06
D144 n145 0 dm1 AREA=9.524e-07
D145 n146 0 dm1 AREA=7.706e-07
D146 n147 0 dm1 AREA=7.518e-07
D147 n148 0 dm1 AREA=1.021e-06
D148 n149 0 dm1 AREA=2.872e-07
D149 n150 0 dm1 AREA=1.280e-06
D150 n151 0 dm1 AREA=7.318e-07
D151 n152 0 dm1 AREA=6.110e-07
D152 n153 0 dm1 AREA=3.461e-07
D153 n154 0 dm1 AREA=1.031e-06
D154 n155 0 dm1 AREA=1.276e-06
D155 n156 0 dm1 AREA=1.061e-06
D156 n157 0 dm1 AREA=1.520e-06
D157 n158 0 dm1 AREA=2.784e-07
D158 n159 0 dm1 AREA=8.815e-07
D159 n160 0 dm1 AREA=1.736e-06
D160 n161 0 dm1 AREA=7.552e-07
D161 n162 0 dm1 AREA=1.031e-06
D162 n163 0 dm1 AREA=9.168e-07
D163 n164 0 dm1 AREA=1.022e-06
D164 n165 0 dm1 AREA=1.863e-06
D165 n166 0 dm1 AREA=1.403e-07
D166 n167 0 dm1 AREA=7.623e-07
D167 n168 0 dm1 AREA=1.116e-06
D168 n169 0 dm1 AREA=6.604e-07
D169 n170 0 dm1 AREA=7.253e-07
D170 n171 0 dm1 AREA=8.543e-07
D171 n172 0 dm1 AREA=8.213e-07
D172 n173 0 dm1 AREA=1.388e-06
D173 n174 0 dm1 AREA=7.550e-07
D174 n1 0 dm1 AREA=3.116e-07
D175 n176 0 dm1 AREA=1.088e-06
D176 n177 0 dm1 AREA=6.280e-07
D177 n178 0 dm1 AREA=8.084e-07
D178 n179 0 dm1 AREA=2.384e-06
D179 n180 0 dm1 AREA=6.449e-07
D180 n181 0 dm1 AREA=6.942e-07
D181 n182 0 dm1 AREA=1.509e-06
D182 n183 0 dm1 AREA=9.229e-07
D183 n184 0 dm1 AREA=1.682e-06
D184 n185 0 dm1 AREA=1.518e-06
D185 n186 0 dm1 AREA=4.404e-07
D186 n187 0 dm1 AREA=6.991e-07
D187 n188 0 dm1 AREA=5.162e-07
D188 n189 0 dm1 AREA=5.656e-07
D189 n190 0 dm1 AREA=8.403e-07
D190 n191 0 dm1 AREA=8.540e-07
D191 n192 0 dm1 AREA=9.868e-07
D192 n193 0 dm1 AREA=8.153e-07
D193 n194 0 dm1 AREA=9.817e-07
D194 n195 0 dm1 AREA=1.354e-06
D195 n196 0 dm1 AREA=7.490e-07
D196 n197 0 dm1 AREA=1.812e-06
D197 n198 0 dm1 AREA=6.654e-07
D198 n199 0 dm1 AREA=7.075e-07
D199 n200 0 dm1 AREA=4.573e-07
D200 n201 0 dm1 AREA=5.507e-07
D201 n202 0 dm1 AREA=8.823e-07
D202 n203 0 dm1 AREA=6.509e-07
D203 n204 0 dm1 AREA=1.134e-06
D204 n205 0 dm1 AREA=9.513e-07
D205 n206 0 dm1 AREA=9.713e-07
D206 n207 0 dm1 AREA=2.493e-07
D207 n208 0 dm1 AREA=6.778e-07
D208 n209 0 dm1 AREA=4.802e-07
D209 n210 0 dm1 AREA=1.116e-06
D210 n211 0 dm1 AREA=6.809e-07
D211 n212 0 dm1 AREA=1.257e-06
D212 n213 0 dm1 AREA=4.486e-07
D213 n214 0 dm1 AREA=6.301e-07
D214 n215 0 dm1 AREA=6.827e-07
D215 n216 0 dm1 AREA=1.134e-06
D216 n217 0 dm1 AREA=5.581e-07
D217 n218 0 dm1 AREA=9.403e-07
D218 n219 0 dm1 AREA=2.426e-06
D219 n220 0 dm1 AREA=1.740e-06
D220 n221 0 dm1 AREA=7.440e-07
D221 n222 0 dm1 AREA=6.907e-07
D222 n223 0 dm1 AREA=7.625e-07
D223 n224 0 dm1 AREA=1.246e-06
D224 n225 0 dm1 AREA=8.199e-07
D225 n226 0 dm1 AREA=2.846e-07
D226 n227 0 dm1 AREA=1.329e-06
D227 n228 0 dm1 AREA=8.607e-07
D228 n229 0 dm1 AREA=4.208e-07
D229 n230 0 dm1 AREA=1.091e-06
D230 n231 0 dm1 AREA=7.345e-07
D231 n1 0 dm1 AREA=5.216e-07
D232 n233 0 dm1 AREA=8.843e-07
D233 n234 0 dm1 AREA=9.722e-07
D234 n235 0 dm1 AREA=5.683e-07
D235 n236 0 dm1 AREA=1.589e-06
D236 n237 0 dm1 AREA=1.701e-06
D237 n238 0 dm1 AREA=6.146e-07
D238 n239 0 dm1 AREA=4.949e-07
D239 n240 0 dm1 AREA=8.789e-07
D240 n241 0 dm1 AREA=5.355e-07
D241 n242 0 dm1 AREA=8.667e-07
D242 n243 0 dm1 AREA=1.357e-06
D243 n244 0 dm1 AREA=1.330e-06
D244 n245 0 dm1 AREA=2.681e-06
D245 n246 0 dm1 AREA=3.731e-07
D246 n247 0 dm1 AREA=4.759e-07
D247 n248 0 dm1 AREA=5.027e-07
D248 n249 0 dm1 AREA=6.673e-07
D249 n250 0 dm1 AREA=6.688e-07
D250 n251 0 dm1 AREA=3.095e-07
D251 n252 0 dm1 AREA=5.354e-07
D252 n253 0 dm1 AREA=1.169e-06
D253 n254 0 dm1 AREA=7.403e-07
D254 n255 0 dm1 AREA=1.281e-06
D255 n256 0 dm1 AREA=1.042e-06
D256 n257 0 dm1 AREA=8.482e-07
D257 n258 0 dm1 AREA=8.679e-07
D258 n259 0 dm1 AREA=8.126e-07
D259 n260 0 dm1 AREA=3.252e-07
D260 n261 0 dm1 AREA=9.272e-07
D261 n262 0 dm1 AREA=1.268e-06
D262 n263 0 dm1 AREA=9.098e-07
D263 n264 0 dm1 AREA=1.573e-06
D264 n265 0 dm1 AREA=7.835e-07
D265 n266 0 dm1 AREA=7.864e-07
D266 n267 0 dm1 AREA=9.937e-07
D267 n268 0 dm1 AREA=7.115e-07
D268 n269 0 dm1 AREA=1.178e-06
D269 n270 0 dm1 AREA=1.136e-06
D270 n271 0 dm1 AREA=6.752e-07
D271 n272 0 dm1 AREA=1.939e-06
D272 n273 0 dm1 AREA=1.347e-06
D273 n274 0 dm1 AREA=3.438e-07
D274 n275 0 dm1 AREA=1.341e-06
D275 n276 0 dm1 AREA=1.514e-06
D276 n277 0 dm1 AREA=2.482e-07
D277 n278 0 dm1 AREA=1.151e-06
D278 n1 0 dm1 AREA=9.026e-07
D279 n280 0 dm1 AREA=1.337e-06
D280 n281 0 dm1 AREA=7.364e-07
D281 n282 0 dm1 AREA=9.972e-07
D282 n283 0 dm1 AREA=1.071e-06
D283 n284 0 dm1 AREA=7.243e-07
D284 n285 0 dm1 AREA=7.236e-07
D285 n286 0 dm1 AREA=1.355e-06
D286 n287 0 dm1 AREA=2.349e-07
D287 n288 0 dm1 AREA=1.070e-06
D288 n289 0 dm1 AREA=8.990e-07
D289 n290 0 dm1 AREA=2.352e-07
D290 n291 0 dm1 AREA=9.428e-07
D291 n292 0 dm1 AREA=6.823e-07
D292 n293 0 dm1 AREA=1.057e-06
D293 n294 0 dm1 AREA=7.779e-07
D294 n295 0 dm1 AREA=6.273e-07
D295 n296 0 dm1 AREA=4.362e-07
D296 n297 0 dm1 AREA=9.841e-07
D297 n298 0 dm1 AREA=1.390e-06
D298 n299 0 dm1 AREA=6.086e-07
D299 n300 0 dm1 AREA=4.720e-07
D300 n301 0 dm1 AREA=4.765e-07
D301 n302 0 dm1 AREA=6.769e-07
D302 n303 0 dm1 AREA=1.955e-06
D303 n304 0 dm1 AREA=4.579e-07
D304 n305 0 dm1 AREA=5.280e-07
D305 n306 0 dm1 AREA=1.382e-06
D306 n307 0 dm1 AREA=5.889e-07
D307 n308 0 dm1 AREA=2.202e-07
D308 n309 0 dm1 AREA=6.689e-07
D309 n310 0 dm1 AREA=9.813e-07
D310 n311 0 dm1 AREA=1.336e-06
D311 n312 0 dm1 AREA=8.846e-07
D312 n313 0 dm1 AREA=7.759e-07
D313 n314 0 dm1 AREA=1.305e-06
D314 n315 0 dm1 AREA=4.139e-07
D315 n1 0 dm1 AREA=7.449e-07
D316 n317 0 dm1 AREA=4.299e-07
D317 n318 0 dm1 AREA=1.609e-06
D318 n319 0 dm1 AREA=7.397e-07
D319 n320 0 dm1 AREA=1.098e-06
D320 n321 0 dm1 AREA=3.681e-07
D321 n322 0 dm1 AREA=6.883e-07
D322 n323 0 dm1 AREA=7.436e-07
D323 n324 0 dm1 AREA=7.772e-07
D324 n325 0 dm1 AREA=1.470e-06
D325 n326 0 dm1 AREA=1.354e-06
D326 n327 0 dm1 AREA=5.480e-07
D327 n328 0 dm1 AREA=2.118e-06
D328 n329 0 dm1 AREA=1.825e-06
D329 n330 0 dm1 AREA=9.061e-07
D330 n331 0 dm1 AREA=1.019e-06
D331 n332 0 dm1 AREA=2.233e-06
D332 n333 0 dm1 AREA=2.277e-06
D333 n334 0 dm1 AREA=1.181e-06
D334 n335 0 dm1 AREA=1.263e-06
D335 n336 0 dm1 AREA=4.404e-07
D336 n337 0 dm1 AREA=1.720e-06
D337 n338 0 dm1 AREA=1.274e-06
D338 n339 0 dm1 AREA=1.582e-06
D339 n340 0 dm1 AREA=1.324e-06
D340 n341 0 dm1 AREA=4.545e-07
D341 n342 0 dm1 AREA=1.200e-06
D342 n343 0 dm1 AREA=1.324e-06
D343 n344 0 dm1 AREA=6.992e-07
D344 n345 0 dm1 AREA=2.438e-07
D345 n346 0 dm1 AREA=4.069e-07
D346 n347 0 dm1 AREA=5.276e-07
D347 n348 0 dm1 AREA=1.262e-06
D348 n349 0 dm1 AREA=1.625e-06
D349 n350 0 dm1 AREA=1.254e-06
D350 n351 0 dm1 AREA=8.401e-07
D351 n352 0 dm1 AREA=1.061e-06
D352 n353 0 dm1 AREA=1.533e-06
D353 n354 0 dm1 AREA=6.102e-07
D354 n355 0 dm1 AREA=1.656e-06
D355 n356 0 dm1 AREA=3.360e-07
D356 n357 0 dm1 AREA=5.933e-07
D357 n358 0 dm1 AREA=3.864e-07
D358 n359 0 dm1 AREA=1.766e-06
D359 n360 0 dm1 AREA=1.469e-06
D360 n361 0 dm1 AREA=7.867e-07
D361 n362 0 dm1 AREA=1.945e-06
D362 n363 0 dm1 AREA=1.010e-06
D363 n364 0 dm1 AREA=8.332e-07
D364 n365 0 dm1 AREA=5.336e-07
D365 n366 0 dm1 AREA=1.826e-06
D366 n367 0 dm1 AREA=2.866e-06
D367 n368 0 dm1 AREA=2.610e-06
D368 n369 0 dm1 AREA=1.125e-06
D369 n370 0 dm1 AREA=1.360e-06
D370 n371 0 dm1 AREA=7.868e-07
D371 n372 0 dm1 AREA=2.445e-06
D372 n373 0 dm1 AREA=9.505e-07
D373 n374 0 dm1 AREA=2.399e-06
D374 n375 0 dm1 AREA=4.883e-07
D375 n376 0 dm1 AREA=1.763e-06
D376 n377 0 dm1 AREA=3.044e-07
D377 n378 0 dm1 AREA=8.654e-07
D378 n379 0 dm1 AREA=6.796e-07
D379 n380 0 dm1 AREA=6.514e-07
D380 n381 0 dm1 AREA=7.339e-07
D381 n382 0 dm1 AREA=2.187e-06
D382 n383 0 dm1 AREA=1.229e-06
D383 n384 0 dm1 AREA=1.327e-06
D384 n385 0 dm1 AREA=3.797e-07
D385 n386 0 dm1 AREA=7.583e-07
D386 n387 0 dm1 AREA=9.801e-07
D387 n388 0 dm1 AREA=3.110e-07
D388 n389 0 dm1 AREA=5.515e-07
D389 n390 0 dm1 AREA=9.278e-07
D390 n391 0 dm1 AREA=9.598e-07
D391 n392 0 dm1 AREA=6.058e-07
D392 n393 0 dm1 AREA=1.298e-06
D393 n394 0 dm1 AREA=1.708e-06
D394 n395 0 dm1 AREA=7.262e-07
D395 n396 0 dm1 AREA=7.621e-07
D396 n397 0 dm1 AREA=7.406e-07
D397 n398 0 dm1 AREA=3.543e-07
D398 n1 0 dm1 AREA=2.022e-06
D399 n400 0 dm1 AREA=9.956e-07
D400 n401 0 dm1 AREA=6.255e-07
D401 n402 0 dm1 AREA=2.440e-06
D402 n403 0 dm1 AREA=1.041e-06
D403 n404 0 dm1 AREA=1.239e-06
D404 n405 0 dm1 AREA=1.294e-06
D405 n406 0 dm1 AREA=5.010e-07
D406 n407 0 dm1 AREA=6.876e-07
D407 n408 0 dm1 AREA=5.898e-07
D408 n409 0 dm1 AREA=7.510e-07
D409 n410 0 dm1 AREA=1.159e-06
D410 n411 0 dm1 AREA=5.910e-07
D411 n412 0 dm1 AREA=9.142e-07
D412 n413 0 dm1 AREA=1.595e-06
D413 n414 0 dm1 AREA=1.823e-07
D414 n415 0 dm1 AREA=1.948e-06
D415 n416 0 dm1 AREA=4.165e-07
D416 n417 0 dm1 AREA=5.817e-07
D417 n418 0 dm1 AREA=8.565e-07
D418 n419 0 dm1 AREA=4.761e-07
D419 n420 0 dm1 AREA=4.035e-07
D420 n421 0 dm1 AREA=1.128e-06
D421 n422 0 dm1 AREA=1.595e-07
D422 n423 0 dm1 AREA=2.733e-06
D423 n424 0 dm1 AREA=2.891e-06
D424 n425 0 dm1 AREA=1.096e-06
D425 n426 0 dm1 AREA=1.094e-06
D426 n427 0 dm1 AREA=7.784e-07
D427 n428 0 dm1 AREA=1.669e-06
D428 n429 0 dm1 AREA=1.020e-06
D429 n430 0 dm1 AREA=1.547e-06
D430 n431 0 dm1 AREA=8.184e-07
D431 n432 0 dm1 AREA=6.470e-07
D432 n433 0 dm1 AREA=6.844e-07
D433 n434 0 dm1 AREA=1.030e-06
D434 n435 0 dm1 AREA=9.088e-07
D435 n436 0 dm1 AREA=1.017e-06
D436 n437 0 dm1 AREA=8.821e-07
D437 n438 0 dm1 AREA=1.395e-06
D438 n439 0 dm1 AREA=5.393e-07
D439 n440 0 dm1 AREA=7.949e-07
D440 n441 0 dm1 AREA=1.985e-06
D441 n442 0 dm1 AREA=1.463e-07
D442 n443 0 dm1 AREA=1.672e-06
D443 n444 0 dm1 AREA=1.318e-06
D444 n445 0 dm1 AREA=1.108e-06
D445 n446 0 dm1 AREA=5.204e-07
D446 n447 0 dm1 AREA=1.397e-06
D447 n448 0 dm1 AREA=1.727e-06
D448 n449 0 dm1 AREA=4.613e-07
D449 n450 0 dm1 AREA=5.923e-07
D450 n451 0 dm1 AREA=1.643e-06
D451 n452 0 dm1 AREA=4.584e-07
D452 n453 0 dm1 AREA=1.333e-06
D453 n454 0 dm1 AREA=9.004e-07
D454 n455 0 dm1 AREA=3.383e-07
D455 n456 0 dm1 AREA=8.690e-07
D456 n457 0 dm1 AREA=1.395e-06
D457 n458 0 dm1 AREA=1.516e-06
D458 n459 0 dm1 AREA=3.992e-07
D459 n460 0 dm1 AREA=1.329e-06
D460 n461 0 dm1 AREA=9.907e-07
D461 n462 0 dm1 AREA=1.011e-06
D462 n463 0 dm1 AREA=2.384e-07
D463 n464 0 dm1 AREA=1.321e-06
D464 n465 0 dm1 AREA=2.070e-07
D465 n466 0 dm1 AREA=8.158e-07
D466 n467 0 dm1 AREA=9.289e-07
D467 n468 0 dm1 AREA=9.012e-07
D468 n469 0 dm1 AREA=8.395e-07
D469 n470 0 dm1 AREA=1.493e-06
D470 n471 0 dm1 AREA=1.527e-06
D471 n472 0 dm1 AREA=1.243e-06
D472 n473 0 dm1 AREA=1.916e-06
D473 n474 0 dm1 AREA=4.917e-07
D474 n475 0 dm1 AREA=5.112e-07
D475 n476 0 dm1 AREA=4.157e-07
D476 n477 0 dm1 AREA=2.187e-06
D477 n478 0 dm1 AREA=8.166e-07
D478 n479 0 dm1 AREA=1.621e-06
D479 n480 0 dm1 AREA=7.468e-07
D480 n481 0 dm1 AREA=4.014e-07
D481 n482 0 dm1 AREA=1.442e-06
D482 n483 0 dm1 AREA=3.818e-07
D483 n1 0 dm1 AREA=1.741e-06
D484 n485 0 dm1 AREA=1.495e-06
D485 n486 0 dm1 AREA=2.334e-06
D486 n487 0 dm1 AREA=6.252e-07
D487 n488 0 dm1 AREA=9.676e-07
D488 n489 0 dm1 AREA=1.114e-06
D489 n490 0 dm1 AREA=1.564e-07
D490 n491 0 dm1 AREA=2.065e-07
D491 n492 0 dm1 AREA=5.031e-07
D492 n493 0 dm1 AREA=2.327e-07
D493 n494 0 dm1 AREA=9.968e-07
D494 n495 0 dm1 AREA=7.256e-07
D495 n496 0 dm1 AREA=8.804e-07
D496 n497 0 dm1 AREA=6.504e-07
D497 n498 0 dm1 AREA=7.260e-07
D498 n499 0 dm1 AREA=5.206e-07
D499 n500 0 dm1 AREA=7.546e-07
D500 n501 0 dm1 AREA=1.110e-06
D501 n502 0 dm1 AREA=5.420e-07
D502 n503 0 dm1 AREA=5.765e-07
D503 n504 0 dm1 AREA=1.127e-06
D504 n505 0 dm1 AREA=1.644e-06
D505 n506 0 dm1 AREA=6.800e-07
D506 n507 0 dm1 AREA=1.084e-06
D507 n508 0 dm1 AREA=8.842e-07
D508 n509 0 dm1 AREA=1.732e-06
D509 n510 0 dm1 AREA=6.401e-07
D510 n511 0 dm1 AREA=1.119e-06
D511 n512 0 dm1 AREA=6.554e-07
D512 n513 0 dm1 AREA=1.146e-06
D513 n514 0 dm1 AREA=5.660e-07
D514 n515 0 dm1 AREA=7.115e-07
D515 n516 0 dm1 AREA=3.132e-07
D516 n517 0 dm1 AREA=7.536e-07
D517 n518 0 dm1 AREA=4.545e-07
D518 n519 0 dm1 AREA=6.963e-07
D519 n520 0 dm1 AREA=1.551e-06
D520 n521 0 dm1 AREA=6.956e-07
D521 n522 0 dm1 AREA=4.249e-07
D522 n523 0 dm1 AREA=2.653e-06
D523 n524 0 dm1 AREA=4.144e-07
D524 n525 0 dm1 AREA=1.132e-06
D525 n526 0 dm1 AREA=4.858e-07
D526 n527 0 dm1 AREA=1.065e-06
D527 n528 0 dm1 AREA=5.348e-07
D528 n529 0 dm1 AREA=1.303e-06
D529 n530 0 dm1 AREA=9.905e-07
D530 n531 0 dm1 AREA=2.518e-06
D531 n532 0 dm1 AREA=3.039e-07
D532 n533 0 dm1 AREA=2.148e-06
D533 n534 0 dm1 AREA=1.418e-06
D534 n535 0 dm1 AREA=3.358e-07
D535 n536 0 dm1 AREA=1.002e-06
D536 n537 0 dm1 AREA=2.771e-06
D537 n538 0 dm1 AREA=1.420e-06
D538 n539 0 dm1 AREA=8.497e-07
D539 n540 0 dm1 AREA=6.195e-07
D540 n541 0 dm1 AREA=7.575e-07
D541 n542 0 dm1 AREA=5.202e-07
D542 n543 0 dm1 AREA=1.725e-06
D543 n544 0 dm1 AREA=1.543e-06
D544 n545 0 dm1 AREA=1.047e-06
D545 n546 0 dm1 AREA=1.214e-06
D546 n547 0 dm1 AREA=7.092e-07
D547 n548 0 dm1 AREA=1.039e-06
D548 n549 0 dm1 AREA=8.370e-07
D549 n550 0 dm1 AREA=1.026e-06
D550 n551 0 dm1 AREA=1.716e-06
D551 n552 0 dm1 AREA=1.060e-06
D552 n553 0 dm1 AREA=1.036e-06
D553 n554 0 dm1 AREA=8.584e-07
D554 n555 0 dm1 AREA=1.142e-06
D555 n556 0 dm1 AREA=2.729e-07
D556 n557 0 dm1 AREA=1.723e-06
D557 n558 0 dm1 AREA=1.134e-06
D558 n559 0 dm1 AREA=8.916e-07
D559 n560 0 dm1 AREA=1.157e-06
D560 n561 0 dm1 AREA=1.700e-06
D561 n562 0 dm1 AREA=5.669e-07
D562 n563 0 dm1 AREA=1.389e-06
D563 n564 0 dm1 AREA=8.302e-07
D564 n565 0 dm1 AREA=3.631e-07
D565 n566 0 dm1 AREA=1.395e-06
D566 n567 0 dm1 AREA=8.817e-07
D567 n568 0 dm1 AREA=1.328e-06
D568 n569 0 dm1 AREA=1.430e-07
D569 n570 0 dm1 AREA=1.166e-06
D570 n571 0 dm1 AREA=3.760e-07
D571 n572 0 dm1 AREA=3.458e-07
D572 n573 0 dm1 AREA=1.021e-06
D573 n574 0 dm1 AREA=1.208e-06
D574 n575 0 dm1 AREA=6.848e-07
D575 n576 0 dm1 AREA=1.041e-06
D576 n577 0 dm1 AREA=1.532e-06
D577 n578 0 dm1 AREA=2.659e-07
D578 n579 0 dm1 AREA=1.078e-06
D579 n580 0 dm1 AREA=1.701e-06
D580 n581 0 dm1 AREA=2.596e-06
D581 n582 0 dm1 AREA=6.833e-07
D582 n583 0 dm1 AREA=1.255e-06
D583 n584 0 dm1 AREA=1.144e-06
D584 n585 0 dm1 AREA=1.042e-06
D585 n586 0 dm1 AREA=9.609e-07
D586 n587 0 dm1 AREA=1.201e-06
D587 n588 0 dm1 AREA=7.061e-07
D588 n589 0 dm1 AREA=4.006e-07
D589 n590 0 dm1 AREA=7.860e-07
D590 n591 0 dm1 AREA=1.772e-06
D591 n592 0 dm1 AREA=2.688e-07
D592 n593 0 dm1 AREA=1.070e-06
D593 n594 0 dm1 AREA=1.358e-06
D594 n595 0 dm1 AREA=1.045e-06
D595 n596 0 dm1 AREA=1.221e-06
D596 n597 0 dm1 AREA=9.846e-07
D597 n598 0 dm1 AREA=8.173e-07
D598 n599 0 dm1 AREA=5.454e-07
D599 n600 0 dm1 AREA=5.407e-07
D600 n601 0 dm1 AREA=7.823e-07
D601 n602 0 dm1 AREA=1.302e-06
D602 n603 0 dm1 AREA=9.015e-07
D603 n604 0 dm1 AREA=3.196e-07
D604 n605 0 dm1 AREA=1.333e-06
D605 n606 0 dm1 AREA=1.468e-06
D606 n607 0 dm1 AREA=1.006e-06
D607 n608 0 dm1 AREA=7.249e-07
D608 n609 0 dm1 AREA=1.080e-06
D609 n610 0 dm1 AREA=5.515e-07
D610 n611 0 dm1 AREA=1.474e-07
D611 n612 0 dm1 AREA=1.182e-06
D612 n613 0 dm1 AREA=8.533e-07
D613 n614 0 dm1 AREA=1.245e-06
D614 n615 0 dm1 AREA=9.486e-07
D615 n616 0 dm1 AREA=4.132e-07
D616 n617 0 dm1 AREA=2.537e-06
D617 n618 0 dm1 AREA=1.319e-06
D618 n619 0 dm1 AREA=1.278e-06
D619 n620 0 dm1 AREA=7.625e-07
D620 n621 0 dm1 AREA=6.512e-07
D621 n622 0 dm1 AREA=4.605e-07
D622 n623 0 dm1 AREA=1.017e-06
D623 n624 0 dm1 AREA=7.482e-07
D624 n625 0 dm1 AREA=6.140e-07
D625 n626 0 dm1 AREA=9.329e-07
D626 n627 0 dm1 AREA=2.441e-07
D627 n628 0 dm1 AREA=6.617e-07
D628 n629 0 dm1 AREA=5.607e-07
D629 n630 0 dm1 AREA=1.689e-06
D630 n631 0 dm1 AREA=4.120e-07
D631 n632 0 dm1 AREA=1.529e-06
D632 n633 0 dm1 AREA=4.789e-07
D633 n634 0 dm1 AREA=6.100e-07
D634 n635 0 dm1 AREA=2.032e-06
D635 n636 0 dm1 AREA=8.097e-07
D636 n637 0 dm1 AREA=4.979e-07
D637 n638 0 dm1 AREA=6.579e-07
D638 n639 0 dm1 AREA=2.312e-06
D639 n640 0 dm1 AREA=8.503e-07
D640 n641 0 dm1 AREA=8.522e-07
D641 n642 0 dm1 AREA=1.832e-06
D642 n643 0 dm1 AREA=6.469e-07
D643 n644 0 dm1 AREA=1.411e-06
D644 n645 0 dm1 AREA=4.632e-07
D645 n646 0 dm1 AREA=4.822e-07
D646 n647 0 dm1 AREA=2.553e-06
D647 n648 0 dm1 AREA=1.207e-06
D648 n649 0 dm1 AREA=1.278e-06
D649 n650 0 dm1 AREA=2.471e-06
D650 n651 0 dm1 AREA=8.734e-07
D651 n652 0 dm1 AREA=8.160e-07
D652 n653 0 dm1 AREA=6.939e-07
D653 n654 0 dm1 AREA=1.272e-06
D654 n655 0 dm1 AREA=8.753e-07
D655 n656 0 dm1 AREA=4.091e-07
D656 n657 0 dm1 AREA=8.357e-07
D657 n658 0 dm1 AREA=4.424e-07
D658 n659 0 dm1 AREA=6.915e-07
D659 n660 0 dm1 AREA=1.832e-06
D660 n661 0 dm1 AREA=1.621e-06
D661 n662 0 dm1 AREA=5.807e-07
D662 n663 0 dm1 AREA=7.805e-07
D663 n664 0 dm1 AREA=5.706e-07
D664 n665 0 dm1 AREA=7.901e-07
D665 n666 0 dm1 AREA=3.967e-07
D666 n667 0 dm1 AREA=1.208e-06
D667 n668 0 dm1 AREA=6.328e-07
D668 n669 0 dm1 AREA=9.679e-07
D669 n670 0 dm1 AREA=1.012e-06
D670 n671 0 dm1 AREA=6.815e-07
D671 n672 0 dm1 AREA=2.757e-06
D672 n673 0 dm1 AREA=1.220e-06
D673 n674 0 dm1 AREA=7.116e-07
D674 n675 0 dm1 AREA=5.721e-07
D675 n676 0 dm1 AREA=7.830e-07
D676 n677 0 dm1 AREA=1.020e-06
D677 n678 0 dm1 AREA=8.388e-07
D678 n679 0 dm1 AREA=6.864e-07
D679 n680 0 dm1 AREA=4.344e-07
D680 n681 0 dm1 AREA=1.602e-06
D681 n682 0 dm1 AREA=7.698e-07
D682 n683 0 dm1 AREA=9.344e-07
D683 n684 0 dm1 AREA=7.830e-07
D684 n685 0 dm1 AREA=2.538e-07
D685 n686 0 dm1 AREA=1.614e-06
D686 n687 0 dm1 AREA=7.077e-07
D687 n688 0 dm1 AREA=2.719e-06
D688 n689 0 dm1 AREA=1.071e-06
D689 n690 0 dm1 AREA=1.302e-06
D690 n691 0 dm1 AREA=9.688e-07
D691 n692 0 dm1 AREA=1.310e-06
D692 n1 0 dm1 AREA=9.627e-07
D693 n694 0 dm1 AREA=8.444e-07
D694 n695 0 dm1 AREA=1.319e-06
D695 n696 0 dm1 AREA=9.658e-07
D696 n697 0 dm1 AREA=5.479e-07
D697 n698 0 dm1 AREA=8.982e-07
D698 n699 0 dm1 AREA=2.068e-06
D699 n700 0 dm1 AREA=1.241e-07
D700 n701 0 dm1 AREA=4.449e-07
D701 n702 0 dm1 AREA=6.839e-07
D702 n703 0 dm1 AREA=8.093e-07
D703 n704 0 dm1 AREA=8.449e-07
D704 n705 0 dm1 AREA=4.703e-07
D705 n706 0 dm1 AREA=1.589e-06
D706 n707 0 dm1 AREA=1.006e-06
D707 n708 0 dm1 AREA=4.137e-07
D708 n709 0 dm1 AREA=2.921e-06
D709 n710 0 dm1 AREA=7.562e-07
D710 n711 0 dm1 AREA=1.619e-06
D711 n712 0 dm1 AREA=1.436e-06
D712 n713 0 dm1 AREA=4.636e-07
D713 n714 0 dm1 AREA=9.167e-07
D714 n715 0 dm1 AREA=1.103e-06
D715 n716 0 dm1 AREA=7.594e-07
D716 n717 0 dm1 AREA=7.290e-07
D717 n718 0 dm1 AREA=5.351e-07
D718 n719 0 dm1 AREA=1.626e-06
D719 n720 0 dm1 AREA=7.818e-07
D720 n721 0 dm1 AREA=9.533e-07
D721 n722 0 dm1 AREA=1.174e-06
D722 n723 0 dm1 AREA=2.427e-07
D723 n724 0 dm1 AREA=3.644e-07
D724 n725 0 dm1 AREA=1.509e-06
D725 n726 0 dm1 AREA=1.380e-06
D726 n727 0 dm1 AREA=1.082e-06
D727 n728 0 dm1 AREA=1.043e-06
D728 n729 0 dm1 AREA=7.722e-07
D729 n730 0 dm1 AREA=1.048e-06
D730 n731 0 dm1 AREA=6.595e-07
D731 n732 0 dm1 AREA=1.301e-06
D732 n733 0 dm1 AREA=4.704e-07
D733 n734 0 dm1 AREA=3.492e-07
D734 n735 0 dm1 AREA=1.642e-06
D735 n736 0 dm1 AREA=9.426e-07
D736 n737 0 dm1 AREA=1.462e-06
D737 n738 0 dm1 AREA=2.224e-06
D738 n739 0 dm1 AREA=1.663e-06
D739 n740 0 dm1 AREA=4.546e-07
D740 n741 0 dm1 AREA=1.365e-06
D741 n742 0 dm1 AREA=8.754e-07
D742 n743 0 dm1 AREA=4.151e-07
D743 n744 0 dm1 AREA=9.681e-07
D744 n745 0 dm1 AREA=7.806e-07
D745 n746 0 dm1 AREA=7.657e-07
D746 n747 0 dm1 AREA=1.069e-06
D747 n748 0 dm1 AREA=8.348e-07
D748 n749 0 dm1 AREA=8.844e-07
D749 n750 0 dm1 AREA=4.445e-07
D750 n751 0 dm1 AREA=1.017e-06
D751 n752 0 dm1 AREA=8.947e-07
D752 n753 0 dm1 AREA=2.024e-06
D753 n754 0 dm1 AREA=1.145e-06
D754 n755 0 dm1 AREA=2.592e-06
D755 n756 0 dm1 AREA=4.768e-07
D756 n757 0 dm1 AREA=5.990e-07
D757 n758 0 dm1 AREA=2.135e-06
D758 n759 0 dm1 AREA=1.491e-06
D759 n760 0 dm1 AREA=6.513e-07
D760 n761 0 dm1 AREA=7.460e-07
D761 n762 0 dm1 AREA=1.779e-06
D762 n763 0 dm1 AREA=2.858e-07
D763 n764 0 dm1 AREA=6.881e-07
D764 n765 0 dm1 AREA=1.110e-06
D765 n766 0 dm1 AREA=8.967e-07
D766 n767 0 dm1 AREA=1.082e-06
D767 n768 0 dm1 AREA=1.366e-06
D768 n769 0 dm1 AREA=1.290e-06
D769 n770 0 dm1 AREA=5.053e-07
D770 n771 0 dm1 AREA=8.371e-07
D771 n772 0 dm1 AREA=3.644e-06
D772 n773 0 dm1 AREA=4.643e-07
D773 n774 0 dm1 AREA=7.137e-07
D774 n775 0 dm1 AREA=8.266e-07
D775 n776 0 dm1 AREA=7.646e-07
D776 n777 0 dm1 AREA=4.175e-07
D777 n778 0 dm1 AREA=8.160e-07
D778 n779 0 dm1 AREA=1.271e-06
D779 n780 0 dm1 AREA=9.448e-07
D780 n781 0 dm1 AREA=1.181e-06
D781 n782 0 dm1 AREA=8.394e-07
D782 n783 0 dm1 AREA=1.034e-06
D783 n784 0 dm1 AREA=1.016e-06
D784 n785 0 dm1 AREA=1.579e-06
D785 n786 0 dm1 AREA=2.905e-07
D786 n787 0 dm1 AREA=8.890e-07
D787 n788 0 dm1 AREA=1.613e-06
D788 n789 0 dm1 AREA=1.568e-06
D789 n790 0 dm1 AREA=6.790e-07
D790 n791 0 dm1 AREA=5.599e-07
D791 n792 0 dm1 AREA=4.254e-07
D792 n793 0 dm1 AREA=1.426e-06
D793 n794 0 dm1 AREA=1.074e-06
D794 n795 0 dm1 AREA=1.205e-06
D795 n796 0 dm1 AREA=2.887e-07
D796 n797 0 dm1 AREA=1.008e-06
D797 n798 0 dm1 AREA=8.800e-07
D798 n799 0 dm1 AREA=1.179e-06
D799 n800 0 dm1 AREA=8.074e-07
D800 n801 0 dm1 AREA=1.492e-06
D801 n802 0 dm1 AREA=2.088e-07
D802 n803 0 dm1 AREA=5.726e-07
D803 n804 0 dm1 AREA=5.478e-07
D804 n805 0 dm1 AREA=4.491e-07
D805 n806 0 dm1 AREA=1.179e-06
D806 n807 0 dm1 AREA=1.456e-06
D807 n808 0 dm1 AREA=1.467e-06
D808 n809 0 dm1 AREA=1.305e-06
D809 n810 0 dm1 AREA=9.733e-07
D810 n811 0 dm1 AREA=6.564e-07
D811 n812 0 dm1 AREA=1.036e-06
D812 n813 0 dm1 AREA=1.277e-06
D813 n814 0 dm1 AREA=1.457e-06
D814 n815 0 dm1 AREA=1.073e-06
D815 n816 0 dm1 AREA=9.696e-07
D816 n817 0 dm1 AREA=1.324e-06
D817 n818 0 dm1 AREA=7.199e-07
D818 n819 0 dm1 AREA=1.143e-06
D819 n820 0 dm1 AREA=5.278e-07
D820 n821 0 dm1 AREA=1.282e-06
D821 n822 0 dm1 AREA=3.693e-07
D822 n823 0 dm1 AREA=1.002e-06
D823 n824 0 dm1 AREA=9.389e-07
D824 n825 0 dm1 AREA=9.990e-07
D825 n826 0 dm1 AREA=8.635e-07
D826 n827 0 dm1 AREA=2.124e-06
D827 n828 0 dm1 AREA=3.769e-07
D828 n829 0 dm1 AREA=1.358e-06
D829 n830 0 dm1 AREA=1.949e-06
D830 n831 0 dm1 AREA=8.666e-07
D831 n832 0 dm1 AREA=1.415e-06
D832 n833 0 dm1 AREA=1.190e-06
D833 n834 0 dm1 AREA=7.378e-07
D834 n835 0 dm1 AREA=1.567e-06
D835 n836 0 dm1 AREA=3.189e-06
D836 n837 0 dm1 AREA=4.309e-07
D837 n838 0 dm1 AREA=1.753e-06
D838 n839 0 dm1 AREA=5.664e-07
D839 n840 0 dm1 AREA=6.919e-07
D840 n841 0 dm1 AREA=1.223e-06
D841 n842 0 dm1 AREA=1.605e-06
D842 n843 0 dm1 AREA=2.555e-07
D843 n844 0 dm1 AREA=1.040e-06
D844 n845 0 dm1 AREA=5.596e-07
D845 n846 0 dm1 AREA=1.171e-06
D846 n847 0 dm1 AREA=6.538e-07
D847 n848 0 dm1 AREA=1.390e-06
D848 n849 0 dm1 AREA=7.676e-07
D849 n850 0 dm1 AREA=7.106e-07
D850 n851 0 dm1 AREA=1.389e-06
D851 n852 0 dm1 AREA=7.680e-07
D852 n853 0 dm1 AREA=1.879e-06
D853 n854 0 dm1 AREA=6.843e-07
D854 n855 0 dm1 AREA=1.364e-06
D855 n856 0 dm1 AREA=9.267e-07
D856 n857 0 dm1 AREA=7.744e-07
D857 n858 0 dm1 AREA=1.019e-06
D858 n859 0 dm1 AREA=3.636e-07
D859 n860 0 dm1 AREA=1.017e-06
D860 n861 0 dm1 AREA=2.092e-06
D861 n862 0 dm1 AREA=2.075e-06
D862 n863 0 dm1 AREA=6.749e-07
D863 n864 0 dm1 AREA=1.304e-06
D864 n865 0 dm1 AREA=8.745e-07
D865 n866 0 dm1 AREA=1.672e-06
D866 n867 0 dm1 AREA=1.071e-06
D867 n868 0 dm1 AREA=2.817e-07
D868 n869 0 dm1 AREA=7.103e-07
D869 n870 0 dm1 AREA=1.391e-06
D870 n871 0 dm1 AREA=1.427e-06
D871 n872 0 dm1 AREA=6.206e-07
D872 n873 0 dm1 AREA=6.815e-07
D873 n874 0 dm1 AREA=1.925e-06
D874 n875 0 dm1 AREA=1.044e-06
D875 n876 0 dm1 AREA=1.427e-06
D876 n877 0 dm1 AREA=5.266e-07
D877 n878 0 dm1 AREA=9.314e-07
D878 n879 0 dm1 AREA=1.726e-06
D879 n880 0 dm1 AREA=6.483e-07
D880 n881 0 dm1 AREA=4.396e-07
D881 n882 0 dm1 AREA=1.986e-06
D882 n883 0 dm1 AREA=5.710e-07
D883 n884 0 dm1 AREA=9.865e-07
D884 n885 0 dm1 AREA=1.026e-06
D885 n886 0 dm1 AREA=1.249e-06
D886 n887 0 dm1 AREA=7.298e-07
D887 n888 0 dm1 AREA=4.309e-07
D888 n889 0 dm1 AREA=2.308e-06
D889 n890 0 dm1 AREA=5.330e-07
D890 n891 0 dm1 AREA=8.695e-07
D891 n892 0 dm1 AREA=7.167e-07
D892 n893 0 dm1 AREA=1.016e-06
D893 n894 0 dm1 AREA=8.941e-07
D894 n895 0 dm1 AREA=7.573e-07
D895 n896 0 dm1 AREA=4.494e-07
D896 n897 0 dm1 AREA=8.369e-07
D897 n1 0 dm1 AREA=3.474e-07
D898 n899 0 dm1 AREA=4.221e-07
D899 n900 0 dm1 AREA=8.044e-07
D900 n901 0 dm1 AREA=2.745e-06
D901 n902 0 dm1 AREA=6.682e-07
D902 n903 0 dm1 AREA=5.532e-07
D903 n904 0 dm1 AREA=1.791e-06
D904 n905 0 dm1 AREA=2.092e-06
D905 n906 0 dm1 AREA=8.343e-07
D906 n907 0 dm1 AREA=1.247e-06
D907 n908 0 dm1 AREA=1.603e-06
D908 n909 0 dm1 AREA=4.201e-07
D909 n910 0 dm1 AREA=6.467e-07
D910 n911 0 dm1 AREA=1.276e-06
D911 n912 0 dm1 AREA=2.583e-07
D912 n913 0 dm1 AREA=5.773e-07
D913 n914 0 dm1 AREA=8.539e-07
D914 n915 0 dm1 AREA=1.703e-06
D915 n916 0 dm1 AREA=4.126e-07
D916 n917 0 dm1 AREA=6.244e-07
D917 n918 0 dm1 AREA=1.805e-06
D918 n919 0 dm1 AREA=6.465e-07
D919 n920 0 dm1 AREA=8.689e-07
D920 n921 0 dm1 AREA=1.794e-06
D921 n922 0 dm1 AREA=1.821e-06
D922 n923 0 dm1 AREA=5.181e-07
D923 n924 0 dm1 AREA=7.770e-07
D924 n925 0 dm1 AREA=5.572e-07
D925 n926 0 dm1 AREA=1.186e-06
D926 n927 0 dm1 AREA=4.811e-07
D927 n928 0 dm1 AREA=5.656e-07
D928 n929 0 dm1 AREA=2.113e-07
D929 n930 0 dm1 AREA=1.283e-06
D930 n931 0 dm1 AREA=7.515e-07
D931 n932 0 dm1 AREA=1.894e-06
D932 n933 0 dm1 AREA=3.893e-07
D933 n934 0 dm1 AREA=1.885e-06
D934 n935 0 dm1 AREA=1.004e-06
D935 n936 0 dm1 AREA=1.174e-07
D936 n937 0 dm1 AREA=8.418e-07
D937 n938 0 dm1 AREA=1.972e-06
D938 n939 0 dm1 AREA=1.454e-06
D939 n940 0 dm1 AREA=6.385e-07
D940 n941 0 dm1 AREA=4.262e-07
D941 n942 0 dm1 AREA=2.533e-07
D942 n943 0 dm1 AREA=3.632e-07
D943 n944 0 dm1 AREA=3.034e-06
D944 n945 0 dm1 AREA=5.936e-07
D945 n946 0 dm1 AREA=1.266e-06
D946 n947 0 dm1 AREA=5.694e-07
D947 n948 0 dm1 AREA=6.230e-07
D948 n949 0 dm1 AREA=9.865e-07
D949 n950 0 dm1 AREA=6.750e-07
D950 n951 0 dm1 AREA=1.849e-06
D951 n952 0 dm1 AREA=4.723e-07
D952 n953 0 dm1 AREA=4.261e-07
D953 n954 0 dm1 AREA=7.252e-07
D954 n955 0 dm1 AREA=6.333e-07
D955 n956 0 dm1 AREA=7.875e-07
D956 n957 0 dm1 AREA=1.393e-06
D957 n958 0 dm1 AREA=1.471e-06
D958 n959 0 dm1 AREA=4.816e-07
D959 n960 0 dm1 AREA=9.772e-07
D960 n961 0 dm1 AREA=9.283e-07
D961 n962 0 dm1 AREA=1.130e-06
D962 n963 0 dm1 AREA=7.910e-07
D963 n964 0 dm1 AREA=1.520e-06
D964 n965 0 dm1 AREA=7.043e-07
D965 n966 0 dm1 AREA=1.570e-06
D966 n967 0 dm1 AREA=4.621e-07
D967 n968 0 dm1 AREA=1.207e-06
D968 n969 0 dm1 AREA=9.323e-07
D969 n970 0 dm1 AREA=3.421e-06
D970 n971 0 dm1 AREA=7.537e-07
D971 n972 0 dm1 AREA=8.525e-07
D972 n973 0 dm1 AREA=1.162e-06
D973 n974 0 dm1 AREA=1.139e-06
D974 n975 0 dm1 AREA=1.602e-06
D975 n976 0 dm1 AREA=4.875e-07
D976 n977 0 dm1 AREA=9.979e-07
D977 n978 0 dm1 AREA=2.139e-06
D978 n979 0 dm1 AREA=5.706e-07
D979 n980 0 dm1 AREA=4.605e-07
D980 n981 0 dm1 AREA=3.420e-07
D981 n982 0 dm1 AREA=1.517e-06
D982 n983 0 dm1 AREA=2.095e-06
D983 n984 0 dm1 AREA=6.055e-07
D984 n985 0 dm1 AREA=9.141e-07
D985 n986 0 dm1 AREA=1.347e-06
D986 n987 0 dm1 AREA=1.205e-07
D987 n988 0 dm1 AREA=1.856e-06
D988 n989 0 dm1 AREA=3.983e-07
D989 n990 0 dm1 AREA=4.008e-07
D990 n991 0 dm1 AREA=1.597e-06
D991 n992 0 dm1 AREA=1.200e-06
D992 n993 0 dm1 AREA=8.942e-07
D993 n994 0 dm1 AREA=9.340e-07
D994 n995 0 dm1 AREA=7.421e-07
D995 n996 0 dm1 AREA=8.892e-07
D996 n997 0 dm1 AREA=7.726e-07
D997 n998 0 dm1 AREA=1.198e-06
D998 n999 0 dm1 AREA=1.302e-06
D999 n1000 0 dm1 AREA=1.729e-06
D1000 n1001 0 dm1 AREA=1.284e-06
D1001 n1002 0 dm1 AREA=5.222e-07
D1002 n1003 0 dm1 AREA=4.123e-07
D1003 n1004 0 dm1 AREA=8.629e-07
D1004 n1005 0 dm1 AREA=7.233e-07
D1005 n1006 0 dm1 AREA=1.454e-06
D1006 n1007 0 dm1 AREA=4.087e-07
D1007 n1008 0 dm1 AREA=5.867e-07
D1008 n1009 0 dm1 AREA=1.072e-06
D1009 n1010 0 dm1 AREA=1.232e-06
D1010 n1011 0 dm1 AREA=7.836e-07
D1011 n1012 0 dm1 AREA=2.219e-07
D1012 n1013 0 dm1 AREA=1.337e-06
D1013 n1014 0 dm1 AREA=6.436e-07
D1014 n1015 0 dm1 AREA=1.038e-06
D1015 n1016 0 dm1 AREA=5.271e-07
D1016 n1017 0 dm1 AREA=8.883e-07
D1017 n1018 0 dm1 AREA=6.726e-07
D1018 n1019 0 dm1 AREA=4.937e-07
D1019 n1020 0 dm1 AREA=9.001e-07
D1020 n1021 0 dm1 AREA=2.020e-06
D1021 n1022 0 dm1 AREA=5.327e-07
D1022 n1023 0 dm1 AREA=4.563e-07
D1023 n1024 0 dm1 AREA=1.484e-06
D1024 n1025 0 dm1 AREA=8.412e-07
D1025 n1026 0 dm1 AREA=1.425e-06
D1026 n1027 0 dm1 AREA=9.694e-07
D1027 n1028 0 dm1 AREA=4.368e-07
D1028 n1029 0 dm1 AREA=4.314e-07
D1029 n1030 0 dm1 AREA=5.495e-07
D1030 n1031 0 dm1 AREA=1.402e-06
D1031 n1032 0 dm1 AREA=3.140e-07
D1032 n1033 0 dm1 AREA=6.079e-07
D1033 n1034 0 dm1 AREA=3.358e-07
D1034 n1035 0 dm1 AREA=9.251e-07
D1035 n1036 0 dm1 AREA=9.467e-07
D1036 n1037 0 dm1 AREA=9.816e-07
D1037 n1038 0 dm1 AREA=2.402e-07
D1038 n1039 0 dm1 AREA=9.594e-07
D1039 n1040 0 dm1 AREA=8.810e-07
D1040 n1041 0 dm1 AREA=1.001e-06
D1041 n1042 0 dm1 AREA=1.579e-06
D1042 n1043 0 dm1 AREA=4.856e-07
D1043 n1044 0 dm1 AREA=1.007e-06
D1044 n1045 0 dm1 AREA=7.230e-07
D1045 n1046 0 dm1 AREA=6.866e-07
D1046 n1047 0 dm1 AREA=1.012e-06
D1047 n1048 0 dm1 AREA=1.467e-06
D1048 n1049 0 dm1 AREA=5.830e-07
D1049 n1050 0 dm1 AREA=7.527e-07
D1050 n1051 0 dm1 AREA=6.642e-07
D1051 n1052 0 dm1 AREA=5.666e-07
D1052 n1053 0 dm1 AREA=9.839e-07
D1053 n1054 0 dm1 AREA=1.556e-06
D1054 n1055 0 dm1 AREA=5.277e-07
D1055 n1056 0 dm1 AREA=1.248e-06
D1056 n1057 0 dm1 AREA=1.159e-06
D1057 n1058 0 dm1 AREA=2.892e-07
D1058 n1059 0 dm1 AREA=3.389e-07
D1059 n1060 0 dm1 AREA=4.291e-07
D1060 n1061 0 dm1 AREA=5.826e-07
D1061 n1062 0 dm1 AREA=1.196e-06
D1062 n1063 0 dm1 AREA=3.238e-07
D1063 n1064 0 dm1 AREA=1.000e-06
D1064 n1065 0 dm1 AREA=1.679e-07
D1065 n1066 0 dm1 AREA=1.662e-06
D1066 n1067 0 dm1 AREA=1.260e-06
D1067 n1068 0 dm1 AREA=2.223e-06
D1068 n1069 0 dm1 AREA=4.112e-07
D1069 n1070 0 dm1 AREA=2.479e-07
D1070 n1071 0 dm1 AREA=1.118e-06
D1071 n1072 0 dm1 AREA=6.374e-07
D1072 n1073 0 dm1 AREA=8.490e-07
D1073 n1074 0 dm1 AREA=1.363e-06
D1074 n1075 0 dm1 AREA=8.383e-07
D1075 n1076 0 dm1 AREA=1.312e-06
D1076 n1077 0 dm1 AREA=8.454e-07
D1077 n1078 0 dm1 AREA=9.880e-07
D1078 n1079 0 dm1 AREA=6.704e-07
D1079 n1080 0 dm1 AREA=1.256e-06
D1080 n1081 0 dm1 AREA=5.184e-07
D1081 n1082 0 dm1 AREA=7.780e-07
D1082 n1083 0 dm1 AREA=1.457e-06
D1083 n1084 0 dm1 AREA=9.524e-07
D1084 n1085 0 dm1 AREA=1.620e-06
D1085 n1086 0 dm1 AREA=4.643e-07
D1086 n1087 0 dm1 AREA=3.534e-07
D1087 n1088 0 dm1 AREA=2.927e-06
D1088 n1089 0 dm1 AREA=9.416e-07
D1089 n1090 0 dm1 AREA=7.030e-07
D1090 n1091 0 dm1 AREA=1.343e-06
D1091 n1092 0 dm1 AREA=5.547e-07
D1092 n1093 0 dm1 AREA=1.104e-06
D1093 n1094 0 dm1 AREA=4.889e-07
D1094 n1095 0 dm1 AREA=1.405e-06
D1095 n1096 0 dm1 AREA=1.881e-06
D1096 n1097 0 dm1 AREA=1.346e-06
D1097 n1098 0 dm1 AREA=4.977e-07
D1098 n1099 0 dm1 AREA=1.340e-06
D1099 n1100 0 dm1 AREA=9.670e-07
D1100 n1101 0 dm1 AREA=5.549e-07
D1101 n1102 0 dm1 AREA=1.047e-06
D1102 n1103 0 dm1 AREA=3.417e-07
D1103 n1104 0 dm1 AREA=2.496e-07
D1104 n1105 0 dm1 AREA=9.603e-07
D1105 n1106 0 dm1 AREA=8.420e-07
D1106 n1107 0 dm1 AREA=7.632e-07
D1107 n1108 0 dm1 AREA=6.593e-07
D1108 n1109 0 dm1 AREA=1.149e-06
D1109 n1110 0 dm1 AREA=9.321e-07
D1110 n1111 0 dm1 AREA=9.308e-07
D1111 n1112 0 dm1 AREA=5.469e-07
D1112 n1113 0 dm1 AREA=4.603e-07
D1113 n1114 0 dm1 AREA=1.602e-06
D1114 n1115 0 dm1 AREA=7.956e-07
D1115 n1116 0 dm1 AREA=1.039e-06
D1116 n1117 0 dm1 AREA=6.046e-07
D1117 n1118 0 dm1 AREA=6.844e-07
D1118 n1119 0 dm1 AREA=1.054e-06
D1119 n1120 0 dm1 AREA=1.216e-06
D1120 n1121 0 dm1 AREA=1.002e-06
D1121 n1122 0 dm1 AREA=1.671e-06
D1122 n1123 0 dm1 AREA=1.216e-06
D1123 n1124 0 dm1 AREA=1.888e-06
D1124 n1125 0 dm1 AREA=5.609e-07
D1125 n1126 0 dm1 AREA=6.535e-07
D1126 n1127 0 dm1 AREA=8.262e-07
D1127 n1128 0 dm1 AREA=7.725e-07
D1128 n1129 0 dm1 AREA=1.012e-06
D1129 n1130 0 dm1 AREA=1.503e-07
D1130 n1131 0 dm1 AREA=1.233e-06
D1131 n1132 0 dm1 AREA=6.558e-07
D1132 n1133 0 dm1 AREA=4.904e-07
D1133 n1134 0 dm1 AREA=1.348e-07
D1134 n1135 0 dm1 AREA=5.693e-07
D1135 n1136 0 dm1 AREA=1.921e-06
D1136 n1137 0 dm1 AREA=6.643e-07
D1137 n1138 0 dm1 AREA=1.544e-06
D1138 n1139 0 dm1 AREA=2.000e-06
D1139 n1140 0 dm1 AREA=9.005e-07
D1140 n1141 0 dm1 AREA=1.078e-06
D1141 n1142 0 dm1 AREA=5.338e-07
D1142 n1143 0 dm1 AREA=1.645e-06
D1143 n1144 0 dm1 AREA=5.375e-07
D1144 n1145 0 dm1 AREA=1.101e-06
D1145 n1146 0 dm1 AREA=5.534e-07
D1146 n1147 0 dm1 AREA=9.812e-07
D1147 n1148 0 dm1 AREA=5.272e-07
D1148 n1149 0 dm1 AREA=1.079e-06
D1149 n1150 0 dm1 AREA=1.069e-06
D1150 n1151 0 dm1 AREA=1.024e-06
D1151 n1152 0 dm1 AREA=1.674e-06
D1152 n1153 0 dm1 AREA=6.382e-07
D1153 n1154 0 dm1 AREA=1.262e-06
D1154 n1 0 dm1 AREA=1.467e-07
D1155 n1156 0 dm1 AREA=3.325e-07
D1156 n1157 0 dm1 AREA=2.280e-06
D1157 n1158 0 dm1 AREA=3.235e-07
D1158 n1159 0 dm1 AREA=6.261e-07
D1159 n1160 0 dm1 AREA=4.874e-07
D1160 n1161 0 dm1 AREA=1.195e-06
D1161 n1162 0 dm1 AREA=2.748e-07
D1162 n1163 0 dm1 AREA=1.147e-06
D1163 n1164 0 dm1 AREA=9.839e-07
D1164 n1165 0 dm1 AREA=8.702e-07
D1165 n1166 0 dm1 AREA=1.089e-06
D1166 n1167 0 dm1 AREA=1.753e-06
D1167 n1168 0 dm1 AREA=1.059e-06
D1168 n1169 0 dm1 AREA=5.824e-07
D1169 n1170 0 dm1 AREA=5.200e-07
D1170 n1171 0 dm1 AREA=4.780e-07
D1171 n1172 0 dm1 AREA=6.333e-07
D1172 n1173 0 dm1 AREA=6.107e-07
D1173 n1174 0 dm1 AREA=1.589e-06
D1174 n1175 0 dm1 AREA=3.762e-07
D1175 n1176 0 dm1 AREA=6.843e-07
D1176 n1177 0 dm1 AREA=1.946e-06
D1177 n1178 0 dm1 AREA=1.198e-06
D1178 n1179 0 dm1 AREA=1.049e-06
D1179 n1 0 dm1 AREA=1.754e-07
D1180 n1181 0 dm1 AREA=1.066e-06
D1181 n1182 0 dm1 AREA=2.980e-06
D1182 n1183 0 dm1 AREA=6.420e-07
D1183 n1184 0 dm1 AREA=1.789e-06
D1184 n1185 0 dm1 AREA=6.495e-07
D1185 n1186 0 dm1 AREA=1.157e-06
D1186 n1187 0 dm1 AREA=3.745e-06
D1187 n1188 0 dm1 AREA=1.505e-06
D1188 n1189 0 dm1 AREA=7.910e-07
D1189 n1190 0 dm1 AREA=3.087e-07
D1190 n1191 0 dm1 AREA=9.167e-07
D1191 n1192 0 dm1 AREA=1.443e-06
D1192 n1193 0 dm1 AREA=9.274e-07
D1193 n1194 0 dm1 AREA=8.541e-07
D1194 n1195 0 dm1 AREA=1.803e-06
D1195 n1196 0 dm1 AREA=9.266e-07
D1196 n1197 0 dm1 AREA=9.330e-07
D1197 n1198 0 dm1 AREA=7.810e-07
D1198 n1199 0 dm1 AREA=1.517e-06
D1199 n1200 0 dm1 AREA=6.532e-07
D1200 n1201 0 dm1 AREA=9.095e-07
D1201 n1 0 dm1 AREA=7.429e-07
D1202 n1203 0 dm1 AREA=1.222e-06
D1203 n1204 0 dm1 AREA=3.085e-07
D1204 n1205 0 dm1 AREA=6.816e-07
D1205 n1206 0 dm1 AREA=1.046e-06
D1206 n1207 0 dm1 AREA=1.549e-06
D1207 n1208 0 dm1 AREA=4.001e-07
D1208 n1209 0 dm1 AREA=3.081e-07
D1209 n1210 0 dm1 AREA=1.452e-06
D1210 n1211 0 dm1 AREA=4.018e-07
D1211 n1212 0 dm1 AREA=8.383e-07
D1212 n1213 0 dm1 AREA=1.097e-06
D1213 n1214 0 dm1 AREA=5.261e-07
D1214 n1215 0 dm1 AREA=1.340e-06
D1215 n1216 0 dm1 AREA=8.519e-07
D1216 n1217 0 dm1 AREA=5.907e-07
D1217 n1218 0 dm1 AREA=4.965e-07
D1218 n1219 0 dm1 AREA=1.076e-06
D1219 n1220 0 dm1 AREA=9.905e-07
D1220 n1221 0 dm1 AREA=1.373e-06
D1221 n1222 0 dm1 AREA=9.037e-07
D1222 n1223 0 dm1 AREA=1.445e-06
D1223 n1224 0 dm1 AREA=1.089e-06
D1224 n1225 0 dm1 AREA=2.026e-06
D1225 n1226 0 dm1 AREA=6.371e-07
D1226 n1227 0 dm1 AREA=1.102e-06
D1227 n1228 0 dm1 AREA=1.423e-06
D1228 n1229 0 dm1 AREA=6.930e-07
D1229 n1230 0 dm1 AREA=5.410e-07
D1230 n1231 0 dm1 AREA=1.181e-06
D1231 n1232 0 dm1 AREA=7.902e-07
D1232 n1233 0 dm1 AREA=1.906e-06
D1233 n1234 0 dm1 AREA=1.627e-06
D1234 n1235 0 dm1 AREA=9.834e-07
D1235 n1236 0 dm1 AREA=7.134e-07
D1236 n1237 0 dm1 AREA=5.238e-07
D1237 n1238 0 dm1 AREA=1.039e-06
D1238 n1239 0 dm1 AREA=4.796e-07
D1239 n1240 0 dm1 AREA=1.231e-06
D1240 n1241 0 dm1 AREA=2.033e-06
D1241 n1242 0 dm1 AREA=1.468e-06
D1242 n1243 0 dm1 AREA=1.187e-06
D1243 n1244 0 dm1 AREA=8.674e-07
D1244 n1245 0 dm1 AREA=1.402e-06
D1245 n1246 0 dm1 AREA=4.845e-07
D1246 n1247 0 dm1 AREA=2.072e-06
D1247 n1248 0 dm1 AREA=1.837e-06
D1248 n1249 0 dm1 AREA=1.429e-06
D1249 n1250 0 dm1 AREA=1.072e-06
D1250 n1251 0 dm1 AREA=2.997e-06
D1251 n1252 0 dm1 AREA=9.704e-07
D1252 n1253 0 dm1 AREA=2.445e-06
D1253 n1254 0 dm1 AREA=5.237e-07
D1254 n1255 0 dm1 AREA=5.501e-07
D1255 n1256 0 dm1 AREA=7.598e-07
D1256 n1257 0 dm1 AREA=3.154e-07
D1257 n1258 0 dm1 AREA=1.677e-06
D1258 n1259 0 dm1 AREA=5.373e-07
D1259 n1260 0 dm1 AREA=2.585e-06
D1260 n1261 0 dm1 AREA=9.400e-07
D1261 n1262 0 dm1 AREA=1.394e-06
D1262 n1263 0 dm1 AREA=6.791e-07
D1263 n1264 0 dm1 AREA=1.149e-06
D1264 n1265 0 dm1 AREA=1.494e-06
D1265 n1266 0 dm1 AREA=1.845e-06
D1266 n1267 0 dm1 AREA=4.265e-07
D1267 n1268 0 dm1 AREA=5.703e-07
D1268 n1269 0 dm1 AREA=6.306e-07
D1269 n1270 0 dm1 AREA=1.273e-06
D1270 n1271 0 dm1 AREA=9.577e-07
D1271 n1 0 dm1 AREA=1.202e-06
D1272 n1273 0 dm1 AREA=7.172e-07
D1273 n1 0 dm1 AREA=1.467e-06
D1274 n1275 0 dm1 AREA=6.894e-07
D1275 n1276 0 dm1 AREA=5.128e-07
D1276 n1277 0 dm1 AREA=6.178e-07
D1277 n1278 0 dm1 AREA=1.030e-06
D1278 n1279 0 dm1 AREA=1.459e-06
D1279 n1280 0 dm1 AREA=1.112e-06
D1280 n1281 0 dm1 AREA=5.704e-07
D1281 n1282 0 dm1 AREA=9.410e-07
D1282 n1283 0 dm1 AREA=5.494e-07
D1283 n1284 0 dm1 AREA=3.777e-07
D1284 n1285 0 dm1 AREA=8.725e-07
D1285 n1286 0 dm1 AREA=8.546e-07
D1286 n1287 0 dm1 AREA=9.583e-07
D1287 n1288 0 dm1 AREA=8.806e-07
D1288 n1289 0 dm1 AREA=1.037e-06
D1289 n1290 0 dm1 AREA=1.736e-06
D1290 n1291 0 dm1 AREA=8.460e-07
D1291 n1292 0 dm1 AREA=1.094e-06
D1292 n1293 0 dm1 AREA=2.990e-07
D1293 n1294 0 dm1 AREA=3.277e-06
D1294 n1295 0 dm1 AREA=8.789e-07
D1295 n1296 0 dm1 AREA=7.119e-07
D1296 n1297 0 dm1 AREA=2.204e-07
D1297 n1298 0 dm1 AREA=5.487e-07
D1298 n1299 0 dm1 AREA=2.187e-06
D1299 n1300 0 dm1 AREA=8.579e-07
D1300 n1301 0 dm1 AREA=4.424e-07
D1301 n1302 0 dm1 AREA=1.099e-06
D1302 n1303 0 dm1 AREA=1.027e-06
D1303 n1304 0 dm1 AREA=9.992e-07
D1304 n1305 0 dm1 AREA=3.724e-07
D1305 n1306 0 dm1 AREA=6.971e-07
D1306 n1307 0 dm1 AREA=6.495e-07
D1307 n1308 0 dm1 AREA=1.654e-06
D1308 n1309 0 dm1 AREA=7.685e-07
D1309 n1310 0 dm1 AREA=2.753e-07
D1310 n1311 0 dm1 AREA=6.639e-07
D1311 n1312 0 dm1 AREA=1.112e-06
D1312 n1313 0 dm1 AREA=9.638e-07
D1313 n1314 0 dm1 AREA=1.336e-06
D1314 n1315 0 dm1 AREA=9.499e-07
D1315 n1316 0 dm1 AREA=7.674e-07
D1316 n1317 0 dm1 AREA=1.118e-06
D1317 n1318 0 dm1 AREA=6.136e-07
D1318 n1319 0 dm1 AREA=8.260e-07
D1319 n1320 0 dm1 AREA=5.301e-07
D1320 n1321 0 dm1 AREA=1.634e-06
D1321 n1322 0 dm1 AREA=1.078e-06
D1322 n1 0 dm1 AREA=8.366e-07
D1323 n1324 0 dm1 AREA=9.161e-07
D1324 n1325 0 dm1 AREA=5.830e-07
D1325 n1326 0 dm1 AREA=7.678e-07
D1326 n1327 0 dm1 AREA=1.152e-06
D1327 n1328 0 dm1 AREA=5.169e-07
D1328 n1329 0 dm1 AREA=1.268e-06
D1329 n1330 0 dm1 AREA=1.589e-06
D1330 n1331 0 dm1 AREA=5.159e-07
D1331 n1332 0 dm1 AREA=1.541e-06
D1332 n1333 0 dm1 AREA=5.760e-07
D1333 n1334 0 dm1 AREA=1.636e-06
D1334 n1335 0 dm1 AREA=6.405e-07
D1335 n1336 0 dm1 AREA=1.263e-06
D1336 n1337 0 dm1 AREA=3.747e-07
D1337 n1338 0 dm1 AREA=1.078e-06
D1338 n1339 0 dm1 AREA=4.879e-07
D1339 n1340 0 dm1 AREA=5.668e-07
D1340 n1341 0 dm1 AREA=6.375e-07
D1341 n1342 0 dm1 AREA=1.525e-06
D1342 n1343 0 dm1 AREA=5.264e-07
D1343 n1344 0 dm1 AREA=1.118e-06
D1344 n1345 0 dm1 AREA=1.133e-06
D1345 n1346 0 dm1 AREA=1.223e-06
D1346 n1347 0 dm1 AREA=9.810e-07
D1347 n1348 0 dm1 AREA=2.095e-07
D1348 n1349 0 dm1 AREA=1.405e-06
D1349 n1350 0 dm1 AREA=1.018e-06
D1350 n1351 0 dm1 AREA=8.551e-07
D1351 n1352 0 dm1 AREA=7.011e-07
D1352 n1353 0 dm1 AREA=1.951e-07
D1353 n1354 0 dm1 AREA=2.472e-06
D1354 n1355 0 dm1 AREA=1.340e-06
D1355 n1356 0 dm1 AREA=5.189e-07
D1356 n1357 0 dm1 AREA=1.393e-06
D1357 n1358 0 dm1 AREA=4.310e-07
D1358 n1359 0 dm1 AREA=6.278e-07
D1359 n1360 0 dm1 AREA=1.474e-06
D1360 n1361 0 dm1 AREA=1.389e-06
D1361 n1362 0 dm1 AREA=1.314e-06
D1362 n1363 0 dm1 AREA=2.150e-07
D1363 n1364 0 dm1 AREA=9.767e-07
D1364 n1365 0 dm1 AREA=1.025e-06
D1365 n1366 0 dm1 AREA=1.153e-06
D1366 n1367 0 dm1 AREA=9.387e-07
D1367 n1368 0 dm1 AREA=1.071e-06
D1368 n1369 0 dm1 AREA=6.779e-07
D1369 n1370 0 dm1 AREA=4.364e-07
D1370 n1371 0 dm1 AREA=2.038e-06
D1371 n1372 0 dm1 AREA=5.232e-07
D1372 n1373 0 dm1 AREA=9.390e-07
D1373 n1374 0 dm1 AREA=1.048e-06
D1374 n1375 0 dm1 AREA=1.848e-06
D1375 n1376 0 dm1 AREA=9.124e-07
D1376 n1377 0 dm1 AREA=3.800e-07
D1377 n1378 0 dm1 AREA=5.474e-07
D1378 n1379 0 dm1 AREA=6.509e-07
D1379 n1380 0 dm1 AREA=6.121e-07
D1380 n1381 0 dm1 AREA=1.382e-06
D1381 n1382 0 dm1 AREA=1.841e-06
D1382 n1383 0 dm1 AREA=1.845e-06
D1383 n1384 0 dm1 AREA=1.273e-06
D1384 n1385 0 dm1 AREA=1.008e-06
D1385 n1386 0 dm1 AREA=8.960e-07
D1386 n1387 0 dm1 AREA=6.383e-07
D1387 n1388 0 dm1 AREA=8.634e-07
D1388 n1389 0 dm1 AREA=6.428e-07
D1389 n1390 0 dm1 AREA=1.337e-06
D1390 n1391 0 dm1 AREA=1.438e-06
D1391 n1392 0 dm1 AREA=1.274e-06
D1392 n1393 0 dm1 AREA=1.400e-06
D1393 n1394 0 dm1 AREA=2.447e-06
D1394 n1395 0 dm1 AREA=3.376e-07
D1395 n1396 0 dm1 AREA=1.658e-06
D1396 n1397 0 dm1 AREA=4.320e-07
D1397 n1398 0 dm1 AREA=2.145e-07
D1398 n1399 0 dm1 AREA=3.584e-07
D1399 n1400 0 dm1 AREA=3.593e-07
D1400 n1401 0 dm1 AREA=1.448e-06
D1401 n1402 0 dm1 AREA=1.679e-07
D1402 n1403 0 dm1 AREA=9.943e-07
D1403 n1404 0 dm1 AREA=6.620e-07
D1404 n1405 0 dm1 AREA=1.620e-06
D1405 n1406 0 dm1 AREA=8.143e-07
D1406 n1407 0 dm1 AREA=1.284e-06
D1407 n1408 0 dm1 AREA=8.231e-07
D1408 n1409 0 dm1 AREA=1.554e-06
D1409 n1410 0 dm1 AREA=2.068e-06
D1410 n1411 0 dm1 AREA=6.382e-07
D1411 n1412 0 dm1 AREA=4.692e-07
D1412 n1413 0 dm1 AREA=1.344e-06
D1413 n1414 0 dm1 AREA=8.122e-07
D1414 n1415 0 dm1 AREA=7.427e-07
D1415 n1416 0 dm1 AREA=1.848e-06
D1416 n1417 0 dm1 AREA=1.176e-06
D1417 n1418 0 dm1 AREA=1.085e-06
D1418 n1419 0 dm1 AREA=5.629e-07
D1419 n1420 0 dm1 AREA=2.393e-07
D1420 n1421 0 dm1 AREA=1.366e-06
D1421 n1422 0 dm1 AREA=1.650e-06
D1422 n1423 0 dm1 AREA=5.174e-07
D1423 n1424 0 dm1 AREA=1.771e-06
D1424 n1425 0 dm1 AREA=5.781e-07
D1425 n1426 0 dm1 AREA=2.063e-07
D1426 n1427 0 dm1 AREA=4.956e-07
D1427 n1428 0 dm1 AREA=1.519e-06
D1428 n1429 0 dm1 AREA=4.957e-07
D1429 n1430 0 dm1 AREA=4.583e-07
D1430 n1431 0 dm1 AREA=1.300e-06
D1431 n1432 0 dm1 AREA=4.333e-07
D1432 n1433 0 dm1 AREA=5.188e-07
D1433 n1434 0 dm1 AREA=2.466e-06
D1434 n1435 0 dm1 AREA=8.620e-07
D1435 n1436 0 dm1 AREA=9.649e-07
D1436 n1437 0 dm1 AREA=5.923e-07
D1437 n1438 0 dm1 AREA=1.521e-06
D1438 n1439 0 dm1 AREA=5.792e-07
D1439 n1440 0 dm1 AREA=1.517e-06
D1440 n1441 0 dm1 AREA=9.445e-07
D1441 n1442 0 dm1 AREA=4.794e-07
D1442 n1443 0 dm1 AREA=1.693e-06
D1443 n1444 0 dm1 AREA=2.112e-06
D1444 n1445 0 dm1 AREA=2.636e-06
D1445 n1446 0 dm1 AREA=6.804e-07
D1446 n1447 0 dm1 AREA=7.208e-07
D1447 n1448 0 dm1 AREA=7.877e-07
D1448 n1449 0 dm1 AREA=8.382e-07
D1449 n1450 0 dm1 AREA=1.134e-06
D1450 n1451 0 dm1 AREA=1.611e-06
D1451 n1452 0 dm1 AREA=1.241e-06
D1452 n1453 0 dm1 AREA=4.432e-07
D1453 n1454 0 dm1 AREA=1.787e-07
D1454 n1455 0 dm1 AREA=1.588e-06
D1455 n1456 0 dm1 AREA=7.620e-07
D1456 n1457 0 dm1 AREA=9.841e-07
D1457 n1458 0 dm1 AREA=1.817e-06
D1458 n1459 0 dm1 AREA=1.642e-06
D1459 n1460 0 dm1 AREA=9.306e-07
D1460 n1461 0 dm1 AREA=3.214e-07
D1461 n1462 0 dm1 AREA=1.567e-06
D1462 n1463 0 dm1 AREA=5.108e-07
D1463 n1464 0 dm1 AREA=6.833e-07
D1464 n1465 0 dm1 AREA=5.559e-07
D1465 n1466 0 dm1 AREA=1.508e-06
D1466 n1467 0 dm1 AREA=2.585e-06
D1467 n1468 0 dm1 AREA=1.476e-06
D1468 n1469 0 dm1 AREA=2.525e-07
D1469 n1470 0 dm1 AREA=7.834e-07
D1470 n1471 0 dm1 AREA=1.247e-06
D1471 n1472 0 dm1 AREA=8.702e-07
D1472 n1473 0 dm1 AREA=6.867e-07
D1473 n1474 0 dm1 AREA=4.001e-07
D1474 n1475 0 dm1 AREA=2.025e-06
D1475 n1476 0 dm1 AREA=1.834e-06
D1476 n1477 0 dm1 AREA=1.915e-06
D1477 n1478 0 dm1 AREA=2.319e-06
D1478 n1479 0 dm1 AREA=6.918e-07
D1479 n1480 0 dm1 AREA=5.841e-07
D1480 n1481 0 dm1 AREA=7.324e-07
D1481 n1482 0 dm1 AREA=4.942e-07
D1482 n1483 0 dm1 AREA=4.433e-07
D1483 n1484 0 dm1 AREA=8.009e-07
D1484 n1 0 dm1 AREA=2.441e-06
D1485 n1486 0 dm1 AREA=1.522e-06
D1486 n1487 0 dm1 AREA=1.151e-06
D1487 n1488 0 dm1 AREA=1.370e-06
D1488 n1489 0 dm1 AREA=6.660e-07
D1489 n1490 0 dm1 AREA=7.215e-07
D1490 n1491 0 dm1 AREA=9.714e-07
D1491 n1492 0 dm1 AREA=7.258e-08
D1492 n1493 0 dm1 AREA=1.252e-06
D1493 n1494 0 dm1 AREA=6.670e-07
D1494 n1495 0 dm1 AREA=1.106e-06
D1495 n1496 0 dm1 AREA=3.938e-07
D1496 n1497 0 dm1 AREA=8.470e-07
D1497 n1498 0 dm1 AREA=6.571e-07
D1498 n1499 0 dm1 AREA=1.482e-07
D1499 n1500 0 dm1 AREA=3.626e-07
D1500 n1501 0 dm1 AREA=1.443e-06
D1501 n1502 0 dm1 AREA=2.580e-07
D1502 n1503 0 dm1 AREA=1.633e-06
D1503 n1504 0 dm1 AREA=4.322e-07
D1504 n1505 0 dm1 AREA=3.472e-07
D1505 n1506 0 dm1 AREA=1.051e-06
D1506 n1507 0 dm1 AREA=8.320e-07
D1507 n1508 0 dm1 AREA=1.092e-06
D1508 n1509 0 dm1 AREA=1.177e-06
D1509 n1510 0 dm1 AREA=1.280e-06
D1510 n1511 0 dm1 AREA=2.356e-06
D1511 n1512 0 dm1 AREA=7.682e-07
D1512 n1513 0 dm1 AREA=1.136e-06
D1513 n1514 0 dm1 AREA=7.346e-07
D1514 n1515 0 dm1 AREA=1.323e-06
D1515 n1516 0 dm1 AREA=8.245e-07
D1516 n1517 0 dm1 AREA=1.191e-06
D1517 n1518 0 dm1 AREA=1.186e-06
D1518 n1519 0 dm1 AREA=1.377e-06
D1519 n1520 0 dm1 AREA=1.207e-06
D1520 n1521 0 dm1 AREA=9.599e-07
D1521 n1522 0 dm1 AREA=8.889e-07
D1522 n1523 0 dm1 AREA=4.371e-07
D1523 n1524 0 dm1 AREA=5.879e-07
D1524 n1525 0 dm1 AREA=2.363e-07
D1525 n1526 0 dm1 AREA=7.867e-07
D1526 n1527 0 dm1 AREA=1.772e-06
D1527 n1528 0 dm1 AREA=3.266e-07
D1528 n1529 0 dm1 AREA=3.685e-07
D1529 n1530 0 dm1 AREA=1.592e-06
D1530 n1531 0 dm1 AREA=5.660e-07
D1531 n1532 0 dm1 AREA=9.475e-07
D1532 n1533 0 dm1 AREA=5.495e-07
D1533 n1534 0 dm1 AREA=1.688e-06
D1534 n1535 0 dm1 AREA=5.259e-07
D1535 n1536 0 dm1 AREA=2.000e-06
D1536 n1537 0 dm1 AREA=6.422e-07
D1537 n1538 0 dm1 AREA=3.411e-07
D1538 n1539 0 dm1 AREA=1.046e-06
D1539 n1540 0 dm1 AREA=8.563e-07
D1540 n1541 0 dm1 AREA=1.542e-06
D1541 n1542 0 dm1 AREA=1.511e-06
D1542 n1543 0 dm1 AREA=1.311e-06
D1543 n1544 0 dm1 AREA=1.150e-06
D1544 n1545 0 dm1 AREA=2.770e-07
D1545 n1546 0 dm1 AREA=2.137e-06
D1546 n1547 0 dm1 AREA=4.020e-07
D1547 n1548 0 dm1 AREA=4.176e-07
D1548 n1549 0 dm1 AREA=5.471e-07
D1549 n1550 0 dm1 AREA=1.423e-06
D1550 n1551 0 dm1 AREA=6.671e-07
D1551 n1552 0 dm1 AREA=1.348e-06
D1552 n1553 0 dm1 AREA=1.624e-06
D1553 n1554 0 dm1 AREA=1.076e-06
D1554 n1555 0 dm1 AREA=8.792e-07
D1555 n1556 0 dm1 AREA=1.050e-06
D1556 n1557 0 dm1 AREA=5.171e-07
D1557 n1558 0 dm1 AREA=1.216e-06
D1558 n1559 0 dm1 AREA=7.760e-07
D1559 n1560 0 dm1 AREA=1.282e-06
D1560 n1561 0 dm1 AREA=1.700e-07
D1561 n1562 0 dm1 AREA=4.044e-07
D1562 n1563 0 dm1 AREA=3.267e-07
D1563 n1564 0 dm1 AREA=7.686e-07
D1564 n1565 0 dm1 AREA=5.320e-07
D1565 n1566 0 dm1 AREA=1.378e-06
D1566 n1567 0 dm1 AREA=1.707e-06
D1567 n1568 0 dm1 AREA=1.455e-06
D1568 n1569 0 dm1 AREA=2.792e-07
D1569 n1570 0 dm1 AREA=1.724e-06
D1570 n1571 0 dm1 AREA=5.279e-07
D1571 n1572 0 dm1 AREA=1.869e-06
D1572 n1573 0 dm1 AREA=3.975e-07
D1573 n1574 0 dm1 AREA=8.179e-07
D1574 n1575 0 dm1 AREA=1.257e-06
D1575 n1576 0 dm1 AREA=8.441e-07
D1576 n1577 0 dm1 AREA=8.631e-07
D1577 n1578 0 dm1 AREA=5.867e-07
D1578 n1579 0 dm1 AREA=1.396e-06
D1579 n1580 0 dm1 AREA=1.290e-06
D1580 n1581 0 dm1 AREA=8.227e-07
D1581 n1582 0 dm1 AREA=4.127e-07
D1582 n1583 0 dm1 AREA=1.042e-06
D1583 n1584 0 dm1 AREA=1.422e-06
D1584 n1585 0 dm1 AREA=5.237e-07
D1585 n1586 0 dm1 AREA=3.643e-07
D1586 n1587 0 dm1 AREA=6.516e-07
D1587 n1588 0 dm1 AREA=1.373e-06
D1588 n1589 0 dm1 AREA=1.645e-06
D1589 n1590 0 dm1 AREA=1.219e-06
D1590 n1591 0 dm1 AREA=3.071e-07
D1591 n1592 0 dm1 AREA=9.230e-07
D1592 n1593 0 dm1 AREA=1.356e-06
D1593 n1594 0 dm1 AREA=1.701e-06
D1594 n1595 0 dm1 AREA=2.293e-06
D1595 n1596 0 dm1 AREA=1.317e-06
D1596 n1597 0 dm1 AREA=5.399e-07
D1597 n1598 0 dm1 AREA=1.530e-06
D1598 n1599 0 dm1 AREA=2.610e-07
D1599 n1600 0 dm1 AREA=2.750e-07
D1600 n1601 0 dm1 AREA=6.347e-07
D1601 n1602 0 dm1 AREA=1.458e-06
D1602 n1603 0 dm1 AREA=1.151e-06
D1603 n1604 0 dm1 AREA=6.874e-07
D1604 n1605 0 dm1 AREA=4.000e-07
D1605 n1606 0 dm1 AREA=1.063e-06
D1606 n1607 0 dm1 AREA=5.919e-07
D1607 n1608 0 dm1 AREA=1.112e-06
D1608 n1609 0 dm1 AREA=4.463e-07
D1609 n1610 0 dm1 AREA=7.720e-07
D1610 n1611 0 dm1 AREA=8.309e-07
D1611 n1612 0 dm1 AREA=1.308e-06
D1612 n1613 0 dm1 AREA=1.858e-07
D1613 n1614 0 dm1 AREA=7.999e-07
D1614 n1615 0 dm1 AREA=4.644e-07
D1615 n1616 0 dm1 AREA=1.214e-06
D1616 n1617 0 dm1 AREA=4.887e-07
D1617 n1618 0 dm1 AREA=2.029e-06
D1618 n1619 0 dm1 AREA=7.213e-07
D1619 n1620 0 dm1 AREA=1.791e-06
D1620 n1621 0 dm1 AREA=9.214e-07
D1621 n1622 0 dm1 AREA=1.473e-06
D1622 n1623 0 dm1 AREA=5.973e-07
D1623 n1624 0 dm1 AREA=6.955e-07
D1624 n1625 0 dm1 AREA=1.976e-06
D1625 n1626 0 dm1 AREA=1.012e-06
D1626 n1627 0 dm1 AREA=9.802e-07
D1627 n1628 0 dm1 AREA=1.100e-06
D1628 n1629 0 dm1 AREA=8.828e-07
D1629 n1630 0 dm1 AREA=1.344e-06
D1630 n1631 0 dm1 AREA=1.563e-06
D1631 n1632 0 dm1 AREA=2.469e-06
D1632 n1633 0 dm1 AREA=4.903e-07
D1633 n1634 0 dm1 AREA=1.271e-06
D1634 n1635 0 dm1 AREA=2.287e-06
D1635 n1636 0 dm1 AREA=1.674e-06
D1636 n1637 0 dm1 AREA=6.028e-07
D1637 n1638 0 dm1 AREA=1.107e-06
D1638 n1639 0 dm1 AREA=7.926e-07
D1639 n1640 0 dm1 AREA=4.163e-07
D1640 n1641 0 dm1 AREA=7.916e-07
D1641 n1642 0 dm1 AREA=4.510e-07
D1642 n1643 0 dm1 AREA=9.843e-07
D1643 n1644 0 dm1 AREA=6.114e-07
D1644 n1645 0 dm1 AREA=1.208e-06
D1645 n1646 0 dm1 AREA=9.548e-07
D1646 n1647 0 dm1 AREA=6.574e-07
D1647 n1648 0 dm1 AREA=1.075e-06
D1648 n1649 0 dm1 AREA=1.077e-06
D1649 n1650 0 dm1 AREA=1.215e-06
D1650 n1651 0 dm1 AREA=1.056e-06
D1651 n1652 0 dm1 AREA=1.607e-06
D1652 n1653 0 dm1 AREA=9.603e-07
D1653 n1654 0 dm1 AREA=5.439e-07
D1654 n1655 0 dm1 AREA=9.337e-07
D1655 n1656 0 dm1 AREA=5.451e-07
D1656 n1657 0 dm1 AREA=1.646e-06
D1657 n1658 0 dm1 AREA=4.881e-07
D1658 n1659 0 dm1 AREA=6.663e-07
D1659 n1660 0 dm1 AREA=7.476e-07
D1660 n1661 0 dm1 AREA=1.675e-06
D1661 n1662 0 dm1 AREA=1.186e-06
D1662 n1663 0 dm1 AREA=6.357e-07
D1663 n1664 0 dm1 AREA=6.737e-07
D1664 n1665 0 dm1 AREA=1.154e-06
D1665 n1666 0 dm1 AREA=9.069e-07
D1666 n1667 0 dm1 AREA=3.178e-07
D1667 n1668 0 dm1 AREA=7.407e-07
D1668 n1669 0 dm1 AREA=9.807e-07
D1669 n1670 0 dm1 AREA=7.755e-07
D1670 n1671 0 dm1 AREA=4.743e-07
D1671 n1672 0 dm1 AREA=5.850e-07
D1672 n1673 0 dm1 AREA=1.202e-06
D1673 n1674 0 dm1 AREA=8.740e-07
D1674 n1675 0 dm1 AREA=1.185e-06
D1675 n1676 0 dm1 AREA=8.754e-07
D1676 n1677 0 dm1 AREA=4.244e-07
D1677 n1678 0 dm1 AREA=1.017e-06
D1678 n1679 0 dm1 AREA=4.769e-07
D1679 n1680 0 dm1 AREA=1.834e-06
D1680 n1681 0 dm1 AREA=7.844e-07
D1681 n1682 0 dm1 AREA=1.285e-06
D1682 n1683 0 dm1 AREA=1.127e-06
D1683 n1684 0 dm1 AREA=9.389e-07
D1684 n1685 0 dm1 AREA=1.079e-06
D1685 n1686 0 dm1 AREA=1.207e-06
D1686 n1687 0 dm1 AREA=2.989e-07
D1687 n1688 0 dm1 AREA=7.529e-07
D1688 n1689 0 dm1 AREA=1.773e-06
D1689 n1690 0 dm1 AREA=7.151e-07
D1690 n1691 0 dm1 AREA=1.445e-06
D1691 n1692 0 dm1 AREA=1.425e-06
D1692 n1693 0 dm1 AREA=4.119e-07
D1693 n1694 0 dm1 AREA=1.584e-06
D1694 n1695 0 dm1 AREA=2.493e-06
D1695 n1696 0 dm1 AREA=7.896e-07
D1696 n1697 0 dm1 AREA=6.651e-07
D1697 n1698 0 dm1 AREA=6.255e-07
D1698 n1699 0 dm1 AREA=6.275e-07
D1699 n1700 0 dm1 AREA=1.346e-06
D1700 n1701 0 dm1 AREA=4.850e-07
D1701 n1702 0 dm1 AREA=5.788e-07
D1702 n1703 0 dm1 AREA=1.174e-06
D1703 n1704 0 dm1 AREA=3.997e-07
D1704 n1705 0 dm1 AREA=2.494e-07
D1705 n1706 0 dm1 AREA=1.732e-06
D1706 n1707 0 dm1 AREA=7.541e-07
D1707 n1708 0 dm1 AREA=8.102e-07
D1708 n1 0 dm1 AREA=1.761e-06
D1709 n1710 0 dm1 AREA=1.113e-06
D1710 n1711 0 dm1 AREA=8.577e-07
D1711 n1712 0 dm1 AREA=5.294e-07
D1712 n1713 0 dm1 AREA=5.657e-07
D1713 n1714 0 dm1 AREA=5.179e-07
D1714 n1715 0 dm1 AREA=7.940e-07
D1715 n1716 0 dm1 AREA=1.025e-06
D1716 n1717 0 dm1 AREA=7.158e-07
D1717 n1718 0 dm1 AREA=8.097e-07
D1718 n1719 0 dm1 AREA=1.363e-06
D1719 n1720 0 dm1 AREA=5.915e-07
D1720 n1721 0 dm1 AREA=5.939e-07
D1721 n1722 0 dm1 AREA=1.247e-06
D1722 n1723 0 dm1 AREA=9.818e-07
D1723 n1724 0 dm1 AREA=9.705e-07
D1724 n1725 0 dm1 AREA=2.419e-07
D1725 n1726 0 dm1 AREA=1.146e-06
D1726 n1727 0 dm1 AREA=1.975e-07
D1727 n1 0 dm1 AREA=1.355e-06
D1728 n1729 0 dm1 AREA=2.292e-07
D1729 n1730 0 dm1 AREA=6.168e-07
D1730 n1731 0 dm1 AREA=6.029e-07
D1731 n1732 0 dm1 AREA=5.500e-07
D1732 n1733 0 dm1 AREA=4.763e-07
D1733 n1734 0 dm1 AREA=4.356e-07
D1734 n1735 0 dm1 AREA=7.707e-07
D1735 n1736 0 dm1 AREA=1.029e-06
D1736 n1737 0 dm1 AREA=5.111e-07
D1737 n1738 0 dm1 AREA=8.900e-07
D1738 n1739 0 dm1 AREA=8.738e-07
D1739 n1740 0 dm1 AREA=1.168e-06
D1740 n1741 0 dm1 AREA=5.439e-07
D1741 n1742 0 dm1 AREA=4.817e-07
D1742 n1743 0 dm1 AREA=1.134e-06
D1743 n1744 0 dm1 AREA=6.644e-07
D1744 n1745 0 dm1 AREA=4.353e-07
D1745 n1746 0 dm1 AREA=1.511e-06
D1746 n1747 0 dm1 AREA=9.676e-07
D1747 n1748 0 dm1 AREA=2.045e-07
D1748 n1749 0 dm1 AREA=1.126e-06
D1749 n1750 0 dm1 AREA=4.397e-07
D1750 n1751 0 dm1 AREA=3.881e-07
D1751 n1752 0 dm1 AREA=6.570e-07
D1752 n1753 0 dm1 AREA=4.137e-07
D1753 n1754 0 dm1 AREA=5.638e-07
D1754 n1755 0 dm1 AREA=8.747e-07
D1755 n1756 0 dm1 AREA=1.916e-06
D1756 n1757 0 dm1 AREA=5.311e-07
D1757 n1758 0 dm1 AREA=7.075e-07
D1758 n1759 0 dm1 AREA=7.066e-07
D1759 n1760 0 dm1 AREA=8.914e-07
D1760 n1761 0 dm1 AREA=2.158e-06
D1761 n1762 0 dm1 AREA=7.873e-07
D1762 n1763 0 dm1 AREA=1.685e-06
D1763 n1764 0 dm1 AREA=8.157e-07
D1764 n1765 0 dm1 AREA=8.651e-07
D1765 n1766 0 dm1 AREA=5.382e-07
D1766 n1767 0 dm1 AREA=7.450e-07
D1767 n1768 0 dm1 AREA=9.319e-07
D1768 n1769 0 dm1 AREA=9.541e-07
D1769 n1770 0 dm1 AREA=1.103e-06
D1770 n1771 0 dm1 AREA=1.572e-06
D1771 n1772 0 dm1 AREA=8.179e-07
D1772 n1773 0 dm1 AREA=6.183e-07
D1773 n1774 0 dm1 AREA=1.322e-06
D1774 n1775 0 dm1 AREA=8.398e-07
D1775 n1776 0 dm1 AREA=1.217e-06
D1776 n1777 0 dm1 AREA=1.311e-06
D1777 n1778 0 dm1 AREA=6.064e-07
D1778 n1779 0 dm1 AREA=8.320e-07
D1779 n1 0 dm1 AREA=8.696e-07
D1780 n1781 0 dm1 AREA=1.507e-06
D1781 n1782 0 dm1 AREA=3.721e-07
D1782 n1783 0 dm1 AREA=3.797e-07
D1783 n1784 0 dm1 AREA=5.793e-07
D1784 n1785 0 dm1 AREA=1.820e-06
D1785 n1786 0 dm1 AREA=1.533e-06
D1786 n1787 0 dm1 AREA=1.111e-06
D1787 n1788 0 dm1 AREA=8.177e-07
D1788 n1789 0 dm1 AREA=1.631e-06
D1789 n1790 0 dm1 AREA=2.270e-07
D1790 n1791 0 dm1 AREA=2.160e-06
D1791 n1792 0 dm1 AREA=6.184e-07
D1792 n1793 0 dm1 AREA=7.211e-07
D1793 n1794 0 dm1 AREA=5.235e-07
D1794 n1795 0 dm1 AREA=3.409e-07
D1795 n1796 0 dm1 AREA=8.828e-07
D1796 n1797 0 dm1 AREA=9.487e-07
D1797 n1798 0 dm1 AREA=1.057e-06
D1798 n1799 0 dm1 AREA=9.554e-07
D1799 n1800 0 dm1 AREA=8.900e-07
D1800 n1801 0 dm1 AREA=1.936e-06
D1801 n1802 0 dm1 AREA=7.800e-07
D1802 n1803 0 dm1 AREA=1.100e-06
D1803 n1804 0 dm1 AREA=1.349e-06
D1804 n1805 0 dm1 AREA=4.342e-07
D1805 n1806 0 dm1 AREA=1.128e-06
D1806 n1807 0 dm1 AREA=1.009e-06
D1807 n1808 0 dm1 AREA=1.054e-06
D1808 n1809 0 dm1 AREA=7.419e-07
D1809 n1810 0 dm1 AREA=1.314e-06
D1810 n1811 0 dm1 AREA=4.422e-07
D1811 n1812 0 dm1 AREA=5.065e-07
D1812 n1813 0 dm1 AREA=2.391e-06
D1813 n1814 0 dm1 AREA=1.926e-07
D1814 n1815 0 dm1 AREA=7.329e-07
D1815 n1816 0 dm1 AREA=1.278e-06
D1816 n1817 0 dm1 AREA=5.955e-07
D1817 n1818 0 dm1 AREA=1.687e-06
D1818 n1819 0 dm1 AREA=3.173e-07
D1819 n1820 0 dm1 AREA=1.580e-06
D1820 n1821 0 dm1 AREA=1.134e-06
D1821 n1822 0 dm1 AREA=1.168e-06
D1822 n1823 0 dm1 AREA=5.286e-07
D1823 n1824 0 dm1 AREA=5.607e-07
D1824 n1825 0 dm1 AREA=5.255e-07
D1825 n1826 0 dm1 AREA=9.545e-07
D1826 n1827 0 dm1 AREA=1.373e-06
D1827 n1828 0 dm1 AREA=1.903e-06
D1828 n1829 0 dm1 AREA=1.101e-06
D1829 n1830 0 dm1 AREA=1.456e-06
D1830 n1831 0 dm1 AREA=7.024e-07
D1831 n1832 0 dm1 AREA=7.832e-07
D1832 n1833 0 dm1 AREA=6.755e-07
D1833 n1834 0 dm1 AREA=1.466e-06
D1834 n1835 0 dm1 AREA=1.033e-06
D1835 n1836 0 dm1 AREA=4.725e-07
D1836 n1837 0 dm1 AREA=9.210e-07
D1837 n1838 0 dm1 AREA=8.962e-07
D1838 n1839 0 dm1 AREA=3.838e-07
D1839 n1 0 dm1 AREA=9.107e-07
D1840 n1841 0 dm1 AREA=5.733e-07
D1841 n1842 0 dm1 AREA=3.929e-07
D1842 n1843 0 dm1 AREA=5.914e-07
D1843 n1844 0 dm1 AREA=1.077e-06
D1844 n1845 0 dm1 AREA=5.239e-07
D1845 n1846 0 dm1 AREA=1.382e-06
D1846 n1847 0 dm1 AREA=6.928e-07
D1847 n1848 0 dm1 AREA=3.247e-07
D1848 n1849 0 dm1 AREA=1.503e-06
D1849 n1850 0 dm1 AREA=2.990e-07
D1850 n1851 0 dm1 AREA=1.144e-06
D1851 n1852 0 dm1 AREA=1.354e-06
D1852 n1853 0 dm1 AREA=2.272e-07
D1853 n1854 0 dm1 AREA=6.682e-07
D1854 n1855 0 dm1 AREA=9.590e-07
D1855 n1856 0 dm1 AREA=1.176e-06
D1856 n1857 0 dm1 AREA=1.351e-06
D1857 n1858 0 dm1 AREA=2.460e-06
D1858 n1859 0 dm1 AREA=3.457e-07
D1859 n1860 0 dm1 AREA=8.739e-07
D1860 n1861 0 dm1 AREA=5.680e-07
D1861 n1862 0 dm1 AREA=1.812e-06
D1862 n1863 0 dm1 AREA=1.108e-06
D1863 n1864 0 dm1 AREA=2.142e-06
D1864 n1865 0 dm1 AREA=1.450e-06
D1865 n1866 0 dm1 AREA=1.452e-06
D1866 n1867 0 dm1 AREA=4.373e-07
D1867 n1868 0 dm1 AREA=3.395e-06
D1868 n1869 0 dm1 AREA=1.463e-06
D1869 n1870 0 dm1 AREA=6.692e-07
D1870 n1871 0 dm1 AREA=7.720e-07
D1871 n1872 0 dm1 AREA=6.258e-07
D1872 n1873 0 dm1 AREA=1.567e-06
D1873 n1874 0 dm1 AREA=5.428e-07
D1874 n1875 0 dm1 AREA=1.265e-06
D1875 n1876 0 dm1 AREA=9.783e-07
D1876 n1877 0 dm1 AREA=3.971e-07
D1877 n1878 0 dm1 AREA=1.812e-07
D1878 n1879 0 dm1 AREA=5.318e-07
D1879 n1880 0 dm1 AREA=1.979e-06
D1880 n1881 0 dm1 AREA=1.549e-06
D1881 n1882 0 dm1 AREA=8.546e-07
D1882 n1883 0 dm1 AREA=7.570e-07
D1883 n1884 0 dm1 AREA=1.481e-06
D1884 n1885 0 dm1 AREA=1.527e-06
D1885 n1886 0 dm1 AREA=5.426e-07
D1886 n1887 0 dm1 AREA=1.632e-06
D1887 n1888 0 dm1 AREA=9.617e-07
D1888 n1889 0 dm1 AREA=1.371e-06
D1889 n1 0 dm1 AREA=1.945e-06
D1890 n1891 0 dm1 AREA=6.287e-07
D1891 n1892 0 dm1 AREA=4.215e-07
D1892 n1893 0 dm1 AREA=1.331e-06
D1893 n1894 0 dm1 AREA=1.685e-06
D1894 n1895 0 dm1 AREA=5.664e-07
D1895 n1896 0 dm1 AREA=1.140e-06
D1896 n1897 0 dm1 AREA=6.472e-07
D1897 n1898 0 dm1 AREA=5.483e-07
D1898 n1899 0 dm1 AREA=2.713e-07
D1899 n1900 0 dm1 AREA=6.003e-07
D1900 n1901 0 dm1 AREA=5.354e-07
D1901 n1902 0 dm1 AREA=1.838e-06
D1902 n1903 0 dm1 AREA=1.767e-06
D1903 n1904 0 dm1 AREA=7.617e-07
D1904 n1905 0 dm1 AREA=1.074e-06
D1905 n1906 0 dm1 AREA=1.049e-06
D1906 n1907 0 dm1 AREA=1.433e-06
D1907 n1908 0 dm1 AREA=9.792e-07
D1908 n1909 0 dm1 AREA=8.329e-07
D1909 n1910 0 dm1 AREA=1.620e-06
D1910 n1911 0 dm1 AREA=9.725e-07
D1911 n1912 0 dm1 AREA=9.399e-07
D1912 n1913 0 dm1 AREA=7.100e-07
D1913 n1914 0 dm1 AREA=8.681e-07
D1914 n1915 0 dm1 AREA=3.674e-07
D1915 n1916 0 dm1 AREA=8.930e-07
D1916 n1917 0 dm1 AREA=1.263e-06
D1917 n1918 0 dm1 AREA=7.159e-07
D1918 n1919 0 dm1 AREA=4.992e-07
D1919 n1920 0 dm1 AREA=2.990e-07
D1920 n1921 0 dm1 AREA=5.317e-07
D1921 n1922 0 dm1 AREA=1.403e-06
D1922 n1923 0 dm1 AREA=1.171e-06
D1923 n1924 0 dm1 AREA=1.828e-06
D1924 n1925 0 dm1 AREA=5.098e-07
D1925 n1926 0 dm1 AREA=8.252e-07
D1926 n1927 0 dm1 AREA=1.780e-06
D1927 n1928 0 dm1 AREA=5.749e-07
D1928 n1929 0 dm1 AREA=1.676e-06
D1929 n1930 0 dm1 AREA=8.815e-07
D1930 n1931 0 dm1 AREA=2.486e-06
D1931 n1932 0 dm1 AREA=7.559e-07
D1932 n1933 0 dm1 AREA=5.553e-07
D1933 n1934 0 dm1 AREA=2.311e-07
D1934 n1935 0 dm1 AREA=1.905e-06
D1935 n1936 0 dm1 AREA=1.660e-06
D1936 n1937 0 dm1 AREA=1.035e-06
D1937 n1938 0 dm1 AREA=1.131e-06
D1938 n1939 0 dm1 AREA=4.850e-07
D1939 n1940 0 dm1 AREA=8.489e-07
D1940 n1941 0 dm1 AREA=5.676e-07
D1941 n1942 0 dm1 AREA=1.102e-06
D1942 n1943 0 dm1 AREA=5.554e-07
D1943 n1944 0 dm1 AREA=1.114e-06
D1944 n1945 0 dm1 AREA=2.621e-07
D1945 n1946 0 dm1 AREA=1.251e-06
D1946 n1947 0 dm1 AREA=1.272e-06
D1947 n1948 0 dm1 AREA=8.436e-07
D1948 n1949 0 dm1 AREA=7.420e-07
D1949 n1950 0 dm1 AREA=2.302e-06
D1950 n1951 0 dm1 AREA=8.677e-07
D1951 n1952 0 dm1 AREA=9.340e-07
D1952 n1953 0 dm1 AREA=7.134e-07
D1953 n1954 0 dm1 AREA=9.262e-07
D1954 n1955 0 dm1 AREA=5.572e-07
D1955 n1956 0 dm1 AREA=5.127e-07
D1956 n1957 0 dm1 AREA=1.276e-06
D1957 n1958 0 dm1 AREA=6.688e-07
D1958 n1959 0 dm1 AREA=1.231e-06
D1959 n1960 0 dm1 AREA=7.938e-07
D1960 n1961 0 dm1 AREA=8.031e-07
D1961 n1962 0 dm1 AREA=8.574e-07
D1962 n1963 0 dm1 AREA=7.206e-07
D1963 n1964 0 dm1 AREA=4.988e-07
D1964 n1965 0 dm1 AREA=3.581e-07
D1965 n1966 0 dm1 AREA=6.842e-07
D1966 n1967 0 dm1 AREA=9.246e-07
D1967 n1968 0 dm1 AREA=4.888e-07
D1968 n1969 0 dm1 AREA=6.645e-07
D1969 n1970 0 dm1 AREA=1.438e-06
D1970 n1971 0 dm1 AREA=6.130e-07
D1971 n1972 0 dm1 AREA=9.062e-07
D1972 n1973 0 dm1 AREA=1.131e-06
D1973 n1974 0 dm1 AREA=9.959e-07
D1974 n1975 0 dm1 AREA=2.902e-07
D1975 n1976 0 dm1 AREA=1.210e-06
D1976 n1977 0 dm1 AREA=6.489e-07
D1977 n1978 0 dm1 AREA=5.623e-07
D1978 n1979 0 dm1 AREA=5.890e-07
D1979 n1980 0 dm1 AREA=9.539e-07
D1980 n1981 0 dm1 AREA=9.019e-07
D1981 n1982 0 dm1 AREA=6.243e-07
D1982 n1983 0 dm1 AREA=2.000e-07
D1983 n1984 0 dm1 AREA=1.057e-06
D1984 n1985 0 dm1 AREA=1.035e-06
D1985 n1986 0 dm1 AREA=2.327e-07
D1986 n1987 0 dm1 AREA=1.612e-06
D1987 n1988 0 dm1 AREA=2.959e-07
D1988 n1989 0 dm1 AREA=9.459e-07
D1989 n1990 0 dm1 AREA=1.021e-06
D1990 n1991 0 dm1 AREA=6.459e-07
D1991 n1992 0 dm1 AREA=1.777e-07
D1992 n1993 0 dm1 AREA=1.181e-06
D1993 n1994 0 dm1 AREA=5.034e-07
D1994 n1995 0 dm1 AREA=3.116e-07
D1995 n1996 0 dm1 AREA=1.757e-06
D1996 n1 0 dm1 AREA=2.182e-07
D1997 n1998 0 dm1 AREA=5.162e-07
D1998 n1999 0 dm1 AREA=9.234e-08
D1999 n2000 0 dm1 AREA=7.823e-07
D2000 n2001 0 dm1 AREA=6.867e-07
D2001 n2002 0 dm1 AREA=6.581e-07
D2002 n2003 0 dm1 AREA=5.059e-07
D2003 n2004 0 dm1 AREA=1.097e-06
D2004 n2005 0 dm1 AREA=1.000e-06
D2005 n2006 0 dm1 AREA=2.263e-06
D2006 n2007 0 dm1 AREA=7.413e-07
D2007 n2008 0 dm1 AREA=3.027e-07
D2008 n2009 0 dm1 AREA=1.505e-06
D2009 n2010 0 dm1 AREA=7.689e-07
D2010 n2011 0 dm1 AREA=1.843e-06
D2011 n2012 0 dm1 AREA=6.532e-07
D2012 n2013 0 dm1 AREA=8.499e-07
D2013 n2014 0 dm1 AREA=1.216e-06
D2014 n2015 0 dm1 AREA=9.929e-07
D2015 n2016 0 dm1 AREA=1.165e-06
D2016 n2017 0 dm1 AREA=9.895e-07
D2017 n2018 0 dm1 AREA=1.855e-06
D2018 n2019 0 dm1 AREA=1.189e-06
D2019 n2020 0 dm1 AREA=1.426e-06
D2020 n2021 0 dm1 AREA=2.278e-07
D2021 n2022 0 dm1 AREA=1.057e-06
D2022 n2023 0 dm1 AREA=5.373e-07
D2023 n2024 0 dm1 AREA=1.290e-06
D2024 n2025 0 dm1 AREA=4.603e-07
D2025 n2026 0 dm1 AREA=3.859e-07
D2026 n2027 0 dm1 AREA=7.638e-07
D2027 n2028 0 dm1 AREA=1.768e-06
D2028 n2029 0 dm1 AREA=1.986e-06
D2029 n2030 0 dm1 AREA=6.722e-07
D2030 n2031 0 dm1 AREA=8.353e-07
D2031 n2032 0 dm1 AREA=8.105e-07
D2032 n2033 0 dm1 AREA=9.030e-07
D2033 n2034 0 dm1 AREA=1.670e-06
D2034 n2035 0 dm1 AREA=8.652e-07
D2035 n2036 0 dm1 AREA=9.608e-07
D2036 n2037 0 dm1 AREA=8.426e-07
D2037 n2038 0 dm1 AREA=2.499e-07
D2038 n2039 0 dm1 AREA=8.031e-07
D2039 n2040 0 dm1 AREA=1.334e-06
D2040 n2041 0 dm1 AREA=9.767e-07
D2041 n2042 0 dm1 AREA=1.655e-06
D2042 n2043 0 dm1 AREA=4.985e-07
D2043 n2044 0 dm1 AREA=8.287e-07
D2044 n2045 0 dm1 AREA=5.938e-07
D2045 n2046 0 dm1 AREA=6.605e-07
D2046 n1 0 dm1 AREA=1.342e-06
D2047 n2048 0 dm1 AREA=8.033e-07
D2048 n2049 0 dm1 AREA=3.635e-07
D2049 n2050 0 dm1 AREA=7.804e-07
D2050 n2051 0 dm1 AREA=1.177e-06
D2051 n2052 0 dm1 AREA=1.547e-06
D2052 n2053 0 dm1 AREA=1.432e-06
D2053 n2054 0 dm1 AREA=8.775e-07
D2054 n2055 0 dm1 AREA=2.473e-06
D2055 n2056 0 dm1 AREA=7.864e-07
D2056 n2057 0 dm1 AREA=6.706e-07
D2057 n2058 0 dm1 AREA=6.701e-07
D2058 n2059 0 dm1 AREA=1.046e-06
D2059 n2060 0 dm1 AREA=5.647e-07
D2060 n2061 0 dm1 AREA=1.498e-06
D2061 n2062 0 dm1 AREA=7.948e-07
D2062 n2063 0 dm1 AREA=3.449e-07
D2063 n1 0 dm1 AREA=1.298e-06
D2064 n2065 0 dm1 AREA=1.233e-06
D2065 n2066 0 dm1 AREA=8.322e-07
D2066 n2067 0 dm1 AREA=9.901e-08
D2067 n2068 0 dm1 AREA=1.405e-06
D2068 n2069 0 dm1 AREA=6.567e-07
D2069 n2070 0 dm1 AREA=6.759e-07
D2070 n2071 0 dm1 AREA=1.327e-06
D2071 n2072 0 dm1 AREA=9.444e-07
D2072 n2073 0 dm1 AREA=7.577e-07
D2073 n2074 0 dm1 AREA=2.917e-06
D2074 n2075 0 dm1 AREA=7.127e-07
D2075 n2076 0 dm1 AREA=8.658e-07
D2076 n2077 0 dm1 AREA=1.321e-06
D2077 n2078 0 dm1 AREA=6.208e-07
D2078 n2079 0 dm1 AREA=1.302e-06
D2079 n2080 0 dm1 AREA=3.437e-07
D2080 n2081 0 dm1 AREA=2.784e-06
D2081 n2082 0 dm1 AREA=9.780e-07
D2082 n2083 0 dm1 AREA=8.265e-07
D2083 n2084 0 dm1 AREA=8.540e-07
D2084 n2085 0 dm1 AREA=7.410e-07
D2085 n2086 0 dm1 AREA=5.644e-07
D2086 n2087 0 dm1 AREA=1.194e-06
D2087 n2088 0 dm1 AREA=1.243e-06
D2088 n2089 0 dm1 AREA=6.347e-07
D2089 n2090 0 dm1 AREA=8.021e-07
D2090 n2091 0 dm1 AREA=6.030e-07
D2091 n1 0 dm1 AREA=7.243e-07
D2092 n2093 0 dm1 AREA=5.088e-07
D2093 n2094 0 dm1 AREA=1.932e-06
D2094 n2095 0 dm1 AREA=2.083e-06
D2095 n2096 0 dm1 AREA=1.405e-06
D2096 n2097 0 dm1 AREA=3.500e-07
D2097 n2098 0 dm1 AREA=6.614e-07
D2098 n2099 0 dm1 AREA=1.235e-06
D2099 n2100 0 dm1 AREA=2.291e-06
D2100 n2101 0 dm1 AREA=1.549e-06
D2101 n2102 0 dm1 AREA=9.375e-07
D2102 n2103 0 dm1 AREA=1.239e-06
D2103 n2104 0 dm1 AREA=6.257e-07
D2104 n2105 0 dm1 AREA=7.990e-07
D2105 n2106 0 dm1 AREA=2.039e-06
D2106 n2107 0 dm1 AREA=1.122e-06
D2107 n2108 0 dm1 AREA=1.017e-06
D2108 n2109 0 dm1 AREA=1.618e-06
D2109 n2110 0 dm1 AREA=6.361e-07
D2110 n2111 0 dm1 AREA=1.836e-06
D2111 n2112 0 dm1 AREA=1.302e-06
D2112 n2113 0 dm1 AREA=7.981e-07
D2113 n2114 0 dm1 AREA=7.469e-07
D2114 n2115 0 dm1 AREA=1.063e-06
D2115 n2116 0 dm1 AREA=1.786e-06
D2116 n2117 0 dm1 AREA=9.167e-07
D2117 n2118 0 dm1 AREA=1.659e-06
D2118 n2119 0 dm1 AREA=1.126e-06
D2119 n2120 0 dm1 AREA=1.783e-06
D2120 n2121 0 dm1 AREA=4.838e-07
D2121 n2122 0 dm1 AREA=1.865e-07
D2122 n2123 0 dm1 AREA=4.438e-07
D2123 n2124 0 dm1 AREA=8.383e-07
D2124 n2125 0 dm1 AREA=7.571e-07
D2125 n2126 0 dm1 AREA=8.509e-07
D2126 n2127 0 dm1 AREA=4.608e-07
D2127 n2128 0 dm1 AREA=5.149e-07
D2128 n2129 0 dm1 AREA=1.741e-06
D2129 n2130 0 dm1 AREA=2.036e-07
D2130 n2131 0 dm1 AREA=4.481e-07
D2131 n2132 0 dm1 AREA=6.967e-07
D2132 n2133 0 dm1 AREA=6.966e-07
D2133 n2134 0 dm1 AREA=4.792e-07
D2134 n2135 0 dm1 AREA=1.373e-06
D2135 n2136 0 dm1 AREA=1.397e-06
D2136 n2137 0 dm1 AREA=3.190e-07
D2137 n2138 0 dm1 AREA=1.173e-06
D2138 n2139 0 dm1 AREA=9.706e-07
D2139 n2140 0 dm1 AREA=6.463e-07
D2140 n2141 0 dm1 AREA=1.744e-06
D2141 n2142 0 dm1 AREA=1.434e-07
D2142 n2143 0 dm1 AREA=9.602e-07
D2143 n2144 0 dm1 AREA=9.740e-07
D2144 n2145 0 dm1 AREA=4.950e-07
D2145 n2146 0 dm1 AREA=6.387e-07
D2146 n2147 0 dm1 AREA=7.913e-07
D2147 n2148 0 dm1 AREA=1.062e-06
D2148 n2149 0 dm1 AREA=7.029e-07
D2149 n2150 0 dm1 AREA=8.487e-07
D2150 n2151 0 dm1 AREA=9.049e-07
D2151 n2152 0 dm1 AREA=4.044e-07
D2152 n2153 0 dm1 AREA=9.971e-07
D2153 n2154 0 dm1 AREA=8.425e-07
D2154 n2155 0 dm1 AREA=2.906e-06
D2155 n2156 0 dm1 AREA=8.577e-07
D2156 n2157 0 dm1 AREA=6.364e-07
D2157 n2158 0 dm1 AREA=1.213e-06
D2158 n2159 0 dm1 AREA=1.787e-06
D2159 n2160 0 dm1 AREA=4.385e-07
D2160 n2161 0 dm1 AREA=1.577e-06
D2161 n2162 0 dm1 AREA=1.406e-07
D2162 n2163 0 dm1 AREA=4.220e-07
D2163 n2164 0 dm1 AREA=2.298e-06
D2164 n2165 0 dm1 AREA=2.135e-06
D2165 n2166 0 dm1 AREA=4.399e-07
D2166 n2167 0 dm1 AREA=1.004e-06
D2167 n2168 0 dm1 AREA=6.744e-07
D2168 n2169 0 dm1 AREA=1.557e-06
D2169 n2170 0 dm1 AREA=9.895e-07
D2170 n2171 0 dm1 AREA=4.565e-07
D2171 n2172 0 dm1 AREA=7.064e-07
D2172 n2173 0 dm1 AREA=2.167e-06
D2173 n2174 0 dm1 AREA=8.865e-07
D2174 n2175 0 dm1 AREA=1.032e-06
D2175 n2176 0 dm1 AREA=5.922e-07
D2176 n2177 0 dm1 AREA=1.342e-06
D2177 n2178 0 dm1 AREA=8.342e-07
D2178 n2179 0 dm1 AREA=8.205e-07
D2179 n2180 0 dm1 AREA=6.534e-07
D2180 n2181 0 dm1 AREA=8.362e-07
D2181 n2182 0 dm1 AREA=8.987e-07
D2182 n2183 0 dm1 AREA=4.565e-07
D2183 n2184 0 dm1 AREA=2.401e-06
D2184 n2185 0 dm1 AREA=9.465e-07
D2185 n2186 0 dm1 AREA=6.285e-07
D2186 n2187 0 dm1 AREA=9.879e-07
D2187 n2188 0 dm1 AREA=7.897e-07
D2188 n2189 0 dm1 AREA=1.046e-06
D2189 n2190 0 dm1 AREA=1.663e-06
D2190 n2191 0 dm1 AREA=4.882e-07
D2191 n2192 0 dm1 AREA=1.737e-06
D2192 n2193 0 dm1 AREA=1.034e-06
D2193 n2194 0 dm1 AREA=1.200e-06
D2194 n2195 0 dm1 AREA=1.549e-06
D2195 n2196 0 dm1 AREA=1.215e-06
D2196 n2197 0 dm1 AREA=2.714e-07
D2197 n2198 0 dm1 AREA=3.861e-07
D2198 n1 0 dm1 AREA=3.887e-07
D2199 n2200 0 dm1 AREA=3.319e-07
D2200 n2201 0 dm1 AREA=2.867e-07
D2201 n2202 0 dm1 AREA=9.656e-07
D2202 n2203 0 dm1 AREA=6.323e-07
D2203 n2204 0 dm1 AREA=6.459e-07
D2204 n2205 0 dm1 AREA=5.207e-07
D2205 n2206 0 dm1 AREA=1.634e-06
D2206 n2207 0 dm1 AREA=1.210e-06
D2207 n2208 0 dm1 AREA=4.689e-07
D2208 n2209 0 dm1 AREA=4.464e-07
D2209 n2210 0 dm1 AREA=8.206e-07
D2210 n2211 0 dm1 AREA=2.393e-07
D2211 n2212 0 dm1 AREA=2.062e-06
D2212 n2213 0 dm1 AREA=7.537e-07
D2213 n2214 0 dm1 AREA=2.761e-06
D2214 n2215 0 dm1 AREA=6.550e-07
D2215 n2216 0 dm1 AREA=8.558e-07
D2216 n2217 0 dm1 AREA=1.511e-06
D2217 n2218 0 dm1 AREA=7.508e-08
D2218 n2219 0 dm1 AREA=5.346e-07
D2219 n2220 0 dm1 AREA=1.361e-06
D2220 n2221 0 dm1 AREA=2.811e-07
D2221 n2222 0 dm1 AREA=9.220e-07
D2222 n2223 0 dm1 AREA=5.009e-07
D2223 n2224 0 dm1 AREA=5.430e-07
D2224 n2225 0 dm1 AREA=6.140e-07
D2225 n2226 0 dm1 AREA=1.192e-06
D2226 n2227 0 dm1 AREA=9.044e-07
D2227 n2228 0 dm1 AREA=1.476e-06
D2228 n2229 0 dm1 AREA=1.875e-06
D2229 n2230 0 dm1 AREA=9.268e-07
D2230 n2231 0 dm1 AREA=2.750e-06
D2231 n2232 0 dm1 AREA=2.554e-06
D2232 n2233 0 dm1 AREA=8.788e-07
D2233 n2234 0 dm1 AREA=1.265e-06
D2234 n2235 0 dm1 AREA=1.327e-06
D2235 n2236 0 dm1 AREA=4.242e-07
D2236 n2237 0 dm1 AREA=4.978e-07
D2237 n2238 0 dm1 AREA=1.125e-06
D2238 n2239 0 dm1 AREA=6.187e-07
D2239 n2240 0 dm1 AREA=7.677e-07
D2240 n2241 0 dm1 AREA=4.882e-07
D2241 n2242 0 dm1 AREA=5.364e-07
D2242 n2243 0 dm1 AREA=7.884e-07
D2243 n2244 0 dm1 AREA=9.529e-07
D2244 n2245 0 dm1 AREA=1.449e-06
D2245 n2246 0 dm1 AREA=7.995e-07
D2246 n2247 0 dm1 AREA=1.856e-07
D2247 n2248 0 dm1 AREA=1.395e-06
D2248 n2249 0 dm1 AREA=4.439e-07
D2249 n2250 0 dm1 AREA=1.138e-06
D2250 n2251 0 dm1 AREA=1.429e-06
D2251 n2252 0 dm1 AREA=8.008e-07
D2252 n2253 0 dm1 AREA=4.394e-07
D2253 n2254 0 dm1 AREA=5.451e-07
D2254 n2255 0 dm1 AREA=6.261e-07
D2255 n2256 0 dm1 AREA=1.005e-06
D2256 n2257 0 dm1 AREA=1.515e-06
D2257 n2258 0 dm1 AREA=1.178e-06
D2258 n2259 0 dm1 AREA=2.041e-06
D2259 n2260 0 dm1 AREA=2.133e-06
D2260 n2261 0 dm1 AREA=4.922e-07
D2261 n2262 0 dm1 AREA=1.363e-06
D2262 n2263 0 dm1 AREA=3.755e-07
D2263 n2264 0 dm1 AREA=1.050e-06
D2264 n2265 0 dm1 AREA=9.658e-07
D2265 n2266 0 dm1 AREA=8.345e-07
D2266 n2267 0 dm1 AREA=5.907e-07
D2267 n2268 0 dm1 AREA=7.686e-07
D2268 n2269 0 dm1 AREA=8.875e-07
D2269 n2270 0 dm1 AREA=5.714e-07
D2270 n2271 0 dm1 AREA=1.160e-06
D2271 n2272 0 dm1 AREA=2.971e-07
D2272 n2273 0 dm1 AREA=5.009e-07
D2273 n2274 0 dm1 AREA=4.281e-07
D2274 n2275 0 dm1 AREA=8.384e-07
D2275 n2276 0 dm1 AREA=1.606e-06
D2276 n2277 0 dm1 AREA=2.624e-06
D2277 n2278 0 dm1 AREA=1.203e-06
D2278 n2279 0 dm1 AREA=5.137e-07
D2279 n2280 0 dm1 AREA=9.832e-07
D2280 n2281 0 dm1 AREA=2.251e-06
D2281 n2282 0 dm1 AREA=3.836e-07
D2282 n2283 0 dm1 AREA=2.938e-07
D2283 n2284 0 dm1 AREA=7.985e-07
D2284 n2285 0 dm1 AREA=1.663e-06
D2285 n2286 0 dm1 AREA=6.374e-07
D2286 n2287 0 dm1 AREA=8.369e-07
D2287 n2288 0 dm1 AREA=9.742e-07
D2288 n2289 0 dm1 AREA=8.272e-07
D2289 n2290 0 dm1 AREA=7.935e-07
D2290 n2291 0 dm1 AREA=1.067e-06
D2291 n2292 0 dm1 AREA=1.255e-06
D2292 n2293 0 dm1 AREA=6.951e-07
D2293 n2294 0 dm1 AREA=9.446e-07
D2294 n2295 0 dm1 AREA=8.201e-07
D2295 n2296 0 dm1 AREA=1.428e-06
D2296 n2297 0 dm1 AREA=2.120e-07
D2297 n2298 0 dm1 AREA=1.543e-06
D2298 n2299 0 dm1 AREA=1.925e-06
D2299 n2300 0 dm1 AREA=7.082e-07
D2300 n2301 0 dm1 AREA=4.028e-07
D2301 n2302 0 dm1 AREA=9.104e-07
D2302 n2303 0 dm1 AREA=2.067e-07
D2303 n2304 0 dm1 AREA=4.619e-07
D2304 n2305 0 dm1 AREA=1.323e-06
D2305 n2306 0 dm1 AREA=7.307e-07
D2306 n2307 0 dm1 AREA=8.662e-07
D2307 n2308 0 dm1 AREA=6.367e-07
D2308 n2309 0 dm1 AREA=2.154e-06
D2309 n2310 0 dm1 AREA=2.136e-07
D2310 n2311 0 dm1 AREA=1.175e-06
D2311 n2312 0 dm1 AREA=8.020e-07
D2312 n2313 0 dm1 AREA=2.294e-06
D2313 n2314 0 dm1 AREA=1.538e-06
D2314 n2315 0 dm1 AREA=5.259e-07
D2315 n2316 0 dm1 AREA=1.132e-06
D2316 n2317 0 dm1 AREA=4.362e-07
D2317 n2318 0 dm1 AREA=2.112e-06
D2318 n2319 0 dm1 AREA=6.480e-07
D2319 n2320 0 dm1 AREA=9.173e-07
D2320 n2321 0 dm1 AREA=3.056e-07
D2321 n2322 0 dm1 AREA=8.414e-07
D2322 n2323 0 dm1 AREA=7.563e-07
D2323 n2324 0 dm1 AREA=1.352e-06
D2324 n2325 0 dm1 AREA=8.671e-07
D2325 n2326 0 dm1 AREA=1.518e-06
D2326 n2327 0 dm1 AREA=1.754e-06
D2327 n2328 0 dm1 AREA=1.782e-06
D2328 n2329 0 dm1 AREA=1.475e-06
D2329 n2330 0 dm1 AREA=9.287e-07
D2330 n2331 0 dm1 AREA=8.393e-07
D2331 n2332 0 dm1 AREA=1.769e-06
D2332 n2333 0 dm1 AREA=1.999e-06
D2333 n2334 0 dm1 AREA=1.345e-06
D2334 n2335 0 dm1 AREA=7.447e-07
D2335 n2336 0 dm1 AREA=4.393e-07
D2336 n2337 0 dm1 AREA=1.258e-06
D2337 n2338 0 dm1 AREA=1.236e-06
D2338 n2339 0 dm1 AREA=1.099e-06
D2339 n2340 0 dm1 AREA=1.862e-06
D2340 n2341 0 dm1 AREA=9.950e-07
D2341 n2342 0 dm1 AREA=1.088e-06
D2342 n2343 0 dm1 AREA=1.170e-06
D2343 n2344 0 dm1 AREA=1.531e-06
D2344 n2345 0 dm1 AREA=8.198e-07
D2345 n2346 0 dm1 AREA=1.329e-06
D2346 n2347 0 dm1 AREA=1.320e-06
D2347 n2348 0 dm1 AREA=7.072e-07
D2348 n2349 0 dm1 AREA=3.952e-07
D2349 n2350 0 dm1 AREA=1.853e-06
D2350 n2351 0 dm1 AREA=7.631e-07
D2351 n2352 0 dm1 AREA=1.628e-06
D2352 n2353 0 dm1 AREA=9.407e-07
D2353 n2354 0 dm1 AREA=8.857e-07
D2354 n2355 0 dm1 AREA=4.743e-07
D2355 n2356 0 dm1 AREA=1.207e-06
D2356 n2357 0 dm1 AREA=6.741e-07
D2357 n2358 0 dm1 AREA=9.194e-07
D2358 n2359 0 dm1 AREA=7.249e-07
D2359 n2360 0 dm1 AREA=1.275e-06
D2360 n2361 0 dm1 AREA=8.858e-07
D2361 n2362 0 dm1 AREA=2.503e-06
D2362 n2363 0 dm1 AREA=5.120e-07
D2363 n2364 0 dm1 AREA=7.487e-07
D2364 n2365 0 dm1 AREA=2.591e-07
D2365 n2366 0 dm1 AREA=2.260e-06
D2366 n2367 0 dm1 AREA=1.291e-06
D2367 n2368 0 dm1 AREA=1.565e-06
D2368 n2369 0 dm1 AREA=7.624e-07
D2369 n2370 0 dm1 AREA=9.977e-07
D2370 n2371 0 dm1 AREA=1.933e-06
D2371 n2372 0 dm1 AREA=1.290e-06
D2372 n2373 0 dm1 AREA=1.131e-06
D2373 n2374 0 dm1 AREA=2.511e-07
D2374 n2375 0 dm1 AREA=9.276e-07
D2375 n2376 0 dm1 AREA=8.498e-07
D2376 n2377 0 dm1 AREA=4.500e-07
D2377 n2378 0 dm1 AREA=3.602e-07
D2378 n2379 0 dm1 AREA=7.984e-07
D2379 n2380 0 dm1 AREA=1.047e-06
D2380 n2381 0 dm1 AREA=1.292e-06
D2381 n2382 0 dm1 AREA=1.629e-06
D2382 n2383 0 dm1 AREA=1.893e-06
D2383 n2384 0 dm1 AREA=1.034e-06
D2384 n2385 0 dm1 AREA=4.862e-07
D2385 n2386 0 dm1 AREA=1.734e-06
D2386 n2387 0 dm1 AREA=4.733e-07
D2387 n2388 0 dm1 AREA=1.608e-06
D2388 n2389 0 dm1 AREA=6.259e-07
D2389 n2390 0 dm1 AREA=7.946e-07
D2390 n2391 0 dm1 AREA=2.454e-06
D2391 n2392 0 dm1 AREA=1.308e-06
D2392 n2393 0 dm1 AREA=1.391e-06
D2393 n2394 0 dm1 AREA=8.803e-07
D2394 n2395 0 dm1 AREA=8.492e-07
D2395 n1 0 dm1 AREA=8.314e-07
D2396 n2397 0 dm1 AREA=1.646e-06
D2397 n2398 0 dm1 AREA=4.386e-07
D2398 n2399 0 dm1 AREA=9.774e-07
D2399 n2400 0 dm1 AREA=7.101e-07
D2400 n2401 0 dm1 AREA=4.350e-07
D2401 n2402 0 dm1 AREA=1.627e-06
D2402 n2403 0 dm1 AREA=1.000e-06
D2403 n2404 0 dm1 AREA=1.339e-06
D2404 n2405 0 dm1 AREA=2.530e-06
D2405 n2406 0 dm1 AREA=1.793e-07
D2406 n2407 0 dm1 AREA=4.290e-07
D2407 n2408 0 dm1 AREA=4.382e-07
D2408 n2409 0 dm1 AREA=5.815e-07
D2409 n2410 0 dm1 AREA=1.024e-06
D2410 n2411 0 dm1 AREA=4.443e-07
D2411 n2412 0 dm1 AREA=7.058e-07
D2412 n2413 0 dm1 AREA=1.171e-06
D2413 n2414 0 dm1 AREA=1.187e-06
D2414 n2415 0 dm1 AREA=1.574e-07
D2415 n2416 0 dm1 AREA=1.912e-06
D2416 n2417 0 dm1 AREA=6.171e-07
D2417 n2418 0 dm1 AREA=7.303e-07
D2418 n2419 0 dm1 AREA=1.452e-06
D2419 n2420 0 dm1 AREA=1.282e-06
D2420 n2421 0 dm1 AREA=1.507e-06
D2421 n2422 0 dm1 AREA=1.140e-06
D2422 n2423 0 dm1 AREA=5.262e-07
D2423 n2424 0 dm1 AREA=1.772e-06
D2424 n2425 0 dm1 AREA=7.328e-07
D2425 n2426 0 dm1 AREA=2.723e-07
D2426 n2427 0 dm1 AREA=5.149e-07
D2427 n2428 0 dm1 AREA=1.037e-06
D2428 n2429 0 dm1 AREA=4.073e-07
D2429 n2430 0 dm1 AREA=6.099e-07
D2430 n2431 0 dm1 AREA=7.608e-07
D2431 n2432 0 dm1 AREA=7.523e-07
D2432 n2433 0 dm1 AREA=2.105e-06
D2433 n2434 0 dm1 AREA=1.661e-06
D2434 n2435 0 dm1 AREA=6.407e-07
D2435 n2436 0 dm1 AREA=1.241e-06
D2436 n2437 0 dm1 AREA=1.334e-06
D2437 n2438 0 dm1 AREA=1.908e-06
D2438 n2439 0 dm1 AREA=9.100e-07
D2439 n1 0 dm1 AREA=8.140e-07
D2440 n2441 0 dm1 AREA=7.192e-07
D2441 n2442 0 dm1 AREA=6.181e-07
D2442 n2443 0 dm1 AREA=9.606e-07
D2443 n2444 0 dm1 AREA=8.612e-07
D2444 n2445 0 dm1 AREA=5.962e-07
D2445 n2446 0 dm1 AREA=5.992e-07
D2446 n1 0 dm1 AREA=6.661e-07
D2447 n2448 0 dm1 AREA=8.987e-07
D2448 n2449 0 dm1 AREA=7.015e-07
D2449 n2450 0 dm1 AREA=8.760e-07
D2450 n2451 0 dm1 AREA=1.185e-06
D2451 n2452 0 dm1 AREA=3.762e-07
D2452 n2453 0 dm1 AREA=8.338e-07
D2453 n2454 0 dm1 AREA=6.166e-07
D2454 n2455 0 dm1 AREA=1.850e-06
D2455 n2456 0 dm1 AREA=3.721e-07
D2456 n2457 0 dm1 AREA=7.840e-07
D2457 n2458 0 dm1 AREA=6.574e-07
D2458 n2459 0 dm1 AREA=1.590e-06
D2459 n2460 0 dm1 AREA=6.168e-07
D2460 n2461 0 dm1 AREA=2.128e-06
D2461 n2462 0 dm1 AREA=2.375e-06
D2462 n2463 0 dm1 AREA=1.184e-06
D2463 n2464 0 dm1 AREA=8.589e-07
D2464 n2465 0 dm1 AREA=8.669e-07
D2465 n2466 0 dm1 AREA=1.448e-06
D2466 n2467 0 dm1 AREA=1.253e-06
D2467 n2468 0 dm1 AREA=1.489e-06
D2468 n2469 0 dm1 AREA=8.677e-07
D2469 n2470 0 dm1 AREA=1.065e-06
D2470 n2471 0 dm1 AREA=8.004e-07
D2471 n2472 0 dm1 AREA=1.796e-06
D2472 n2473 0 dm1 AREA=7.839e-07
D2473 n2474 0 dm1 AREA=1.183e-06
D2474 n2475 0 dm1 AREA=1.400e-06
D2475 n2476 0 dm1 AREA=1.799e-06
D2476 n2477 0 dm1 AREA=1.019e-06
D2477 n2478 0 dm1 AREA=6.991e-07
D2478 n2479 0 dm1 AREA=3.040e-07
D2479 n2480 0 dm1 AREA=2.283e-07
D2480 n2481 0 dm1 AREA=6.262e-07
D2481 n2482 0 dm1 AREA=7.751e-07
D2482 n2483 0 dm1 AREA=1.470e-06
D2483 n2484 0 dm1 AREA=9.797e-07
D2484 n2485 0 dm1 AREA=1.165e-06
D2485 n2486 0 dm1 AREA=1.458e-06
D2486 n2487 0 dm1 AREA=7.819e-07
D2487 n2488 0 dm1 AREA=2.581e-06
D2488 n2489 0 dm1 AREA=1.565e-06
D2489 n2490 0 dm1 AREA=1.010e-06
D2490 n2491 0 dm1 AREA=1.366e-06
D2491 n2492 0 dm1 AREA=1.218e-06
D2492 n2493 0 dm1 AREA=2.969e-07
D2493 n2494 0 dm1 AREA=1.901e-06
D2494 n2495 0 dm1 AREA=6.021e-07
D2495 n2496 0 dm1 AREA=2.527e-06
D2496 n2497 0 dm1 AREA=3.817e-07
D2497 n2498 0 dm1 AREA=1.268e-06
D2498 n2499 0 dm1 AREA=1.553e-06
D2499 n2500 0 dm1 AREA=1.166e-06
D2500 n2501 0 dm1 AREA=1.164e-06
D2501 n2502 0 dm1 AREA=3.794e-07
D2502 n2503 0 dm1 AREA=2.255e-07
D2503 n2504 0 dm1 AREA=1.341e-06
D2504 n2505 0 dm1 AREA=2.153e-06
D2505 n2506 0 dm1 AREA=8.914e-07
D2506 n2507 0 dm1 AREA=5.773e-07
D2507 n2508 0 dm1 AREA=8.529e-07
D2508 n2509 0 dm1 AREA=2.473e-06
D2509 n2510 0 dm1 AREA=5.346e-07
D2510 n2511 0 dm1 AREA=7.277e-07
D2511 n2512 0 dm1 AREA=6.381e-07
D2512 n2513 0 dm1 AREA=2.244e-06
D2513 n2514 0 dm1 AREA=8.029e-07
D2514 n2515 0 dm1 AREA=1.078e-06
D2515 n2516 0 dm1 AREA=9.418e-07
D2516 n2517 0 dm1 AREA=9.086e-07
D2517 n2518 0 dm1 AREA=2.688e-07
D2518 n2519 0 dm1 AREA=7.714e-07
D2519 n2520 0 dm1 AREA=3.710e-07
D2520 n2521 0 dm1 AREA=8.298e-07
D2521 n2522 0 dm1 AREA=7.694e-07
D2522 n2523 0 dm1 AREA=5.372e-07
D2523 n2524 0 dm1 AREA=1.260e-06
D2524 n2525 0 dm1 AREA=1.470e-07
D2525 n2526 0 dm1 AREA=1.162e-06
D2526 n2527 0 dm1 AREA=3.333e-07
D2527 n2528 0 dm1 AREA=3.868e-07
D2528 n2529 0 dm1 AREA=1.221e-06
D2529 n2530 0 dm1 AREA=5.357e-07
D2530 n2531 0 dm1 AREA=3.518e-07
D2531 n2532 0 dm1 AREA=6.841e-07
D2532 n2533 0 dm1 AREA=9.216e-07
D2533 n2534 0 dm1 AREA=1.469e-06
D2534 n2535 0 dm1 AREA=5.862e-07
D2535 n2536 0 dm1 AREA=8.243e-07
D2536 n2537 0 dm1 AREA=1.433e-06
D2537 n2538 0 dm1 AREA=5.693e-07
D2538 n2539 0 dm1 AREA=8.337e-07
D2539 n2540 0 dm1 AREA=1.421e-06
D2540 n2541 0 dm1 AREA=4.370e-07
D2541 n2542 0 dm1 AREA=5.394e-07
D2542 n2543 0 dm1 AREA=3.093e-07
D2543 n2544 0 dm1 AREA=2.746e-07
D2544 n2545 0 dm1 AREA=2.135e-06
D2545 n2546 0 dm1 AREA=6.211e-07
D2546 n2547 0 dm1 AREA=4.799e-07
D2547 n2548 0 dm1 AREA=6.559e-07
D2548 n2549 0 dm1 AREA=3.161e-07
D2549 n2550 0 dm1 AREA=1.393e-06
D2550 n2551 0 dm1 AREA=1.157e-06
D2551 n2552 0 dm1 AREA=8.334e-07
D2552 n2553 0 dm1 AREA=6.920e-07
D2553 n2554 0 dm1 AREA=5.610e-07
D2554 n2555 0 dm1 AREA=6.037e-07
D2555 n2556 0 dm1 AREA=1.416e-06
D2556 n2557 0 dm1 AREA=1.097e-06
D2557 n2558 0 dm1 AREA=5.185e-07
D2558 n2559 0 dm1 AREA=5.197e-07
D2559 n2560 0 dm1 AREA=5.407e-07
D2560 n2561 0 dm1 AREA=6.848e-07
D2561 n2562 0 dm1 AREA=1.812e-06
D2562 n2563 0 dm1 AREA=1.781e-06
D2563 n2564 0 dm1 AREA=1.069e-06
D2564 n2565 0 dm1 AREA=1.635e-06
D2565 n2566 0 dm1 AREA=1.360e-06
D2566 n2567 0 dm1 AREA=5.008e-07
D2567 n2568 0 dm1 AREA=1.106e-06
D2568 n2569 0 dm1 AREA=1.779e-06
D2569 n2570 0 dm1 AREA=6.979e-07
D2570 n2571 0 dm1 AREA=9.677e-07
D2571 n1 0 dm1 AREA=9.258e-07
D2572 n2573 0 dm1 AREA=5.622e-07
D2573 n2574 0 dm1 AREA=2.028e-07
D2574 n2575 0 dm1 AREA=1.268e-06
D2575 n2576 0 dm1 AREA=9.871e-07
D2576 n2577 0 dm1 AREA=1.046e-06
D2577 n2578 0 dm1 AREA=1.007e-06
D2578 n2579 0 dm1 AREA=6.481e-07
D2579 n2580 0 dm1 AREA=7.577e-07
D2580 n2581 0 dm1 AREA=3.136e-07
D2581 n2582 0 dm1 AREA=9.670e-07
D2582 n2583 0 dm1 AREA=5.466e-07
D2583 n2584 0 dm1 AREA=1.964e-06
D2584 n2585 0 dm1 AREA=3.953e-07
D2585 n2586 0 dm1 AREA=1.016e-06
D2586 n2587 0 dm1 AREA=6.430e-07
D2587 n2588 0 dm1 AREA=7.140e-07
D2588 n2589 0 dm1 AREA=9.229e-07
D2589 n2590 0 dm1 AREA=5.621e-07
D2590 n2591 0 dm1 AREA=5.487e-07
D2591 n2592 0 dm1 AREA=1.060e-06
D2592 n2593 0 dm1 AREA=1.065e-06
D2593 n2594 0 dm1 AREA=6.890e-07
D2594 n2595 0 dm1 AREA=8.534e-07
D2595 n2596 0 dm1 AREA=1.902e-06
D2596 n2597 0 dm1 AREA=9.030e-07
D2597 n2598 0 dm1 AREA=4.148e-07
D2598 n2599 0 dm1 AREA=4.005e-07
D2599 n2600 0 dm1 AREA=1.358e-06
D2600 n2601 0 dm1 AREA=2.236e-07
D2601 n2602 0 dm1 AREA=9.544e-07
D2602 n2603 0 dm1 AREA=2.660e-07
D2603 n2604 0 dm1 AREA=7.735e-07
D2604 n2605 0 dm1 AREA=1.077e-06
D2605 n2606 0 dm1 AREA=7.866e-07
D2606 n2607 0 dm1 AREA=8.451e-07
D2607 n2608 0 dm1 AREA=1.112e-07
D2608 n2609 0 dm1 AREA=1.086e-06
D2609 n2610 0 dm1 AREA=2.092e-07
D2610 n1 0 dm1 AREA=1.060e-06
D2611 n2612 0 dm1 AREA=1.952e-07
D2612 n2613 0 dm1 AREA=1.601e-06
D2613 n2614 0 dm1 AREA=6.157e-07
D2614 n2615 0 dm1 AREA=9.849e-07
D2615 n2616 0 dm1 AREA=5.728e-07
D2616 n2617 0 dm1 AREA=9.350e-07
D2617 n2618 0 dm1 AREA=2.005e-06
D2618 n2619 0 dm1 AREA=6.181e-07
D2619 n2620 0 dm1 AREA=1.636e-06
D2620 n2621 0 dm1 AREA=6.408e-07
D2621 n2622 0 dm1 AREA=4.041e-07
D2622 n2623 0 dm1 AREA=6.394e-07
D2623 n2624 0 dm1 AREA=6.523e-07
D2624 n2625 0 dm1 AREA=1.576e-06
D2625 n2626 0 dm1 AREA=7.881e-07
D2626 n2627 0 dm1 AREA=1.539e-06
D2627 n2628 0 dm1 AREA=4.961e-07
D2628 n2629 0 dm1 AREA=5.368e-07
D2629 n2630 0 dm1 AREA=6.427e-07
D2630 n2631 0 dm1 AREA=1.276e-06
D2631 n2632 0 dm1 AREA=6.877e-07
D2632 n2633 0 dm1 AREA=5.634e-07
D2633 n2634 0 dm1 AREA=1.264e-06
D2634 n2635 0 dm1 AREA=1.887e-06
D2635 n2636 0 dm1 AREA=2.043e-06
D2636 n2637 0 dm1 AREA=1.443e-06
D2637 n2638 0 dm1 AREA=4.173e-07
D2638 n2639 0 dm1 AREA=6.590e-07
D2639 n2640 0 dm1 AREA=2.518e-06
D2640 n2641 0 dm1 AREA=8.809e-07
D2641 n2642 0 dm1 AREA=1.543e-06
D2642 n2643 0 dm1 AREA=5.506e-07
D2643 n2644 0 dm1 AREA=1.446e-06
D2644 n2645 0 dm1 AREA=1.418e-06
D2645 n2646 0 dm1 AREA=1.815e-07
D2646 n2647 0 dm1 AREA=4.567e-07
D2647 n2648 0 dm1 AREA=9.418e-07
D2648 n2649 0 dm1 AREA=7.747e-07
D2649 n2650 0 dm1 AREA=3.421e-07
D2650 n2651 0 dm1 AREA=9.129e-07
D2651 n2652 0 dm1 AREA=2.070e-06
D2652 n2653 0 dm1 AREA=1.154e-06
D2653 n2654 0 dm1 AREA=3.262e-07
D2654 n2655 0 dm1 AREA=1.212e-06
D2655 n2656 0 dm1 AREA=7.641e-07
D2656 n2657 0 dm1 AREA=6.564e-07
D2657 n2658 0 dm1 AREA=2.673e-06
D2658 n2659 0 dm1 AREA=1.233e-06
D2659 n2660 0 dm1 AREA=7.925e-07
D2660 n2661 0 dm1 AREA=1.174e-06
D2661 n2662 0 dm1 AREA=2.343e-06
D2662 n2663 0 dm1 AREA=3.245e-07
D2663 n2664 0 dm1 AREA=4.950e-07
D2664 n2665 0 dm1 AREA=8.129e-07
D2665 n2666 0 dm1 AREA=1.073e-06
D2666 n2667 0 dm1 AREA=7.750e-07
D2667 n2668 0 dm1 AREA=2.695e-06
D2668 n2669 0 dm1 AREA=1.210e-06
D2669 n2670 0 dm1 AREA=3.770e-07
D2670 n2671 0 dm1 AREA=1.155e-06
D2671 n2672 0 dm1 AREA=6.021e-07
D2672 n2673 0 dm1 AREA=1.269e-06
D2673 n2674 0 dm1 AREA=1.171e-06
D2674 n2675 0 dm1 AREA=7.859e-07
D2675 n2676 0 dm1 AREA=3.980e-07
D2676 n2677 0 dm1 AREA=7.305e-07
D2677 n2678 0 dm1 AREA=7.919e-07
D2678 n2679 0 dm1 AREA=1.797e-06
D2679 n2680 0 dm1 AREA=9.168e-07
D2680 n2681 0 dm1 AREA=9.091e-07
D2681 n2682 0 dm1 AREA=9.946e-07
D2682 n2683 0 dm1 AREA=6.996e-07
D2683 n2684 0 dm1 AREA=1.247e-06
D2684 n2685 0 dm1 AREA=6.130e-07
D2685 n2686 0 dm1 AREA=7.127e-07
D2686 n2687 0 dm1 AREA=1.634e-06
D2687 n2688 0 dm1 AREA=1.062e-06
D2688 n2689 0 dm1 AREA=1.684e-06
D2689 n2690 0 dm1 AREA=6.999e-07
D2690 n2691 0 dm1 AREA=9.522e-07
D2691 n2692 0 dm1 AREA=1.317e-06
D2692 n2693 0 dm1 AREA=9.925e-07
D2693 n2694 0 dm1 AREA=7.051e-07
D2694 n2695 0 dm1 AREA=4.137e-07
D2695 n2696 0 dm1 AREA=2.306e-06
D2696 n2697 0 dm1 AREA=9.962e-07
D2697 n2698 0 dm1 AREA=7.819e-07
D2698 n2699 0 dm1 AREA=4.075e-07
D2699 n2700 0 dm1 AREA=9.080e-07
D2700 n2701 0 dm1 AREA=7.656e-07
D2701 n2702 0 dm1 AREA=1.282e-06
D2702 n2703 0 dm1 AREA=8.332e-07
D2703 n2704 0 dm1 AREA=8.778e-07
D2704 n2705 0 dm1 AREA=4.092e-07
D2705 n2706 0 dm1 AREA=1.038e-06
D2706 n2707 0 dm1 AREA=6.395e-07
D2707 n2708 0 dm1 AREA=1.412e-06
D2708 n2709 0 dm1 AREA=1.192e-06
D2709 n2710 0 dm1 AREA=1.638e-06
D2710 n2711 0 dm1 AREA=5.842e-07
D2711 n2712 0 dm1 AREA=1.452e-06
D2712 n2713 0 dm1 AREA=3.241e-07
D2713 n2714 0 dm1 AREA=1.218e-06
D2714 n2715 0 dm1 AREA=6.326e-07
D2715 n2716 0 dm1 AREA=1.707e-06
D2716 n2717 0 dm1 AREA=2.573e-06
D2717 n2718 0 dm1 AREA=8.477e-07
D2718 n2719 0 dm1 AREA=1.034e-06
D2719 n2720 0 dm1 AREA=1.845e-06
D2720 n2721 0 dm1 AREA=1.609e-06
D2721 n2722 0 dm1 AREA=3.801e-07
D2722 n2723 0 dm1 AREA=1.482e-07
D2723 n2724 0 dm1 AREA=6.670e-07
D2724 n2725 0 dm1 AREA=2.078e-06
D2725 n2726 0 dm1 AREA=7.247e-07
D2726 n2727 0 dm1 AREA=7.174e-07
D2727 n2728 0 dm1 AREA=4.640e-07
D2728 n2729 0 dm1 AREA=6.898e-07
D2729 n2730 0 dm1 AREA=1.095e-06
D2730 n2731 0 dm1 AREA=1.210e-06
D2731 n2732 0 dm1 AREA=1.050e-06
D2732 n2733 0 dm1 AREA=8.959e-07
D2733 n2734 0 dm1 AREA=1.628e-06
D2734 n2735 0 dm1 AREA=1.478e-06
D2735 n2736 0 dm1 AREA=1.184e-06
D2736 n2737 0 dm1 AREA=1.030e-06
D2737 n2738 0 dm1 AREA=1.347e-06
D2738 n2739 0 dm1 AREA=1.891e-06
D2739 n2740 0 dm1 AREA=8.545e-07
D2740 n2741 0 dm1 AREA=1.286e-06
D2741 n2742 0 dm1 AREA=1.030e-07
D2742 n2743 0 dm1 AREA=1.137e-06
D2743 n2744 0 dm1 AREA=1.062e-06
D2744 n2745 0 dm1 AREA=9.689e-07
D2745 n2746 0 dm1 AREA=8.505e-07
D2746 n2747 0 dm1 AREA=1.003e-06
D2747 n1 0 dm1 AREA=1.052e-06
D2748 n2749 0 dm1 AREA=1.481e-06
D2749 n2750 0 dm1 AREA=1.538e-06
D2750 n2751 0 dm1 AREA=7.363e-07
D2751 n2752 0 dm1 AREA=1.575e-06
D2752 n2753 0 dm1 AREA=1.107e-06
D2753 n2754 0 dm1 AREA=1.266e-06
D2754 n2755 0 dm1 AREA=1.026e-06
D2755 n2756 0 dm1 AREA=1.430e-06
D2756 n2757 0 dm1 AREA=1.048e-06
D2757 n2758 0 dm1 AREA=1.748e-06
D2758 n2759 0 dm1 AREA=1.931e-06
D2759 n2760 0 dm1 AREA=8.461e-07
D2760 n2761 0 dm1 AREA=7.410e-07
D2761 n2762 0 dm1 AREA=2.027e-06
D2762 n2763 0 dm1 AREA=1.547e-06
D2763 n2764 0 dm1 AREA=1.144e-06
D2764 n2765 0 dm1 AREA=3.119e-07
D2765 n2766 0 dm1 AREA=8.726e-07
D2766 n2767 0 dm1 AREA=1.141e-06
D2767 n2768 0 dm1 AREA=1.207e-06
D2768 n2769 0 dm1 AREA=1.103e-06
D2769 n2770 0 dm1 AREA=1.084e-06
D2770 n2771 0 dm1 AREA=1.061e-06
D2771 n2772 0 dm1 AREA=1.300e-06
D2772 n2773 0 dm1 AREA=8.614e-08
D2773 n2774 0 dm1 AREA=1.022e-06
D2774 n2775 0 dm1 AREA=2.185e-07
D2775 n2776 0 dm1 AREA=1.037e-06
D2776 n2777 0 dm1 AREA=3.077e-07
D2777 n2778 0 dm1 AREA=9.192e-07
D2778 n2779 0 dm1 AREA=1.286e-06
D2779 n2780 0 dm1 AREA=7.662e-07
D2780 n2781 0 dm1 AREA=1.831e-06
D2781 n2782 0 dm1 AREA=1.630e-06
D2782 n2783 0 dm1 AREA=5.734e-07
D2783 n2784 0 dm1 AREA=1.090e-06
D2784 n2785 0 dm1 AREA=1.100e-06
D2785 n2786 0 dm1 AREA=1.105e-06
D2786 n2787 0 dm1 AREA=7.726e-07
D2787 n2788 0 dm1 AREA=1.031e-06
D2788 n2789 0 dm1 AREA=7.063e-07
D2789 n2790 0 dm1 AREA=1.642e-06
D2790 n2791 0 dm1 AREA=1.397e-06
D2791 n2792 0 dm1 AREA=6.917e-07
D2792 n2793 0 dm1 AREA=4.373e-07
D2793 n2794 0 dm1 AREA=5.513e-07
D2794 n2795 0 dm1 AREA=1.522e-06
D2795 n2796 0 dm1 AREA=1.663e-06
D2796 n2797 0 dm1 AREA=1.144e-06
D2797 n2798 0 dm1 AREA=4.594e-07
D2798 n2799 0 dm1 AREA=8.332e-07
D2799 n2800 0 dm1 AREA=4.595e-07
D2800 n2801 0 dm1 AREA=4.474e-07
D2801 n2802 0 dm1 AREA=9.438e-07
D2802 n2803 0 dm1 AREA=8.881e-07
D2803 n2804 0 dm1 AREA=4.215e-07
D2804 n2805 0 dm1 AREA=2.336e-07
D2805 n2806 0 dm1 AREA=1.539e-06
D2806 n2807 0 dm1 AREA=2.331e-07
D2807 n2808 0 dm1 AREA=1.814e-06
D2808 n2809 0 dm1 AREA=8.649e-07
D2809 n2810 0 dm1 AREA=1.279e-06
D2810 n2811 0 dm1 AREA=3.409e-07
D2811 n2812 0 dm1 AREA=1.205e-06
D2812 n2813 0 dm1 AREA=1.839e-06
D2813 n2814 0 dm1 AREA=5.285e-07
D2814 n2815 0 dm1 AREA=5.084e-07
D2815 n2816 0 dm1 AREA=1.545e-06
D2816 n2817 0 dm1 AREA=1.845e-06
D2817 n2818 0 dm1 AREA=4.437e-07
D2818 n2819 0 dm1 AREA=1.622e-06
D2819 n2820 0 dm1 AREA=6.849e-07
D2820 n2821 0 dm1 AREA=4.758e-07
D2821 n2822 0 dm1 AREA=1.257e-06
D2822 n2823 0 dm1 AREA=7.162e-07
D2823 n2824 0 dm1 AREA=8.013e-07
D2824 n2825 0 dm1 AREA=2.403e-06
D2825 n2826 0 dm1 AREA=6.093e-07
D2826 n2827 0 dm1 AREA=6.514e-07
D2827 n2828 0 dm1 AREA=9.764e-07
D2828 n2829 0 dm1 AREA=1.580e-06
D2829 n2830 0 dm1 AREA=7.741e-07
D2830 n2831 0 dm1 AREA=7.442e-07
D2831 n2832 0 dm1 AREA=2.872e-06
D2832 n2833 0 dm1 AREA=1.100e-06
D2833 n2834 0 dm1 AREA=1.373e-06
D2834 n2835 0 dm1 AREA=1.425e-06
D2835 n2836 0 dm1 AREA=4.089e-07
D2836 n2837 0 dm1 AREA=1.432e-06
D2837 n2838 0 dm1 AREA=9.954e-07
D2838 n2839 0 dm1 AREA=1.586e-06
D2839 n2840 0 dm1 AREA=1.250e-06
D2840 n2841 0 dm1 AREA=9.772e-07
D2841 n2842 0 dm1 AREA=5.573e-07
D2842 n2843 0 dm1 AREA=1.189e-06
D2843 n2844 0 dm1 AREA=1.699e-06
D2844 n2845 0 dm1 AREA=1.263e-06
D2845 n2846 0 dm1 AREA=5.649e-07
D2846 n2847 0 dm1 AREA=1.424e-06
D2847 n2848 0 dm1 AREA=1.232e-06
D2848 n2849 0 dm1 AREA=8.870e-07
D2849 n2850 0 dm1 AREA=1.305e-06
D2850 n1 0 dm1 AREA=1.992e-06
D2851 n2852 0 dm1 AREA=8.638e-07
D2852 n2853 0 dm1 AREA=6.221e-07
D2853 n2854 0 dm1 AREA=1.188e-06
D2854 n2855 0 dm1 AREA=1.505e-06
D2855 n2856 0 dm1 AREA=1.845e-06
D2856 n2857 0 dm1 AREA=2.093e-06
D2857 n2858 0 dm1 AREA=1.880e-06
D2858 n2859 0 dm1 AREA=1.558e-06
D2859 n2860 0 dm1 AREA=6.558e-07
D2860 n2861 0 dm1 AREA=6.821e-07
D2861 n2862 0 dm1 AREA=7.736e-07
D2862 n2863 0 dm1 AREA=1.094e-06
D2863 n2864 0 dm1 AREA=8.240e-07
D2864 n2865 0 dm1 AREA=1.115e-06
D2865 n2866 0 dm1 AREA=6.941e-07
D2866 n2867 0 dm1 AREA=9.778e-07
D2867 n2868 0 dm1 AREA=1.121e-06
D2868 n2869 0 dm1 AREA=4.851e-07
D2869 n1 0 dm1 AREA=3.150e-07
D2870 n2871 0 dm1 AREA=1.657e-06
D2871 n2872 0 dm1 AREA=1.210e-06
D2872 n2873 0 dm1 AREA=6.970e-07
D2873 n2874 0 dm1 AREA=2.248e-06
D2874 n2875 0 dm1 AREA=6.349e-07
D2875 n2876 0 dm1 AREA=8.074e-07
D2876 n2877 0 dm1 AREA=6.018e-07
D2877 n2878 0 dm1 AREA=1.024e-06
D2878 n2879 0 dm1 AREA=6.078e-07
D2879 n2880 0 dm1 AREA=6.619e-07
D2880 n2881 0 dm1 AREA=8.128e-07
D2881 n2882 0 dm1 AREA=6.642e-07
D2882 n2883 0 dm1 AREA=1.042e-06
D2883 n2884 0 dm1 AREA=7.542e-07
D2884 n2885 0 dm1 AREA=1.413e-06
D2885 n2886 0 dm1 AREA=6.335e-07
D2886 n2887 0 dm1 AREA=1.152e-06
D2887 n2888 0 dm1 AREA=3.106e-07
D2888 n2889 0 dm1 AREA=1.306e-06
D2889 n2890 0 dm1 AREA=1.311e-06
D2890 n2891 0 dm1 AREA=7.706e-07
D2891 n2892 0 dm1 AREA=8.970e-07
D2892 n2893 0 dm1 AREA=1.658e-06
D2893 n2894 0 dm1 AREA=7.981e-07
D2894 n2895 0 dm1 AREA=9.583e-07
D2895 n2896 0 dm1 AREA=5.051e-07
D2896 n2897 0 dm1 AREA=9.950e-07
D2897 n2898 0 dm1 AREA=1.876e-06
D2898 n2899 0 dm1 AREA=1.258e-06
D2899 n2900 0 dm1 AREA=1.429e-06
D2900 n1 0 dm1 AREA=8.099e-07
D2901 n2902 0 dm1 AREA=1.261e-06
D2902 n2903 0 dm1 AREA=7.333e-07
D2903 n2904 0 dm1 AREA=5.524e-07
D2904 n2905 0 dm1 AREA=1.059e-06
D2905 n2906 0 dm1 AREA=4.484e-07
D2906 n2907 0 dm1 AREA=1.928e-06
D2907 n2908 0 dm1 AREA=8.942e-07
D2908 n2909 0 dm1 AREA=7.699e-07
D2909 n2910 0 dm1 AREA=2.160e-06
D2910 n2911 0 dm1 AREA=1.768e-06
D2911 n2912 0 dm1 AREA=7.927e-07
D2912 n2913 0 dm1 AREA=1.526e-06
D2913 n2914 0 dm1 AREA=1.288e-06
D2914 n2915 0 dm1 AREA=1.345e-07
D2915 n2916 0 dm1 AREA=1.103e-06
D2916 n2917 0 dm1 AREA=1.096e-06
D2917 n2918 0 dm1 AREA=8.873e-07
D2918 n2919 0 dm1 AREA=1.102e-06
D2919 n2920 0 dm1 AREA=8.306e-07
D2920 n2921 0 dm1 AREA=8.841e-07
D2921 n2922 0 dm1 AREA=1.040e-06
D2922 n2923 0 dm1 AREA=1.748e-06
D2923 n2924 0 dm1 AREA=4.302e-07
D2924 n2925 0 dm1 AREA=6.497e-07
D2925 n2926 0 dm1 AREA=2.193e-06
D2926 n2927 0 dm1 AREA=1.190e-06
D2927 n2928 0 dm1 AREA=1.074e-06
D2928 n2929 0 dm1 AREA=1.288e-06
D2929 n2930 0 dm1 AREA=6.538e-07
D2930 n2931 0 dm1 AREA=3.487e-07
D2931 n2932 0 dm1 AREA=7.912e-07
D2932 n2933 0 dm1 AREA=6.743e-07
D2933 n2934 0 dm1 AREA=1.114e-06
D2934 n2935 0 dm1 AREA=1.387e-06
D2935 n2936 0 dm1 AREA=6.331e-07
D2936 n2937 0 dm1 AREA=1.018e-06
D2937 n2938 0 dm1 AREA=1.276e-06
D2938 n2939 0 dm1 AREA=1.048e-06
D2939 n2940 0 dm1 AREA=7.280e-07
D2940 n2941 0 dm1 AREA=3.393e-07
D2941 n2942 0 dm1 AREA=3.274e-07
D2942 n2943 0 dm1 AREA=1.059e-06
D2943 n1 0 dm1 AREA=4.512e-07
D2944 n2945 0 dm1 AREA=1.567e-06
D2945 n2946 0 dm1 AREA=1.507e-06
D2946 n2947 0 dm1 AREA=1.287e-06
D2947 n2948 0 dm1 AREA=2.124e-06
D2948 n2949 0 dm1 AREA=8.761e-07
D2949 n2950 0 dm1 AREA=2.327e-06
D2950 n2951 0 dm1 AREA=9.287e-07
D2951 n2952 0 dm1 AREA=1.378e-06
D2952 n2953 0 dm1 AREA=6.255e-07
D2953 n2954 0 dm1 AREA=7.248e-07
D2954 n2955 0 dm1 AREA=8.598e-07
D2955 n2956 0 dm1 AREA=4.687e-07
D2956 n2957 0 dm1 AREA=3.026e-07
D2957 n2958 0 dm1 AREA=8.844e-07
D2958 n2959 0 dm1 AREA=1.487e-06
D2959 n2960 0 dm1 AREA=5.238e-07
D2960 n2961 0 dm1 AREA=1.042e-06
D2961 n2962 0 dm1 AREA=1.072e-07
D2962 n2963 0 dm1 AREA=1.044e-06
D2963 n2964 0 dm1 AREA=1.201e-06
D2964 n2965 0 dm1 AREA=4.328e-07
D2965 n2966 0 dm1 AREA=1.173e-06
D2966 n2967 0 dm1 AREA=1.057e-06
D2967 n2968 0 dm1 AREA=1.363e-06
D2968 n2969 0 dm1 AREA=1.354e-06
D2969 n2970 0 dm1 AREA=4.780e-07
D2970 n2971 0 dm1 AREA=3.578e-07
D2971 n2972 0 dm1 AREA=7.403e-07
D2972 n2973 0 dm1 AREA=7.584e-07
D2973 n2974 0 dm1 AREA=7.201e-07
D2974 n2975 0 dm1 AREA=2.446e-07
D2975 n2976 0 dm1 AREA=1.103e-06
D2976 n2977 0 dm1 AREA=1.933e-07
D2977 n2978 0 dm1 AREA=1.871e-06
D2978 n2979 0 dm1 AREA=8.287e-07
D2979 n2980 0 dm1 AREA=6.050e-07
D2980 n2981 0 dm1 AREA=6.873e-07
D2981 n2982 0 dm1 AREA=6.928e-07
D2982 n2983 0 dm1 AREA=9.135e-07
D2983 n2984 0 dm1 AREA=5.239e-07
D2984 n2985 0 dm1 AREA=8.435e-07
D2985 n2986 0 dm1 AREA=2.620e-07
D2986 n2987 0 dm1 AREA=6.226e-07
D2987 n2988 0 dm1 AREA=5.507e-07
D2988 n2989 0 dm1 AREA=7.369e-07
D2989 n2990 0 dm1 AREA=1.231e-06
D2990 n2991 0 dm1 AREA=2.365e-06
D2991 n2992 0 dm1 AREA=3.884e-07
D2992 n2993 0 dm1 AREA=1.951e-07
D2993 n2994 0 dm1 AREA=5.448e-07
D2994 n2995 0 dm1 AREA=8.526e-07
D2995 n2996 0 dm1 AREA=4.551e-07
D2996 n2997 0 dm1 AREA=1.071e-06
D2997 n2998 0 dm1 AREA=9.658e-07
D2998 n2999 0 dm1 AREA=5.638e-07
D2999 n3000 0 dm1 AREA=4.506e-07
D3000 n3001 0 dm1 AREA=1.210e-06
D3001 n3002 0 dm1 AREA=6.687e-07
D3002 n3003 0 dm1 AREA=6.748e-07
D3003 n3004 0 dm1 AREA=1.244e-06
D3004 n3005 0 dm1 AREA=4.963e-07
D3005 n3006 0 dm1 AREA=1.479e-06
D3006 n3007 0 dm1 AREA=1.400e-06
D3007 n3008 0 dm1 AREA=5.122e-07
D3008 n3009 0 dm1 AREA=7.978e-07
D3009 n3010 0 dm1 AREA=9.648e-07
D3010 n3011 0 dm1 AREA=1.890e-07
D3011 n3012 0 dm1 AREA=1.283e-06
D3012 n3013 0 dm1 AREA=3.545e-07
D3013 n3014 0 dm1 AREA=1.704e-06
D3014 n3015 0 dm1 AREA=6.319e-07
D3015 n3016 0 dm1 AREA=6.229e-07
D3016 n3017 0 dm1 AREA=9.590e-07
D3017 n3018 0 dm1 AREA=6.316e-07
D3018 n3019 0 dm1 AREA=4.826e-07
D3019 n3020 0 dm1 AREA=1.352e-06
D3020 n3021 0 dm1 AREA=5.110e-07
D3021 n3022 0 dm1 AREA=7.575e-07
D3022 n3023 0 dm1 AREA=1.141e-06
D3023 n3024 0 dm1 AREA=6.584e-07
D3024 n3025 0 dm1 AREA=1.370e-06
D3025 n3026 0 dm1 AREA=1.519e-06
D3026 n3027 0 dm1 AREA=6.546e-07
D3027 n3028 0 dm1 AREA=8.026e-07
D3028 n3029 0 dm1 AREA=7.483e-07
D3029 n3030 0 dm1 AREA=1.624e-06
D3030 n3031 0 dm1 AREA=1.389e-06
D3031 n3032 0 dm1 AREA=1.423e-06
D3032 n3033 0 dm1 AREA=1.145e-06
D3033 n3034 0 dm1 AREA=1.934e-06
D3034 n3035 0 dm1 AREA=9.968e-07
D3035 n3036 0 dm1 AREA=5.329e-07
D3036 n3037 0 dm1 AREA=2.795e-07
D3037 n3038 0 dm1 AREA=1.496e-06
D3038 n3039 0 dm1 AREA=2.314e-06
D3039 n1 0 dm1 AREA=8.598e-07
D3040 n3041 0 dm1 AREA=1.105e-06
D3041 n3042 0 dm1 AREA=6.260e-07
D3042 n3043 0 dm1 AREA=1.045e-06
D3043 n3044 0 dm1 AREA=1.040e-06
D3044 n3045 0 dm1 AREA=5.659e-07
D3045 n3046 0 dm1 AREA=6.913e-07
D3046 n3047 0 dm1 AREA=3.177e-07
D3047 n3048 0 dm1 AREA=2.671e-06
D3048 n3049 0 dm1 AREA=1.763e-07
D3049 n3050 0 dm1 AREA=1.509e-06
D3050 n3051 0 dm1 AREA=1.236e-06
D3051 n3052 0 dm1 AREA=1.944e-06
D3052 n3053 0 dm1 AREA=7.637e-07
D3053 n3054 0 dm1 AREA=4.088e-07
D3054 n3055 0 dm1 AREA=1.767e-06
D3055 n3056 0 dm1 AREA=9.397e-07
D3056 n3057 0 dm1 AREA=9.379e-07
D3057 n3058 0 dm1 AREA=4.370e-07
D3058 n3059 0 dm1 AREA=2.346e-06
D3059 n3060 0 dm1 AREA=1.004e-06
D3060 n3061 0 dm1 AREA=7.516e-07
D3061 n3062 0 dm1 AREA=1.238e-06
D3062 n3063 0 dm1 AREA=8.882e-07
D3063 n3064 0 dm1 AREA=6.832e-07
D3064 n3065 0 dm1 AREA=1.197e-06
D3065 n3066 0 dm1 AREA=7.290e-07
D3066 n3067 0 dm1 AREA=5.046e-07
D3067 n3068 0 dm1 AREA=6.312e-07
D3068 n3069 0 dm1 AREA=9.035e-07
D3069 n3070 0 dm1 AREA=2.501e-07
D3070 n3071 0 dm1 AREA=1.431e-06
D3071 n3072 0 dm1 AREA=7.918e-07
D3072 n3073 0 dm1 AREA=2.383e-07
D3073 n3074 0 dm1 AREA=8.397e-07
D3074 n3075 0 dm1 AREA=1.009e-06
D3075 n3076 0 dm1 AREA=7.869e-07
D3076 n3077 0 dm1 AREA=3.836e-07
D3077 n3078 0 dm1 AREA=1.171e-06
D3078 n3079 0 dm1 AREA=7.467e-07
D3079 n3080 0 dm1 AREA=5.089e-07
D3080 n3081 0 dm1 AREA=7.583e-07
D3081 n3082 0 dm1 AREA=1.043e-06
D3082 n3083 0 dm1 AREA=9.499e-07
D3083 n3084 0 dm1 AREA=7.259e-07
D3084 n3085 0 dm1 AREA=1.292e-06
D3085 n3086 0 dm1 AREA=3.168e-06
D3086 n3087 0 dm1 AREA=9.293e-07
D3087 n3088 0 dm1 AREA=7.963e-07
D3088 n3089 0 dm1 AREA=6.874e-07
D3089 n3090 0 dm1 AREA=5.622e-07
D3090 n3091 0 dm1 AREA=1.168e-06
D3091 n3092 0 dm1 AREA=3.077e-07
D3092 n3093 0 dm1 AREA=8.051e-07
D3093 n3094 0 dm1 AREA=7.781e-07
D3094 n3095 0 dm1 AREA=1.969e-06
D3095 n3096 0 dm1 AREA=5.864e-07
D3096 n3097 0 dm1 AREA=1.170e-06
D3097 n1 0 dm1 AREA=8.112e-07
D3098 n3099 0 dm1 AREA=9.582e-07
D3099 n3100 0 dm1 AREA=7.084e-07
D3100 n3101 0 dm1 AREA=1.219e-06
D3101 n3102 0 dm1 AREA=9.306e-07
D3102 n3103 0 dm1 AREA=1.219e-06
D3103 n3104 0 dm1 AREA=6.750e-07
D3104 n3105 0 dm1 AREA=6.249e-07
D3105 n3106 0 dm1 AREA=9.499e-07
D3106 n3107 0 dm1 AREA=1.793e-06
D3107 n3108 0 dm1 AREA=1.068e-06
D3108 n3109 0 dm1 AREA=1.819e-06
D3109 n3110 0 dm1 AREA=2.095e-06
D3110 n3111 0 dm1 AREA=2.091e-07
D3111 n1 0 dm1 AREA=6.818e-07
D3112 n3113 0 dm1 AREA=8.972e-07
D3113 n3114 0 dm1 AREA=9.313e-07
D3114 n3115 0 dm1 AREA=8.400e-07
D3115 n3116 0 dm1 AREA=2.551e-06
D3116 n3117 0 dm1 AREA=9.038e-07
D3117 n3118 0 dm1 AREA=1.205e-06
D3118 n3119 0 dm1 AREA=6.252e-07
D3119 n3120 0 dm1 AREA=1.306e-06
D3120 n3121 0 dm1 AREA=1.133e-06
D3121 n3122 0 dm1 AREA=2.951e-07
D3122 n3123 0 dm1 AREA=1.065e-06
D3123 n3124 0 dm1 AREA=3.100e-07
D3124 n3125 0 dm1 AREA=2.477e-06
D3125 n3126 0 dm1 AREA=9.202e-07
D3126 n3127 0 dm1 AREA=8.589e-07
D3127 n3128 0 dm1 AREA=8.086e-07
D3128 n3129 0 dm1 AREA=1.199e-06
D3129 n3130 0 dm1 AREA=2.096e-07
D3130 n3131 0 dm1 AREA=7.131e-07
D3131 n3132 0 dm1 AREA=5.885e-07
D3132 n3133 0 dm1 AREA=6.421e-07
D3133 n3134 0 dm1 AREA=1.557e-06
D3134 n3135 0 dm1 AREA=1.333e-06
D3135 n3136 0 dm1 AREA=4.375e-07
D3136 n3137 0 dm1 AREA=1.842e-06
D3137 n3138 0 dm1 AREA=7.350e-07
D3138 n3139 0 dm1 AREA=8.150e-07
D3139 n3140 0 dm1 AREA=3.884e-07
D3140 n3141 0 dm1 AREA=1.122e-06
D3141 n3142 0 dm1 AREA=1.264e-06
D3142 n3143 0 dm1 AREA=1.698e-06
D3143 n3144 0 dm1 AREA=9.457e-07
D3144 n3145 0 dm1 AREA=3.199e-07
D3145 n3146 0 dm1 AREA=9.039e-07
D3146 n3147 0 dm1 AREA=5.886e-07
D3147 n3148 0 dm1 AREA=1.837e-07
D3148 n3149 0 dm1 AREA=7.564e-07
D3149 n3150 0 dm1 AREA=1.911e-06
D3150 n3151 0 dm1 AREA=3.866e-07
D3151 n3152 0 dm1 AREA=5.437e-07
D3152 n3153 0 dm1 AREA=2.471e-06
D3153 n3154 0 dm1 AREA=1.527e-06
D3154 n3155 0 dm1 AREA=9.242e-07
D3155 n3156 0 dm1 AREA=2.815e-07
D3156 n3157 0 dm1 AREA=4.096e-07
D3157 n3158 0 dm1 AREA=1.195e-06
D3158 n3159 0 dm1 AREA=3.585e-07
D3159 n3160 0 dm1 AREA=1.427e-06
D3160 n3161 0 dm1 AREA=6.595e-07
D3161 n3162 0 dm1 AREA=3.674e-07
D3162 n3163 0 dm1 AREA=5.909e-07
D3163 n3164 0 dm1 AREA=1.406e-06
D3164 n3165 0 dm1 AREA=8.995e-07
D3165 n3166 0 dm1 AREA=1.434e-06
D3166 n3167 0 dm1 AREA=9.021e-07
D3167 n3168 0 dm1 AREA=4.819e-07
D3168 n1 0 dm1 AREA=5.590e-07
D3169 n3170 0 dm1 AREA=6.624e-07
D3170 n3171 0 dm1 AREA=1.604e-06
D3171 n3172 0 dm1 AREA=7.385e-07
D3172 n3173 0 dm1 AREA=1.737e-06
D3173 n3174 0 dm1 AREA=4.944e-07
D3174 n3175 0 dm1 AREA=1.518e-06
D3175 n3176 0 dm1 AREA=1.206e-06
D3176 n3177 0 dm1 AREA=9.571e-07
D3177 n3178 0 dm1 AREA=5.500e-07
D3178 n3179 0 dm1 AREA=2.243e-06
D3179 n3180 0 dm1 AREA=2.543e-06
D3180 n3181 0 dm1 AREA=1.555e-06
D3181 n3182 0 dm1 AREA=1.292e-06
D3182 n3183 0 dm1 AREA=7.488e-07
D3183 n3184 0 dm1 AREA=9.221e-07
D3184 n3185 0 dm1 AREA=1.035e-06
D3185 n3186 0 dm1 AREA=8.766e-07
D3186 n3187 0 dm1 AREA=7.471e-07
D3187 n3188 0 dm1 AREA=7.138e-07
D3188 n3189 0 dm1 AREA=1.063e-06
D3189 n3190 0 dm1 AREA=1.673e-06
D3190 n3191 0 dm1 AREA=2.002e-06
D3191 n3192 0 dm1 AREA=1.573e-06
D3192 n3193 0 dm1 AREA=5.667e-07
D3193 n3194 0 dm1 AREA=9.128e-07
D3194 n3195 0 dm1 AREA=1.175e-06
D3195 n3196 0 dm1 AREA=4.331e-07
D3196 n3197 0 dm1 AREA=4.904e-07
D3197 n3198 0 dm1 AREA=1.337e-06
D3198 n3199 0 dm1 AREA=5.878e-07
D3199 n3200 0 dm1 AREA=6.193e-07
D3200 n3201 0 dm1 AREA=9.687e-07
D3201 n3202 0 dm1 AREA=5.935e-07
D3202 n3203 0 dm1 AREA=1.650e-06
D3203 n3204 0 dm1 AREA=8.513e-07
D3204 n3205 0 dm1 AREA=3.276e-06
D3205 n3206 0 dm1 AREA=9.200e-07
D3206 n3207 0 dm1 AREA=2.237e-07
D3207 n3208 0 dm1 AREA=1.623e-06
D3208 n3209 0 dm1 AREA=2.144e-06
D3209 n3210 0 dm1 AREA=7.932e-07
D3210 n3211 0 dm1 AREA=5.045e-07
D3211 n3212 0 dm1 AREA=1.642e-06
D3212 n3213 0 dm1 AREA=1.706e-06
D3213 n3214 0 dm1 AREA=1.646e-06
D3214 n3215 0 dm1 AREA=7.743e-07
D3215 n3216 0 dm1 AREA=1.050e-06
D3216 n3217 0 dm1 AREA=6.950e-07
D3217 n3218 0 dm1 AREA=1.650e-06
D3218 n3219 0 dm1 AREA=9.950e-07
D3219 n3220 0 dm1 AREA=7.357e-07
D3220 n3221 0 dm1 AREA=9.130e-07
D3221 n3222 0 dm1 AREA=1.256e-06
D3222 n3223 0 dm1 AREA=9.531e-07
D3223 n1 0 dm1 AREA=1.541e-06
D3224 n3225 0 dm1 AREA=1.068e-06
D3225 n3226 0 dm1 AREA=1.586e-06
D3226 n3227 0 dm1 AREA=3.361e-07
D3227 n3228 0 dm1 AREA=1.186e-06
D3228 n3229 0 dm1 AREA=4.805e-07
D3229 n3230 0 dm1 AREA=1.298e-06
D3230 n3231 0 dm1 AREA=1.017e-06
D3231 n3232 0 dm1 AREA=3.678e-07
D3232 n3233 0 dm1 AREA=1.294e-06
D3233 n3234 0 dm1 AREA=6.979e-07
D3234 n3235 0 dm1 AREA=5.370e-07
D3235 n3236 0 dm1 AREA=2.337e-06
D3236 n3237 0 dm1 AREA=9.499e-07
D3237 n3238 0 dm1 AREA=1.205e-06
D3238 n3239 0 dm1 AREA=3.072e-07
D3239 n3240 0 dm1 AREA=1.185e-06
D3240 n3241 0 dm1 AREA=5.544e-07
D3241 n3242 0 dm1 AREA=1.182e-06
D3242 n3243 0 dm1 AREA=1.484e-06
D3243 n3244 0 dm1 AREA=4.547e-07
D3244 n3245 0 dm1 AREA=1.330e-06
D3245 n3246 0 dm1 AREA=1.250e-06
D3246 n3247 0 dm1 AREA=6.190e-07
D3247 n3248 0 dm1 AREA=1.735e-06
D3248 n3249 0 dm1 AREA=8.484e-07
D3249 n3250 0 dm1 AREA=8.984e-07
D3250 n3251 0 dm1 AREA=1.075e-06
D3251 n3252 0 dm1 AREA=1.981e-06
D3252 n3253 0 dm1 AREA=2.834e-07
D3253 n3254 0 dm1 AREA=7.942e-07
D3254 n3255 0 dm1 AREA=1.821e-06
D3255 n3256 0 dm1 AREA=1.178e-06
D3256 n3257 0 dm1 AREA=1.245e-06
D3257 n3258 0 dm1 AREA=1.262e-06
D3258 n3259 0 dm1 AREA=6.216e-07
D3259 n3260 0 dm1 AREA=1.317e-06
D3260 n3261 0 dm1 AREA=1.943e-06
D3261 n3262 0 dm1 AREA=1.014e-06
D3262 n3263 0 dm1 AREA=7.745e-07
D3263 n3264 0 dm1 AREA=8.424e-07
D3264 n3265 0 dm1 AREA=1.671e-06
D3265 n3266 0 dm1 AREA=9.595e-07
D3266 n3267 0 dm1 AREA=1.811e-06
D3267 n3268 0 dm1 AREA=3.827e-07
D3268 n3269 0 dm1 AREA=9.709e-07
D3269 n3270 0 dm1 AREA=8.924e-07
D3270 n3271 0 dm1 AREA=1.354e-06
D3271 n3272 0 dm1 AREA=1.102e-06
D3272 n3273 0 dm1 AREA=4.783e-07
D3273 n3274 0 dm1 AREA=1.675e-06
D3274 n3275 0 dm1 AREA=3.001e-07
D3275 n3276 0 dm1 AREA=1.166e-06
D3276 n3277 0 dm1 AREA=1.204e-06
D3277 n3278 0 dm1 AREA=1.913e-06
D3278 n3279 0 dm1 AREA=1.475e-06
D3279 n3280 0 dm1 AREA=5.593e-07
D3280 n3281 0 dm1 AREA=3.517e-07
D3281 n3282 0 dm1 AREA=4.707e-07
D3282 n3283 0 dm1 AREA=1.963e-06
D3283 n3284 0 dm1 AREA=8.975e-07
D3284 n3285 0 dm1 AREA=1.219e-06
D3285 n3286 0 dm1 AREA=8.695e-07
D3286 n3287 0 dm1 AREA=1.220e-06
D3287 n3288 0 dm1 AREA=1.005e-06
D3288 n3289 0 dm1 AREA=1.195e-06
D3289 n3290 0 dm1 AREA=1.116e-06
D3290 n3291 0 dm1 AREA=3.205e-07
D3291 n3292 0 dm1 AREA=3.278e-07
D3292 n3293 0 dm1 AREA=4.874e-07
D3293 n3294 0 dm1 AREA=8.093e-07
D3294 n3295 0 dm1 AREA=6.401e-07
D3295 n3296 0 dm1 AREA=1.014e-06
D3296 n3297 0 dm1 AREA=4.697e-07
D3297 n3298 0 dm1 AREA=9.805e-07
D3298 n3299 0 dm1 AREA=2.225e-07
D3299 n3300 0 dm1 AREA=1.319e-06
D3300 n3301 0 dm1 AREA=1.168e-06
D3301 n3302 0 dm1 AREA=1.077e-06
D3302 n3303 0 dm1 AREA=8.574e-07
D3303 n3304 0 dm1 AREA=1.037e-06
D3304 n3305 0 dm1 AREA=9.708e-07
D3305 n3306 0 dm1 AREA=8.413e-07
D3306 n3307 0 dm1 AREA=6.561e-07
D3307 n3308 0 dm1 AREA=1.410e-06
D3308 n1 0 dm1 AREA=4.512e-07
D3309 n3310 0 dm1 AREA=3.962e-07
D3310 n3311 0 dm1 AREA=1.168e-06
D3311 n3312 0 dm1 AREA=1.559e-06
D3312 n3313 0 dm1 AREA=1.205e-06
D3313 n3314 0 dm1 AREA=6.442e-07
D3314 n3315 0 dm1 AREA=9.995e-07
D3315 n3316 0 dm1 AREA=7.204e-07
D3316 n3317 0 dm1 AREA=1.118e-06
D3317 n3318 0 dm1 AREA=8.018e-07
D3318 n3319 0 dm1 AREA=1.487e-06
D3319 n3320 0 dm1 AREA=1.948e-07
D3320 n3321 0 dm1 AREA=1.329e-06
D3321 n3322 0 dm1 AREA=1.658e-06
D3322 n3323 0 dm1 AREA=3.894e-07
D3323 n3324 0 dm1 AREA=1.165e-06
D3324 n3325 0 dm1 AREA=7.764e-07
D3325 n3326 0 dm1 AREA=2.292e-06
D3326 n3327 0 dm1 AREA=1.103e-06
D3327 n3328 0 dm1 AREA=6.603e-07
D3328 n3329 0 dm1 AREA=3.853e-07
D3329 n3330 0 dm1 AREA=5.541e-07
D3330 n3331 0 dm1 AREA=7.181e-07
D3331 n3332 0 dm1 AREA=1.374e-06
D3332 n3333 0 dm1 AREA=6.538e-07
D3333 n3334 0 dm1 AREA=1.214e-06
D3334 n3335 0 dm1 AREA=1.400e-06
D3335 n3336 0 dm1 AREA=1.720e-07
D3336 n3337 0 dm1 AREA=7.276e-07
D3337 n3338 0 dm1 AREA=6.675e-07
D3338 n3339 0 dm1 AREA=1.317e-06
D3339 n3340 0 dm1 AREA=4.944e-07
D3340 n3341 0 dm1 AREA=2.774e-07
D3341 n3342 0 dm1 AREA=1.085e-06
D3342 n3343 0 dm1 AREA=5.248e-07
D3343 n3344 0 dm1 AREA=1.442e-06
D3344 n3345 0 dm1 AREA=7.903e-07
D3345 n3346 0 dm1 AREA=8.975e-07
D3346 n3347 0 dm1 AREA=3.263e-07
D3347 n3348 0 dm1 AREA=8.164e-07
D3348 n3349 0 dm1 AREA=1.577e-06
D3349 n3350 0 dm1 AREA=1.438e-06
D3350 n3351 0 dm1 AREA=1.158e-06
D3351 n3352 0 dm1 AREA=1.738e-06
D3352 n3353 0 dm1 AREA=2.105e-06
D3353 n3354 0 dm1 AREA=1.195e-06
D3354 n3355 0 dm1 AREA=8.934e-07
D3355 n3356 0 dm1 AREA=6.286e-07
D3356 n3357 0 dm1 AREA=1.577e-06
D3357 n3358 0 dm1 AREA=1.255e-06
D3358 n3359 0 dm1 AREA=1.531e-06
D3359 n3360 0 dm1 AREA=1.168e-06
D3360 n3361 0 dm1 AREA=6.232e-07
D3361 n3362 0 dm1 AREA=6.038e-07
D3362 n3363 0 dm1 AREA=2.118e-07
D3363 n3364 0 dm1 AREA=4.762e-07
D3364 n3365 0 dm1 AREA=3.399e-06
D3365 n3366 0 dm1 AREA=7.991e-07
D3366 n3367 0 dm1 AREA=7.441e-07
D3367 n3368 0 dm1 AREA=1.105e-06
D3368 n3369 0 dm1 AREA=6.136e-07
D3369 n3370 0 dm1 AREA=9.790e-07
D3370 n3371 0 dm1 AREA=1.709e-06
D3371 n3372 0 dm1 AREA=1.329e-06
D3372 n3373 0 dm1 AREA=5.898e-07
D3373 n3374 0 dm1 AREA=6.460e-07
D3374 n3375 0 dm1 AREA=9.353e-07
D3375 n3376 0 dm1 AREA=4.603e-07
D3376 n3377 0 dm1 AREA=4.813e-07
D3377 n3378 0 dm1 AREA=1.112e-06
D3378 n3379 0 dm1 AREA=5.421e-07
D3379 n3380 0 dm1 AREA=9.532e-07
D3380 n3381 0 dm1 AREA=9.892e-07
D3381 n3382 0 dm1 AREA=1.011e-06
D3382 n3383 0 dm1 AREA=5.068e-07
D3383 n3384 0 dm1 AREA=8.408e-07
D3384 n3385 0 dm1 AREA=1.070e-06
D3385 n3386 0 dm1 AREA=2.150e-06
D3386 n3387 0 dm1 AREA=2.400e-06
D3387 n3388 0 dm1 AREA=1.893e-06
D3388 n3389 0 dm1 AREA=2.107e-07
D3389 n1 0 dm1 AREA=1.303e-06
D3390 n3391 0 dm1 AREA=8.001e-07
D3391 n3392 0 dm1 AREA=8.373e-07
D3392 n3393 0 dm1 AREA=4.289e-07
D3393 n3394 0 dm1 AREA=8.073e-07
D3394 n3395 0 dm1 AREA=5.557e-07
D3395 n3396 0 dm1 AREA=4.272e-07
D3396 n3397 0 dm1 AREA=9.078e-07
D3397 n3398 0 dm1 AREA=1.197e-06
D3398 n3399 0 dm1 AREA=1.134e-06
D3399 n3400 0 dm1 AREA=9.934e-07
D3400 n3401 0 dm1 AREA=7.343e-07
D3401 n3402 0 dm1 AREA=6.339e-07
D3402 n3403 0 dm1 AREA=1.073e-06
D3403 n3404 0 dm1 AREA=5.057e-07
D3404 n3405 0 dm1 AREA=4.601e-07
D3405 n3406 0 dm1 AREA=4.014e-07
D3406 n3407 0 dm1 AREA=1.278e-06
D3407 n3408 0 dm1 AREA=6.991e-07
D3408 n3409 0 dm1 AREA=5.256e-07
D3409 n3410 0 dm1 AREA=4.602e-07
D3410 n3411 0 dm1 AREA=6.855e-07
D3411 n3412 0 dm1 AREA=8.425e-07
D3412 n3413 0 dm1 AREA=1.047e-06
D3413 n3414 0 dm1 AREA=6.204e-07
D3414 n3415 0 dm1 AREA=5.029e-07
D3415 n3416 0 dm1 AREA=9.759e-07
D3416 n3417 0 dm1 AREA=2.203e-06
D3417 n3418 0 dm1 AREA=2.839e-06
D3418 n3419 0 dm1 AREA=9.128e-07
D3419 n3420 0 dm1 AREA=6.342e-07
D3420 n3421 0 dm1 AREA=9.046e-07
D3421 n3422 0 dm1 AREA=1.046e-06
D3422 n3423 0 dm1 AREA=1.956e-06
D3423 n3424 0 dm1 AREA=5.614e-07
D3424 n3425 0 dm1 AREA=8.055e-07
D3425 n3426 0 dm1 AREA=6.947e-07
D3426 n3427 0 dm1 AREA=8.997e-07
D3427 n3428 0 dm1 AREA=8.377e-07
D3428 n3429 0 dm1 AREA=6.291e-07
D3429 n3430 0 dm1 AREA=9.511e-07
D3430 n3431 0 dm1 AREA=6.853e-07
D3431 n3432 0 dm1 AREA=4.940e-07
D3432 n3433 0 dm1 AREA=9.948e-07
D3433 n3434 0 dm1 AREA=1.039e-06
D3434 n3435 0 dm1 AREA=6.267e-07
D3435 n3436 0 dm1 AREA=9.085e-07
D3436 n3437 0 dm1 AREA=1.018e-06
D3437 n3438 0 dm1 AREA=1.868e-06
D3438 n3439 0 dm1 AREA=1.389e-06
D3439 n3440 0 dm1 AREA=1.234e-06
D3440 n3441 0 dm1 AREA=1.280e-06
D3441 n3442 0 dm1 AREA=5.854e-07
D3442 n3443 0 dm1 AREA=3.899e-07
D3443 n3444 0 dm1 AREA=8.201e-07
D3444 n3445 0 dm1 AREA=2.094e-06
D3445 n3446 0 dm1 AREA=1.419e-06
D3446 n3447 0 dm1 AREA=1.547e-06
D3447 n3448 0 dm1 AREA=6.824e-07
D3448 n3449 0 dm1 AREA=1.199e-06
D3449 n3450 0 dm1 AREA=1.235e-06
D3450 n3451 0 dm1 AREA=1.154e-06
D3451 n3452 0 dm1 AREA=1.001e-06
D3452 n3453 0 dm1 AREA=1.270e-06
D3453 n3454 0 dm1 AREA=1.179e-06
D3454 n3455 0 dm1 AREA=1.038e-06
D3455 n3456 0 dm1 AREA=8.039e-07
D3456 n3457 0 dm1 AREA=1.072e-06
D3457 n3458 0 dm1 AREA=1.196e-06
D3458 n3459 0 dm1 AREA=6.508e-07
D3459 n3460 0 dm1 AREA=1.262e-06
D3460 n3461 0 dm1 AREA=1.130e-06
D3461 n3462 0 dm1 AREA=1.067e-06
D3462 n3463 0 dm1 AREA=2.235e-07
D3463 n3464 0 dm1 AREA=9.599e-07
D3464 n3465 0 dm1 AREA=1.863e-06
D3465 n3466 0 dm1 AREA=1.197e-06
D3466 n3467 0 dm1 AREA=5.227e-07
D3467 n3468 0 dm1 AREA=1.373e-06
D3468 n3469 0 dm1 AREA=1.440e-06
D3469 n3470 0 dm1 AREA=1.922e-06
D3470 n3471 0 dm1 AREA=1.047e-06
D3471 n3472 0 dm1 AREA=9.311e-07
D3472 n3473 0 dm1 AREA=5.262e-07
D3473 n3474 0 dm1 AREA=5.634e-07
D3474 n3475 0 dm1 AREA=4.553e-07
D3475 n3476 0 dm1 AREA=6.511e-07
D3476 n3477 0 dm1 AREA=8.479e-07
D3477 n3478 0 dm1 AREA=4.146e-07
D3478 n3479 0 dm1 AREA=3.726e-07
D3479 n3480 0 dm1 AREA=1.159e-06
D3480 n3481 0 dm1 AREA=4.782e-07
D3481 n3482 0 dm1 AREA=2.054e-06
D3482 n3483 0 dm1 AREA=1.548e-06
D3483 n3484 0 dm1 AREA=1.712e-07
D3484 n3485 0 dm1 AREA=1.472e-07
D3485 n3486 0 dm1 AREA=7.066e-07
D3486 n3487 0 dm1 AREA=1.656e-06
D3487 n3488 0 dm1 AREA=1.123e-06
D3488 n3489 0 dm1 AREA=6.639e-07
D3489 n3490 0 dm1 AREA=1.095e-06
D3490 n3491 0 dm1 AREA=1.486e-06
D3491 n3492 0 dm1 AREA=1.221e-06
D3492 n1 0 dm1 AREA=8.609e-07
D3493 n3494 0 dm1 AREA=1.991e-06
D3494 n3495 0 dm1 AREA=3.499e-07
D3495 n3496 0 dm1 AREA=6.659e-07
D3496 n3497 0 dm1 AREA=1.197e-06
D3497 n3498 0 dm1 AREA=7.153e-07
D3498 n3499 0 dm1 AREA=4.466e-07
D3499 n3500 0 dm1 AREA=9.738e-07
D3500 n3501 0 dm1 AREA=1.068e-06
D3501 n3502 0 dm1 AREA=6.088e-07
D3502 n3503 0 dm1 AREA=1.255e-06
D3503 n3504 0 dm1 AREA=1.329e-06
D3504 n3505 0 dm1 AREA=1.168e-06
D3505 n3506 0 dm1 AREA=4.340e-07
D3506 n3507 0 dm1 AREA=5.992e-07
D3507 n3508 0 dm1 AREA=1.200e-06
D3508 n3509 0 dm1 AREA=1.564e-06
D3509 n3510 0 dm1 AREA=7.002e-07
D3510 n3511 0 dm1 AREA=1.360e-06
D3511 n3512 0 dm1 AREA=1.663e-07
D3512 n3513 0 dm1 AREA=8.436e-07
D3513 n3514 0 dm1 AREA=1.075e-06
D3514 n3515 0 dm1 AREA=1.701e-06
D3515 n3516 0 dm1 AREA=1.102e-06
D3516 n3517 0 dm1 AREA=1.729e-06
D3517 n3518 0 dm1 AREA=1.079e-06
D3518 n3519 0 dm1 AREA=8.206e-07
D3519 n3520 0 dm1 AREA=4.018e-07
D3520 n3521 0 dm1 AREA=4.024e-07
D3521 n3522 0 dm1 AREA=9.371e-07
D3522 n3523 0 dm1 AREA=1.169e-06
D3523 n3524 0 dm1 AREA=5.914e-07
D3524 n3525 0 dm1 AREA=8.012e-07
D3525 n3526 0 dm1 AREA=6.652e-07
D3526 n3527 0 dm1 AREA=6.790e-07
D3527 n3528 0 dm1 AREA=1.091e-06
D3528 n3529 0 dm1 AREA=1.311e-06
D3529 n3530 0 dm1 AREA=1.367e-06
D3530 n3531 0 dm1 AREA=1.117e-06
D3531 n3532 0 dm1 AREA=6.338e-07
D3532 n3533 0 dm1 AREA=4.755e-07
D3533 n3534 0 dm1 AREA=1.025e-06
D3534 n3535 0 dm1 AREA=1.193e-06
D3535 n3536 0 dm1 AREA=1.101e-06
D3536 n3537 0 dm1 AREA=1.503e-06
D3537 n3538 0 dm1 AREA=5.089e-07
D3538 n3539 0 dm1 AREA=1.694e-06
D3539 n3540 0 dm1 AREA=5.611e-07
D3540 n3541 0 dm1 AREA=9.565e-07
D3541 n3542 0 dm1 AREA=3.052e-07
D3542 n3543 0 dm1 AREA=1.661e-06
D3543 n3544 0 dm1 AREA=4.717e-07
D3544 n3545 0 dm1 AREA=5.777e-07
D3545 n3546 0 dm1 AREA=1.097e-06
D3546 n3547 0 dm1 AREA=1.057e-06
D3547 n3548 0 dm1 AREA=1.149e-06
D3548 n3549 0 dm1 AREA=8.004e-07
D3549 n3550 0 dm1 AREA=3.880e-07
D3550 n3551 0 dm1 AREA=8.372e-07
D3551 n3552 0 dm1 AREA=1.303e-06
D3552 n3553 0 dm1 AREA=9.362e-07
D3553 n3554 0 dm1 AREA=1.474e-06
D3554 n3555 0 dm1 AREA=9.057e-07
D3555 n3556 0 dm1 AREA=1.265e-06
D3556 n3557 0 dm1 AREA=1.295e-06
D3557 n3558 0 dm1 AREA=1.297e-06
D3558 n3559 0 dm1 AREA=8.131e-07
D3559 n3560 0 dm1 AREA=5.561e-07
D3560 n3561 0 dm1 AREA=9.633e-07
D3561 n3562 0 dm1 AREA=1.347e-06
D3562 n3563 0 dm1 AREA=3.811e-07
D3563 n3564 0 dm1 AREA=1.004e-06
D3564 n3565 0 dm1 AREA=1.225e-06
D3565 n3566 0 dm1 AREA=6.895e-07
D3566 n3567 0 dm1 AREA=9.378e-07
D3567 n3568 0 dm1 AREA=8.345e-07
D3568 n3569 0 dm1 AREA=6.322e-07
D3569 n3570 0 dm1 AREA=1.114e-06
D3570 n3571 0 dm1 AREA=1.205e-06
D3571 n3572 0 dm1 AREA=1.251e-06
D3572 n3573 0 dm1 AREA=2.637e-07
D3573 n3574 0 dm1 AREA=4.824e-07
D3574 n3575 0 dm1 AREA=6.628e-07
D3575 n3576 0 dm1 AREA=9.062e-07
D3576 n3577 0 dm1 AREA=9.680e-07
D3577 n3578 0 dm1 AREA=6.220e-07
D3578 n3579 0 dm1 AREA=1.318e-06
D3579 n3580 0 dm1 AREA=1.269e-06
D3580 n3581 0 dm1 AREA=8.664e-07
D3581 n3582 0 dm1 AREA=9.764e-07
D3582 n3583 0 dm1 AREA=2.039e-07
D3583 n3584 0 dm1 AREA=1.362e-06
D3584 n3585 0 dm1 AREA=1.858e-06
D3585 n3586 0 dm1 AREA=6.656e-07
D3586 n3587 0 dm1 AREA=8.165e-07
D3587 n3588 0 dm1 AREA=7.933e-07
D3588 n3589 0 dm1 AREA=1.183e-06
D3589 n3590 0 dm1 AREA=1.706e-06
D3590 n3591 0 dm1 AREA=1.444e-06
D3591 n3592 0 dm1 AREA=1.495e-06
D3592 n3593 0 dm1 AREA=1.759e-06
D3593 n3594 0 dm1 AREA=1.413e-06
D3594 n3595 0 dm1 AREA=4.286e-07
D3595 n3596 0 dm1 AREA=1.285e-06
D3596 n3597 0 dm1 AREA=2.806e-06
D3597 n3598 0 dm1 AREA=8.495e-07
D3598 n3599 0 dm1 AREA=1.073e-06
D3599 n3600 0 dm1 AREA=8.035e-07
D3600 n3601 0 dm1 AREA=6.542e-07
D3601 n3602 0 dm1 AREA=6.276e-07
D3602 n3603 0 dm1 AREA=1.561e-06
D3603 n3604 0 dm1 AREA=9.641e-07
D3604 n3605 0 dm1 AREA=8.403e-07
D3605 n3606 0 dm1 AREA=1.072e-06
D3606 n3607 0 dm1 AREA=1.011e-06
D3607 n3608 0 dm1 AREA=8.701e-07
D3608 n3609 0 dm1 AREA=1.191e-06
D3609 n3610 0 dm1 AREA=8.743e-07
D3610 n3611 0 dm1 AREA=2.543e-07
D3611 n3612 0 dm1 AREA=1.302e-06
D3612 n3613 0 dm1 AREA=4.432e-07
D3613 n3614 0 dm1 AREA=1.542e-07
D3614 n3615 0 dm1 AREA=2.613e-06
D3615 n3616 0 dm1 AREA=3.373e-07
D3616 n3617 0 dm1 AREA=6.871e-07
D3617 n3618 0 dm1 AREA=7.901e-07
D3618 n3619 0 dm1 AREA=1.175e-06
D3619 n3620 0 dm1 AREA=5.834e-07
D3620 n3621 0 dm1 AREA=5.379e-07
D3621 n3622 0 dm1 AREA=6.775e-07
D3622 n3623 0 dm1 AREA=6.263e-07
D3623 n3624 0 dm1 AREA=1.496e-06
D3624 n3625 0 dm1 AREA=1.579e-06
D3625 n3626 0 dm1 AREA=2.819e-07
D3626 n3627 0 dm1 AREA=1.627e-06
D3627 n3628 0 dm1 AREA=3.135e-07
D3628 n3629 0 dm1 AREA=3.588e-07
D3629 n3630 0 dm1 AREA=6.379e-07
D3630 n3631 0 dm1 AREA=5.745e-07
D3631 n3632 0 dm1 AREA=3.903e-07
D3632 n3633 0 dm1 AREA=1.052e-06
D3633 n3634 0 dm1 AREA=2.176e-06
D3634 n3635 0 dm1 AREA=1.286e-06
D3635 n3636 0 dm1 AREA=9.360e-07
D3636 n3637 0 dm1 AREA=5.289e-07
D3637 n3638 0 dm1 AREA=9.777e-07
D3638 n3639 0 dm1 AREA=1.263e-06
D3639 n3640 0 dm1 AREA=6.518e-07
D3640 n3641 0 dm1 AREA=1.013e-06
D3641 n3642 0 dm1 AREA=9.030e-07
D3642 n3643 0 dm1 AREA=1.000e-06
D3643 n3644 0 dm1 AREA=1.066e-06
D3644 n3645 0 dm1 AREA=9.494e-07
D3645 n3646 0 dm1 AREA=8.755e-07
D3646 n3647 0 dm1 AREA=1.094e-06
D3647 n3648 0 dm1 AREA=1.267e-06
D3648 n3649 0 dm1 AREA=7.411e-07
D3649 n3650 0 dm1 AREA=8.164e-07
D3650 n3651 0 dm1 AREA=1.320e-06
D3651 n3652 0 dm1 AREA=9.501e-07
D3652 n3653 0 dm1 AREA=8.165e-07
D3653 n3654 0 dm1 AREA=5.036e-07
D3654 n3655 0 dm1 AREA=8.015e-07
D3655 n3656 0 dm1 AREA=1.366e-06
D3656 n3657 0 dm1 AREA=8.999e-07
D3657 n3658 0 dm1 AREA=5.180e-07
D3658 n3659 0 dm1 AREA=3.751e-07
D3659 n3660 0 dm1 AREA=4.227e-07
D3660 n3661 0 dm1 AREA=4.283e-07
D3661 n3662 0 dm1 AREA=1.656e-06
D3662 n3663 0 dm1 AREA=5.555e-07
D3663 n3664 0 dm1 AREA=1.055e-06
D3664 n3665 0 dm1 AREA=9.698e-07
D3665 n3666 0 dm1 AREA=7.029e-07
D3666 n3667 0 dm1 AREA=2.396e-06
D3667 n3668 0 dm1 AREA=8.458e-07
D3668 n3669 0 dm1 AREA=1.745e-06
D3669 n3670 0 dm1 AREA=9.766e-07
D3670 n3671 0 dm1 AREA=1.787e-06
D3671 n3672 0 dm1 AREA=5.659e-07
D3672 n3673 0 dm1 AREA=1.170e-06
D3673 n3674 0 dm1 AREA=7.940e-07
D3674 n3675 0 dm1 AREA=8.162e-07
D3675 n3676 0 dm1 AREA=8.300e-07
D3676 n3677 0 dm1 AREA=7.528e-07
D3677 n3678 0 dm1 AREA=1.633e-06
D3678 n3679 0 dm1 AREA=8.258e-07
D3679 n3680 0 dm1 AREA=1.171e-06
D3680 n3681 0 dm1 AREA=6.355e-07
D3681 n3682 0 dm1 AREA=3.364e-07
D3682 n3683 0 dm1 AREA=2.264e-07
D3683 n3684 0 dm1 AREA=7.555e-07
D3684 n3685 0 dm1 AREA=1.155e-06
D3685 n3686 0 dm1 AREA=2.897e-07
D3686 n3687 0 dm1 AREA=6.324e-07
D3687 n3688 0 dm1 AREA=2.077e-07
D3688 n3689 0 dm1 AREA=1.111e-06
D3689 n3690 0 dm1 AREA=8.593e-07
D3690 n3691 0 dm1 AREA=1.691e-06
D3691 n3692 0 dm1 AREA=3.398e-07
D3692 n3693 0 dm1 AREA=1.509e-06
D3693 n3694 0 dm1 AREA=8.456e-07
D3694 n3695 0 dm1 AREA=1.476e-06
D3695 n3696 0 dm1 AREA=2.403e-06
D3696 n3697 0 dm1 AREA=1.030e-06
D3697 n3698 0 dm1 AREA=2.367e-07
D3698 n3699 0 dm1 AREA=9.434e-07
D3699 n3700 0 dm1 AREA=7.311e-07
D3700 n3701 0 dm1 AREA=8.188e-07
D3701 n3702 0 dm1 AREA=4.997e-07
D3702 n3703 0 dm1 AREA=1.271e-06
D3703 n3704 0 dm1 AREA=6.334e-07
D3704 n3705 0 dm1 AREA=1.029e-06
D3705 n3706 0 dm1 AREA=3.424e-07
D3706 n3707 0 dm1 AREA=8.759e-07
D3707 n3708 0 dm1 AREA=6.741e-07
D3708 n3709 0 dm1 AREA=2.050e-06
D3709 n3710 0 dm1 AREA=8.945e-07
D3710 n3711 0 dm1 AREA=9.582e-07
D3711 n3712 0 dm1 AREA=8.029e-07
D3712 n3713 0 dm1 AREA=1.159e-06
D3713 n3714 0 dm1 AREA=5.949e-07
D3714 n3715 0 dm1 AREA=2.587e-06
D3715 n3716 0 dm1 AREA=1.456e-06
D3716 n3717 0 dm1 AREA=2.625e-07
D3717 n3718 0 dm1 AREA=2.430e-06
D3718 n3719 0 dm1 AREA=7.714e-07
D3719 n3720 0 dm1 AREA=8.536e-07
D3720 n3721 0 dm1 AREA=2.497e-06
D3721 n3722 0 dm1 AREA=5.500e-07
D3722 n3723 0 dm1 AREA=1.118e-06
D3723 n3724 0 dm1 AREA=1.922e-06
D3724 n3725 0 dm1 AREA=4.843e-07
D3725 n3726 0 dm1 AREA=1.442e-06
D3726 n3727 0 dm1 AREA=1.487e-06
D3727 n3728 0 dm1 AREA=4.958e-07
D3728 n3729 0 dm1 AREA=8.478e-07
D3729 n3730 0 dm1 AREA=7.523e-07
D3730 n3731 0 dm1 AREA=1.085e-06
D3731 n3732 0 dm1 AREA=6.988e-07
D3732 n3733 0 dm1 AREA=6.509e-07
D3733 n3734 0 dm1 AREA=2.483e-06
D3734 n3735 0 dm1 AREA=1.758e-06
D3735 n3736 0 dm1 AREA=9.130e-07
D3736 n3737 0 dm1 AREA=4.440e-07
D3737 n3738 0 dm1 AREA=9.703e-07
D3738 n3739 0 dm1 AREA=6.794e-07
D3739 n3740 0 dm1 AREA=5.190e-07
D3740 n3741 0 dm1 AREA=1.230e-06
D3741 n3742 0 dm1 AREA=1.347e-06
D3742 n3743 0 dm1 AREA=2.322e-07
D3743 n3744 0 dm1 AREA=3.729e-07
D3744 n3745 0 dm1 AREA=7.807e-07
D3745 n3746 0 dm1 AREA=5.555e-07
D3746 n3747 0 dm1 AREA=1.194e-06
D3747 n3748 0 dm1 AREA=1.160e-06
D3748 n3749 0 dm1 AREA=2.453e-06
D3749 n3750 0 dm1 AREA=6.547e-07
D3750 n3751 0 dm1 AREA=1.437e-07
D3751 n3752 0 dm1 AREA=1.727e-06
D3752 n3753 0 dm1 AREA=1.105e-06
D3753 n3754 0 dm1 AREA=1.151e-06
D3754 n3755 0 dm1 AREA=7.075e-07
D3755 n3756 0 dm1 AREA=4.709e-07
D3756 n3757 0 dm1 AREA=6.466e-07
D3757 n3758 0 dm1 AREA=9.032e-07
D3758 n3759 0 dm1 AREA=1.097e-06
D3759 n3760 0 dm1 AREA=4.878e-07
D3760 n3761 0 dm1 AREA=1.006e-06
D3761 n3762 0 dm1 AREA=6.838e-07
D3762 n3763 0 dm1 AREA=1.582e-06
D3763 n3764 0 dm1 AREA=7.305e-07
D3764 n3765 0 dm1 AREA=3.445e-07
D3765 n3766 0 dm1 AREA=3.228e-07
D3766 n3767 0 dm1 AREA=1.579e-06
D3767 n3768 0 dm1 AREA=1.870e-06
D3768 n3769 0 dm1 AREA=1.546e-06
D3769 n3770 0 dm1 AREA=1.247e-06
D3770 n3771 0 dm1 AREA=5.771e-07
D3771 n3772 0 dm1 AREA=8.279e-07
D3772 n3773 0 dm1 AREA=6.017e-07
D3773 n3774 0 dm1 AREA=1.147e-06
D3774 n3775 0 dm1 AREA=2.479e-06
D3775 n3776 0 dm1 AREA=1.225e-06
D3776 n3777 0 dm1 AREA=3.666e-06
D3777 n3778 0 dm1 AREA=1.502e-06
D3778 n3779 0 dm1 AREA=4.181e-07
D3779 n3780 0 dm1 AREA=1.308e-06
D3780 n3781 0 dm1 AREA=2.553e-06
D3781 n3782 0 dm1 AREA=1.705e-06
D3782 n3783 0 dm1 AREA=6.911e-07
D3783 n3784 0 dm1 AREA=1.318e-06
D3784 n3785 0 dm1 AREA=1.251e-06
D3785 n3786 0 dm1 AREA=1.960e-06
D3786 n3787 0 dm1 AREA=2.378e-06
D3787 n3788 0 dm1 AREA=8.510e-07
D3788 n3789 0 dm1 AREA=7.216e-07
D3789 n3790 0 dm1 AREA=1.877e-07
D3790 n3791 0 dm1 AREA=4.995e-07
D3791 n3792 0 dm1 AREA=2.938e-06
D3792 n3793 0 dm1 AREA=1.545e-06
D3793 n3794 0 dm1 AREA=1.158e-06
D3794 n3795 0 dm1 AREA=9.355e-07
D3795 n3796 0 dm1 AREA=7.078e-07
D3796 n3797 0 dm1 AREA=1.438e-06
D3797 n3798 0 dm1 AREA=9.696e-07
D3798 n3799 0 dm1 AREA=2.716e-06
D3799 n3800 0 dm1 AREA=1.022e-06
D3800 n3801 0 dm1 AREA=1.447e-06
D3801 n3802 0 dm1 AREA=7.202e-07
D3802 n3803 0 dm1 AREA=1.342e-06
D3803 n3804 0 dm1 AREA=1.302e-06
D3804 n3805 0 dm1 AREA=5.343e-07
D3805 n3806 0 dm1 AREA=1.045e-07
D3806 n3807 0 dm1 AREA=1.800e-06
D3807 n3808 0 dm1 AREA=1.811e-06
D3808 n3809 0 dm1 AREA=3.795e-07
D3809 n3810 0 dm1 AREA=1.179e-06
D3810 n3811 0 dm1 AREA=1.098e-06
D3811 n3812 0 dm1 AREA=7.647e-07
D3812 n3813 0 dm1 AREA=5.347e-07
D3813 n3814 0 dm1 AREA=1.030e-06
D3814 n3815 0 dm1 AREA=1.066e-06
D3815 n3816 0 dm1 AREA=2.039e-07
D3816 n3817 0 dm1 AREA=4.828e-07
D3817 n3818 0 dm1 AREA=2.026e-06
D3818 n3819 0 dm1 AREA=1.570e-06
D3819 n3820 0 dm1 AREA=8.063e-07
D3820 n3821 0 dm1 AREA=1.157e-06
D3821 n3822 0 dm1 AREA=4.548e-07
D3822 n3823 0 dm1 AREA=4.584e-07
D3823 n3824 0 dm1 AREA=2.085e-06
D3824 n3825 0 dm1 AREA=1.605e-06
D3825 n3826 0 dm1 AREA=4.210e-07
D3826 n3827 0 dm1 AREA=9.730e-07
D3827 n3828 0 dm1 AREA=8.246e-07
D3828 n3829 0 dm1 AREA=9.755e-07
D3829 n3830 0 dm1 AREA=9.656e-07
D3830 n3831 0 dm1 AREA=8.125e-07
D3831 n3832 0 dm1 AREA=1.443e-06
D3832 n3833 0 dm1 AREA=6.724e-07
D3833 n3834 0 dm1 AREA=3.696e-07
D3834 n3835 0 dm1 AREA=8.609e-07
D3835 n3836 0 dm1 AREA=1.286e-06
D3836 n3837 0 dm1 AREA=1.003e-06
D3837 n3838 0 dm1 AREA=1.209e-06
D3838 n3839 0 dm1 AREA=5.160e-07
D3839 n3840 0 dm1 AREA=9.438e-07
D3840 n3841 0 dm1 AREA=5.285e-07
D3841 n3842 0 dm1 AREA=9.412e-07
D3842 n3843 0 dm1 AREA=5.619e-07
D3843 n3844 0 dm1 AREA=6.681e-07
D3844 n3845 0 dm1 AREA=7.623e-07
D3845 n3846 0 dm1 AREA=3.175e-07
D3846 n3847 0 dm1 AREA=1.671e-06
D3847 n3848 0 dm1 AREA=8.044e-07
D3848 n3849 0 dm1 AREA=1.320e-06
D3849 n3850 0 dm1 AREA=1.322e-06
D3850 n3851 0 dm1 AREA=1.278e-06
D3851 n3852 0 dm1 AREA=3.744e-07
D3852 n3853 0 dm1 AREA=8.123e-07
D3853 n3854 0 dm1 AREA=1.884e-06
D3854 n3855 0 dm1 AREA=1.474e-06
D3855 n3856 0 dm1 AREA=5.409e-07
D3856 n3857 0 dm1 AREA=9.930e-07
D3857 n3858 0 dm1 AREA=6.365e-07
D3858 n3859 0 dm1 AREA=3.776e-08
D3859 n3860 0 dm1 AREA=3.613e-07
D3860 n3861 0 dm1 AREA=8.328e-07
D3861 n3862 0 dm1 AREA=1.127e-06
D3862 n3863 0 dm1 AREA=2.099e-07
D3863 n3864 0 dm1 AREA=5.383e-07
D3864 n3865 0 dm1 AREA=1.315e-06
D3865 n3866 0 dm1 AREA=1.629e-06
D3866 n3867 0 dm1 AREA=3.564e-07
D3867 n3868 0 dm1 AREA=1.356e-06
D3868 n3869 0 dm1 AREA=1.950e-06
D3869 n3870 0 dm1 AREA=9.083e-07
D3870 n3871 0 dm1 AREA=9.430e-07
D3871 n3872 0 dm1 AREA=2.075e-06
D3872 n3873 0 dm1 AREA=1.049e-06
D3873 n3874 0 dm1 AREA=1.628e-06
D3874 n3875 0 dm1 AREA=8.192e-07
D3875 n3876 0 dm1 AREA=1.089e-06
D3876 n3877 0 dm1 AREA=9.792e-07
D3877 n3878 0 dm1 AREA=8.124e-07
D3878 n3879 0 dm1 AREA=6.025e-07
D3879 n3880 0 dm1 AREA=8.938e-07
D3880 n3881 0 dm1 AREA=7.428e-07
D3881 n3882 0 dm1 AREA=7.821e-07
D3882 n3883 0 dm1 AREA=1.380e-06
D3883 n3884 0 dm1 AREA=1.034e-06
D3884 n3885 0 dm1 AREA=2.630e-07
D3885 n3886 0 dm1 AREA=1.012e-06
D3886 n3887 0 dm1 AREA=6.967e-07
D3887 n3888 0 dm1 AREA=4.540e-07
D3888 n3889 0 dm1 AREA=6.820e-07
D3889 n3890 0 dm1 AREA=4.847e-07
D3890 n3891 0 dm1 AREA=1.088e-06
D3891 n3892 0 dm1 AREA=7.831e-07
D3892 n3893 0 dm1 AREA=7.094e-07
D3893 n3894 0 dm1 AREA=6.013e-07
D3894 n3895 0 dm1 AREA=5.032e-07
D3895 n3896 0 dm1 AREA=1.083e-06
D3896 n3897 0 dm1 AREA=6.876e-07
D3897 n3898 0 dm1 AREA=9.702e-07
D3898 n3899 0 dm1 AREA=1.018e-06
D3899 n3900 0 dm1 AREA=1.779e-06
D3900 n3901 0 dm1 AREA=1.252e-06
D3901 n3902 0 dm1 AREA=1.160e-06
D3902 n3903 0 dm1 AREA=1.187e-06
D3903 n3904 0 dm1 AREA=1.442e-06
D3904 n3905 0 dm1 AREA=2.253e-07
D3905 n3906 0 dm1 AREA=7.124e-07
D3906 n3907 0 dm1 AREA=3.710e-07
D3907 n3908 0 dm1 AREA=9.550e-07
D3908 n3909 0 dm1 AREA=5.417e-07
D3909 n3910 0 dm1 AREA=6.207e-07
D3910 n3911 0 dm1 AREA=5.088e-07
D3911 n3912 0 dm1 AREA=7.641e-07
D3912 n3913 0 dm1 AREA=2.786e-07
D3913 n3914 0 dm1 AREA=6.048e-07
D3914 n3915 0 dm1 AREA=5.120e-07
D3915 n3916 0 dm1 AREA=2.000e-06
D3916 n3917 0 dm1 AREA=9.889e-07
D3917 n3918 0 dm1 AREA=9.928e-07
D3918 n3919 0 dm1 AREA=7.103e-07
D3919 n3920 0 dm1 AREA=1.135e-06
D3920 n3921 0 dm1 AREA=6.284e-07
D3921 n3922 0 dm1 AREA=1.019e-06
D3922 n3923 0 dm1 AREA=8.489e-07
D3923 n3924 0 dm1 AREA=1.004e-06
D3924 n3925 0 dm1 AREA=1.484e-06
D3925 n3926 0 dm1 AREA=8.006e-07
D3926 n3927 0 dm1 AREA=6.419e-07
D3927 n3928 0 dm1 AREA=3.753e-07
D3928 n3929 0 dm1 AREA=5.239e-07
D3929 n3930 0 dm1 AREA=2.094e-06
D3930 n3931 0 dm1 AREA=9.051e-07
D3931 n3932 0 dm1 AREA=3.897e-07
D3932 n3933 0 dm1 AREA=2.878e-06
D3933 n3934 0 dm1 AREA=1.507e-06
D3934 n3935 0 dm1 AREA=9.366e-07
D3935 n3936 0 dm1 AREA=6.612e-07
D3936 n3937 0 dm1 AREA=1.956e-06
D3937 n3938 0 dm1 AREA=1.135e-06
D3938 n3939 0 dm1 AREA=1.520e-07
D3939 n3940 0 dm1 AREA=1.601e-06
D3940 n3941 0 dm1 AREA=8.622e-07
D3941 n3942 0 dm1 AREA=1.365e-06
D3942 n3943 0 dm1 AREA=4.352e-07
D3943 n3944 0 dm1 AREA=1.051e-06
D3944 n3945 0 dm1 AREA=9.823e-07
D3945 n3946 0 dm1 AREA=2.581e-06
D3946 n3947 0 dm1 AREA=7.096e-07
D3947 n3948 0 dm1 AREA=1.792e-06
D3948 n3949 0 dm1 AREA=3.447e-07
D3949 n3950 0 dm1 AREA=2.303e-06
D3950 n3951 0 dm1 AREA=1.836e-07
D3951 n1 0 dm1 AREA=1.134e-06
D3952 n3953 0 dm1 AREA=1.525e-06
D3953 n3954 0 dm1 AREA=1.255e-06
D3954 n3955 0 dm1 AREA=8.089e-07
D3955 n3956 0 dm1 AREA=1.139e-06
D3956 n3957 0 dm1 AREA=1.695e-06
D3957 n3958 0 dm1 AREA=9.380e-07
D3958 n3959 0 dm1 AREA=1.450e-06
D3959 n3960 0 dm1 AREA=1.646e-06
D3960 n3961 0 dm1 AREA=4.707e-07
D3961 n3962 0 dm1 AREA=1.263e-06
D3962 n3963 0 dm1 AREA=1.187e-06
D3963 n3964 0 dm1 AREA=9.064e-07
D3964 n3965 0 dm1 AREA=1.630e-06
D3965 n3966 0 dm1 AREA=5.200e-07
D3966 n3967 0 dm1 AREA=1.685e-06
D3967 n3968 0 dm1 AREA=8.600e-07
D3968 n3969 0 dm1 AREA=7.040e-07
D3969 n3970 0 dm1 AREA=2.497e-06
D3970 n3971 0 dm1 AREA=8.638e-07
D3971 n3972 0 dm1 AREA=1.522e-06
D3972 n3973 0 dm1 AREA=7.603e-07
D3973 n3974 0 dm1 AREA=1.736e-06
D3974 n3975 0 dm1 AREA=1.195e-06
D3975 n3976 0 dm1 AREA=9.135e-07
D3976 n3977 0 dm1 AREA=3.964e-07
D3977 n3978 0 dm1 AREA=1.853e-07
D3978 n3979 0 dm1 AREA=1.893e-06
D3979 n3980 0 dm1 AREA=5.427e-07
D3980 n3981 0 dm1 AREA=4.704e-07
D3981 n3982 0 dm1 AREA=1.044e-06
D3982 n3983 0 dm1 AREA=5.805e-07
D3983 n3984 0 dm1 AREA=2.422e-06
D3984 n3985 0 dm1 AREA=9.561e-07
D3985 n3986 0 dm1 AREA=6.093e-07
D3986 n3987 0 dm1 AREA=2.702e-06
D3987 n3988 0 dm1 AREA=7.391e-07
D3988 n3989 0 dm1 AREA=6.121e-07
D3989 n3990 0 dm1 AREA=7.973e-07
D3990 n3991 0 dm1 AREA=7.523e-07
D3991 n3992 0 dm1 AREA=9.225e-07
D3992 n3993 0 dm1 AREA=7.699e-07
D3993 n3994 0 dm1 AREA=1.148e-07
D3994 n3995 0 dm1 AREA=6.335e-07
D3995 n3996 0 dm1 AREA=1.372e-06
D3996 n3997 0 dm1 AREA=2.198e-06
D3997 n3998 0 dm1 AREA=1.528e-06
D3998 n3999 0 dm1 AREA=1.140e-06
D3999 n4000 0 dm1 AREA=6.874e-07
D4000 n4001 0 dm1 AREA=2.002e-07
D4001 n4002 0 dm1 AREA=1.476e-06
D4002 n4003 0 dm1 AREA=1.080e-06
D4003 n4004 0 dm1 AREA=6.948e-07
D4004 n4005 0 dm1 AREA=5.536e-07
D4005 n4006 0 dm1 AREA=8.652e-07
D4006 n4007 0 dm1 AREA=9.365e-07
D4007 n4008 0 dm1 AREA=1.385e-06
D4008 n4009 0 dm1 AREA=5.870e-07
D4009 n4010 0 dm1 AREA=5.456e-07
D4010 n4011 0 dm1 AREA=6.999e-07
D4011 n4012 0 dm1 AREA=1.250e-06
D4012 n4013 0 dm1 AREA=1.096e-06
D4013 n4014 0 dm1 AREA=8.570e-07
D4014 n4015 0 dm1 AREA=1.494e-06
D4015 n4016 0 dm1 AREA=1.832e-06
D4016 n4017 0 dm1 AREA=9.298e-07
D4017 n4018 0 dm1 AREA=8.067e-07
D4018 n4019 0 dm1 AREA=2.317e-07
D4019 n4020 0 dm1 AREA=4.479e-07
D4020 n4021 0 dm1 AREA=2.360e-06
D4021 n4022 0 dm1 AREA=3.218e-06
D4022 n4023 0 dm1 AREA=1.064e-06
D4023 n4024 0 dm1 AREA=2.398e-06
D4024 n4025 0 dm1 AREA=5.349e-07
D4025 n4026 0 dm1 AREA=1.218e-06
D4026 n4027 0 dm1 AREA=1.275e-06
D4027 n4028 0 dm1 AREA=8.261e-07
D4028 n4029 0 dm1 AREA=6.988e-07
D4029 n4030 0 dm1 AREA=1.148e-06
D4030 n4031 0 dm1 AREA=8.716e-07
D4031 n4032 0 dm1 AREA=1.038e-06
D4032 n4033 0 dm1 AREA=1.060e-06
D4033 n4034 0 dm1 AREA=1.181e-06
D4034 n4035 0 dm1 AREA=8.606e-07
D4035 n4036 0 dm1 AREA=8.316e-07
D4036 n4037 0 dm1 AREA=1.266e-06
D4037 n4038 0 dm1 AREA=1.049e-06
D4038 n4039 0 dm1 AREA=4.756e-07
D4039 n4040 0 dm1 AREA=8.496e-07
D4040 n4041 0 dm1 AREA=1.079e-06
D4041 n4042 0 dm1 AREA=1.177e-06
D4042 n4043 0 dm1 AREA=1.955e-06
D4043 n4044 0 dm1 AREA=2.842e-07
D4044 n4045 0 dm1 AREA=1.350e-06
D4045 n4046 0 dm1 AREA=2.084e-06
D4046 n4047 0 dm1 AREA=3.935e-07
D4047 n4048 0 dm1 AREA=2.813e-06
D4048 n4049 0 dm1 AREA=3.126e-07
D4049 n4050 0 dm1 AREA=3.708e-07
D4050 n4051 0 dm1 AREA=5.874e-07
D4051 n4052 0 dm1 AREA=9.194e-07
D4052 n4053 0 dm1 AREA=1.671e-06
D4053 n4054 0 dm1 AREA=9.562e-07
D4054 n4055 0 dm1 AREA=1.271e-06
D4055 n4056 0 dm1 AREA=1.213e-06
D4056 n4057 0 dm1 AREA=1.055e-06
D4057 n4058 0 dm1 AREA=6.047e-07
D4058 n4059 0 dm1 AREA=2.382e-06
D4059 n4060 0 dm1 AREA=6.332e-07
D4060 n4061 0 dm1 AREA=8.426e-07
D4061 n4062 0 dm1 AREA=1.200e-06
D4062 n4063 0 dm1 AREA=6.048e-07
D4063 n4064 0 dm1 AREA=1.559e-06
D4064 n4065 0 dm1 AREA=3.125e-07
D4065 n4066 0 dm1 AREA=6.412e-07
D4066 n4067 0 dm1 AREA=2.975e-07
D4067 n4068 0 dm1 AREA=2.566e-06
D4068 n4069 0 dm1 AREA=6.065e-07
D4069 n4070 0 dm1 AREA=8.303e-07
D4070 n4071 0 dm1 AREA=9.999e-07
D4071 n4072 0 dm1 AREA=7.605e-07
D4072 n4073 0 dm1 AREA=1.195e-06
D4073 n4074 0 dm1 AREA=4.947e-07
D4074 n4075 0 dm1 AREA=9.973e-07
D4075 n4076 0 dm1 AREA=8.370e-07
D4076 n4077 0 dm1 AREA=6.294e-07
D4077 n4078 0 dm1 AREA=3.909e-07
D4078 n4079 0 dm1 AREA=2.546e-06
D4079 n4080 0 dm1 AREA=1.590e-06
D4080 n4081 0 dm1 AREA=5.466e-07
D4081 n4082 0 dm1 AREA=1.393e-06
D4082 n4083 0 dm1 AREA=8.094e-07
D4083 n4084 0 dm1 AREA=1.023e-06
D4084 n4085 0 dm1 AREA=7.720e-07
D4085 n4086 0 dm1 AREA=3.493e-07
D4086 n4087 0 dm1 AREA=4.234e-07
D4087 n4088 0 dm1 AREA=4.867e-07
D4088 n4089 0 dm1 AREA=1.985e-06
D4089 n4090 0 dm1 AREA=8.145e-07
D4090 n4091 0 dm1 AREA=8.285e-07
D4091 n4092 0 dm1 AREA=8.436e-07
D4092 n4093 0 dm1 AREA=1.694e-06
D4093 n4094 0 dm1 AREA=1.266e-06
D4094 n4095 0 dm1 AREA=1.175e-06
D4095 n4096 0 dm1 AREA=1.059e-06
D4096 n4097 0 dm1 AREA=2.293e-06
D4097 n4098 0 dm1 AREA=9.917e-07
D4098 n4099 0 dm1 AREA=7.242e-07
D4099 n4100 0 dm1 AREA=5.620e-07
D4100 n4101 0 dm1 AREA=1.446e-06
D4101 n4102 0 dm1 AREA=4.386e-07
D4102 n4103 0 dm1 AREA=1.455e-06
D4103 n4104 0 dm1 AREA=3.738e-07
D4104 n4105 0 dm1 AREA=1.385e-06
D4105 n4106 0 dm1 AREA=2.057e-06
D4106 n4107 0 dm1 AREA=1.107e-06
D4107 n4108 0 dm1 AREA=1.026e-06
D4108 n4109 0 dm1 AREA=7.103e-07
D4109 n4110 0 dm1 AREA=1.404e-06
D4110 n4111 0 dm1 AREA=3.599e-07
D4111 n4112 0 dm1 AREA=1.140e-06
D4112 n4113 0 dm1 AREA=7.060e-07
D4113 n4114 0 dm1 AREA=1.449e-06
D4114 n4115 0 dm1 AREA=1.106e-06
D4115 n4116 0 dm1 AREA=1.291e-06
D4116 n4117 0 dm1 AREA=1.313e-06
D4117 n4118 0 dm1 AREA=3.748e-07
D4118 n4119 0 dm1 AREA=3.540e-07
D4119 n4120 0 dm1 AREA=1.944e-06
D4120 n4121 0 dm1 AREA=1.339e-06
D4121 n4122 0 dm1 AREA=4.032e-07
D4122 n4123 0 dm1 AREA=1.115e-06
D4123 n4124 0 dm1 AREA=3.487e-07
D4124 n4125 0 dm1 AREA=1.120e-06
D4125 n4126 0 dm1 AREA=1.135e-06
D4126 n4127 0 dm1 AREA=4.728e-07
D4127 n4128 0 dm1 AREA=8.735e-07
D4128 n4129 0 dm1 AREA=1.837e-06
D4129 n4130 0 dm1 AREA=2.166e-06
D4130 n4131 0 dm1 AREA=1.690e-06
D4131 n4132 0 dm1 AREA=5.911e-07
D4132 n4133 0 dm1 AREA=3.983e-07
D4133 n4134 0 dm1 AREA=7.826e-07
D4134 n4135 0 dm1 AREA=1.827e-06
D4135 n4136 0 dm1 AREA=3.929e-07
D4136 n4137 0 dm1 AREA=1.211e-06
D4137 n4138 0 dm1 AREA=2.087e-06
D4138 n4139 0 dm1 AREA=2.578e-06
D4139 n4140 0 dm1 AREA=4.896e-07
D4140 n4141 0 dm1 AREA=1.103e-06
D4141 n4142 0 dm1 AREA=7.332e-07
D4142 n4143 0 dm1 AREA=1.459e-06
D4143 n4144 0 dm1 AREA=2.489e-06
D4144 n4145 0 dm1 AREA=5.223e-07
D4145 n4146 0 dm1 AREA=5.902e-07
D4146 n4147 0 dm1 AREA=1.363e-06
D4147 n4148 0 dm1 AREA=1.919e-06
D4148 n4149 0 dm1 AREA=6.256e-07
D4149 n4150 0 dm1 AREA=1.422e-06
D4150 n4151 0 dm1 AREA=1.244e-06
D4151 n4152 0 dm1 AREA=6.705e-07
D4152 n4153 0 dm1 AREA=1.623e-06
D4153 n4154 0 dm1 AREA=8.136e-07
D4154 n4155 0 dm1 AREA=1.255e-06
D4155 n4156 0 dm1 AREA=6.143e-07
D4156 n4157 0 dm1 AREA=9.150e-07
D4157 n4158 0 dm1 AREA=9.773e-07
D4158 n4159 0 dm1 AREA=1.884e-06
D4159 n4160 0 dm1 AREA=2.920e-07
D4160 n4161 0 dm1 AREA=5.072e-07
D4161 n4162 0 dm1 AREA=5.440e-07
D4162 n4163 0 dm1 AREA=1.707e-06
D4163 n4164 0 dm1 AREA=7.917e-07
D4164 n4165 0 dm1 AREA=2.480e-06
D4165 n4166 0 dm1 AREA=7.679e-07
D4166 n4167 0 dm1 AREA=8.071e-07
D4167 n4168 0 dm1 AREA=5.845e-07
D4168 n4169 0 dm1 AREA=1.159e-06
D4169 n4170 0 dm1 AREA=7.948e-07
D4170 n4171 0 dm1 AREA=9.418e-07
D4171 n4172 0 dm1 AREA=1.059e-06
D4172 n4173 0 dm1 AREA=6.433e-07
D4173 n4174 0 dm1 AREA=9.255e-07
D4174 n4175 0 dm1 AREA=1.313e-06
D4175 n4176 0 dm1 AREA=9.170e-07
D4176 n4177 0 dm1 AREA=7.866e-07
D4177 n4178 0 dm1 AREA=8.215e-07
D4178 n4179 0 dm1 AREA=1.591e-06
D4179 n4180 0 dm1 AREA=3.525e-07
D4180 n4181 0 dm1 AREA=8.303e-07
D4181 n4182 0 dm1 AREA=4.523e-07
D4182 n4183 0 dm1 AREA=4.228e-07
D4183 n4184 0 dm1 AREA=9.439e-07
D4184 n4185 0 dm1 AREA=1.109e-06
D4185 n4186 0 dm1 AREA=5.079e-07
D4186 n4187 0 dm1 AREA=8.967e-07
D4187 n4188 0 dm1 AREA=8.215e-07
D4188 n4189 0 dm1 AREA=6.405e-07
D4189 n1 0 dm1 AREA=1.048e-06
D4190 n4191 0 dm1 AREA=9.232e-07
D4191 n4192 0 dm1 AREA=1.488e-06
D4192 n4193 0 dm1 AREA=1.138e-06
D4193 n4194 0 dm1 AREA=1.069e-06
D4194 n4195 0 dm1 AREA=1.183e-07
D4195 n4196 0 dm1 AREA=2.495e-06
D4196 n4197 0 dm1 AREA=4.611e-07
D4197 n4198 0 dm1 AREA=5.078e-07
D4198 n4199 0 dm1 AREA=1.599e-06
D4199 n4200 0 dm1 AREA=8.638e-07
D4200 n4201 0 dm1 AREA=6.423e-07
D4201 n4202 0 dm1 AREA=6.893e-07
D4202 n4203 0 dm1 AREA=7.532e-07
D4203 n4204 0 dm1 AREA=5.643e-07
D4204 n4205 0 dm1 AREA=1.390e-06
D4205 n4206 0 dm1 AREA=4.057e-07
D4206 n4207 0 dm1 AREA=5.832e-07
D4207 n4208 0 dm1 AREA=4.457e-07
D4208 n4209 0 dm1 AREA=2.666e-07
D4209 n4210 0 dm1 AREA=9.526e-07
D4210 n4211 0 dm1 AREA=2.191e-06
D4211 n4212 0 dm1 AREA=1.060e-06
D4212 n4213 0 dm1 AREA=7.373e-07
D4213 n4214 0 dm1 AREA=4.472e-07
D4214 n4215 0 dm1 AREA=3.838e-07
D4215 n4216 0 dm1 AREA=2.414e-06
D4216 n4217 0 dm1 AREA=8.533e-07
D4217 n4218 0 dm1 AREA=7.939e-07
D4218 n4219 0 dm1 AREA=1.650e-06
D4219 n4220 0 dm1 AREA=6.948e-07
D4220 n4221 0 dm1 AREA=5.896e-07
D4221 n4222 0 dm1 AREA=9.310e-07
D4222 n4223 0 dm1 AREA=3.161e-07
D4223 n4224 0 dm1 AREA=5.248e-07
D4224 n4225 0 dm1 AREA=1.365e-06
D4225 n4226 0 dm1 AREA=6.717e-07
D4226 n4227 0 dm1 AREA=1.635e-07
D4227 n4228 0 dm1 AREA=9.423e-07
D4228 n4229 0 dm1 AREA=7.847e-07
D4229 n4230 0 dm1 AREA=1.110e-06
D4230 n4231 0 dm1 AREA=8.525e-07
D4231 n4232 0 dm1 AREA=1.025e-06
D4232 n4233 0 dm1 AREA=4.814e-07
D4233 n4234 0 dm1 AREA=4.058e-07
D4234 n4235 0 dm1 AREA=1.738e-06
D4235 n4236 0 dm1 AREA=8.729e-07
D4236 n4237 0 dm1 AREA=6.838e-07
D4237 n4238 0 dm1 AREA=2.495e-06
D4238 n4239 0 dm1 AREA=8.585e-07
D4239 n4240 0 dm1 AREA=1.069e-06
D4240 n4241 0 dm1 AREA=1.140e-06
D4241 n4242 0 dm1 AREA=8.617e-07
D4242 n4243 0 dm1 AREA=2.667e-07
D4243 n4244 0 dm1 AREA=3.775e-07
D4244 n4245 0 dm1 AREA=8.489e-07
D4245 n4246 0 dm1 AREA=8.519e-07
D4246 n4247 0 dm1 AREA=8.189e-07
D4247 n4248 0 dm1 AREA=6.930e-07
D4248 n4249 0 dm1 AREA=1.373e-06
D4249 n4250 0 dm1 AREA=8.628e-07
D4250 n4251 0 dm1 AREA=9.185e-07
D4251 n4252 0 dm1 AREA=1.102e-06
D4252 n4253 0 dm1 AREA=4.924e-07
D4253 n4254 0 dm1 AREA=5.864e-07
D4254 n4255 0 dm1 AREA=1.413e-06
D4255 n4256 0 dm1 AREA=1.292e-06
D4256 n4257 0 dm1 AREA=4.708e-07
D4257 n4258 0 dm1 AREA=7.233e-07
D4258 n4259 0 dm1 AREA=1.170e-06
D4259 n4260 0 dm1 AREA=9.257e-07
D4260 n4261 0 dm1 AREA=1.796e-06
D4261 n4262 0 dm1 AREA=1.851e-06
D4262 n4263 0 dm1 AREA=1.084e-06
D4263 n4264 0 dm1 AREA=6.369e-07
D4264 n4265 0 dm1 AREA=7.541e-07
D4265 n4266 0 dm1 AREA=1.747e-06
D4266 n4267 0 dm1 AREA=1.829e-07
D4267 n4268 0 dm1 AREA=6.147e-07
D4268 n4269 0 dm1 AREA=1.382e-06
D4269 n4270 0 dm1 AREA=1.043e-06
D4270 n4271 0 dm1 AREA=6.632e-07
D4271 n4272 0 dm1 AREA=2.035e-06
D4272 n4273 0 dm1 AREA=8.499e-07
D4273 n4274 0 dm1 AREA=1.730e-06
D4274 n4275 0 dm1 AREA=1.061e-06
D4275 n4276 0 dm1 AREA=3.174e-07
D4276 n4277 0 dm1 AREA=9.379e-07
D4277 n4278 0 dm1 AREA=1.003e-06
D4278 n4279 0 dm1 AREA=1.464e-06
D4279 n4280 0 dm1 AREA=7.483e-07
D4280 n4281 0 dm1 AREA=1.687e-06
D4281 n4282 0 dm1 AREA=1.092e-06
D4282 n4283 0 dm1 AREA=8.773e-07
D4283 n4284 0 dm1 AREA=9.578e-07
D4284 n4285 0 dm1 AREA=1.307e-06
D4285 n4286 0 dm1 AREA=3.727e-07
D4286 n4287 0 dm1 AREA=2.431e-07
D4287 n4288 0 dm1 AREA=1.487e-06
D4288 n4289 0 dm1 AREA=3.472e-07
D4289 n4290 0 dm1 AREA=8.070e-07
D4290 n4291 0 dm1 AREA=1.004e-06
D4291 n4292 0 dm1 AREA=1.109e-06
D4292 n4293 0 dm1 AREA=1.617e-06
D4293 n4294 0 dm1 AREA=3.929e-07
D4294 n4295 0 dm1 AREA=1.030e-06
D4295 n4296 0 dm1 AREA=9.951e-07
D4296 n4297 0 dm1 AREA=3.791e-07
D4297 n4298 0 dm1 AREA=5.411e-07
D4298 n4299 0 dm1 AREA=3.892e-07
D4299 n4300 0 dm1 AREA=1.971e-06
D4300 n4301 0 dm1 AREA=1.276e-06
D4301 n4302 0 dm1 AREA=1.726e-06
D4302 n4303 0 dm1 AREA=1.181e-06
D4303 n4304 0 dm1 AREA=1.665e-06
D4304 n4305 0 dm1 AREA=1.452e-06
D4305 n4306 0 dm1 AREA=2.394e-07
D4306 n4307 0 dm1 AREA=5.411e-07
D4307 n4308 0 dm1 AREA=8.108e-07
D4308 n4309 0 dm1 AREA=5.124e-07
D4309 n4310 0 dm1 AREA=1.016e-06
D4310 n4311 0 dm1 AREA=1.096e-06
D4311 n4312 0 dm1 AREA=7.745e-07
D4312 n4313 0 dm1 AREA=1.343e-06
D4313 n4314 0 dm1 AREA=1.650e-06
D4314 n4315 0 dm1 AREA=2.876e-06
D4315 n4316 0 dm1 AREA=1.062e-06
D4316 n4317 0 dm1 AREA=6.877e-07
D4317 n4318 0 dm1 AREA=5.937e-07
D4318 n4319 0 dm1 AREA=7.740e-07
D4319 n4320 0 dm1 AREA=6.598e-07
D4320 n4321 0 dm1 AREA=3.790e-07
D4321 n4322 0 dm1 AREA=5.738e-07
D4322 n4323 0 dm1 AREA=2.108e-06
D4323 n4324 0 dm1 AREA=5.369e-07
D4324 n4325 0 dm1 AREA=1.344e-06
D4325 n4326 0 dm1 AREA=8.138e-07
D4326 n4327 0 dm1 AREA=1.313e-06
D4327 n4328 0 dm1 AREA=8.785e-07
D4328 n4329 0 dm1 AREA=7.887e-07
D4329 n4330 0 dm1 AREA=1.709e-06
D4330 n1 0 dm1 AREA=4.818e-07
D4331 n1 0 dm1 AREA=8.180e-07
D4332 n4333 0 dm1 AREA=6.799e-07
D4333 n4334 0 dm1 AREA=1.051e-06
D4334 n4335 0 dm1 AREA=5.873e-07
D4335 n4336 0 dm1 AREA=1.073e-06
D4336 n4337 0 dm1 AREA=7.384e-07
D4337 n4338 0 dm1 AREA=1.312e-06
D4338 n1 0 dm1 AREA=7.876e-07
D4339 n4340 0 dm1 AREA=5.262e-07
D4340 n4341 0 dm1 AREA=7.622e-07
D4341 n4342 0 dm1 AREA=4.644e-07
D4342 n4343 0 dm1 AREA=2.045e-06
D4343 n4344 0 dm1 AREA=3.291e-06
D4344 n4345 0 dm1 AREA=1.273e-06
D4345 n4346 0 dm1 AREA=1.505e-06
D4346 n4347 0 dm1 AREA=9.687e-07
D4347 n4348 0 dm1 AREA=3.825e-07
D4348 n4349 0 dm1 AREA=6.595e-07
D4349 n4350 0 dm1 AREA=3.473e-07
D4350 n4351 0 dm1 AREA=8.975e-07
D4351 n4352 0 dm1 AREA=1.182e-06
D4352 n4353 0 dm1 AREA=1.262e-06
D4353 n4354 0 dm1 AREA=2.211e-06
D4354 n4355 0 dm1 AREA=2.060e-06
D4355 n4356 0 dm1 AREA=3.707e-07
D4356 n4357 0 dm1 AREA=8.471e-07
D4357 n4358 0 dm1 AREA=7.446e-07
D4358 n4359 0 dm1 AREA=5.947e-07
D4359 n4360 0 dm1 AREA=1.389e-06
D4360 n4361 0 dm1 AREA=1.093e-06
D4361 n4362 0 dm1 AREA=8.821e-07
D4362 n4363 0 dm1 AREA=2.226e-06
D4363 n4364 0 dm1 AREA=2.440e-06
D4364 n4365 0 dm1 AREA=8.322e-07
D4365 n4366 0 dm1 AREA=6.755e-07
D4366 n4367 0 dm1 AREA=1.184e-06
D4367 n4368 0 dm1 AREA=1.377e-06
D4368 n4369 0 dm1 AREA=4.658e-07
D4369 n4370 0 dm1 AREA=9.097e-07
D4370 n4371 0 dm1 AREA=6.594e-07
D4371 n4372 0 dm1 AREA=6.060e-07
D4372 n4373 0 dm1 AREA=1.410e-06
D4373 n4374 0 dm1 AREA=6.746e-07
D4374 n4375 0 dm1 AREA=1.179e-06
D4375 n4376 0 dm1 AREA=1.530e-06
D4376 n4377 0 dm1 AREA=2.051e-07
D4377 n4378 0 dm1 AREA=8.812e-07
D4378 n4379 0 dm1 AREA=2.603e-06
D4379 n4380 0 dm1 AREA=4.134e-07
D4380 n4381 0 dm1 AREA=1.151e-06
D4381 n4382 0 dm1 AREA=7.858e-07
D4382 n4383 0 dm1 AREA=8.157e-07
D4383 n4384 0 dm1 AREA=1.006e-06
D4384 n4385 0 dm1 AREA=7.641e-07
D4385 n1 0 dm1 AREA=7.157e-07
D4386 n4387 0 dm1 AREA=1.172e-06
D4387 n4388 0 dm1 AREA=7.395e-07
D4388 n4389 0 dm1 AREA=7.918e-07
D4389 n4390 0 dm1 AREA=1.484e-06
D4390 n4391 0 dm1 AREA=1.088e-06
D4391 n4392 0 dm1 AREA=2.196e-06
D4392 n4393 0 dm1 AREA=2.890e-06
D4393 n4394 0 dm1 AREA=1.694e-06
D4394 n4395 0 dm1 AREA=4.613e-07
D4395 n4396 0 dm1 AREA=6.283e-07
D4396 n4397 0 dm1 AREA=6.655e-07
D4397 n4398 0 dm1 AREA=2.150e-06
D4398 n4399 0 dm1 AREA=2.153e-06
D4399 n4400 0 dm1 AREA=1.474e-06
D4400 n4401 0 dm1 AREA=8.503e-07
D4401 n4402 0 dm1 AREA=1.852e-06
D4402 n4403 0 dm1 AREA=1.347e-06
D4403 n4404 0 dm1 AREA=3.539e-07
D4404 n4405 0 dm1 AREA=3.538e-07
D4405 n4406 0 dm1 AREA=6.409e-07
D4406 n4407 0 dm1 AREA=9.869e-07
D4407 n4408 0 dm1 AREA=6.869e-07
D4408 n4409 0 dm1 AREA=1.075e-06
D4409 n4410 0 dm1 AREA=1.377e-06
D4410 n4411 0 dm1 AREA=3.502e-07
D4411 n4412 0 dm1 AREA=3.620e-07
D4412 n4413 0 dm1 AREA=1.201e-06
D4413 n4414 0 dm1 AREA=7.283e-07
D4414 n4415 0 dm1 AREA=1.257e-06
D4415 n4416 0 dm1 AREA=5.114e-07
D4416 n4417 0 dm1 AREA=9.447e-07
D4417 n4418 0 dm1 AREA=1.026e-06
D4418 n4419 0 dm1 AREA=1.807e-07
D4419 n4420 0 dm1 AREA=1.168e-06
D4420 n4421 0 dm1 AREA=9.629e-07
D4421 n4422 0 dm1 AREA=3.128e-06
D4422 n4423 0 dm1 AREA=6.792e-07
D4423 n4424 0 dm1 AREA=5.093e-07
D4424 n4425 0 dm1 AREA=5.670e-07
D4425 n4426 0 dm1 AREA=1.612e-06
D4426 n4427 0 dm1 AREA=1.621e-07
D4427 n4428 0 dm1 AREA=3.540e-07
D4428 n4429 0 dm1 AREA=4.925e-07
D4429 n4430 0 dm1 AREA=8.668e-07
D4430 n4431 0 dm1 AREA=1.126e-06
D4431 n4432 0 dm1 AREA=2.066e-07
D4432 n4433 0 dm1 AREA=9.135e-07
D4433 n4434 0 dm1 AREA=1.220e-06
D4434 n4435 0 dm1 AREA=1.255e-06
D4435 n4436 0 dm1 AREA=7.393e-07
D4436 n4437 0 dm1 AREA=1.668e-07
D4437 n4438 0 dm1 AREA=1.809e-06
D4438 n4439 0 dm1 AREA=7.077e-07
D4439 n4440 0 dm1 AREA=1.328e-06
D4440 n4441 0 dm1 AREA=4.566e-07
D4441 n4442 0 dm1 AREA=3.957e-07
D4442 n4443 0 dm1 AREA=7.970e-07
D4443 n4444 0 dm1 AREA=1.316e-06
D4444 n4445 0 dm1 AREA=1.205e-06
D4445 n4446 0 dm1 AREA=1.257e-06
D4446 n4447 0 dm1 AREA=6.599e-07
D4447 n4448 0 dm1 AREA=5.796e-07
D4448 n4449 0 dm1 AREA=8.215e-07
D4449 n4450 0 dm1 AREA=3.691e-07
D4450 n4451 0 dm1 AREA=2.042e-06
D4451 n4452 0 dm1 AREA=1.088e-06
D4452 n4453 0 dm1 AREA=7.657e-07
D4453 n4454 0 dm1 AREA=4.744e-07
D4454 n4455 0 dm1 AREA=1.649e-06
D4455 n4456 0 dm1 AREA=1.778e-07
D4456 n4457 0 dm1 AREA=2.251e-07
D4457 n4458 0 dm1 AREA=9.499e-07
D4458 n4459 0 dm1 AREA=8.332e-07
D4459 n4460 0 dm1 AREA=1.340e-06
D4460 n4461 0 dm1 AREA=1.050e-06
D4461 n4462 0 dm1 AREA=3.449e-07
D4462 n4463 0 dm1 AREA=1.620e-06
D4463 n4464 0 dm1 AREA=1.048e-06
D4464 n4465 0 dm1 AREA=1.069e-06
D4465 n4466 0 dm1 AREA=9.725e-07
D4466 n4467 0 dm1 AREA=2.680e-07
D4467 n4468 0 dm1 AREA=6.168e-07
D4468 n4469 0 dm1 AREA=5.317e-07
D4469 n4470 0 dm1 AREA=1.215e-06
D4470 n4471 0 dm1 AREA=9.827e-07
D4471 n4472 0 dm1 AREA=7.004e-07
D4472 n4473 0 dm1 AREA=2.665e-06
D4473 n4474 0 dm1 AREA=8.190e-07
D4474 n4475 0 dm1 AREA=9.317e-07
D4475 n4476 0 dm1 AREA=5.397e-07
D4476 n4477 0 dm1 AREA=4.978e-07
D4477 n4478 0 dm1 AREA=8.607e-07
D4478 n4479 0 dm1 AREA=1.070e-06
D4479 n4480 0 dm1 AREA=1.575e-06
D4480 n4481 0 dm1 AREA=4.924e-07
D4481 n4482 0 dm1 AREA=5.499e-07
D4482 n4483 0 dm1 AREA=1.463e-06
D4483 n4484 0 dm1 AREA=8.438e-07
D4484 n4485 0 dm1 AREA=7.316e-07
D4485 n4486 0 dm1 AREA=2.182e-06
D4486 n4487 0 dm1 AREA=1.050e-06
D4487 n4488 0 dm1 AREA=7.267e-07
D4488 n4489 0 dm1 AREA=9.928e-07
D4489 n4490 0 dm1 AREA=4.149e-07
D4490 n4491 0 dm1 AREA=9.077e-07
D4491 n4492 0 dm1 AREA=9.199e-07
D4492 n4493 0 dm1 AREA=6.912e-07
D4493 n4494 0 dm1 AREA=4.884e-07
D4494 n4495 0 dm1 AREA=1.855e-06
D4495 n4496 0 dm1 AREA=8.807e-07
D4496 n4497 0 dm1 AREA=5.235e-07
D4497 n4498 0 dm1 AREA=1.913e-06
D4498 n4499 0 dm1 AREA=7.979e-07
D4499 n4500 0 dm1 AREA=1.572e-06
D4500 n4501 0 dm1 AREA=1.324e-06
D4501 n4502 0 dm1 AREA=1.156e-06
D4502 n4503 0 dm1 AREA=2.222e-07
D4503 n4504 0 dm1 AREA=1.514e-06
D4504 n4505 0 dm1 AREA=5.984e-07
D4505 n4506 0 dm1 AREA=7.083e-07
D4506 n4507 0 dm1 AREA=1.454e-06
D4507 n4508 0 dm1 AREA=7.352e-07
D4508 n4509 0 dm1 AREA=6.859e-07
D4509 n4510 0 dm1 AREA=1.279e-06
D4510 n4511 0 dm1 AREA=1.580e-06
D4511 n4512 0 dm1 AREA=6.058e-07
D4512 n4513 0 dm1 AREA=5.350e-07
D4513 n4514 0 dm1 AREA=5.929e-07
D4514 n4515 0 dm1 AREA=1.549e-06
D4515 n4516 0 dm1 AREA=7.770e-07
D4516 n4517 0 dm1 AREA=6.097e-07
D4517 n4518 0 dm1 AREA=5.069e-07
D4518 n4519 0 dm1 AREA=1.736e-06
D4519 n4520 0 dm1 AREA=8.891e-07
D4520 n4521 0 dm1 AREA=1.903e-06
D4521 n4522 0 dm1 AREA=4.467e-07
D4522 n4523 0 dm1 AREA=9.193e-07
D4523 n4524 0 dm1 AREA=6.443e-07
D4524 n4525 0 dm1 AREA=1.203e-06
D4525 n4526 0 dm1 AREA=7.676e-07
D4526 n4527 0 dm1 AREA=2.064e-06
D4527 n4528 0 dm1 AREA=8.549e-07
D4528 n4529 0 dm1 AREA=1.221e-06
D4529 n4530 0 dm1 AREA=1.613e-06
D4530 n1 0 dm1 AREA=1.208e-06
D4531 n4532 0 dm1 AREA=9.056e-07
D4532 n4533 0 dm1 AREA=1.742e-06
D4533 n4534 0 dm1 AREA=6.537e-07
D4534 n4535 0 dm1 AREA=9.614e-07
D4535 n4536 0 dm1 AREA=1.760e-07
D4536 n4537 0 dm1 AREA=7.775e-07
D4537 n4538 0 dm1 AREA=7.564e-07
D4538 n4539 0 dm1 AREA=7.788e-07
D4539 n4540 0 dm1 AREA=4.542e-07
D4540 n4541 0 dm1 AREA=1.293e-06
D4541 n4542 0 dm1 AREA=4.628e-07
D4542 n4543 0 dm1 AREA=2.408e-06
D4543 n4544 0 dm1 AREA=3.579e-07
D4544 n4545 0 dm1 AREA=1.453e-06
D4545 n4546 0 dm1 AREA=1.020e-06
D4546 n4547 0 dm1 AREA=9.347e-07
D4547 n4548 0 dm1 AREA=9.275e-07
D4548 n4549 0 dm1 AREA=3.829e-07
D4549 n4550 0 dm1 AREA=1.124e-06
D4550 n4551 0 dm1 AREA=1.254e-06
D4551 n4552 0 dm1 AREA=5.122e-07
D4552 n4553 0 dm1 AREA=1.770e-06
D4553 n4554 0 dm1 AREA=1.185e-06
D4554 n4555 0 dm1 AREA=9.783e-07
D4555 n4556 0 dm1 AREA=6.685e-07
D4556 n4557 0 dm1 AREA=8.692e-07
D4557 n4558 0 dm1 AREA=1.194e-06
D4558 n4559 0 dm1 AREA=3.357e-07
D4559 n4560 0 dm1 AREA=1.472e-06
D4560 n4561 0 dm1 AREA=8.490e-07
D4561 n4562 0 dm1 AREA=2.437e-07
D4562 n4563 0 dm1 AREA=6.516e-07
D4563 n4564 0 dm1 AREA=5.830e-07
D4564 n4565 0 dm1 AREA=8.914e-07
D4565 n4566 0 dm1 AREA=7.273e-07
D4566 n4567 0 dm1 AREA=1.239e-06
D4567 n4568 0 dm1 AREA=1.076e-06
D4568 n4569 0 dm1 AREA=7.158e-07
D4569 n4570 0 dm1 AREA=3.087e-07
D4570 n4571 0 dm1 AREA=9.207e-07
D4571 n4572 0 dm1 AREA=2.711e-06
D4572 n4573 0 dm1 AREA=1.258e-06
D4573 n4574 0 dm1 AREA=1.109e-06
D4574 n4575 0 dm1 AREA=6.088e-07
D4575 n4576 0 dm1 AREA=8.902e-07
D4576 n4577 0 dm1 AREA=1.519e-06
D4577 n4578 0 dm1 AREA=8.457e-07
D4578 n4579 0 dm1 AREA=1.119e-06
D4579 n4580 0 dm1 AREA=2.124e-06
D4580 n4581 0 dm1 AREA=5.874e-07
D4581 n4582 0 dm1 AREA=7.023e-07
D4582 n4583 0 dm1 AREA=4.113e-07
D4583 n4584 0 dm1 AREA=9.607e-07
D4584 n4585 0 dm1 AREA=1.556e-06
D4585 n4586 0 dm1 AREA=1.891e-06
D4586 n4587 0 dm1 AREA=8.939e-07
D4587 n4588 0 dm1 AREA=1.253e-06
D4588 n4589 0 dm1 AREA=4.110e-07
D4589 n4590 0 dm1 AREA=7.043e-07
D4590 n4591 0 dm1 AREA=8.203e-07
D4591 n4592 0 dm1 AREA=9.205e-07
D4592 n4593 0 dm1 AREA=1.545e-06
D4593 n4594 0 dm1 AREA=1.177e-06
D4594 n4595 0 dm1 AREA=2.002e-06
D4595 n4596 0 dm1 AREA=1.137e-06
D4596 n4597 0 dm1 AREA=1.442e-06
D4597 n4598 0 dm1 AREA=9.858e-07
D4598 n4599 0 dm1 AREA=6.698e-07
D4599 n4600 0 dm1 AREA=1.468e-06
D4600 n4601 0 dm1 AREA=1.743e-07
D4601 n4602 0 dm1 AREA=1.156e-06
D4602 n4603 0 dm1 AREA=6.210e-07
D4603 n4604 0 dm1 AREA=1.724e-06
D4604 n4605 0 dm1 AREA=8.507e-07
D4605 n4606 0 dm1 AREA=2.574e-06
D4606 n4607 0 dm1 AREA=1.073e-06
D4607 n4608 0 dm1 AREA=8.583e-07
D4608 n4609 0 dm1 AREA=5.222e-07
D4609 n1 0 dm1 AREA=1.412e-06
D4610 n4611 0 dm1 AREA=1.053e-06
D4611 n4612 0 dm1 AREA=1.019e-06
D4612 n4613 0 dm1 AREA=1.371e-06
D4613 n4614 0 dm1 AREA=1.233e-06
D4614 n4615 0 dm1 AREA=9.963e-07
D4615 n4616 0 dm1 AREA=2.111e-06
D4616 n4617 0 dm1 AREA=7.486e-07
D4617 n4618 0 dm1 AREA=2.933e-07
D4618 n4619 0 dm1 AREA=1.033e-06
D4619 n4620 0 dm1 AREA=5.758e-07
D4620 n4621 0 dm1 AREA=4.930e-07
D4621 n4622 0 dm1 AREA=1.230e-06
D4622 n4623 0 dm1 AREA=8.840e-07
D4623 n4624 0 dm1 AREA=5.672e-07
D4624 n4625 0 dm1 AREA=1.028e-06
D4625 n4626 0 dm1 AREA=7.985e-07
D4626 n4627 0 dm1 AREA=2.937e-07
D4627 n4628 0 dm1 AREA=7.059e-07
D4628 n4629 0 dm1 AREA=9.912e-07
D4629 n4630 0 dm1 AREA=8.790e-07
D4630 n4631 0 dm1 AREA=1.360e-06
D4631 n4632 0 dm1 AREA=7.005e-07
D4632 n4633 0 dm1 AREA=1.428e-06
D4633 n4634 0 dm1 AREA=4.700e-07
D4634 n4635 0 dm1 AREA=1.087e-06
D4635 n4636 0 dm1 AREA=7.478e-07
D4636 n4637 0 dm1 AREA=9.424e-07
D4637 n4638 0 dm1 AREA=3.143e-07
D4638 n4639 0 dm1 AREA=5.717e-07
D4639 n4640 0 dm1 AREA=1.499e-06
D4640 n4641 0 dm1 AREA=4.347e-07
D4641 n4642 0 dm1 AREA=3.311e-07
D4642 n4643 0 dm1 AREA=7.428e-07
D4643 n4644 0 dm1 AREA=2.913e-07
D4644 n4645 0 dm1 AREA=4.348e-07
D4645 n4646 0 dm1 AREA=9.540e-07
D4646 n4647 0 dm1 AREA=1.716e-06
D4647 n4648 0 dm1 AREA=9.178e-07
D4648 n4649 0 dm1 AREA=9.487e-07
D4649 n4650 0 dm1 AREA=1.302e-06
D4650 n4651 0 dm1 AREA=4.838e-07
D4651 n4652 0 dm1 AREA=1.122e-06
D4652 n4653 0 dm1 AREA=1.279e-06
D4653 n4654 0 dm1 AREA=1.907e-06
D4654 n4655 0 dm1 AREA=7.492e-07
D4655 n4656 0 dm1 AREA=6.288e-07
D4656 n4657 0 dm1 AREA=5.471e-07
D4657 n4658 0 dm1 AREA=3.988e-07
D4658 n4659 0 dm1 AREA=7.652e-07
D4659 n4660 0 dm1 AREA=4.826e-07
D4660 n4661 0 dm1 AREA=8.577e-07
D4661 n4662 0 dm1 AREA=2.752e-06
D4662 n4663 0 dm1 AREA=9.810e-07
D4663 n4664 0 dm1 AREA=8.048e-07
D4664 n4665 0 dm1 AREA=1.123e-06
D4665 n4666 0 dm1 AREA=6.877e-07
D4666 n1 0 dm1 AREA=9.757e-07
D4667 n4668 0 dm1 AREA=6.223e-07
D4668 n4669 0 dm1 AREA=7.155e-07
D4669 n4670 0 dm1 AREA=1.219e-06
D4670 n4671 0 dm1 AREA=1.008e-06
D4671 n4672 0 dm1 AREA=7.146e-07
D4672 n4673 0 dm1 AREA=1.044e-06
D4673 n4674 0 dm1 AREA=1.735e-06
D4674 n4675 0 dm1 AREA=1.954e-06
D4675 n4676 0 dm1 AREA=9.395e-07
D4676 n4677 0 dm1 AREA=1.526e-06
D4677 n4678 0 dm1 AREA=7.287e-07
D4678 n4679 0 dm1 AREA=1.134e-07
D4679 n4680 0 dm1 AREA=7.958e-07
D4680 n4681 0 dm1 AREA=5.796e-07
D4681 n4682 0 dm1 AREA=6.636e-07
D4682 n4683 0 dm1 AREA=1.229e-06
D4683 n4684 0 dm1 AREA=1.500e-06
D4684 n4685 0 dm1 AREA=4.386e-07
D4685 n4686 0 dm1 AREA=1.869e-06
D4686 n4687 0 dm1 AREA=6.567e-07
D4687 n4688 0 dm1 AREA=1.977e-06
D4688 n4689 0 dm1 AREA=1.656e-06
D4689 n4690 0 dm1 AREA=6.939e-07
D4690 n4691 0 dm1 AREA=9.286e-07
D4691 n4692 0 dm1 AREA=4.328e-07
D4692 n4693 0 dm1 AREA=7.343e-07
D4693 n4694 0 dm1 AREA=7.578e-07
D4694 n4695 0 dm1 AREA=1.324e-06
D4695 n4696 0 dm1 AREA=1.295e-06
D4696 n4697 0 dm1 AREA=6.542e-07
D4697 n4698 0 dm1 AREA=6.369e-07
D4698 n4699 0 dm1 AREA=7.161e-07
D4699 n4700 0 dm1 AREA=1.447e-06
D4700 n4701 0 dm1 AREA=1.370e-06
D4701 n4702 0 dm1 AREA=9.511e-07
D4702 n4703 0 dm1 AREA=1.542e-06
D4703 n4704 0 dm1 AREA=2.137e-06
D4704 n4705 0 dm1 AREA=2.028e-06
D4705 n4706 0 dm1 AREA=5.523e-07
D4706 n4707 0 dm1 AREA=1.684e-06
D4707 n4708 0 dm1 AREA=1.570e-06
D4708 n4709 0 dm1 AREA=1.682e-06
D4709 n4710 0 dm1 AREA=1.677e-06
D4710 n4711 0 dm1 AREA=1.370e-06
D4711 n4712 0 dm1 AREA=1.467e-06
D4712 n4713 0 dm1 AREA=4.934e-07
D4713 n4714 0 dm1 AREA=1.247e-06
D4714 n4715 0 dm1 AREA=1.500e-06
D4715 n4716 0 dm1 AREA=7.945e-07
D4716 n4717 0 dm1 AREA=6.502e-07
D4717 n4718 0 dm1 AREA=1.149e-06
D4718 n4719 0 dm1 AREA=1.093e-06
D4719 n4720 0 dm1 AREA=3.755e-07
D4720 n4721 0 dm1 AREA=4.603e-07
D4721 n4722 0 dm1 AREA=1.188e-06
D4722 n4723 0 dm1 AREA=6.627e-07
D4723 n4724 0 dm1 AREA=7.543e-07
D4724 n4725 0 dm1 AREA=1.142e-06
D4725 n4726 0 dm1 AREA=2.414e-07
D4726 n4727 0 dm1 AREA=1.151e-06
D4727 n4728 0 dm1 AREA=5.673e-07
D4728 n4729 0 dm1 AREA=8.875e-07
D4729 n4730 0 dm1 AREA=1.231e-06
D4730 n4731 0 dm1 AREA=1.127e-06
D4731 n4732 0 dm1 AREA=6.826e-07
D4732 n4733 0 dm1 AREA=9.684e-07
D4733 n4734 0 dm1 AREA=1.642e-06
D4734 n4735 0 dm1 AREA=1.130e-06
D4735 n4736 0 dm1 AREA=2.138e-07
D4736 n4737 0 dm1 AREA=7.361e-07
D4737 n4738 0 dm1 AREA=8.079e-07
D4738 n4739 0 dm1 AREA=1.245e-06
D4739 n4740 0 dm1 AREA=6.017e-07
D4740 n4741 0 dm1 AREA=1.173e-06
D4741 n4742 0 dm1 AREA=5.031e-07
D4742 n4743 0 dm1 AREA=1.444e-06
D4743 n4744 0 dm1 AREA=6.538e-07
D4744 n4745 0 dm1 AREA=1.676e-06
D4745 n4746 0 dm1 AREA=4.110e-07
D4746 n4747 0 dm1 AREA=1.522e-06
D4747 n4748 0 dm1 AREA=8.666e-07
D4748 n4749 0 dm1 AREA=9.732e-07
D4749 n4750 0 dm1 AREA=3.532e-07
D4750 n4751 0 dm1 AREA=1.222e-06
D4751 n4752 0 dm1 AREA=2.170e-06
D4752 n4753 0 dm1 AREA=1.017e-06
D4753 n4754 0 dm1 AREA=3.766e-07
D4754 n4755 0 dm1 AREA=4.555e-07
D4755 n4756 0 dm1 AREA=1.118e-06
D4756 n4757 0 dm1 AREA=1.612e-06
D4757 n4758 0 dm1 AREA=8.456e-07
D4758 n4759 0 dm1 AREA=1.280e-06
D4759 n4760 0 dm1 AREA=3.538e-07
D4760 n4761 0 dm1 AREA=9.195e-07
D4761 n4762 0 dm1 AREA=1.634e-06
D4762 n4763 0 dm1 AREA=1.337e-06
D4763 n4764 0 dm1 AREA=3.890e-07
D4764 n4765 0 dm1 AREA=1.657e-06
D4765 n4766 0 dm1 AREA=7.270e-07
D4766 n4767 0 dm1 AREA=6.937e-07
D4767 n4768 0 dm1 AREA=3.200e-07
D4768 n4769 0 dm1 AREA=1.337e-06
D4769 n4770 0 dm1 AREA=1.345e-06
D4770 n4771 0 dm1 AREA=8.278e-07
D4771 n4772 0 dm1 AREA=1.066e-06
D4772 n4773 0 dm1 AREA=1.140e-06
D4773 n4774 0 dm1 AREA=7.059e-07
D4774 n4775 0 dm1 AREA=1.059e-06
D4775 n4776 0 dm1 AREA=1.313e-06
D4776 n4777 0 dm1 AREA=1.440e-06
D4777 n4778 0 dm1 AREA=4.035e-07
D4778 n1 0 dm1 AREA=3.751e-07
D4779 n4780 0 dm1 AREA=1.271e-06
D4780 n4781 0 dm1 AREA=7.076e-07
D4781 n4782 0 dm1 AREA=7.602e-07
D4782 n4783 0 dm1 AREA=9.778e-07
D4783 n4784 0 dm1 AREA=9.722e-07
D4784 n4785 0 dm1 AREA=7.447e-07
D4785 n4786 0 dm1 AREA=5.884e-07
D4786 n4787 0 dm1 AREA=4.085e-07
D4787 n4788 0 dm1 AREA=8.302e-07
D4788 n4789 0 dm1 AREA=2.072e-06
D4789 n4790 0 dm1 AREA=8.547e-07
D4790 n4791 0 dm1 AREA=1.188e-06
D4791 n4792 0 dm1 AREA=2.215e-06
D4792 n4793 0 dm1 AREA=2.420e-07
D4793 n4794 0 dm1 AREA=1.245e-06
D4794 n4795 0 dm1 AREA=4.390e-07
D4795 n4796 0 dm1 AREA=4.431e-07
D4796 n4797 0 dm1 AREA=1.104e-06
D4797 n4798 0 dm1 AREA=1.274e-06
D4798 n4799 0 dm1 AREA=2.887e-07
D4799 n4800 0 dm1 AREA=2.443e-06
D4800 n4801 0 dm1 AREA=6.392e-07
D4801 n4802 0 dm1 AREA=1.761e-06
D4802 n4803 0 dm1 AREA=2.469e-06
D4803 n4804 0 dm1 AREA=7.483e-07
D4804 n4805 0 dm1 AREA=1.412e-06
D4805 n4806 0 dm1 AREA=1.193e-06
D4806 n4807 0 dm1 AREA=1.771e-06
D4807 n1 0 dm1 AREA=9.124e-07
D4808 n4809 0 dm1 AREA=1.379e-06
D4809 n4810 0 dm1 AREA=5.655e-07
D4810 n4811 0 dm1 AREA=9.968e-07
D4811 n4812 0 dm1 AREA=6.343e-07
D4812 n4813 0 dm1 AREA=8.651e-07
D4813 n4814 0 dm1 AREA=1.783e-06
D4814 n4815 0 dm1 AREA=8.734e-07
D4815 n4816 0 dm1 AREA=5.766e-07
D4816 n4817 0 dm1 AREA=2.751e-07
D4817 n4818 0 dm1 AREA=6.912e-07
D4818 n4819 0 dm1 AREA=9.673e-07
D4819 n4820 0 dm1 AREA=6.823e-07
D4820 n4821 0 dm1 AREA=4.447e-07
D4821 n4822 0 dm1 AREA=1.560e-06
D4822 n4823 0 dm1 AREA=1.925e-06
D4823 n4824 0 dm1 AREA=7.476e-07
D4824 n4825 0 dm1 AREA=4.740e-07
D4825 n4826 0 dm1 AREA=3.363e-07
D4826 n4827 0 dm1 AREA=1.751e-06
D4827 n4828 0 dm1 AREA=6.548e-07
D4828 n4829 0 dm1 AREA=1.872e-07
D4829 n4830 0 dm1 AREA=7.444e-07
D4830 n4831 0 dm1 AREA=1.209e-06
D4831 n4832 0 dm1 AREA=1.146e-06
D4832 n4833 0 dm1 AREA=8.973e-07
D4833 n4834 0 dm1 AREA=1.226e-06
D4834 n4835 0 dm1 AREA=3.120e-07
D4835 n4836 0 dm1 AREA=7.289e-07
D4836 n4837 0 dm1 AREA=3.702e-07
D4837 n4838 0 dm1 AREA=9.609e-07
D4838 n4839 0 dm1 AREA=5.808e-07
D4839 n4840 0 dm1 AREA=3.344e-07
D4840 n4841 0 dm1 AREA=1.399e-06
D4841 n4842 0 dm1 AREA=1.547e-06
D4842 n4843 0 dm1 AREA=1.143e-06
D4843 n4844 0 dm1 AREA=3.111e-07
D4844 n4845 0 dm1 AREA=1.063e-06
D4845 n4846 0 dm1 AREA=6.490e-07
D4846 n4847 0 dm1 AREA=9.578e-07
D4847 n4848 0 dm2 AREA=1.046e-06
D4848 n4849 0 dm2 AREA=7.614e-07
D4849 n4850 0 dm2 AREA=1.053e-06
D4850 n4851 0 dm2 AREA=1.328e-06
D4851 n4852 0 dm2 AREA=4.409e-07
D4852 n4853 0 dm2 AREA=1.204e-06
D4853 n4854 0 dm2 AREA=8.714e-07
D4854 n4855 0 dm2 AREA=3.476e-07
D4855 n4856 0 dm2 AREA=7.279e-07
D4856 n4857 0 dm2 AREA=4.012e-06
D4857 n4858 0 dm2 AREA=1.837e-06
D4858 n4859 0 dm2 AREA=9.303e-07
D4859 n4860 0 dm2 AREA=2.686e-07
D4860 n4861 0 dm2 AREA=8.868e-07
D4861 n4862 0 dm2 AREA=2.902e-07
D4862 n4863 0 dm2 AREA=5.308e-07
D4863 n4864 0 dm2 AREA=1.422e-06
D4864 n4865 0 dm2 AREA=9.156e-07
D4865 n4866 0 dm2 AREA=9.049e-07
D4866 n4867 0 dm2 AREA=1.857e-06
D4867 n4868 0 dm2 AREA=8.523e-07
D4868 n4869 0 dm2 AREA=9.346e-07
D4869 n4870 0 dm2 AREA=7.523e-07
D4870 n4871 0 dm2 AREA=1.171e-06
D4871 n4872 0 dm2 AREA=4.187e-07
D4872 n4873 0 dm2 AREA=9.190e-07
D4873 n4874 0 dm2 AREA=1.169e-06
D4874 n4875 0 dm2 AREA=4.616e-07
D4875 n4876 0 dm2 AREA=8.934e-07
D4876 n4877 0 dm2 AREA=1.450e-06
D4877 n4878 0 dm2 AREA=2.544e-07
D4878 n4879 0 dm2 AREA=1.144e-06
D4879 n4880 0 dm2 AREA=9.680e-07
D4880 n4881 0 dm2 AREA=6.387e-07
D4881 n4882 0 dm2 AREA=9.759e-07
D4882 n4883 0 dm2 AREA=7.238e-07
D4883 n4884 0 dm2 AREA=1.043e-06
D4884 n4885 0 dm2 AREA=3.366e-07
D4885 n4886 0 dm2 AREA=4.044e-07
D4886 n4887 0 dm2 AREA=1.745e-06
D4887 n4888 0 dm2 AREA=1.804e-06
D4888 n4889 0 dm2 AREA=1.170e-06
D4889 n4890 0 dm2 AREA=6.821e-07
D4890 n4891 0 dm2 AREA=2.558e-07
D4891 n4892 0 dm2 AREA=3.185e-07
D4892 n4893 0 dm2 AREA=7.170e-07
D4893 n4894 0 dm2 AREA=1.118e-06
D4894 n4895 0 dm2 AREA=5.745e-07
D4895 n4896 0 dm2 AREA=4.835e-07
D4896 n4897 0 dm2 AREA=6.224e-07
D4897 n4898 0 dm2 AREA=7.356e-07
D4898 n4899 0 dm2 AREA=8.107e-07
D4899 n4900 0 dm2 AREA=7.691e-07
D4900 n4901 0 dm2 AREA=8.602e-07
D4901 n4902 0 dm2 AREA=7.421e-07
D4902 n4903 0 dm2 AREA=1.344e-06
D4903 n4904 0 dm2 AREA=1.542e-06
D4904 n4905 0 dm2 AREA=6.035e-07
D4905 n4906 0 dm2 AREA=5.768e-07
D4906 n4907 0 dm2 AREA=6.036e-07
D4907 n4908 0 dm2 AREA=1.652e-06
D4908 n4909 0 dm2 AREA=2.023e-06
D4909 n4910 0 dm2 AREA=5.563e-07
D4910 n4911 0 dm2 AREA=5.590e-07
D4911 n4912 0 dm2 AREA=6.625e-07
D4912 n4913 0 dm2 AREA=2.097e-06
D4913 n4914 0 dm2 AREA=1.607e-06
D4914 n4915 0 dm2 AREA=3.663e-07
D4915 n4916 0 dm2 AREA=1.284e-06
D4916 n4917 0 dm2 AREA=6.208e-07
D4917 n4918 0 dm2 AREA=1.487e-06
D4918 n4919 0 dm2 AREA=8.912e-07
D4919 n1 0 dm2 AREA=3.125e-07
D4920 n4921 0 dm2 AREA=2.055e-06
D4921 n4922 0 dm2 AREA=8.014e-07
D4922 n4923 0 dm2 AREA=1.056e-06
D4923 n4924 0 dm2 AREA=1.310e-06
D4924 n4925 0 dm2 AREA=7.943e-07
D4925 n4926 0 dm2 AREA=5.858e-07
D4926 n4927 0 dm2 AREA=7.364e-07
D4927 n4928 0 dm2 AREA=8.525e-07
D4928 n4929 0 dm2 AREA=7.454e-07
D4929 n4930 0 dm2 AREA=1.269e-06
D4930 n4931 0 dm2 AREA=2.875e-06
D4931 n4932 0 dm2 AREA=1.105e-06
D4932 n4933 0 dm2 AREA=1.558e-07
D4933 n4934 0 dm2 AREA=1.888e-07
D4934 n4935 0 dm2 AREA=6.545e-07
D4935 n4936 0 dm2 AREA=6.274e-07
D4936 n4937 0 dm2 AREA=2.607e-06
D4937 n4938 0 dm2 AREA=1.343e-06
D4938 n4939 0 dm2 AREA=1.062e-06
D4939 n4940 0 dm2 AREA=6.856e-07
D4940 n4941 0 dm2 AREA=1.025e-06
D4941 n4942 0 dm2 AREA=1.246e-06
D4942 n4943 0 dm2 AREA=1.295e-06
D4943 n4944 0 dm2 AREA=1.016e-06
D4944 n4945 0 dm2 AREA=9.476e-07
D4945 n4946 0 dm2 AREA=2.738e-07
D4946 n4947 0 dm2 AREA=4.281e-07
D4947 n4948 0 dm2 AREA=4.377e-07
D4948 n4949 0 dm2 AREA=2.578e-06
D4949 n4950 0 dm2 AREA=5.885e-07
D4950 n4951 0 dm2 AREA=7.572e-07
D4951 n4952 0 dm2 AREA=9.881e-07
D4952 n4953 0 dm2 AREA=1.886e-06
D4953 n4954 0 dm2 AREA=3.354e-07
D4954 n4955 0 dm2 AREA=1.720e-06
D4955 n4956 0 dm2 AREA=7.478e-07
D4956 n4957 0 dm2 AREA=2.388e-06
D4957 n4958 0 dm2 AREA=7.157e-07
D4958 n4959 0 dm2 AREA=8.521e-07
D4959 n4960 0 dm2 AREA=3.183e-07
D4960 n4961 0 dm2 AREA=4.207e-07
D4961 n4962 0 dm2 AREA=1.446e-06
D4962 n4963 0 dm2 AREA=3.635e-07
D4963 n4964 0 dm2 AREA=8.401e-07
D4964 n4965 0 dm2 AREA=2.220e-07
D4965 n4966 0 dm2 AREA=1.910e-06
D4966 n4967 0 dm2 AREA=1.832e-06
D4967 n4968 0 dm2 AREA=1.112e-06
D4968 n4969 0 dm2 AREA=1.503e-06
D4969 n4970 0 dm2 AREA=8.235e-07
D4970 n4971 0 dm2 AREA=3.260e-07
D4971 n4972 0 dm2 AREA=8.690e-07
D4972 n4973 0 dm2 AREA=8.397e-07
D4973 n4974 0 dm2 AREA=9.962e-07
D4974 n4975 0 dm2 AREA=1.055e-06
D4975 n4976 0 dm2 AREA=9.329e-07
D4976 n4977 0 dm2 AREA=5.377e-07
D4977 n4978 0 dm2 AREA=1.724e-06
D4978 n4979 0 dm2 AREA=1.343e-06
D4979 n4980 0 dm2 AREA=1.334e-06
D4980 n4981 0 dm2 AREA=1.202e-06
D4981 n4982 0 dm2 AREA=2.907e-06
D4982 n4983 0 dm2 AREA=8.334e-07
D4983 n4984 0 dm2 AREA=1.427e-06
D4984 n4985 0 dm2 AREA=3.703e-07
D4985 n4986 0 dm2 AREA=9.487e-07
D4986 n4987 0 dm2 AREA=1.121e-06
D4987 n4988 0 dm2 AREA=2.594e-06
D4988 n4989 0 dm2 AREA=7.244e-07
D4989 n4990 0 dm2 AREA=9.051e-07
D4990 n4991 0 dm2 AREA=1.321e-06
D4991 n4992 0 dm2 AREA=1.421e-06
D4992 n4993 0 dm2 AREA=2.648e-06
D4993 n4994 0 dm2 AREA=1.101e-06
D4994 n4995 0 dm2 AREA=9.097e-07
D4995 n4996 0 dm2 AREA=1.831e-06
D4996 n1 0 dm2 AREA=1.000e-06
D4997 n4998 0 dm2 AREA=9.628e-07
D4998 n4999 0 dm2 AREA=1.485e-06
D4999 n5000 0 dm2 AREA=5.188e-07
D5000 n5001 0 dm2 AREA=2.183e-06
D5001 n5002 0 dm2 AREA=1.446e-06
D5002 n5003 0 dm2 AREA=2.108e-06
D5003 n5004 0 dm2 AREA=1.618e-06
D5004 n5005 0 dm2 AREA=6.537e-07
D5005 n5006 0 dm2 AREA=6.469e-07
D5006 n5007 0 dm2 AREA=2.414e-06
D5007 n5008 0 dm2 AREA=1.031e-06
D5008 n5009 0 dm2 AREA=4.610e-07
D5009 n5010 0 dm2 AREA=5.483e-07
D5010 n5011 0 dm2 AREA=1.326e-06
D5011 n5012 0 dm2 AREA=5.782e-07
D5012 n5013 0 dm2 AREA=1.350e-06
D5013 n5014 0 dm2 AREA=1.034e-06
D5014 n5015 0 dm2 AREA=2.047e-06
D5015 n5016 0 dm2 AREA=9.660e-07
D5016 n5017 0 dm2 AREA=4.306e-07
D5017 n5018 0 dm2 AREA=6.264e-07
D5018 n5019 0 dm2 AREA=8.126e-07
D5019 n5020 0 dm2 AREA=8.900e-07
D5020 n5021 0 dm2 AREA=7.378e-07
D5021 n5022 0 dm2 AREA=1.700e-07
D5022 n5023 0 dm2 AREA=5.695e-07
D5023 n5024 0 dm2 AREA=1.557e-06
D5024 n5025 0 dm2 AREA=3.888e-07
D5025 n5026 0 dm2 AREA=5.091e-07
D5026 n5027 0 dm2 AREA=6.649e-07
D5027 n5028 0 dm2 AREA=7.829e-07
D5028 n5029 0 dm2 AREA=6.270e-07
D5029 n5030 0 dm2 AREA=5.877e-07
D5030 n5031 0 dm2 AREA=1.155e-06
D5031 n5032 0 dm2 AREA=6.314e-07
D5032 n5033 0 dm2 AREA=3.843e-07
D5033 n5034 0 dm2 AREA=3.390e-07
D5034 n5035 0 dm2 AREA=2.038e-06
D5035 n5036 0 dm2 AREA=9.973e-07
D5036 n5037 0 dm2 AREA=1.184e-06
D5037 n5038 0 dm2 AREA=1.340e-06
D5038 n5039 0 dm2 AREA=1.651e-07
D5039 n5040 0 dm2 AREA=7.603e-07
D5040 n5041 0 dm2 AREA=7.741e-07
D5041 n5042 0 dm2 AREA=7.156e-07
D5042 n5043 0 dm2 AREA=1.331e-06
D5043 n5044 0 dm2 AREA=2.924e-07
D5044 n5045 0 dm2 AREA=1.390e-06
D5045 n5046 0 dm2 AREA=3.589e-07
D5046 n5047 0 dm2 AREA=4.495e-07
D5047 n5048 0 dm2 AREA=7.244e-07
D5048 n5049 0 dm2 AREA=1.151e-06
D5049 n5050 0 dm2 AREA=9.764e-07
D5050 n5051 0 dm2 AREA=3.893e-07
D5051 n5052 0 dm2 AREA=1.686e-06
D5052 n5053 0 dm2 AREA=9.205e-07
D5053 n5054 0 dm2 AREA=8.258e-07
D5054 n5055 0 dm2 AREA=1.018e-06
D5055 n5056 0 dm2 AREA=1.325e-06
D5056 n5057 0 dm2 AREA=9.168e-07
D5057 n5058 0 dm2 AREA=1.206e-06
D5058 n5059 0 dm2 AREA=9.646e-07
D5059 n5060 0 dm2 AREA=8.015e-07
D5060 n5061 0 dm2 AREA=2.013e-06
D5061 n5062 0 dm2 AREA=4.647e-07
D5062 n5063 0 dm2 AREA=6.884e-07
D5063 n5064 0 dm2 AREA=1.189e-06
D5064 n5065 0 dm2 AREA=1.534e-06
D5065 n5066 0 dm2 AREA=8.549e-07
D5066 n5067 0 dm2 AREA=5.895e-07
D5067 n5068 0 dm2 AREA=5.794e-07
D5068 n5069 0 dm2 AREA=6.845e-07
D5069 n5070 0 dm2 AREA=1.537e-06
D5070 n5071 0 dm2 AREA=5.793e-07
D5071 n5072 0 dm2 AREA=1.932e-06
D5072 n5073 0 dm2 AREA=1.390e-06
D5073 n5074 0 dm2 AREA=1.135e-06
D5074 n5075 0 dm2 AREA=8.154e-07
D5075 n5076 0 dm2 AREA=4.848e-07
D5076 n5077 0 dm2 AREA=2.621e-07
D5077 n5078 0 dm2 AREA=5.245e-07
D5078 n5079 0 dm2 AREA=1.344e-06
D5079 n5080 0 dm2 AREA=1.082e-06
D5080 n5081 0 dm2 AREA=1.265e-06
D5081 n5082 0 dm2 AREA=1.383e-06
D5082 n5083 0 dm2 AREA=1.251e-06
D5083 n5084 0 dm2 AREA=8.326e-07
D5084 n5085 0 dm2 AREA=1.623e-06
D5085 n5086 0 dm2 AREA=1.991e-06
D5086 n5087 0 dm2 AREA=6.515e-07
D5087 n5088 0 dm2 AREA=1.032e-06
D5088 n5089 0 dm2 AREA=5.068e-07
D5089 n5090 0 dm2 AREA=6.705e-07
D5090 n5091 0 dm2 AREA=1.734e-06
D5091 n5092 0 dm2 AREA=1.420e-06
D5092 n5093 0 dm2 AREA=7.939e-07
D5093 n5094 0 dm2 AREA=3.395e-07
D5094 n1 0 dm2 AREA=4.032e-07
D5095 n5096 0 dm2 AREA=8.039e-07
D5096 n5097 0 dm2 AREA=3.698e-07
D5097 n5098 0 dm2 AREA=4.993e-07
D5098 n5099 0 dm2 AREA=1.188e-06
D5099 n5100 0 dm2 AREA=1.595e-06
D5100 n5101 0 dm2 AREA=1.940e-06
D5101 n5102 0 dm2 AREA=9.582e-07
D5102 n5103 0 dm2 AREA=1.187e-06
D5103 n5104 0 dm2 AREA=6.970e-07
D5104 n5105 0 dm2 AREA=1.021e-06
D5105 n5106 0 dm2 AREA=6.657e-07
D5106 n5107 0 dm2 AREA=7.126e-07
D5107 n5108 0 dm2 AREA=1.190e-06
D5108 n5109 0 dm2 AREA=5.948e-07
D5109 n5110 0 dm2 AREA=5.510e-07
D5110 n5111 0 dm2 AREA=1.929e-06
D5111 n5112 0 dm2 AREA=3.678e-07
D5112 n5113 0 dm2 AREA=9.511e-07
D5113 n5114 0 dm2 AREA=1.214e-06
D5114 n5115 0 dm2 AREA=8.266e-07
D5115 n5116 0 dm2 AREA=7.226e-07
D5116 n5117 0 dm2 AREA=4.822e-07
D5117 n5118 0 dm2 AREA=8.821e-07
D5118 n5119 0 dm2 AREA=1.099e-06
D5119 n5120 0 dm2 AREA=3.654e-07
D5120 n5121 0 dm2 AREA=1.129e-06
D5121 n5122 0 dm2 AREA=8.076e-07
D5122 n5123 0 dm2 AREA=1.746e-06
D5123 n5124 0 dm2 AREA=1.308e-06
D5124 n5125 0 dm2 AREA=8.004e-07
D5125 n5126 0 dm2 AREA=2.776e-07
D5126 n5127 0 dm2 AREA=1.133e-06
D5127 n5128 0 dm2 AREA=1.324e-06
D5128 n5129 0 dm2 AREA=1.443e-06
D5129 n5130 0 dm2 AREA=7.094e-07
D5130 n5131 0 dm2 AREA=8.073e-07
D5131 n5132 0 dm2 AREA=1.303e-06
D5132 n5133 0 dm2 AREA=1.423e-06
D5133 n5134 0 dm2 AREA=9.717e-07
D5134 n5135 0 dm2 AREA=2.361e-07
D5135 n5136 0 dm2 AREA=2.498e-07
D5136 n5137 0 dm2 AREA=7.545e-07
D5137 n5138 0 dm2 AREA=1.070e-06
D5138 n5139 0 dm2 AREA=7.045e-07
D5139 n5140 0 dm2 AREA=6.116e-07
D5140 n5141 0 dm2 AREA=4.974e-07
D5141 n5142 0 dm2 AREA=1.427e-06
D5142 n5143 0 dm2 AREA=8.906e-07
D5143 n5144 0 dm2 AREA=1.208e-06
D5144 n5145 0 dm2 AREA=9.229e-07
D5145 n5146 0 dm2 AREA=1.438e-06
D5146 n5147 0 dm2 AREA=1.562e-06
D5147 n5148 0 dm2 AREA=1.409e-07
D5148 n5149 0 dm2 AREA=1.176e-06
D5149 n5150 0 dm2 AREA=9.290e-07
D5150 n5151 0 dm2 AREA=2.235e-06
D5151 n5152 0 dm2 AREA=1.107e-06
D5152 n5153 0 dm2 AREA=4.809e-07
D5153 n5154 0 dm2 AREA=1.253e-06
D5154 n5155 0 dm2 AREA=2.488e-07
D5155 n5156 0 dm2 AREA=1.777e-06
D5156 n5157 0 dm2 AREA=7.559e-07
D5157 n5158 0 dm2 AREA=1.003e-06
D5158 n5159 0 dm2 AREA=6.154e-07
D5159 n5160 0 dm2 AREA=5.843e-07
D5160 n5161 0 dm2 AREA=4.649e-07
D5161 n5162 0 dm2 AREA=4.749e-07
D5162 n5163 0 dm2 AREA=8.593e-07
D5163 n5164 0 dm2 AREA=1.167e-06
D5164 n5165 0 dm2 AREA=1.137e-06
D5165 n5166 0 dm2 AREA=3.195e-07
D5166 n5167 0 dm2 AREA=8.925e-07
D5167 n5168 0 dm2 AREA=5.451e-07
D5168 n5169 0 dm2 AREA=1.183e-06
D5169 n5170 0 dm2 AREA=1.144e-06
D5170 n5171 0 dm2 AREA=3.620e-07
D5171 n5172 0 dm2 AREA=4.163e-07
D5172 n5173 0 dm2 AREA=9.836e-07
D5173 n5174 0 dm2 AREA=7.003e-07
D5174 n5175 0 dm2 AREA=6.543e-07
D5175 n5176 0 dm2 AREA=1.220e-06
D5176 n5177 0 dm2 AREA=3.973e-07
D5177 n5178 0 dm2 AREA=5.614e-07
D5178 n5179 0 dm2 AREA=4.510e-07
D5179 n5180 0 dm2 AREA=1.485e-06
D5180 n5181 0 dm2 AREA=1.469e-06
D5181 n5182 0 dm2 AREA=9.666e-07
D5182 n5183 0 dm2 AREA=6.918e-07
D5183 n5184 0 dm2 AREA=1.922e-07
D5184 n5185 0 dm2 AREA=7.631e-07
D5185 n5186 0 dm2 AREA=1.296e-06
D5186 n5187 0 dm2 AREA=1.404e-06
D5187 n5188 0 dm2 AREA=8.764e-07
D5188 n5189 0 dm2 AREA=3.220e-07
D5189 n5190 0 dm2 AREA=1.118e-06
D5190 n5191 0 dm2 AREA=3.030e-07
D5191 n5192 0 dm2 AREA=7.597e-07
D5192 n5193 0 dm2 AREA=3.521e-07
D5193 n5194 0 dm2 AREA=1.369e-06
D5194 n5195 0 dm2 AREA=4.260e-07
D5195 n5196 0 dm2 AREA=1.192e-06
D5196 n5197 0 dm2 AREA=1.150e-06
D5197 n5198 0 dm2 AREA=2.148e-07
D5198 n5199 0 dm2 AREA=2.094e-06
D5199 n5200 0 dm2 AREA=3.264e-07
D5200 n5201 0 dm2 AREA=4.653e-07
D5201 n5202 0 dm2 AREA=6.667e-07
D5202 n5203 0 dm2 AREA=2.075e-07
D5203 n5204 0 dm2 AREA=1.607e-06
D5204 n5205 0 dm2 AREA=1.069e-06
D5205 n5206 0 dm2 AREA=8.965e-07
D5206 n5207 0 dm2 AREA=7.218e-07
D5207 n5208 0 dm2 AREA=1.173e-06
D5208 n5209 0 dm2 AREA=1.344e-06
D5209 n1 0 dm2 AREA=6.978e-07
D5210 n5211 0 dm2 AREA=2.867e-06
D5211 n5212 0 dm2 AREA=7.528e-07
D5212 n5213 0 dm2 AREA=1.022e-06
D5213 n5214 0 dm2 AREA=1.075e-06
D5214 n5215 0 dm2 AREA=1.349e-06
D5215 n5216 0 dm2 AREA=6.489e-07
D5216 n5217 0 dm2 AREA=5.055e-07
D5217 n5218 0 dm2 AREA=8.185e-07
D5218 n5219 0 dm2 AREA=1.035e-06
D5219 n5220 0 dm2 AREA=1.269e-06
D5220 n5221 0 dm2 AREA=1.299e-06
D5221 n5222 0 dm2 AREA=5.758e-07
D5222 n5223 0 dm2 AREA=1.769e-06
D5223 n5224 0 dm2 AREA=3.758e-07
D5224 n5225 0 dm2 AREA=1.199e-06
D5225 n5226 0 dm2 AREA=1.646e-07
D5226 n5227 0 dm2 AREA=4.583e-07
D5227 n5228 0 dm2 AREA=1.012e-06
D5228 n5229 0 dm2 AREA=8.616e-07
D5229 n5230 0 dm2 AREA=1.763e-07
D5230 n5231 0 dm2 AREA=5.722e-07
D5231 n5232 0 dm2 AREA=1.305e-07
D5232 n5233 0 dm2 AREA=9.308e-07
D5233 n5234 0 dm2 AREA=9.161e-07
D5234 n5235 0 dm2 AREA=6.711e-07
D5235 n5236 0 dm2 AREA=5.345e-07
D5236 n5237 0 dm2 AREA=2.724e-07
D5237 n5238 0 dm2 AREA=1.684e-06
D5238 n5239 0 dm2 AREA=7.514e-07
D5239 n5240 0 dm2 AREA=1.442e-06
D5240 n5241 0 dm2 AREA=5.889e-07
D5241 n5242 0 dm2 AREA=8.515e-07
D5242 n5243 0 dm2 AREA=3.208e-07
D5243 n1 0 dm2 AREA=1.390e-06
D5244 n5245 0 dm2 AREA=4.197e-07
D5245 n5246 0 dm2 AREA=2.239e-06
D5246 n5247 0 dm2 AREA=1.161e-06
D5247 n5248 0 dm2 AREA=7.479e-07
D5248 n5249 0 dm2 AREA=5.327e-07
D5249 n5250 0 dm2 AREA=6.708e-07
D5250 n5251 0 dm2 AREA=1.242e-06
D5251 n5252 0 dm2 AREA=2.784e-07
D5252 n5253 0 dm2 AREA=2.420e-07
D5253 n5254 0 dm2 AREA=1.748e-06
D5254 n5255 0 dm2 AREA=1.052e-06
D5255 n5256 0 dm2 AREA=2.003e-06
D5256 n5257 0 dm2 AREA=1.570e-06
D5257 n5258 0 dm2 AREA=7.546e-07
D5258 n5259 0 dm2 AREA=4.515e-07
D5259 n5260 0 dm2 AREA=1.214e-06
D5260 n5261 0 dm2 AREA=8.871e-07
D5261 n5262 0 dm2 AREA=6.020e-07
D5262 n5263 0 dm2 AREA=1.205e-06
D5263 n5264 0 dm2 AREA=4.606e-07
D5264 n5265 0 dm2 AREA=1.702e-06
D5265 n5266 0 dm2 AREA=6.798e-07
D5266 n5267 0 dm2 AREA=6.368e-07
D5267 n5268 0 dm2 AREA=2.154e-07
D5268 n5269 0 dm2 AREA=2.515e-07
D5269 n5270 0 dm2 AREA=1.283e-06
D5270 n5271 0 dm2 AREA=8.802e-07
D5271 n5272 0 dm2 AREA=3.179e-07
D5272 n5273 0 dm2 AREA=2.547e-07
D5273 n5274 0 dm2 AREA=1.325e-06
D5274 n5275 0 dm2 AREA=1.716e-06
D5275 n5276 0 dm2 AREA=3.952e-07
D5276 n5277 0 dm2 AREA=1.055e-06
D5277 n5278 0 dm2 AREA=1.097e-06
D5278 n5279 0 dm2 AREA=1.306e-06
D5279 n5280 0 dm2 AREA=1.798e-06
D5280 n5281 0 dm2 AREA=5.670e-07
D5281 n5282 0 dm2 AREA=8.507e-07
D5282 n5283 0 dm2 AREA=9.775e-07
D5283 n5284 0 dm2 AREA=2.364e-07
D5284 n5285 0 dm2 AREA=9.483e-07
D5285 n5286 0 dm2 AREA=1.045e-06
D5286 n5287 0 dm2 AREA=8.461e-07
D5287 n5288 0 dm2 AREA=5.995e-07
D5288 n5289 0 dm2 AREA=7.001e-07
D5289 n5290 0 dm2 AREA=2.833e-07
D5290 n5291 0 dm2 AREA=1.314e-06
D5291 n5292 0 dm2 AREA=1.332e-06
D5292 n5293 0 dm2 AREA=1.404e-06
D5293 n5294 0 dm2 AREA=1.043e-06
D5294 n5295 0 dm2 AREA=9.204e-07
D5295 n5296 0 dm2 AREA=1.416e-06
D5296 n5297 0 dm2 AREA=2.117e-06
D5297 n5298 0 dm2 AREA=2.144e-07
D5298 n5299 0 dm2 AREA=7.369e-07
D5299 n5300 0 dm2 AREA=9.461e-07
D5300 n5301 0 dm2 AREA=5.026e-07
D5301 n5302 0 dm2 AREA=5.388e-07
D5302 n5303 0 dm2 AREA=2.453e-07
D5303 n5304 0 dm2 AREA=5.823e-07
D5304 n5305 0 dm2 AREA=6.598e-07
D5305 n5306 0 dm2 AREA=3.787e-07
D5306 n5307 0 dm2 AREA=9.436e-07
D5307 n5308 0 dm2 AREA=6.058e-07
D5308 n5309 0 dm2 AREA=2.696e-07
D5309 n5310 0 dm2 AREA=8.503e-07
D5310 n5311 0 dm2 AREA=1.564e-06
D5311 n5312 0 dm2 AREA=1.801e-06
D5312 n5313 0 dm2 AREA=7.214e-07
D5313 n5314 0 dm2 AREA=1.308e-06
D5314 n5315 0 dm2 AREA=5.606e-07
D5315 n5316 0 dm2 AREA=6.878e-07
D5316 n5317 0 dm2 AREA=6.703e-07
D5317 n5318 0 dm2 AREA=1.387e-06
D5318 n5319 0 dm2 AREA=1.089e-06
D5319 n5320 0 dm2 AREA=4.618e-07
D5320 n5321 0 dm2 AREA=2.499e-07
D5321 n5322 0 dm2 AREA=7.210e-07
D5322 n5323 0 dm2 AREA=7.848e-07
D5323 n5324 0 dm2 AREA=1.477e-06
D5324 n5325 0 dm2 AREA=8.349e-07
D5325 n5326 0 dm2 AREA=3.935e-07
D5326 n5327 0 dm2 AREA=1.227e-06
D5327 n5328 0 dm2 AREA=2.139e-06
D5328 n5329 0 dm2 AREA=3.723e-07
D5329 n5330 0 dm2 AREA=1.248e-06
D5330 n5331 0 dm2 AREA=9.141e-07
D5331 n5332 0 dm2 AREA=5.783e-07
D5332 n5333 0 dm2 AREA=2.254e-06
D5333 n5334 0 dm2 AREA=3.276e-07
D5334 n5335 0 dm2 AREA=1.578e-06
D5335 n5336 0 dm2 AREA=3.298e-07
D5336 n5337 0 dm2 AREA=1.061e-06
D5337 n5338 0 dm2 AREA=9.671e-07
D5338 n5339 0 dm2 AREA=1.295e-06
D5339 n5340 0 dm2 AREA=1.299e-06
D5340 n5341 0 dm2 AREA=1.155e-06
D5341 n5342 0 dm2 AREA=7.233e-07
D5342 n5343 0 dm2 AREA=5.343e-07
D5343 n5344 0 dm2 AREA=4.430e-07
D5344 n5345 0 dm2 AREA=7.275e-07
D5345 n5346 0 dm2 AREA=9.684e-07
D5346 n5347 0 dm2 AREA=8.046e-07
D5347 n5348 0 dm2 AREA=1.688e-07
D5348 n5349 0 dm2 AREA=9.796e-07
D5349 n5350 0 dm2 AREA=1.060e-06
D5350 n5351 0 dm2 AREA=8.965e-07
D5351 n5352 0 dm2 AREA=2.814e-07
D5352 n5353 0 dm2 AREA=4.814e-07
D5353 n5354 0 dm2 AREA=8.295e-07
D5354 n5355 0 dm2 AREA=1.094e-06
D5355 n5356 0 dm2 AREA=9.000e-07
D5356 n5357 0 dm2 AREA=4.412e-07
D5357 n5358 0 dm2 AREA=1.352e-06
D5358 n5359 0 dm2 AREA=1.342e-06
D5359 n5360 0 dm2 AREA=4.872e-07
D5360 n5361 0 dm2 AREA=1.045e-06
D5361 n5362 0 dm2 AREA=9.111e-07
D5362 n5363 0 dm2 AREA=1.313e-06
D5363 n5364 0 dm2 AREA=1.540e-06
D5364 n5365 0 dm2 AREA=1.236e-06
D5365 n5366 0 dm2 AREA=2.400e-06
D5366 n5367 0 dm2 AREA=1.760e-06
D5367 n5368 0 dm2 AREA=6.904e-08
D5368 n5369 0 dm2 AREA=1.772e-07
D5369 n5370 0 dm2 AREA=8.096e-07
D5370 n5371 0 dm2 AREA=2.098e-06
D5371 n5372 0 dm2 AREA=8.861e-07
D5372 n5373 0 dm2 AREA=1.494e-06
D5373 n5374 0 dm2 AREA=6.265e-07
D5374 n5375 0 dm2 AREA=2.348e-06
D5375 n5376 0 dm2 AREA=5.884e-07
D5376 n5377 0 dm2 AREA=1.762e-07
D5377 n5378 0 dm2 AREA=5.182e-07
D5378 n5379 0 dm2 AREA=8.774e-07
D5379 n5380 0 dm2 AREA=1.027e-06
D5380 n5381 0 dm2 AREA=4.558e-07
D5381 n5382 0 dm2 AREA=7.521e-07
D5382 n5383 0 dm2 AREA=6.567e-07
D5383 n5384 0 dm2 AREA=9.371e-07
D5384 n5385 0 dm2 AREA=2.434e-06
D5385 n5386 0 dm2 AREA=7.716e-07
D5386 n5387 0 dm2 AREA=6.949e-07
D5387 n5388 0 dm2 AREA=1.036e-06
D5388 n5389 0 dm2 AREA=9.503e-07
D5389 n5390 0 dm2 AREA=7.684e-07
D5390 n5391 0 dm2 AREA=2.349e-06
D5391 n5392 0 dm2 AREA=9.470e-07
D5392 n5393 0 dm2 AREA=4.759e-07
D5393 n5394 0 dm2 AREA=6.734e-07
D5394 n5395 0 dm2 AREA=5.288e-07
D5395 n5396 0 dm2 AREA=7.910e-07
D5396 n5397 0 dm2 AREA=5.639e-07
D5397 n5398 0 dm2 AREA=8.941e-07
D5398 n5399 0 dm2 AREA=3.689e-07
D5399 n5400 0 dm2 AREA=9.194e-07
D5400 n5401 0 dm2 AREA=1.105e-06
D5401 n5402 0 dm2 AREA=2.506e-06
D5402 n5403 0 dm2 AREA=2.284e-06
D5403 n5404 0 dm2 AREA=1.371e-06
D5404 n5405 0 dm2 AREA=5.407e-07
D5405 n5406 0 dm2 AREA=1.207e-06
D5406 n5407 0 dm2 AREA=1.161e-06
D5407 n5408 0 dm2 AREA=7.868e-07
D5408 n5409 0 dm2 AREA=8.129e-07
D5409 n5410 0 dm2 AREA=1.307e-06
D5410 n5411 0 dm2 AREA=1.326e-06
D5411 n5412 0 dm2 AREA=1.189e-06
D5412 n5413 0 dm2 AREA=3.866e-07
D5413 n5414 0 dm2 AREA=1.176e-06
D5414 n5415 0 dm2 AREA=1.427e-06
D5415 n5416 0 dm2 AREA=1.846e-07
D5416 n5417 0 dm2 AREA=7.639e-07
D5417 n5418 0 dm2 AREA=7.399e-07
D5418 n5419 0 dm2 AREA=2.045e-06
D5419 n5420 0 dm2 AREA=1.555e-06
D5420 n5421 0 dm2 AREA=8.036e-07
D5421 n5422 0 dm2 AREA=4.920e-07
D5422 n5423 0 dm2 AREA=5.411e-07
D5423 n5424 0 dm2 AREA=7.185e-07
D5424 n5425 0 dm2 AREA=4.957e-07
D5425 n5426 0 dm2 AREA=5.996e-07
D5426 n5427 0 dm2 AREA=1.281e-06
D5427 n5428 0 dm2 AREA=1.467e-06
D5428 n5429 0 dm2 AREA=9.382e-07
D5429 n5430 0 dm2 AREA=6.983e-07
D5430 n5431 0 dm2 AREA=1.168e-06
D5431 n5432 0 dm2 AREA=1.242e-06
D5432 n5433 0 dm2 AREA=1.219e-06
D5433 n5434 0 dm2 AREA=1.208e-06
D5434 n5435 0 dm2 AREA=5.811e-07
D5435 n5436 0 dm2 AREA=8.932e-07
D5436 n5437 0 dm2 AREA=1.111e-06
D5437 n5438 0 dm2 AREA=1.640e-06
D5438 n5439 0 dm2 AREA=5.352e-07
D5439 n5440 0 dm2 AREA=2.452e-06
D5440 n5441 0 dm2 AREA=3.886e-07
D5441 n5442 0 dm2 AREA=9.856e-07
D5442 n5443 0 dm2 AREA=1.556e-06
D5443 n5444 0 dm2 AREA=1.191e-06
D5444 n5445 0 dm2 AREA=4.370e-07
D5445 n5446 0 dm2 AREA=8.786e-07
D5446 n5447 0 dm2 AREA=8.432e-07
D5447 n5448 0 dm2 AREA=6.067e-07
D5448 n5449 0 dm2 AREA=1.462e-06
D5449 n5450 0 dm2 AREA=7.166e-07
D5450 n5451 0 dm2 AREA=3.072e-07
D5451 n5452 0 dm2 AREA=1.574e-06
D5452 n5453 0 dm2 AREA=9.093e-07
D5453 n5454 0 dm2 AREA=2.891e-06
D5454 n5455 0 dm2 AREA=7.072e-07
D5455 n5456 0 dm2 AREA=1.291e-06
D5456 n5457 0 dm2 AREA=1.569e-06
D5457 n5458 0 dm2 AREA=1.815e-06
D5458 n5459 0 dm2 AREA=1.368e-06
D5459 n5460 0 dm2 AREA=6.825e-07
D5460 n5461 0 dm2 AREA=5.995e-07
D5461 n5462 0 dm2 AREA=1.598e-06
D5462 n1 0 dm2 AREA=7.589e-07
D5463 n5464 0 dm2 AREA=1.031e-06
D5464 n5465 0 dm2 AREA=8.655e-07
D5465 n5466 0 dm2 AREA=7.245e-07
D5466 n5467 0 dm2 AREA=1.012e-06
D5467 n5468 0 dm2 AREA=1.103e-06
D5468 n5469 0 dm2 AREA=1.143e-06
D5469 n5470 0 dm2 AREA=8.380e-07
D5470 n5471 0 dm2 AREA=1.209e-06
D5471 n5472 0 dm2 AREA=3.073e-07
D5472 n5473 0 dm2 AREA=9.071e-07
D5473 n5474 0 dm2 AREA=4.829e-07
D5474 n5475 0 dm2 AREA=3.433e-07
D5475 n5476 0 dm2 AREA=4.926e-07
D5476 n5477 0 dm2 AREA=5.980e-07
D5477 n5478 0 dm2 AREA=1.149e-06
D5478 n5479 0 dm2 AREA=8.801e-07
D5479 n5480 0 dm2 AREA=5.020e-07
D5480 n5481 0 dm2 AREA=9.801e-07
D5481 n5482 0 dm2 AREA=1.056e-06
D5482 n5483 0 dm2 AREA=1.001e-06
D5483 n5484 0 dm2 AREA=1.369e-06
D5484 n5485 0 dm2 AREA=9.767e-07
D5485 n5486 0 dm2 AREA=5.177e-07
D5486 n5487 0 dm2 AREA=6.527e-07
D5487 n5488 0 dm2 AREA=1.491e-06
D5488 n5489 0 dm2 AREA=1.394e-06
D5489 n5490 0 dm2 AREA=1.196e-06
D5490 n5491 0 dm2 AREA=7.104e-07
D5491 n5492 0 dm2 AREA=1.188e-06
D5492 n5493 0 dm2 AREA=3.055e-07
D5493 n5494 0 dm2 AREA=5.677e-07
D5494 n5495 0 dm2 AREA=1.255e-06
D5495 n5496 0 dm2 AREA=3.502e-07
D5496 n5497 0 dm2 AREA=9.397e-07
D5497 n5498 0 dm2 AREA=1.303e-06
D5498 n5499 0 dm2 AREA=3.181e-06
D5499 n5500 0 dm2 AREA=1.434e-06
D5500 n5501 0 dm2 AREA=9.352e-07
D5501 n5502 0 dm2 AREA=4.204e-07
D5502 n5503 0 dm2 AREA=8.260e-07
D5503 n1 0 dm2 AREA=5.417e-07
D5504 n5505 0 dm2 AREA=2.153e-06
D5505 n5506 0 dm2 AREA=2.956e-07
D5506 n5507 0 dm2 AREA=1.670e-06
D5507 n5508 0 dm2 AREA=7.773e-07
D5508 n5509 0 dm2 AREA=7.023e-07
D5509 n5510 0 dm2 AREA=4.563e-07
D5510 n5511 0 dm2 AREA=8.592e-07
D5511 n5512 0 dm2 AREA=5.534e-07
D5512 n5513 0 dm2 AREA=6.994e-07
D5513 n5514 0 dm2 AREA=1.165e-06
D5514 n5515 0 dm2 AREA=1.376e-06
D5515 n5516 0 dm2 AREA=2.477e-06
D5516 n5517 0 dm2 AREA=6.183e-07
D5517 n5518 0 dm2 AREA=6.515e-07
D5518 n5519 0 dm2 AREA=7.284e-07
D5519 n5520 0 dm2 AREA=1.541e-06
D5520 n5521 0 dm2 AREA=1.510e-06
D5521 n5522 0 dm2 AREA=1.160e-06
D5522 n5523 0 dm2 AREA=8.133e-07
D5523 n1 0 dm2 AREA=3.191e-07
D5524 n5525 0 dm2 AREA=7.955e-07
D5525 n5526 0 dm2 AREA=6.398e-07
D5526 n5527 0 dm2 AREA=2.069e-06
D5527 n5528 0 dm2 AREA=1.124e-06
D5528 n5529 0 dm2 AREA=6.838e-07
D5529 n5530 0 dm2 AREA=5.466e-07
D5530 n5531 0 dm2 AREA=5.453e-07
D5531 n5532 0 dm2 AREA=2.404e-06
D5532 n5533 0 dm2 AREA=1.018e-06
D5533 n5534 0 dm2 AREA=6.538e-07
D5534 n5535 0 dm2 AREA=9.133e-07
D5535 n5536 0 dm2 AREA=6.155e-07
D5536 n5537 0 dm2 AREA=6.219e-07
D5537 n5538 0 dm2 AREA=6.797e-07
D5538 n5539 0 dm2 AREA=4.600e-07
D5539 n5540 0 dm2 AREA=8.972e-07
D5540 n5541 0 dm2 AREA=6.791e-07
D5541 n5542 0 dm2 AREA=9.833e-07
D5542 n5543 0 dm2 AREA=1.333e-06
D5543 n5544 0 dm2 AREA=9.160e-07
D5544 n5545 0 dm2 AREA=1.663e-06
D5545 n5546 0 dm2 AREA=1.809e-06
D5546 n5547 0 dm2 AREA=1.387e-06
D5547 n5548 0 dm2 AREA=1.445e-06
D5548 n5549 0 dm2 AREA=1.045e-06
D5549 n5550 0 dm2 AREA=4.297e-07
D5550 n5551 0 dm2 AREA=1.577e-06
D5551 n5552 0 dm2 AREA=6.999e-07
D5552 n5553 0 dm2 AREA=1.385e-06
D5553 n5554 0 dm2 AREA=1.104e-06
D5554 n5555 0 dm2 AREA=1.336e-06
D5555 n5556 0 dm2 AREA=7.614e-07
D5556 n5557 0 dm2 AREA=9.728e-07
D5557 n5558 0 dm2 AREA=2.814e-06
D5558 n5559 0 dm2 AREA=8.780e-07
D5559 n5560 0 dm2 AREA=1.331e-06
D5560 n5561 0 dm2 AREA=5.211e-07
D5561 n5562 0 dm2 AREA=5.382e-07
D5562 n5563 0 dm2 AREA=1.141e-06
D5563 n5564 0 dm2 AREA=1.846e-06
D5564 n5565 0 dm2 AREA=1.577e-06
D5565 n5566 0 dm2 AREA=5.229e-07
D5566 n5567 0 dm2 AREA=6.791e-07
D5567 n5568 0 dm2 AREA=4.545e-07
D5568 n5569 0 dm2 AREA=6.619e-07
D5569 n5570 0 dm2 AREA=8.432e-07
D5570 n1 0 dm2 AREA=2.994e-07
D5571 n5572 0 dm2 AREA=1.733e-06
D5572 n5573 0 dm2 AREA=1.706e-06
D5573 n5574 0 dm2 AREA=8.488e-07
D5574 n5575 0 dm2 AREA=1.342e-06
D5575 n5576 0 dm2 AREA=1.296e-06
D5576 n5577 0 dm2 AREA=1.460e-06
D5577 n5578 0 dm2 AREA=7.540e-07
D5578 n5579 0 dm2 AREA=5.345e-07
D5579 n5580 0 dm2 AREA=5.001e-07
D5580 n5581 0 dm2 AREA=1.115e-06
D5581 n5582 0 dm2 AREA=7.876e-07
D5582 n5583 0 dm2 AREA=1.537e-06
D5583 n5584 0 dm2 AREA=4.665e-07
D5584 n5585 0 dm2 AREA=1.319e-06
D5585 n5586 0 dm2 AREA=8.413e-07
D5586 n5587 0 dm2 AREA=1.448e-06
D5587 n5588 0 dm2 AREA=7.847e-07
D5588 n5589 0 dm2 AREA=2.008e-06
D5589 n5590 0 dm2 AREA=6.705e-07
D5590 n5591 0 dm2 AREA=1.168e-06
D5591 n5592 0 dm2 AREA=1.038e-06
D5592 n5593 0 dm2 AREA=1.961e-06
D5593 n5594 0 dm2 AREA=1.069e-06
D5594 n5595 0 dm2 AREA=1.100e-06
D5595 n5596 0 dm2 AREA=4.956e-07
D5596 n5597 0 dm2 AREA=3.639e-07
D5597 n5598 0 dm2 AREA=1.180e-06
D5598 n5599 0 dm2 AREA=9.677e-07
D5599 n5600 0 dm2 AREA=1.276e-06
D5600 n5601 0 dm2 AREA=1.326e-06
D5601 n5602 0 dm2 AREA=4.969e-07
D5602 n1 0 dm2 AREA=1.445e-06
D5603 n5604 0 dm2 AREA=8.921e-07
D5604 n5605 0 dm2 AREA=3.784e-07
D5605 n5606 0 dm2 AREA=6.814e-07
D5606 n5607 0 dm2 AREA=1.066e-06
D5607 n5608 0 dm2 AREA=9.867e-07
D5608 n5609 0 dm2 AREA=7.303e-07
D5609 n5610 0 dm2 AREA=6.324e-07
D5610 n5611 0 dm2 AREA=2.216e-06
D5611 n5612 0 dm2 AREA=7.338e-07
D5612 n5613 0 dm2 AREA=1.517e-07
D5613 n5614 0 dm2 AREA=8.546e-07
D5614 n5615 0 dm2 AREA=4.042e-07
D5615 n5616 0 dm2 AREA=6.246e-07
D5616 n5617 0 dm2 AREA=1.352e-06
D5617 n5618 0 dm2 AREA=6.086e-07
D5618 n5619 0 dm2 AREA=1.441e-06
D5619 n5620 0 dm2 AREA=9.208e-07
D5620 n5621 0 dm2 AREA=8.983e-07
D5621 n5622 0 dm2 AREA=4.745e-07
D5622 n5623 0 dm2 AREA=8.279e-07
D5623 n5624 0 dm2 AREA=9.148e-07
D5624 n5625 0 dm2 AREA=7.702e-07
D5625 n5626 0 dm2 AREA=3.516e-07
D5626 n5627 0 dm2 AREA=4.677e-07
D5627 n5628 0 dm2 AREA=1.352e-06
D5628 n5629 0 dm2 AREA=1.309e-06
D5629 n5630 0 dm2 AREA=1.005e-06
D5630 n5631 0 dm2 AREA=6.823e-07
D5631 n5632 0 dm2 AREA=2.502e-07
D5632 n5633 0 dm2 AREA=8.812e-07
D5633 n5634 0 dm2 AREA=1.249e-06
D5634 n5635 0 dm2 AREA=1.814e-06
D5635 n5636 0 dm2 AREA=9.676e-07
D5636 n5637 0 dm2 AREA=1.484e-06
D5637 n5638 0 dm2 AREA=3.627e-07
D5638 n5639 0 dm2 AREA=9.678e-07
D5639 n5640 0 dm2 AREA=6.474e-07
D5640 n5641 0 dm2 AREA=9.367e-07
D5641 n5642 0 dm2 AREA=7.925e-07
D5642 n5643 0 dm2 AREA=1.395e-06
D5643 n5644 0 dm2 AREA=1.065e-06
D5644 n5645 0 dm2 AREA=4.934e-07
D5645 n5646 0 dm2 AREA=3.291e-07
D5646 n5647 0 dm2 AREA=2.310e-07
D5647 n5648 0 dm2 AREA=4.196e-07
D5648 n5649 0 dm2 AREA=5.361e-07
D5649 n5650 0 dm2 AREA=1.717e-06
D5650 n5651 0 dm2 AREA=7.728e-07
D5651 n5652 0 dm2 AREA=5.324e-07
D5652 n5653 0 dm2 AREA=7.774e-07
D5653 n5654 0 dm2 AREA=7.579e-07
D5654 n5655 0 dm2 AREA=7.718e-07
D5655 n5656 0 dm2 AREA=5.293e-07
D5656 n5657 0 dm2 AREA=2.018e-06
D5657 n5658 0 dm2 AREA=1.589e-06
D5658 n5659 0 dm2 AREA=8.850e-07
D5659 n5660 0 dm2 AREA=1.835e-06
D5660 n5661 0 dm2 AREA=2.302e-06
D5661 n5662 0 dm2 AREA=1.110e-06
D5662 n5663 0 dm2 AREA=4.376e-07
D5663 n5664 0 dm2 AREA=9.806e-07
D5664 n5665 0 dm2 AREA=1.523e-06
D5665 n5666 0 dm2 AREA=1.196e-06
D5666 n5667 0 dm2 AREA=1.091e-06
D5667 n5668 0 dm2 AREA=6.100e-07
D5668 n5669 0 dm2 AREA=1.634e-06
D5669 n5670 0 dm2 AREA=1.471e-06
D5670 n5671 0 dm2 AREA=9.254e-07
D5671 n5672 0 dm2 AREA=5.075e-07
D5672 n5673 0 dm2 AREA=8.763e-07
D5673 n5674 0 dm2 AREA=9.733e-07
D5674 n5675 0 dm2 AREA=1.407e-06
D5675 n5676 0 dm2 AREA=9.768e-07
D5676 n5677 0 dm2 AREA=5.402e-07
D5677 n5678 0 dm2 AREA=1.343e-06
D5678 n5679 0 dm2 AREA=9.556e-07
D5679 n5680 0 dm2 AREA=6.862e-07
D5680 n5681 0 dm2 AREA=8.392e-07
D5681 n5682 0 dm2 AREA=7.882e-07
D5682 n5683 0 dm2 AREA=7.303e-07
D5683 n5684 0 dm2 AREA=2.869e-07
D5684 n5685 0 dm2 AREA=1.136e-06
D5685 n5686 0 dm2 AREA=1.802e-07
D5686 n5687 0 dm2 AREA=2.626e-06
D5687 n5688 0 dm2 AREA=4.972e-07
D5688 n5689 0 dm2 AREA=2.957e-07
D5689 n5690 0 dm2 AREA=2.744e-06
D5690 n5691 0 dm2 AREA=6.076e-07
D5691 n5692 0 dm2 AREA=7.112e-07
D5692 n5693 0 dm2 AREA=5.852e-07
D5693 n5694 0 dm2 AREA=1.536e-06
D5694 n5695 0 dm2 AREA=1.087e-06
D5695 n5696 0 dm2 AREA=7.048e-07
D5696 n5697 0 dm2 AREA=3.201e-07
D5697 n5698 0 dm2 AREA=6.198e-07
D5698 n5699 0 dm2 AREA=8.441e-07
D5699 n5700 0 dm2 AREA=1.756e-06
D5700 n5701 0 dm2 AREA=1.599e-06
D5701 n5702 0 dm2 AREA=1.222e-06
D5702 n5703 0 dm2 AREA=2.066e-06
D5703 n5704 0 dm2 AREA=6.806e-07
D5704 n5705 0 dm2 AREA=5.343e-07
D5705 n5706 0 dm2 AREA=3.088e-07
D5706 n5707 0 dm2 AREA=1.571e-06
D5707 n1 0 dm2 AREA=3.653e-07
D5708 n5709 0 dm2 AREA=4.882e-07
D5709 n5710 0 dm2 AREA=1.516e-06
D5710 n5711 0 dm2 AREA=2.485e-07
D5711 n5712 0 dm2 AREA=4.497e-07
D5712 n5713 0 dm2 AREA=1.633e-06
D5713 n5714 0 dm2 AREA=1.865e-06
D5714 n5715 0 dm2 AREA=1.613e-06
D5715 n5716 0 dm2 AREA=6.100e-07
D5716 n5717 0 dm2 AREA=9.517e-07
D5717 n5718 0 dm2 AREA=6.287e-07
D5718 n5719 0 dm2 AREA=1.092e-06
D5719 n5720 0 dm2 AREA=3.753e-07
D5720 n5721 0 dm2 AREA=9.269e-07
D5721 n5722 0 dm2 AREA=8.185e-07
D5722 n5723 0 dm2 AREA=1.600e-06
D5723 n5724 0 dm2 AREA=7.491e-08
D5724 n5725 0 dm2 AREA=8.243e-07
D5725 n5726 0 dm2 AREA=9.301e-07
D5726 n5727 0 dm2 AREA=2.606e-07
D5727 n5728 0 dm2 AREA=5.763e-07
D5728 n5729 0 dm2 AREA=1.192e-06
D5729 n5730 0 dm2 AREA=1.084e-06
D5730 n5731 0 dm2 AREA=8.984e-07
D5731 n5732 0 dm2 AREA=2.472e-07
D5732 n5733 0 dm2 AREA=8.375e-07
D5733 n5734 0 dm2 AREA=5.209e-07
D5734 n5735 0 dm2 AREA=7.979e-07
D5735 n5736 0 dm2 AREA=1.354e-06
D5736 n5737 0 dm2 AREA=1.391e-06
D5737 n5738 0 dm2 AREA=1.469e-06
D5738 n5739 0 dm2 AREA=5.304e-07
D5739 n5740 0 dm2 AREA=4.282e-07
D5740 n5741 0 dm2 AREA=1.202e-06
D5741 n5742 0 dm2 AREA=5.365e-07
D5742 n5743 0 dm2 AREA=8.106e-07
D5743 n5744 0 dm2 AREA=1.441e-06
D5744 n5745 0 dm2 AREA=4.367e-07
D5745 n5746 0 dm2 AREA=1.802e-06
D5746 n5747 0 dm2 AREA=2.020e-06
D5747 n5748 0 dm2 AREA=9.502e-07
D5748 n5749 0 dm2 AREA=1.548e-06
D5749 n5750 0 dm2 AREA=5.643e-07
D5750 n5751 0 dm2 AREA=4.087e-07
D5751 n5752 0 dm2 AREA=1.127e-06
D5752 n5753 0 dm2 AREA=5.888e-07
D5753 n5754 0 dm2 AREA=1.886e-06
D5754 n5755 0 dm2 AREA=2.997e-07
D5755 n5756 0 dm2 AREA=7.040e-07
D5756 n5757 0 dm2 AREA=1.480e-06
D5757 n5758 0 dm2 AREA=9.274e-07
D5758 n5759 0 dm2 AREA=1.091e-06
D5759 n5760 0 dm2 AREA=9.908e-07
D5760 n5761 0 dm2 AREA=7.545e-07
D5761 n5762 0 dm2 AREA=2.226e-06
D5762 n5763 0 dm2 AREA=6.223e-07
D5763 n5764 0 dm2 AREA=5.412e-07
D5764 n5765 0 dm2 AREA=1.073e-07
D5765 n5766 0 dm2 AREA=7.808e-07
D5766 n5767 0 dm2 AREA=9.668e-07
D5767 n5768 0 dm2 AREA=2.168e-07
D5768 n5769 0 dm2 AREA=3.047e-07
D5769 n5770 0 dm2 AREA=1.494e-06
D5770 n5771 0 dm2 AREA=1.696e-06
D5771 n5772 0 dm2 AREA=1.032e-06
D5772 n5773 0 dm2 AREA=6.535e-07
D5773 n5774 0 dm2 AREA=7.477e-07
D5774 n5775 0 dm2 AREA=2.059e-07
D5775 n5776 0 dm2 AREA=5.453e-07
D5776 n5777 0 dm2 AREA=3.987e-07
D5777 n5778 0 dm2 AREA=1.159e-06
D5778 n5779 0 dm2 AREA=1.162e-06
D5779 n5780 0 dm2 AREA=3.714e-07
D5780 n5781 0 dm2 AREA=4.329e-07
D5781 n5782 0 dm2 AREA=5.782e-07
D5782 n5783 0 dm2 AREA=3.619e-07
D5783 n5784 0 dm2 AREA=1.104e-06
D5784 n5785 0 dm2 AREA=9.505e-07
D5785 n5786 0 dm2 AREA=1.170e-06
D5786 n5787 0 dm2 AREA=1.532e-06
D5787 n5788 0 dm2 AREA=8.691e-07
D5788 n5789 0 dm2 AREA=1.754e-06
D5789 n5790 0 dm2 AREA=9.321e-07
D5790 n5791 0 dm2 AREA=1.749e-06
D5791 n5792 0 dm2 AREA=1.051e-06
D5792 n5793 0 dm2 AREA=6.825e-07
D5793 n5794 0 dm2 AREA=1.389e-06
D5794 n5795 0 dm2 AREA=1.418e-06
D5795 n5796 0 dm2 AREA=9.042e-07
D5796 n5797 0 dm2 AREA=1.181e-06
D5797 n5798 0 dm2 AREA=2.137e-06
D5798 n5799 0 dm2 AREA=8.245e-07
D5799 n5800 0 dm2 AREA=1.181e-06
D5800 n5801 0 dm2 AREA=5.116e-07
D5801 n5802 0 dm2 AREA=5.745e-07
D5802 n5803 0 dm2 AREA=4.088e-07
D5803 n5804 0 dm2 AREA=7.103e-07
D5804 n5805 0 dm2 AREA=1.962e-06
D5805 n5806 0 dm2 AREA=1.530e-06
D5806 n5807 0 dm2 AREA=1.520e-06
D5807 n5808 0 dm2 AREA=1.107e-06
D5808 n5809 0 dm2 AREA=1.366e-06
D5809 n5810 0 dm2 AREA=4.332e-07
D5810 n5811 0 dm2 AREA=4.474e-07
D5811 n5812 0 dm2 AREA=8.070e-07
D5812 n5813 0 dm2 AREA=3.197e-07
D5813 n5814 0 dm2 AREA=6.854e-07
D5814 n5815 0 dm2 AREA=6.664e-07
D5815 n5816 0 dm2 AREA=4.168e-07
D5816 n5817 0 dm2 AREA=1.405e-06
D5817 n5818 0 dm2 AREA=1.825e-06
D5818 n5819 0 dm2 AREA=1.978e-06
D5819 n5820 0 dm2 AREA=1.613e-06
D5820 n5821 0 dm2 AREA=1.039e-06
D5821 n5822 0 dm2 AREA=1.048e-06
D5822 n5823 0 dm2 AREA=7.762e-07
D5823 n5824 0 dm2 AREA=5.464e-07
D5824 n5825 0 dm2 AREA=2.096e-06
D5825 n5826 0 dm2 AREA=2.287e-07
D5826 n5827 0 dm2 AREA=1.415e-06
D5827 n5828 0 dm2 AREA=9.594e-07
D5828 n5829 0 dm2 AREA=8.186e-07
D5829 n5830 0 dm2 AREA=1.723e-06
D5830 n5831 0 dm2 AREA=2.427e-07
D5831 n5832 0 dm2 AREA=1.653e-06
D5832 n5833 0 dm2 AREA=1.894e-06
D5833 n5834 0 dm2 AREA=2.374e-06
D5834 n5835 0 dm2 AREA=3.895e-07
D5835 n5836 0 dm2 AREA=5.180e-07
D5836 n5837 0 dm2 AREA=9.015e-07
D5837 n5838 0 dm2 AREA=6.468e-07
D5838 n5839 0 dm2 AREA=1.327e-06
D5839 n5840 0 dm2 AREA=9.656e-07
D5840 n5841 0 dm2 AREA=5.730e-07
D5841 n5842 0 dm2 AREA=1.673e-06
D5842 n5843 0 dm2 AREA=1.038e-06
D5843 n5844 0 dm2 AREA=1.590e-06
D5844 n5845 0 dm2 AREA=1.027e-06
D5845 n5846 0 dm2 AREA=1.815e-06
D5846 n5847 0 dm2 AREA=1.006e-06
D5847 n5848 0 dm2 AREA=1.988e-06
D5848 n5849 0 dm2 AREA=9.804e-07
D5849 n5850 0 dm2 AREA=1.605e-06
D5850 n5851 0 dm2 AREA=8.210e-07
D5851 n5852 0 dm2 AREA=1.379e-06
D5852 n5853 0 dm2 AREA=1.937e-07
D5853 n5854 0 dm2 AREA=1.036e-06
D5854 n5855 0 dm2 AREA=1.080e-06
D5855 n5856 0 dm2 AREA=4.808e-07
D5856 n5857 0 dm2 AREA=9.662e-07
D5857 n5858 0 dm2 AREA=1.009e-06
D5858 n5859 0 dm2 AREA=1.559e-06
D5859 n5860 0 dm2 AREA=8.079e-08
D5860 n5861 0 dm2 AREA=8.616e-07
D5861 n5862 0 dm2 AREA=1.090e-06
D5862 n5863 0 dm2 AREA=1.590e-06
D5863 n5864 0 dm2 AREA=2.496e-06
D5864 n5865 0 dm2 AREA=1.683e-06
D5865 n5866 0 dm2 AREA=1.304e-06
D5866 n5867 0 dm2 AREA=2.170e-06
D5867 n5868 0 dm2 AREA=9.652e-07
D5868 n5869 0 dm2 AREA=7.275e-07
D5869 n5870 0 dm2 AREA=1.672e-06
D5870 n5871 0 dm2 AREA=8.758e-07
D5871 n5872 0 dm2 AREA=4.816e-07
D5872 n5873 0 dm2 AREA=4.797e-07
D5873 n5874 0 dm2 AREA=7.951e-07
D5874 n5875 0 dm2 AREA=9.659e-07
D5875 n5876 0 dm2 AREA=9.033e-07
D5876 n5877 0 dm2 AREA=7.426e-07
D5877 n5878 0 dm2 AREA=4.183e-07
D5878 n5879 0 dm2 AREA=4.619e-07
D5879 n5880 0 dm2 AREA=1.668e-06
D5880 n5881 0 dm2 AREA=9.980e-07
D5881 n5882 0 dm2 AREA=1.551e-06
D5882 n5883 0 dm2 AREA=1.524e-06
D5883 n5884 0 dm2 AREA=4.383e-07
D5884 n5885 0 dm2 AREA=7.039e-07
D5885 n5886 0 dm2 AREA=8.816e-07
D5886 n5887 0 dm2 AREA=9.779e-07
D5887 n5888 0 dm2 AREA=8.115e-07
D5888 n5889 0 dm2 AREA=6.475e-07
D5889 n5890 0 dm2 AREA=1.237e-06
D5890 n5891 0 dm2 AREA=3.868e-07
D5891 n5892 0 dm2 AREA=9.896e-07
D5892 n5893 0 dm2 AREA=1.110e-06
D5893 n5894 0 dm2 AREA=5.005e-07
D5894 n5895 0 dm2 AREA=1.536e-06
D5895 n5896 0 dm2 AREA=1.293e-06
D5896 n5897 0 dm2 AREA=1.555e-06
D5897 n5898 0 dm2 AREA=7.891e-07
D5898 n5899 0 dm2 AREA=3.538e-07
D5899 n5900 0 dm2 AREA=8.610e-07
D5900 n5901 0 dm2 AREA=9.009e-07
D5901 n5902 0 dm2 AREA=3.957e-07
D5902 n5903 0 dm2 AREA=6.258e-07
D5903 n5904 0 dm2 AREA=1.578e-06
D5904 n5905 0 dm2 AREA=7.278e-07
D5905 n5906 0 dm2 AREA=2.015e-07
D5906 n5907 0 dm2 AREA=2.207e-06
D5907 n5908 0 dm2 AREA=9.813e-07
D5908 n5909 0 dm2 AREA=7.120e-07
D5909 n1 0 dm2 AREA=1.027e-06
D5910 n5911 0 dm2 AREA=1.136e-06
D5911 n5912 0 dm2 AREA=5.802e-08
D5912 n5913 0 dm2 AREA=7.248e-07
D5913 n5914 0 dm2 AREA=1.781e-06
D5914 n5915 0 dm2 AREA=1.388e-06
D5915 n5916 0 dm2 AREA=8.736e-07
D5916 n5917 0 dm2 AREA=2.169e-06
D5917 n5918 0 dm2 AREA=8.338e-07
D5918 n5919 0 dm2 AREA=1.016e-06
D5919 n5920 0 dm2 AREA=1.279e-06
D5920 n5921 0 dm2 AREA=8.514e-07
D5921 n5922 0 dm2 AREA=1.455e-06
D5922 n5923 0 dm2 AREA=5.314e-07
D5923 n5924 0 dm2 AREA=4.059e-07
D5924 n5925 0 dm2 AREA=6.819e-07
D5925 n5926 0 dm2 AREA=9.849e-07
D5926 n5927 0 dm2 AREA=1.376e-06
D5927 n5928 0 dm2 AREA=3.215e-07
D5928 n5929 0 dm2 AREA=6.784e-07
D5929 n5930 0 dm2 AREA=2.686e-07
D5930 n5931 0 dm2 AREA=1.146e-06
D5931 n5932 0 dm2 AREA=1.684e-06
D5932 n1 0 dm2 AREA=1.412e-06
D5933 n5934 0 dm2 AREA=8.425e-07
D5934 n5935 0 dm2 AREA=1.325e-06
D5935 n5936 0 dm2 AREA=4.340e-07
D5936 n5937 0 dm2 AREA=1.190e-06
D5937 n5938 0 dm2 AREA=1.778e-06
D5938 n5939 0 dm2 AREA=4.648e-07
D5939 n5940 0 dm2 AREA=1.469e-06
D5940 n5941 0 dm2 AREA=6.708e-07
D5941 n5942 0 dm2 AREA=4.447e-07
D5942 n5943 0 dm2 AREA=7.645e-07
D5943 n5944 0 dm2 AREA=1.066e-06
D5944 n5945 0 dm2 AREA=1.030e-06
D5945 n5946 0 dm2 AREA=1.649e-06
D5946 n5947 0 dm2 AREA=7.442e-07
D5947 n5948 0 dm2 AREA=6.225e-07
D5948 n5949 0 dm2 AREA=8.243e-07
D5949 n5950 0 dm2 AREA=1.135e-06
D5950 n5951 0 dm2 AREA=1.636e-06
D5951 n5952 0 dm2 AREA=7.468e-07
D5952 n5953 0 dm2 AREA=1.659e-06
D5953 n5954 0 dm2 AREA=6.575e-07
D5954 n5955 0 dm2 AREA=8.868e-07
D5955 n5956 0 dm2 AREA=5.622e-07
D5956 n5957 0 dm2 AREA=1.438e-06
D5957 n5958 0 dm2 AREA=1.240e-06
D5958 n5959 0 dm2 AREA=1.266e-06
D5959 n5960 0 dm2 AREA=7.156e-07
D5960 n5961 0 dm2 AREA=4.957e-07
D5961 n5962 0 dm2 AREA=3.352e-06
D5962 n5963 0 dm2 AREA=1.554e-06
D5963 n5964 0 dm2 AREA=1.513e-06
D5964 n5965 0 dm2 AREA=7.027e-07
D5965 n5966 0 dm2 AREA=3.919e-07
D5966 n5967 0 dm2 AREA=1.350e-06
D5967 n5968 0 dm2 AREA=7.114e-07
D5968 n5969 0 dm2 AREA=3.768e-07
D5969 n5970 0 dm2 AREA=1.258e-06
D5970 n5971 0 dm2 AREA=9.144e-07
D5971 n5972 0 dm2 AREA=2.857e-06
D5972 n5973 0 dm2 AREA=6.271e-07
D5973 n5974 0 dm2 AREA=6.788e-07
D5974 n5975 0 dm2 AREA=8.066e-07
D5975 n5976 0 dm2 AREA=9.573e-07
D5976 n5977 0 dm2 AREA=9.825e-07
D5977 n5978 0 dm2 AREA=4.999e-07
D5978 n5979 0 dm2 AREA=5.826e-07
D5979 n5980 0 dm2 AREA=2.104e-06
D5980 n5981 0 dm2 AREA=6.339e-07
D5981 n5982 0 dm2 AREA=9.897e-07
D5982 n5983 0 dm2 AREA=1.049e-06
D5983 n5984 0 dm2 AREA=7.634e-07
D5984 n5985 0 dm2 AREA=1.385e-06
D5985 n5986 0 dm2 AREA=5.255e-07
D5986 n5987 0 dm2 AREA=1.235e-06
D5987 n5988 0 dm2 AREA=4.323e-07
D5988 n5989 0 dm2 AREA=6.926e-07
D5989 n5990 0 dm2 AREA=6.565e-07
D5990 n5991 0 dm2 AREA=9.406e-07
D5991 n5992 0 dm2 AREA=2.549e-07
D5992 n5993 0 dm2 AREA=2.837e-07
D5993 n5994 0 dm2 AREA=9.192e-07
D5994 n5995 0 dm2 AREA=1.246e-06
D5995 n5996 0 dm2 AREA=5.610e-07
D5996 n5997 0 dm2 AREA=1.129e-06
D5997 n5998 0 dm2 AREA=5.633e-07
D5998 n5999 0 dm2 AREA=5.025e-07
D5999 n6000 0 dm2 AREA=1.026e-06
D6000 n6001 0 dm2 AREA=1.889e-06
D6001 n6002 0 dm2 AREA=1.249e-06
D6002 n6003 0 dm2 AREA=6.767e-07
D6003 n6004 0 dm2 AREA=1.042e-06
D6004 n6005 0 dm2 AREA=5.617e-07
D6005 n6006 0 dm2 AREA=8.100e-07
D6006 n6007 0 dm2 AREA=1.126e-06
D6007 n6008 0 dm2 AREA=6.967e-07
D6008 n6009 0 dm2 AREA=1.172e-07
D6009 n6010 0 dm2 AREA=1.187e-06
D6010 n6011 0 dm2 AREA=5.798e-07
D6011 n6012 0 dm2 AREA=8.565e-07
D6012 n6013 0 dm2 AREA=1.379e-06
D6013 n6014 0 dm2 AREA=1.316e-06
D6014 n6015 0 dm2 AREA=1.868e-06
D6015 n6016 0 dm2 AREA=6.620e-07
D6016 n6017 0 dm2 AREA=2.196e-07
D6017 n6018 0 dm2 AREA=1.411e-06
D6018 n6019 0 dm2 AREA=1.418e-06
D6019 n6020 0 dm2 AREA=9.521e-07
D6020 n6021 0 dm2 AREA=6.190e-07
D6021 n6022 0 dm2 AREA=3.840e-07
D6022 n6023 0 dm2 AREA=2.041e-06
D6023 n6024 0 dm2 AREA=9.165e-07
D6024 n6025 0 dm2 AREA=8.202e-07
D6025 n6026 0 dm2 AREA=1.388e-07
D6026 n6027 0 dm2 AREA=8.540e-07
D6027 n6028 0 dm2 AREA=1.570e-06
D6028 n6029 0 dm2 AREA=9.443e-07
D6029 n6030 0 dm2 AREA=1.631e-06
D6030 n6031 0 dm2 AREA=3.222e-07
D6031 n6032 0 dm2 AREA=2.519e-06
D6032 n6033 0 dm2 AREA=4.803e-07
D6033 n6034 0 dm2 AREA=1.230e-06
D6034 n6035 0 dm2 AREA=4.788e-07
D6035 n6036 0 dm2 AREA=4.684e-07
D6036 n6037 0 dm2 AREA=7.227e-07
D6037 n6038 0 dm2 AREA=4.136e-07
D6038 n6039 0 dm2 AREA=1.142e-06
D6039 n6040 0 dm2 AREA=1.114e-06
D6040 n6041 0 dm2 AREA=2.065e-06
D6041 n1 0 dm2 AREA=8.357e-07
D6042 n6043 0 dm2 AREA=1.373e-06
D6043 n6044 0 dm2 AREA=3.447e-07
D6044 n6045 0 dm2 AREA=1.635e-06
D6045 n6046 0 dm2 AREA=2.996e-06
D6046 n6047 0 dm2 AREA=1.065e-06
D6047 n6048 0 dm2 AREA=6.173e-07
D6048 n6049 0 dm2 AREA=1.036e-06
D6049 n6050 0 dm2 AREA=2.196e-06
D6050 n6051 0 dm2 AREA=9.337e-07
D6051 n6052 0 dm2 AREA=6.564e-07
D6052 n6053 0 dm2 AREA=5.446e-07
D6053 n6054 0 dm2 AREA=2.421e-06
D6054 n6055 0 dm2 AREA=7.790e-07
D6055 n6056 0 dm2 AREA=3.390e-06
D6056 n6057 0 dm2 AREA=1.084e-06
D6057 n6058 0 dm2 AREA=1.258e-06
D6058 n6059 0 dm2 AREA=7.069e-07
D6059 n6060 0 dm2 AREA=8.453e-07
D6060 n6061 0 dm2 AREA=9.155e-07
D6061 n6062 0 dm2 AREA=1.425e-06
D6062 n6063 0 dm2 AREA=1.001e-06
D6063 n6064 0 dm2 AREA=1.081e-06
D6064 n6065 0 dm2 AREA=9.849e-07
D6065 n6066 0 dm2 AREA=8.879e-07
D6066 n6067 0 dm2 AREA=1.224e-06
D6067 n6068 0 dm2 AREA=6.146e-07
D6068 n6069 0 dm2 AREA=4.282e-07
D6069 n6070 0 dm2 AREA=5.767e-07
D6070 n6071 0 dm2 AREA=5.539e-07
D6071 n6072 0 dm2 AREA=3.303e-07
D6072 n6073 0 dm2 AREA=2.834e-07
D6073 n6074 0 dm2 AREA=8.939e-07
D6074 n6075 0 dm2 AREA=6.740e-07
D6075 n6076 0 dm2 AREA=1.740e-06
D6076 n6077 0 dm2 AREA=5.105e-07
D6077 n6078 0 dm2 AREA=1.300e-06
D6078 n6079 0 dm2 AREA=9.511e-07
D6079 n6080 0 dm2 AREA=8.584e-07
D6080 n6081 0 dm2 AREA=7.585e-07
D6081 n6082 0 dm2 AREA=1.507e-06
D6082 n6083 0 dm2 AREA=3.761e-07
D6083 n6084 0 dm2 AREA=4.884e-07
D6084 n6085 0 dm2 AREA=3.524e-07
D6085 n6086 0 dm2 AREA=6.899e-07
D6086 n6087 0 dm2 AREA=1.593e-07
D6087 n6088 0 dm2 AREA=1.010e-06
D6088 n6089 0 dm2 AREA=8.431e-07
D6089 n6090 0 dm2 AREA=7.542e-07
D6090 n6091 0 dm2 AREA=1.059e-06
D6091 n6092 0 dm2 AREA=9.565e-07
D6092 n6093 0 dm2 AREA=1.870e-06
D6093 n6094 0 dm2 AREA=5.695e-07
D6094 n6095 0 dm2 AREA=8.721e-07
D6095 n6096 0 dm2 AREA=1.934e-06
D6096 n6097 0 dm2 AREA=9.766e-07
D6097 n6098 0 dm2 AREA=9.305e-07
D6098 n6099 0 dm2 AREA=1.063e-06
D6099 n6100 0 dm2 AREA=6.594e-07
D6100 n6101 0 dm2 AREA=8.897e-07
D6101 n6102 0 dm2 AREA=3.187e-07
D6102 n6103 0 dm2 AREA=1.136e-06
D6103 n6104 0 dm2 AREA=1.429e-06
D6104 n6105 0 dm2 AREA=8.522e-07
D6105 n6106 0 dm2 AREA=4.150e-07
D6106 n6107 0 dm2 AREA=4.474e-07
D6107 n6108 0 dm2 AREA=4.624e-07
D6108 n6109 0 dm2 AREA=1.302e-06
D6109 n6110 0 dm2 AREA=8.057e-07
D6110 n6111 0 dm2 AREA=1.223e-07
D6111 n6112 0 dm2 AREA=1.637e-06
D6112 n6113 0 dm2 AREA=1.714e-06
D6113 n6114 0 dm2 AREA=7.786e-07
D6114 n6115 0 dm2 AREA=7.114e-07
D6115 n6116 0 dm2 AREA=2.549e-07
D6116 n6117 0 dm2 AREA=1.735e-06
D6117 n6118 0 dm2 AREA=5.700e-07
D6118 n6119 0 dm2 AREA=8.047e-07
D6119 n1 0 dm2 AREA=1.593e-06
D6120 n6121 0 dm2 AREA=7.764e-07
D6121 n6122 0 dm2 AREA=8.460e-07
D6122 n6123 0 dm2 AREA=8.480e-07
D6123 n6124 0 dm2 AREA=1.723e-06
D6124 n6125 0 dm2 AREA=2.619e-07
D6125 n6126 0 dm2 AREA=5.305e-07
D6126 n6127 0 dm2 AREA=1.785e-06
D6127 n6128 0 dm2 AREA=1.733e-06
D6128 n6129 0 dm2 AREA=1.160e-06
D6129 n6130 0 dm2 AREA=9.293e-07
D6130 n6131 0 dm2 AREA=1.993e-06
D6131 n6132 0 dm2 AREA=1.290e-06
D6132 n6133 0 dm2 AREA=3.094e-06
D6133 n6134 0 dm2 AREA=1.524e-06
D6134 n6135 0 dm2 AREA=1.491e-06
D6135 n6136 0 dm2 AREA=9.753e-07
D6136 n6137 0 dm2 AREA=1.288e-06
D6137 n6138 0 dm2 AREA=1.510e-06
D6138 n6139 0 dm2 AREA=1.088e-06
D6139 n6140 0 dm2 AREA=5.954e-07
D6140 n6141 0 dm2 AREA=6.073e-07
D6141 n6142 0 dm2 AREA=9.430e-07
D6142 n6143 0 dm2 AREA=1.319e-06
D6143 n6144 0 dm2 AREA=2.496e-07
D6144 n6145 0 dm2 AREA=2.484e-07
D6145 n6146 0 dm2 AREA=8.105e-07
D6146 n6147 0 dm2 AREA=1.172e-06
D6147 n6148 0 dm2 AREA=1.108e-06
D6148 n6149 0 dm2 AREA=6.767e-07
D6149 n6150 0 dm2 AREA=4.744e-07
D6150 n6151 0 dm2 AREA=8.493e-07
D6151 n6152 0 dm2 AREA=7.010e-07
D6152 n6153 0 dm2 AREA=3.023e-07
D6153 n6154 0 dm2 AREA=1.622e-06
D6154 n6155 0 dm2 AREA=2.300e-06
D6155 n6156 0 dm2 AREA=7.398e-07
D6156 n6157 0 dm2 AREA=9.660e-07
D6157 n6158 0 dm2 AREA=1.347e-06
D6158 n6159 0 dm2 AREA=1.372e-06
D6159 n6160 0 dm2 AREA=8.318e-07
D6160 n6161 0 dm2 AREA=1.561e-06
D6161 n6162 0 dm2 AREA=1.505e-06
D6162 n6163 0 dm2 AREA=4.520e-07
D6163 n6164 0 dm2 AREA=7.555e-07
D6164 n6165 0 dm2 AREA=6.706e-07
D6165 n6166 0 dm2 AREA=1.544e-06
D6166 n6167 0 dm2 AREA=7.001e-07
D6167 n6168 0 dm2 AREA=9.994e-07
D6168 n6169 0 dm2 AREA=1.313e-06
D6169 n6170 0 dm2 AREA=7.440e-07
D6170 n6171 0 dm2 AREA=8.998e-07
D6171 n6172 0 dm2 AREA=1.667e-06
D6172 n6173 0 dm2 AREA=1.813e-06
D6173 n6174 0 dm2 AREA=6.986e-07
D6174 n1 0 dm2 AREA=6.605e-07
D6175 n6176 0 dm2 AREA=5.889e-07
D6176 n6177 0 dm2 AREA=6.479e-07
D6177 n6178 0 dm2 AREA=9.661e-07
D6178 n6179 0 dm2 AREA=1.413e-06
D6179 n6180 0 dm2 AREA=6.165e-07
D6180 n6181 0 dm2 AREA=4.764e-07
D6181 n6182 0 dm2 AREA=7.710e-07
D6182 n6183 0 dm2 AREA=6.853e-07
D6183 n6184 0 dm2 AREA=6.425e-07
D6184 n6185 0 dm2 AREA=1.322e-06
D6185 n6186 0 dm2 AREA=1.497e-06
D6186 n6187 0 dm2 AREA=1.239e-06
D6187 n6188 0 dm2 AREA=9.959e-07
D6188 n6189 0 dm2 AREA=1.967e-06
D6189 n6190 0 dm2 AREA=1.549e-07
D6190 n6191 0 dm2 AREA=6.373e-07
D6191 n6192 0 dm2 AREA=2.731e-07
D6192 n6193 0 dm2 AREA=1.261e-06
D6193 n6194 0 dm2 AREA=1.641e-06
D6194 n6195 0 dm2 AREA=2.120e-07
D6195 n6196 0 dm2 AREA=3.348e-07
D6196 n6197 0 dm2 AREA=4.663e-07
D6197 n6198 0 dm2 AREA=1.368e-06
D6198 n6199 0 dm2 AREA=1.099e-06
D6199 n6200 0 dm2 AREA=6.262e-07
D6200 n6201 0 dm2 AREA=9.603e-07
D6201 n6202 0 dm2 AREA=7.031e-07
D6202 n6203 0 dm2 AREA=6.485e-07
D6203 n6204 0 dm2 AREA=7.716e-07
D6204 n6205 0 dm2 AREA=1.424e-06
D6205 n6206 0 dm2 AREA=5.646e-07
D6206 n6207 0 dm2 AREA=1.587e-06
D6207 n6208 0 dm2 AREA=1.205e-06
D6208 n6209 0 dm2 AREA=1.291e-06
D6209 n6210 0 dm2 AREA=4.979e-07
D6210 n6211 0 dm2 AREA=1.328e-06
D6211 n6212 0 dm2 AREA=1.404e-07
D6212 n6213 0 dm2 AREA=8.239e-07
D6213 n6214 0 dm2 AREA=1.014e-06
D6214 n6215 0 dm2 AREA=6.344e-08
D6215 n6216 0 dm2 AREA=2.822e-07
D6216 n6217 0 dm2 AREA=1.748e-06
D6217 n6218 0 dm2 AREA=2.595e-07
D6218 n6219 0 dm2 AREA=1.665e-06
D6219 n6220 0 dm2 AREA=8.980e-07
D6220 n6221 0 dm2 AREA=1.583e-06
D6221 n6222 0 dm2 AREA=4.543e-07
D6222 n6223 0 dm2 AREA=8.112e-07
D6223 n6224 0 dm2 AREA=1.561e-06
D6224 n6225 0 dm2 AREA=1.577e-06
D6225 n6226 0 dm2 AREA=1.181e-06
D6226 n6227 0 dm2 AREA=1.170e-06
D6227 n6228 0 dm2 AREA=1.299e-06
D6228 n6229 0 dm2 AREA=5.158e-07
D6229 n6230 0 dm2 AREA=1.768e-06
D6230 n6231 0 dm2 AREA=4.372e-07
D6231 n6232 0 dm2 AREA=2.532e-07
D6232 n6233 0 dm2 AREA=1.042e-06
D6233 n6234 0 dm2 AREA=1.838e-06
D6234 n6235 0 dm2 AREA=1.381e-06
D6235 n6236 0 dm2 AREA=4.102e-07
D6236 n6237 0 dm2 AREA=6.637e-07
D6237 n6238 0 dm2 AREA=1.692e-06
D6238 n6239 0 dm2 AREA=1.408e-06
D6239 n6240 0 dm2 AREA=6.966e-07
D6240 n6241 0 dm2 AREA=1.802e-06
D6241 n6242 0 dm2 AREA=1.082e-06
D6242 n6243 0 dm2 AREA=1.553e-06
D6243 n6244 0 dm2 AREA=1.064e-06
D6244 n6245 0 dm2 AREA=1.128e-06
D6245 n6246 0 dm2 AREA=1.169e-06
D6246 n6247 0 dm2 AREA=1.388e-06
D6247 n6248 0 dm2 AREA=1.154e-06
D6248 n6249 0 dm2 AREA=8.186e-07
D6249 n6250 0 dm2 AREA=8.047e-07
D6250 n6251 0 dm2 AREA=1.177e-06
D6251 n6252 0 dm2 AREA=2.321e-06
D6252 n6253 0 dm2 AREA=2.161e-06
D6253 n6254 0 dm2 AREA=1.361e-06
D6254 n6255 0 dm2 AREA=1.595e-06
D6255 n6256 0 dm2 AREA=1.536e-06
D6256 n6257 0 dm2 AREA=5.306e-07
D6257 n6258 0 dm2 AREA=9.960e-07
D6258 n6259 0 dm2 AREA=1.342e-06
D6259 n6260 0 dm2 AREA=1.720e-06
D6260 n6261 0 dm2 AREA=8.745e-07
D6261 n6262 0 dm2 AREA=6.743e-07
D6262 n6263 0 dm2 AREA=1.887e-06
D6263 n6264 0 dm2 AREA=1.165e-06
D6264 n6265 0 dm2 AREA=6.028e-07
D6265 n6266 0 dm2 AREA=8.434e-07
D6266 n6267 0 dm2 AREA=1.225e-06
D6267 n6268 0 dm2 AREA=1.150e-06
D6268 n6269 0 dm2 AREA=4.561e-07
D6269 n6270 0 dm2 AREA=7.159e-07
D6270 n6271 0 dm2 AREA=9.907e-07
D6271 n6272 0 dm2 AREA=1.057e-06
D6272 n6273 0 dm2 AREA=1.247e-06
D6273 n6274 0 dm2 AREA=1.319e-06
D6274 n6275 0 dm2 AREA=5.935e-07
D6275 n6276 0 dm2 AREA=8.640e-07
D6276 n6277 0 dm2 AREA=1.415e-06
D6277 n6278 0 dm2 AREA=1.595e-07
D6278 n6279 0 dm2 AREA=8.679e-07
D6279 n6280 0 dm2 AREA=8.710e-07
D6280 n6281 0 dm2 AREA=1.268e-06
D6281 n6282 0 dm2 AREA=5.187e-07
D6282 n6283 0 dm2 AREA=6.978e-07
D6283 n6284 0 dm2 AREA=2.658e-07
D6284 n6285 0 dm2 AREA=1.202e-06
D6285 n6286 0 dm2 AREA=8.817e-07
D6286 n6287 0 dm2 AREA=1.033e-06
D6287 n6288 0 dm2 AREA=6.443e-07
D6288 n6289 0 dm2 AREA=1.495e-06
D6289 n6290 0 dm2 AREA=1.090e-06
D6290 n6291 0 dm2 AREA=3.304e-07
D6291 n6292 0 dm2 AREA=2.475e-06
D6292 n6293 0 dm2 AREA=9.661e-07
D6293 n6294 0 dm2 AREA=1.310e-06
D6294 n6295 0 dm2 AREA=1.608e-06
D6295 n6296 0 dm2 AREA=4.479e-07
D6296 n6297 0 dm2 AREA=8.873e-07
D6297 n6298 0 dm2 AREA=1.355e-06
D6298 n6299 0 dm2 AREA=1.626e-06
D6299 n6300 0 dm2 AREA=7.928e-07
D6300 n6301 0 dm2 AREA=5.500e-07
D6301 n6302 0 dm2 AREA=6.839e-07
D6302 n6303 0 dm2 AREA=1.515e-06
D6303 n6304 0 dm2 AREA=2.581e-06
D6304 n6305 0 dm2 AREA=3.297e-07
D6305 n6306 0 dm2 AREA=8.101e-07
D6306 n6307 0 dm2 AREA=1.722e-06
D6307 n6308 0 dm2 AREA=9.768e-07
D6308 n6309 0 dm2 AREA=4.683e-07
D6309 n6310 0 dm2 AREA=1.379e-06
D6310 n6311 0 dm2 AREA=1.545e-07
D6311 n6312 0 dm2 AREA=9.597e-07
D6312 n6313 0 dm2 AREA=2.889e-07
D6313 n6314 0 dm2 AREA=1.479e-06
D6314 n6315 0 dm2 AREA=1.266e-06
D6315 n6316 0 dm2 AREA=1.122e-06
D6316 n6317 0 dm2 AREA=9.791e-07
D6317 n6318 0 dm2 AREA=1.115e-06
D6318 n6319 0 dm2 AREA=1.448e-06
D6319 n6320 0 dm2 AREA=9.281e-07
D6320 n6321 0 dm2 AREA=1.212e-06
D6321 n6322 0 dm2 AREA=1.793e-06
D6322 n6323 0 dm2 AREA=1.809e-06
D6323 n6324 0 dm2 AREA=6.341e-07
D6324 n6325 0 dm2 AREA=1.094e-06
D6325 n6326 0 dm2 AREA=1.128e-06
D6326 n6327 0 dm2 AREA=8.110e-07
D6327 n6328 0 dm2 AREA=8.565e-07
D6328 n6329 0 dm2 AREA=1.816e-06
D6329 n6330 0 dm2 AREA=1.558e-06
D6330 n6331 0 dm2 AREA=9.532e-07
D6331 n6332 0 dm2 AREA=5.541e-07
D6332 n6333 0 dm2 AREA=9.980e-07
D6333 n6334 0 dm2 AREA=2.334e-07
D6334 n6335 0 dm2 AREA=1.111e-06
D6335 n6336 0 dm2 AREA=1.168e-06
D6336 n6337 0 dm2 AREA=7.384e-07
D6337 n6338 0 dm2 AREA=3.182e-07
D6338 n6339 0 dm2 AREA=1.190e-06
D6339 n6340 0 dm2 AREA=7.563e-07
D6340 n6341 0 dm2 AREA=2.392e-06
D6341 n6342 0 dm2 AREA=1.482e-06
D6342 n1 0 dm2 AREA=1.145e-06
D6343 n6344 0 dm2 AREA=9.208e-07
D6344 n6345 0 dm2 AREA=6.689e-07
D6345 n6346 0 dm2 AREA=5.136e-07
D6346 n6347 0 dm2 AREA=2.520e-06
D6347 n6348 0 dm2 AREA=7.361e-07
D6348 n6349 0 dm2 AREA=1.121e-06
D6349 n6350 0 dm2 AREA=1.058e-06
D6350 n6351 0 dm2 AREA=9.083e-07
D6351 n6352 0 dm2 AREA=9.816e-07
D6352 n6353 0 dm2 AREA=1.221e-06
D6353 n6354 0 dm2 AREA=4.309e-07
D6354 n6355 0 dm2 AREA=4.629e-07
D6355 n6356 0 dm2 AREA=1.481e-06
D6356 n6357 0 dm2 AREA=2.264e-06
D6357 n6358 0 dm2 AREA=1.075e-06
D6358 n6359 0 dm2 AREA=6.103e-07
D6359 n6360 0 dm2 AREA=1.155e-06
D6360 n6361 0 dm2 AREA=1.139e-06
D6361 n6362 0 dm2 AREA=1.133e-06
D6362 n6363 0 dm2 AREA=1.509e-06
D6363 n6364 0 dm2 AREA=1.010e-06
D6364 n6365 0 dm2 AREA=8.119e-07
D6365 n6366 0 dm2 AREA=4.466e-07
D6366 n6367 0 dm2 AREA=7.454e-07
D6367 n6368 0 dm2 AREA=1.536e-06
D6368 n6369 0 dm2 AREA=1.667e-06
D6369 n6370 0 dm2 AREA=2.094e-06
D6370 n6371 0 dm2 AREA=1.110e-06
D6371 n6372 0 dm2 AREA=1.012e-06
D6372 n6373 0 dm2 AREA=1.167e-06
D6373 n6374 0 dm2 AREA=9.281e-07
D6374 n6375 0 dm2 AREA=1.079e-06
D6375 n6376 0 dm2 AREA=8.413e-07
D6376 n6377 0 dm2 AREA=1.485e-06
D6377 n6378 0 dm2 AREA=2.556e-07
D6378 n6379 0 dm2 AREA=3.278e-07
D6379 n6380 0 dm2 AREA=2.121e-06
D6380 n6381 0 dm2 AREA=1.135e-06
D6381 n6382 0 dm2 AREA=9.497e-07
D6382 n6383 0 dm2 AREA=6.847e-07
D6383 n6384 0 dm2 AREA=5.834e-07
D6384 n6385 0 dm2 AREA=8.812e-07
D6385 n6386 0 dm2 AREA=6.801e-07
D6386 n6387 0 dm2 AREA=8.076e-07
D6387 n6388 0 dm2 AREA=1.256e-06
D6388 n6389 0 dm2 AREA=1.872e-06
D6389 n6390 0 dm2 AREA=8.114e-07
D6390 n6391 0 dm2 AREA=7.371e-07
D6391 n6392 0 dm2 AREA=8.133e-07
D6392 n6393 0 dm2 AREA=3.980e-07
D6393 n6394 0 dm2 AREA=7.114e-07
D6394 n6395 0 dm2 AREA=8.750e-07
D6395 n6396 0 dm2 AREA=1.263e-06
D6396 n6397 0 dm2 AREA=1.317e-06
D6397 n6398 0 dm2 AREA=1.237e-06
D6398 n6399 0 dm2 AREA=5.676e-07
D6399 n6400 0 dm2 AREA=5.533e-07
D6400 n6401 0 dm2 AREA=4.578e-07
D6401 n6402 0 dm2 AREA=6.405e-07
D6402 n6403 0 dm2 AREA=1.461e-06
D6403 n6404 0 dm2 AREA=2.800e-07
D6404 n6405 0 dm2 AREA=1.059e-06
D6405 n6406 0 dm2 AREA=1.987e-06
D6406 n6407 0 dm2 AREA=1.999e-06
D6407 n6408 0 dm2 AREA=2.123e-06
D6408 n6409 0 dm2 AREA=1.184e-06
D6409 n6410 0 dm2 AREA=9.703e-07
D6410 n6411 0 dm2 AREA=9.881e-07
D6411 n6412 0 dm2 AREA=7.483e-07
D6412 n6413 0 dm2 AREA=5.563e-07
D6413 n6414 0 dm2 AREA=1.327e-06
D6414 n6415 0 dm2 AREA=2.124e-07
D6415 n6416 0 dm2 AREA=4.599e-07
D6416 n6417 0 dm2 AREA=3.359e-07
D6417 n6418 0 dm2 AREA=1.189e-06
D6418 n6419 0 dm2 AREA=8.087e-07
D6419 n6420 0 dm2 AREA=6.376e-07
D6420 n6421 0 dm2 AREA=3.815e-07
D6421 n6422 0 dm2 AREA=1.080e-06
D6422 n6423 0 dm2 AREA=5.153e-07
D6423 n6424 0 dm2 AREA=9.426e-07
D6424 n6425 0 dm2 AREA=4.241e-07
D6425 n6426 0 dm2 AREA=2.259e-07
D6426 n6427 0 dm2 AREA=1.924e-06
D6427 n6428 0 dm2 AREA=1.140e-06
D6428 n6429 0 dm2 AREA=1.666e-06
D6429 n6430 0 dm2 AREA=9.277e-07
D6430 n6431 0 dm2 AREA=1.106e-06
D6431 n6432 0 dm2 AREA=6.130e-07
D6432 n6433 0 dm2 AREA=8.986e-07
D6433 n6434 0 dm2 AREA=1.146e-06
D6434 n6435 0 dm2 AREA=1.061e-06
D6435 n6436 0 dm2 AREA=1.356e-07
D6436 n6437 0 dm2 AREA=1.674e-06
D6437 n6438 0 dm2 AREA=7.925e-07
D6438 n6439 0 dm2 AREA=6.762e-07
D6439 n6440 0 dm2 AREA=5.100e-07
D6440 n6441 0 dm2 AREA=6.300e-07
D6441 n6442 0 dm2 AREA=1.332e-06
D6442 n6443 0 dm2 AREA=2.293e-06
D6443 n6444 0 dm2 AREA=7.740e-07
D6444 n6445 0 dm2 AREA=9.385e-07
D6445 n6446 0 dm2 AREA=7.981e-07
D6446 n6447 0 dm2 AREA=6.534e-07
D6447 n6448 0 dm2 AREA=1.156e-06
D6448 n6449 0 dm2 AREA=8.883e-07
D6449 n6450 0 dm2 AREA=2.438e-06
D6450 n6451 0 dm2 AREA=1.242e-06
D6451 n6452 0 dm2 AREA=7.908e-07
D6452 n6453 0 dm2 AREA=1.806e-06
D6453 n6454 0 dm2 AREA=4.154e-07
D6454 n6455 0 dm2 AREA=1.064e-06
D6455 n6456 0 dm2 AREA=1.200e-06
D6456 n6457 0 dm2 AREA=8.263e-07
D6457 n6458 0 dm2 AREA=4.122e-07
D6458 n6459 0 dm2 AREA=1.861e-06
D6459 n6460 0 dm2 AREA=3.327e-07
D6460 n6461 0 dm2 AREA=1.120e-06
D6461 n6462 0 dm2 AREA=2.261e-07
D6462 n6463 0 dm2 AREA=1.999e-06
D6463 n6464 0 dm2 AREA=4.307e-07
D6464 n6465 0 dm2 AREA=2.762e-06
D6465 n6466 0 dm2 AREA=7.413e-07
D6466 n6467 0 dm2 AREA=9.771e-07
D6467 n6468 0 dm2 AREA=1.227e-06
D6468 n6469 0 dm2 AREA=8.842e-07
D6469 n1 0 dm2 AREA=2.747e-07
D6470 n6471 0 dm2 AREA=1.024e-06
D6471 n6472 0 dm2 AREA=5.212e-07
D6472 n6473 0 dm2 AREA=6.349e-07
D6473 n6474 0 dm2 AREA=6.778e-07
D6474 n6475 0 dm2 AREA=1.037e-06
D6475 n6476 0 dm2 AREA=7.276e-07
D6476 n6477 0 dm2 AREA=1.093e-06
D6477 n6478 0 dm2 AREA=8.051e-07
D6478 n6479 0 dm2 AREA=6.204e-07
D6479 n6480 0 dm2 AREA=1.091e-06
D6480 n6481 0 dm2 AREA=1.048e-06
D6481 n6482 0 dm2 AREA=1.069e-06
D6482 n6483 0 dm2 AREA=6.810e-07
D6483 n6484 0 dm2 AREA=1.056e-06
D6484 n6485 0 dm2 AREA=1.640e-06
D6485 n6486 0 dm2 AREA=1.016e-06
D6486 n6487 0 dm2 AREA=1.003e-06
D6487 n6488 0 dm2 AREA=5.766e-07
D6488 n6489 0 dm2 AREA=1.590e-06
D6489 n6490 0 dm2 AREA=1.674e-06
D6490 n6491 0 dm2 AREA=1.010e-06
D6491 n6492 0 dm2 AREA=8.331e-07
D6492 n6493 0 dm2 AREA=1.652e-06
D6493 n6494 0 dm2 AREA=8.447e-07
D6494 n6495 0 dm2 AREA=1.957e-06
D6495 n6496 0 dm2 AREA=5.733e-07
D6496 n6497 0 dm2 AREA=8.672e-07
D6497 n6498 0 dm2 AREA=8.244e-07
D6498 n6499 0 dm2 AREA=2.311e-07
D6499 n6500 0 dm2 AREA=2.042e-06
D6500 n6501 0 dm2 AREA=7.595e-07
D6501 n6502 0 dm2 AREA=4.144e-07
D6502 n6503 0 dm2 AREA=6.993e-07
D6503 n6504 0 dm2 AREA=1.634e-06
D6504 n6505 0 dm2 AREA=6.438e-07
D6505 n6506 0 dm2 AREA=5.892e-07
D6506 n6507 0 dm2 AREA=1.091e-06
D6507 n6508 0 dm2 AREA=8.508e-07
D6508 n6509 0 dm2 AREA=9.457e-07
D6509 n6510 0 dm2 AREA=1.879e-06
D6510 n6511 0 dm2 AREA=1.312e-06
D6511 n6512 0 dm2 AREA=5.262e-07
D6512 n6513 0 dm2 AREA=1.528e-06
D6513 n6514 0 dm2 AREA=1.136e-06
D6514 n6515 0 dm2 AREA=1.012e-06
D6515 n6516 0 dm2 AREA=1.378e-06
D6516 n6517 0 dm2 AREA=8.884e-07
D6517 n6518 0 dm2 AREA=5.982e-07
D6518 n6519 0 dm2 AREA=1.064e-06
D6519 n6520 0 dm2 AREA=5.608e-07
D6520 n6521 0 dm2 AREA=7.260e-07
D6521 n6522 0 dm2 AREA=1.008e-06
D6522 n6523 0 dm2 AREA=1.735e-06
D6523 n6524 0 dm2 AREA=1.548e-06
D6524 n6525 0 dm2 AREA=1.206e-06
D6525 n6526 0 dm2 AREA=2.079e-06
D6526 n6527 0 dm2 AREA=7.247e-07
D6527 n6528 0 dm2 AREA=1.478e-06
D6528 n6529 0 dm2 AREA=8.107e-07
D6529 n6530 0 dm2 AREA=1.993e-06
D6530 n6531 0 dm2 AREA=1.922e-06
D6531 n6532 0 dm2 AREA=4.763e-07
D6532 n6533 0 dm2 AREA=4.632e-07
D6533 n6534 0 dm2 AREA=9.854e-07
D6534 n6535 0 dm2 AREA=8.199e-07
D6535 n6536 0 dm2 AREA=1.049e-06
D6536 n6537 0 dm2 AREA=1.509e-06
D6537 n6538 0 dm2 AREA=9.350e-07
D6538 n6539 0 dm2 AREA=7.016e-07
D6539 n6540 0 dm2 AREA=1.952e-06
D6540 n6541 0 dm2 AREA=7.957e-07
D6541 n6542 0 dm2 AREA=5.938e-07
D6542 n6543 0 dm2 AREA=8.415e-07
D6543 n6544 0 dm2 AREA=2.354e-06
D6544 n6545 0 dm2 AREA=5.064e-07
D6545 n6546 0 dm2 AREA=2.355e-07
D6546 n6547 0 dm2 AREA=4.938e-07
D6547 n6548 0 dm2 AREA=9.645e-07
D6548 n6549 0 dm2 AREA=6.352e-07
D6549 n6550 0 dm2 AREA=3.310e-07
D6550 n6551 0 dm2 AREA=3.600e-07
D6551 n6552 0 dm2 AREA=1.338e-06
D6552 n6553 0 dm2 AREA=1.315e-06
D6553 n6554 0 dm2 AREA=2.537e-07
D6554 n6555 0 dm2 AREA=9.237e-07
D6555 n6556 0 dm2 AREA=5.346e-07
D6556 n6557 0 dm2 AREA=3.800e-07
D6557 n6558 0 dm2 AREA=4.212e-07
D6558 n6559 0 dm2 AREA=1.640e-06
D6559 n6560 0 dm2 AREA=5.836e-07
D6560 n6561 0 dm2 AREA=3.608e-07
D6561 n6562 0 dm2 AREA=6.380e-07
D6562 n6563 0 dm2 AREA=7.754e-07
D6563 n6564 0 dm2 AREA=1.438e-06
D6564 n6565 0 dm2 AREA=9.009e-07
D6565 n6566 0 dm2 AREA=5.848e-07
D6566 n6567 0 dm2 AREA=1.382e-06
D6567 n6568 0 dm2 AREA=1.364e-06
D6568 n6569 0 dm2 AREA=1.527e-06
D6569 n6570 0 dm2 AREA=1.320e-06
D6570 n6571 0 dm2 AREA=8.526e-07
D6571 n6572 0 dm2 AREA=6.696e-07
D6572 n6573 0 dm2 AREA=1.099e-06
D6573 n6574 0 dm2 AREA=3.481e-07
D6574 n6575 0 dm2 AREA=1.292e-06
D6575 n6576 0 dm2 AREA=1.105e-06
D6576 n6577 0 dm2 AREA=1.010e-06
D6577 n6578 0 dm2 AREA=4.838e-07
D6578 n6579 0 dm2 AREA=1.665e-06
D6579 n6580 0 dm2 AREA=8.200e-07
D6580 n6581 0 dm2 AREA=2.524e-07
D6581 n6582 0 dm2 AREA=5.716e-07
D6582 n6583 0 dm2 AREA=5.987e-07
D6583 n6584 0 dm2 AREA=4.369e-07
D6584 n6585 0 dm2 AREA=1.191e-06
D6585 n6586 0 dm2 AREA=5.611e-07
D6586 n6587 0 dm2 AREA=2.965e-07
D6587 n6588 0 dm2 AREA=1.717e-06
D6588 n6589 0 dm2 AREA=1.250e-06
D6589 n6590 0 dm2 AREA=4.345e-07
D6590 n6591 0 dm2 AREA=4.866e-07
D6591 n6592 0 dm2 AREA=1.360e-06
D6592 n6593 0 dm2 AREA=1.015e-06
D6593 n6594 0 dm2 AREA=6.801e-07
D6594 n6595 0 dm2 AREA=4.848e-07
D6595 n6596 0 dm2 AREA=2.477e-06
D6596 n6597 0 dm2 AREA=1.879e-06
D6597 n6598 0 dm2 AREA=1.157e-06
D6598 n6599 0 dm2 AREA=1.052e-06
D6599 n6600 0 dm2 AREA=1.528e-06
D6600 n6601 0 dm2 AREA=1.170e-06
D6601 n6602 0 dm2 AREA=1.585e-06
D6602 n6603 0 dm2 AREA=1.138e-06
D6603 n6604 0 dm2 AREA=1.942e-06
D6604 n6605 0 dm2 AREA=6.837e-07
D6605 n6606 0 dm2 AREA=5.664e-07
D6606 n6607 0 dm2 AREA=6.266e-07
D6607 n6608 0 dm2 AREA=5.565e-07
D6608 n6609 0 dm2 AREA=5.505e-07
D6609 n6610 0 dm2 AREA=4.797e-07
D6610 n6611 0 dm2 AREA=4.086e-07
D6611 n6612 0 dm2 AREA=8.390e-07
D6612 n6613 0 dm2 AREA=7.562e-07
D6613 n6614 0 dm2 AREA=1.470e-06
D6614 n6615 0 dm2 AREA=1.054e-06
D6615 n6616 0 dm2 AREA=6.917e-07
D6616 n6617 0 dm2 AREA=9.748e-07
D6617 n6618 0 dm2 AREA=3.851e-07
D6618 n6619 0 dm2 AREA=1.581e-06
D6619 n6620 0 dm2 AREA=8.485e-07
D6620 n6621 0 dm2 AREA=9.538e-07
D6621 n6622 0 dm2 AREA=1.966e-07
D6622 n6623 0 dm2 AREA=4.653e-07
D6623 n6624 0 dm2 AREA=9.217e-07
D6624 n6625 0 dm2 AREA=9.486e-07
D6625 n6626 0 dm2 AREA=1.258e-06
D6626 n6627 0 dm2 AREA=6.009e-07
D6627 n6628 0 dm2 AREA=6.427e-07
D6628 n6629 0 dm2 AREA=5.126e-07
D6629 n6630 0 dm2 AREA=1.440e-06
D6630 n6631 0 dm2 AREA=5.035e-07
D6631 n6632 0 dm2 AREA=6.530e-07
D6632 n6633 0 dm2 AREA=1.885e-06
D6633 n6634 0 dm2 AREA=1.873e-06
D6634 n6635 0 dm2 AREA=2.481e-07
D6635 n6636 0 dm2 AREA=1.997e-06
D6636 n6637 0 dm2 AREA=6.767e-07
D6637 n6638 0 dm2 AREA=1.538e-06
D6638 n6639 0 dm2 AREA=4.616e-07
D6639 n6640 0 dm2 AREA=2.700e-07
D6640 n6641 0 dm2 AREA=1.593e-06
D6641 n6642 0 dm2 AREA=1.938e-06
D6642 n6643 0 dm2 AREA=2.000e-06
D6643 n6644 0 dm2 AREA=1.227e-06
D6644 n6645 0 dm2 AREA=1.065e-06
D6645 n6646 0 dm2 AREA=1.081e-06
D6646 n1 0 dm2 AREA=5.536e-07
D6647 n6648 0 dm2 AREA=1.252e-06
D6648 n6649 0 dm2 AREA=8.564e-07
D6649 n6650 0 dm2 AREA=1.150e-06
D6650 n6651 0 dm2 AREA=1.717e-06
D6651 n6652 0 dm2 AREA=2.947e-06
D6652 n6653 0 dm2 AREA=5.658e-07
D6653 n6654 0 dm2 AREA=1.269e-06
D6654 n6655 0 dm2 AREA=7.774e-07
D6655 n6656 0 dm2 AREA=1.496e-06
D6656 n6657 0 dm2 AREA=7.571e-07
D6657 n6658 0 dm2 AREA=1.200e-06
D6658 n6659 0 dm2 AREA=3.567e-07
D6659 n6660 0 dm2 AREA=2.503e-06
D6660 n6661 0 dm2 AREA=1.417e-06
D6661 n6662 0 dm2 AREA=1.034e-06
D6662 n6663 0 dm2 AREA=1.457e-06
D6663 n6664 0 dm2 AREA=1.057e-06
D6664 n6665 0 dm2 AREA=4.464e-07
D6665 n6666 0 dm2 AREA=1.548e-06
D6666 n6667 0 dm2 AREA=1.083e-06
D6667 n6668 0 dm2 AREA=1.007e-06
D6668 n6669 0 dm2 AREA=2.258e-06
D6669 n6670 0 dm2 AREA=4.813e-07
D6670 n6671 0 dm2 AREA=9.900e-07
D6671 n6672 0 dm2 AREA=6.013e-07
D6672 n6673 0 dm2 AREA=4.423e-07
D6673 n6674 0 dm2 AREA=2.703e-06
D6674 n6675 0 dm2 AREA=1.750e-06
D6675 n6676 0 dm2 AREA=7.992e-07
D6676 n6677 0 dm2 AREA=5.602e-07
D6677 n6678 0 dm2 AREA=1.699e-06
D6678 n6679 0 dm2 AREA=1.861e-06
D6679 n6680 0 dm2 AREA=9.573e-07
D6680 n6681 0 dm2 AREA=5.364e-07
D6681 n6682 0 dm2 AREA=9.004e-07
D6682 n6683 0 dm2 AREA=8.500e-07
D6683 n6684 0 dm2 AREA=4.327e-07
D6684 n6685 0 dm2 AREA=2.130e-07
D6685 n6686 0 dm2 AREA=7.854e-07
D6686 n6687 0 dm2 AREA=7.085e-07
D6687 n6688 0 dm2 AREA=2.551e-06
D6688 n6689 0 dm2 AREA=1.386e-06
D6689 n6690 0 dm2 AREA=9.354e-07
D6690 n6691 0 dm2 AREA=1.202e-07
D6691 n6692 0 dm2 AREA=8.412e-07
D6692 n6693 0 dm2 AREA=7.471e-07
D6693 n6694 0 dm2 AREA=1.902e-06
D6694 n6695 0 dm2 AREA=1.375e-06
D6695 n6696 0 dm2 AREA=4.524e-07
D6696 n6697 0 dm2 AREA=8.529e-07
D6697 n6698 0 dm2 AREA=1.991e-06
D6698 n6699 0 dm2 AREA=8.797e-07
D6699 n6700 0 dm2 AREA=3.279e-07
D6700 n6701 0 dm2 AREA=6.935e-07
D6701 n6702 0 dm2 AREA=4.993e-07
D6702 n6703 0 dm2 AREA=5.364e-07
D6703 n6704 0 dm2 AREA=5.881e-07
D6704 n6705 0 dm2 AREA=8.583e-07
D6705 n6706 0 dm2 AREA=2.827e-06
D6706 n6707 0 dm2 AREA=8.344e-07
D6707 n6708 0 dm2 AREA=6.138e-07
D6708 n6709 0 dm2 AREA=1.999e-06
D6709 n6710 0 dm2 AREA=1.247e-06
D6710 n6711 0 dm2 AREA=1.482e-06
D6711 n6712 0 dm2 AREA=6.313e-07
D6712 n6713 0 dm2 AREA=1.742e-06
D6713 n6714 0 dm2 AREA=1.448e-06
D6714 n6715 0 dm2 AREA=8.041e-07
D6715 n6716 0 dm2 AREA=1.071e-06
D6716 n6717 0 dm2 AREA=2.937e-07
D6717 n6718 0 dm2 AREA=1.688e-07
D6718 n6719 0 dm2 AREA=4.896e-07
D6719 n6720 0 dm2 AREA=5.290e-07
D6720 n6721 0 dm2 AREA=7.135e-07
D6721 n6722 0 dm2 AREA=6.118e-07
D6722 n6723 0 dm2 AREA=7.680e-07
D6723 n6724 0 dm2 AREA=2.670e-06
D6724 n6725 0 dm2 AREA=6.224e-07
D6725 n6726 0 dm2 AREA=6.563e-07
D6726 n6727 0 dm2 AREA=5.911e-07
D6727 n6728 0 dm2 AREA=7.429e-07
D6728 n6729 0 dm2 AREA=8.701e-07
D6729 n6730 0 dm2 AREA=1.141e-06
D6730 n6731 0 dm2 AREA=1.554e-06
D6731 n6732 0 dm2 AREA=8.146e-07
D6732 n6733 0 dm2 AREA=7.921e-07
D6733 n6734 0 dm2 AREA=1.223e-06
D6734 n6735 0 dm2 AREA=7.561e-07
D6735 n6736 0 dm2 AREA=4.134e-07
D6736 n6737 0 dm2 AREA=3.686e-07
D6737 n6738 0 dm2 AREA=6.335e-07
D6738 n6739 0 dm2 AREA=3.718e-07
D6739 n6740 0 dm2 AREA=1.189e-06
D6740 n6741 0 dm2 AREA=8.153e-07
D6741 n6742 0 dm2 AREA=7.430e-07
D6742 n6743 0 dm2 AREA=1.129e-06
D6743 n6744 0 dm2 AREA=9.255e-07
D6744 n6745 0 dm2 AREA=5.497e-07
D6745 n6746 0 dm2 AREA=6.985e-07
D6746 n6747 0 dm2 AREA=1.098e-06
D6747 n6748 0 dm2 AREA=4.024e-07
D6748 n6749 0 dm2 AREA=9.304e-07
D6749 n6750 0 dm2 AREA=8.235e-07
D6750 n6751 0 dm2 AREA=1.855e-06
D6751 n6752 0 dm2 AREA=2.591e-07
D6752 n6753 0 dm2 AREA=8.525e-07
D6753 n6754 0 dm2 AREA=3.428e-07
D6754 n6755 0 dm2 AREA=5.755e-07
D6755 n6756 0 dm2 AREA=4.975e-07
D6756 n6757 0 dm2 AREA=8.460e-07
D6757 n6758 0 dm2 AREA=7.740e-07
D6758 n6759 0 dm2 AREA=9.007e-07
D6759 n6760 0 dm2 AREA=1.117e-06
D6760 n6761 0 dm2 AREA=5.144e-07
D6761 n6762 0 dm2 AREA=7.848e-07
D6762 n6763 0 dm2 AREA=8.832e-07
D6763 n6764 0 dm2 AREA=1.253e-06
D6764 n6765 0 dm2 AREA=1.653e-06
D6765 n6766 0 dm2 AREA=5.606e-07
D6766 n6767 0 dm2 AREA=9.906e-07
D6767 n6768 0 dm2 AREA=8.795e-07
D6768 n6769 0 dm2 AREA=1.351e-06
D6769 n6770 0 dm2 AREA=1.423e-06
D6770 n6771 0 dm2 AREA=8.477e-07
D6771 n6772 0 dm2 AREA=6.827e-07
D6772 n6773 0 dm2 AREA=9.882e-07
D6773 n6774 0 dm2 AREA=7.507e-07
D6774 n6775 0 dm2 AREA=7.080e-07
D6775 n6776 0 dm2 AREA=8.368e-07
D6776 n6777 0 dm2 AREA=9.572e-07
D6777 n6778 0 dm2 AREA=8.325e-07
D6778 n6779 0 dm2 AREA=1.366e-06
D6779 n6780 0 dm2 AREA=1.513e-06
D6780 n6781 0 dm2 AREA=9.063e-07
D6781 n6782 0 dm2 AREA=2.042e-07
D6782 n6783 0 dm2 AREA=7.354e-07
D6783 n6784 0 dm2 AREA=2.516e-06
D6784 n6785 0 dm2 AREA=5.206e-07
D6785 n6786 0 dm2 AREA=1.300e-07
D6786 n6787 0 dm2 AREA=4.601e-07
D6787 n6788 0 dm2 AREA=4.960e-07
D6788 n6789 0 dm2 AREA=1.991e-06
D6789 n6790 0 dm2 AREA=9.159e-07
D6790 n6791 0 dm2 AREA=1.384e-06
D6791 n6792 0 dm2 AREA=2.237e-06
D6792 n6793 0 dm2 AREA=7.658e-07
D6793 n6794 0 dm2 AREA=8.507e-07
D6794 n6795 0 dm2 AREA=1.354e-06
D6795 n6796 0 dm2 AREA=8.910e-07
D6796 n6797 0 dm2 AREA=1.462e-07
D6797 n6798 0 dm2 AREA=5.764e-07
D6798 n6799 0 dm2 AREA=3.318e-07
D6799 n6800 0 dm2 AREA=8.248e-07
D6800 n6801 0 dm2 AREA=7.684e-07
D6801 n6802 0 dm2 AREA=1.244e-06
D6802 n6803 0 dm2 AREA=1.062e-06
D6803 n6804 0 dm2 AREA=1.513e-06
D6804 n6805 0 dm2 AREA=1.310e-06
D6805 n6806 0 dm2 AREA=2.320e-06
D6806 n6807 0 dm2 AREA=8.625e-07
D6807 n6808 0 dm2 AREA=6.042e-07
D6808 n6809 0 dm2 AREA=5.931e-07
D6809 n6810 0 dm2 AREA=1.007e-06
D6810 n6811 0 dm2 AREA=1.314e-06
D6811 n6812 0 dm2 AREA=2.274e-06
D6812 n6813 0 dm2 AREA=6.624e-07
D6813 n6814 0 dm2 AREA=1.207e-06
D6814 n6815 0 dm2 AREA=1.091e-06
D6815 n6816 0 dm2 AREA=2.120e-07
D6816 n6817 0 dm2 AREA=8.122e-07
D6817 n6818 0 dm2 AREA=5.828e-07
D6818 n6819 0 dm2 AREA=5.995e-07
D6819 n6820 0 dm2 AREA=6.214e-07
D6820 n6821 0 dm2 AREA=1.437e-06
D6821 n6822 0 dm2 AREA=1.465e-06
D6822 n6823 0 dm2 AREA=3.887e-07
D6823 n6824 0 dm2 AREA=1.526e-06
D6824 n6825 0 dm2 AREA=9.028e-07
D6825 n6826 0 dm2 AREA=1.032e-06
D6826 n6827 0 dm2 AREA=6.258e-07
D6827 n6828 0 dm2 AREA=6.318e-07
D6828 n6829 0 dm2 AREA=8.051e-07
D6829 n6830 0 dm2 AREA=1.034e-06
D6830 n6831 0 dm2 AREA=8.445e-07
D6831 n6832 0 dm2 AREA=2.865e-07
D6832 n6833 0 dm2 AREA=1.209e-06
D6833 n6834 0 dm2 AREA=1.522e-06
D6834 n6835 0 dm2 AREA=8.150e-07
D6835 n6836 0 dm2 AREA=4.158e-07
D6836 n6837 0 dm2 AREA=1.098e-06
D6837 n6838 0 dm2 AREA=1.197e-06
D6838 n6839 0 dm2 AREA=1.194e-06
D6839 n6840 0 dm2 AREA=1.814e-06
D6840 n6841 0 dm2 AREA=1.090e-06
D6841 n6842 0 dm2 AREA=1.495e-06
D6842 n6843 0 dm2 AREA=1.121e-06
D6843 n6844 0 dm2 AREA=4.681e-07
D6844 n6845 0 dm2 AREA=4.058e-07
D6845 n6846 0 dm2 AREA=1.167e-06
D6846 n6847 0 dm2 AREA=1.236e-06
D6847 n6848 0 dm2 AREA=1.140e-06
D6848 n6849 0 dm2 AREA=1.801e-07
D6849 n6850 0 dm2 AREA=7.520e-07
D6850 n6851 0 dm2 AREA=5.091e-07
D6851 n6852 0 dm2 AREA=3.926e-07
D6852 n6853 0 dm2 AREA=9.244e-07
D6853 n6854 0 dm2 AREA=3.374e-06
D6854 n6855 0 dm2 AREA=7.713e-07
D6855 n6856 0 dm2 AREA=1.424e-06
D6856 n6857 0 dm2 AREA=1.650e-06
D6857 n6858 0 dm2 AREA=1.404e-06
D6858 n6859 0 dm2 AREA=1.038e-06
D6859 n6860 0 dm2 AREA=9.372e-07
D6860 n6861 0 dm2 AREA=1.914e-06
D6861 n6862 0 dm2 AREA=5.576e-07
D6862 n6863 0 dm2 AREA=9.290e-07
D6863 n6864 0 dm2 AREA=5.137e-07
D6864 n6865 0 dm2 AREA=7.042e-08
D6865 n6866 0 dm2 AREA=4.628e-07
D6866 n6867 0 dm2 AREA=6.348e-07
D6867 n6868 0 dm2 AREA=1.329e-06
D6868 n6869 0 dm2 AREA=2.812e-06
D6869 n6870 0 dm2 AREA=5.195e-07
D6870 n6871 0 dm2 AREA=3.099e-07
D6871 n6872 0 dm2 AREA=7.729e-07
D6872 n6873 0 dm2 AREA=1.243e-06
D6873 n6874 0 dm2 AREA=8.202e-07
D6874 n6875 0 dm2 AREA=5.241e-07
D6875 n6876 0 dm2 AREA=1.061e-06
D6876 n6877 0 dm2 AREA=7.334e-07
D6877 n6878 0 dm2 AREA=7.541e-07
D6878 n6879 0 dm2 AREA=1.136e-06
D6879 n6880 0 dm2 AREA=1.182e-06
D6880 n6881 0 dm2 AREA=4.630e-07
D6881 n6882 0 dm2 AREA=8.095e-07
D6882 n6883 0 dm2 AREA=4.492e-07
D6883 n6884 0 dm2 AREA=7.642e-07
D6884 n6885 0 dm2 AREA=2.118e-06
D6885 n6886 0 dm2 AREA=1.326e-06
D6886 n6887 0 dm2 AREA=7.498e-07
D6887 n6888 0 dm2 AREA=1.483e-06
D6888 n6889 0 dm2 AREA=1.071e-06
D6889 n6890 0 dm2 AREA=6.602e-07
D6890 n6891 0 dm2 AREA=1.185e-06
D6891 n6892 0 dm2 AREA=2.535e-06
D6892 n6893 0 dm2 AREA=3.702e-07
D6893 n6894 0 dm2 AREA=8.358e-07
D6894 n6895 0 dm2 AREA=8.962e-07
D6895 n6896 0 dm2 AREA=8.031e-07
D6896 n6897 0 dm2 AREA=2.255e-07
D6897 n6898 0 dm2 AREA=2.504e-07
D6898 n6899 0 dm2 AREA=5.770e-07
D6899 n6900 0 dm2 AREA=6.353e-07
D6900 n6901 0 dm2 AREA=7.280e-07
D6901 n6902 0 dm2 AREA=2.172e-06
D6902 n6903 0 dm2 AREA=8.278e-07
D6903 n6904 0 dm2 AREA=8.967e-07
D6904 n6905 0 dm2 AREA=1.500e-06
D6905 n6906 0 dm2 AREA=7.494e-07
D6906 n6907 0 dm2 AREA=1.143e-06
D6907 n6908 0 dm2 AREA=1.431e-06
D6908 n6909 0 dm2 AREA=1.183e-06
D6909 n6910 0 dm2 AREA=1.159e-06
D6910 n6911 0 dm2 AREA=7.997e-07
D6911 n6912 0 dm2 AREA=1.849e-06
D6912 n6913 0 dm2 AREA=2.945e-06
D6913 n6914 0 dm2 AREA=1.238e-06
D6914 n6915 0 dm2 AREA=1.489e-06
D6915 n6916 0 dm2 AREA=9.382e-07
D6916 n6917 0 dm2 AREA=7.988e-07
D6917 n6918 0 dm2 AREA=3.017e-07
D6918 n6919 0 dm2 AREA=1.063e-06
D6919 n6920 0 dm2 AREA=7.082e-07
D6920 n6921 0 dm2 AREA=1.545e-06
D6921 n6922 0 dm2 AREA=4.670e-07
D6922 n6923 0 dm2 AREA=1.002e-06
D6923 n6924 0 dm2 AREA=8.202e-07
D6924 n6925 0 dm2 AREA=1.161e-06
D6925 n6926 0 dm2 AREA=1.543e-07
D6926 n6927 0 dm2 AREA=4.467e-07
D6927 n6928 0 dm2 AREA=5.007e-07
D6928 n6929 0 dm2 AREA=1.435e-06
D6929 n6930 0 dm2 AREA=3.219e-07
D6930 n6931 0 dm2 AREA=1.438e-06
D6931 n6932 0 dm2 AREA=6.053e-07
D6932 n6933 0 dm2 AREA=2.308e-07
D6933 n6934 0 dm2 AREA=2.245e-06
D6934 n6935 0 dm2 AREA=1.206e-07
D6935 n6936 0 dm2 AREA=5.972e-07
D6936 n6937 0 dm2 AREA=1.300e-06
D6937 n6938 0 dm2 AREA=1.481e-06
D6938 n6939 0 dm2 AREA=1.486e-06
D6939 n6940 0 dm2 AREA=1.263e-06
D6940 n6941 0 dm2 AREA=7.115e-07
D6941 n6942 0 dm2 AREA=3.629e-07
D6942 n6943 0 dm2 AREA=1.258e-06
D6943 n6944 0 dm2 AREA=5.553e-07
D6944 n6945 0 dm2 AREA=7.323e-07
D6945 n6946 0 dm2 AREA=1.418e-06
D6946 n6947 0 dm2 AREA=6.412e-07
D6947 n6948 0 dm2 AREA=5.113e-07
D6948 n6949 0 dm2 AREA=1.235e-06
D6949 n6950 0 dm2 AREA=7.348e-07
D6950 n6951 0 dm2 AREA=7.974e-07
D6951 n6952 0 dm2 AREA=4.211e-07
D6952 n6953 0 dm2 AREA=2.143e-06
D6953 n6954 0 dm2 AREA=5.467e-07
D6954 n6955 0 dm2 AREA=1.097e-06
D6955 n6956 0 dm2 AREA=1.490e-06
D6956 n6957 0 dm2 AREA=1.288e-06
D6957 n6958 0 dm2 AREA=6.000e-07
D6958 n6959 0 dm2 AREA=6.940e-07
D6959 n6960 0 dm2 AREA=1.335e-06
D6960 n6961 0 dm2 AREA=1.461e-06
D6961 n6962 0 dm2 AREA=9.446e-07
D6962 n6963 0 dm2 AREA=3.583e-06
D6963 n6964 0 dm2 AREA=8.129e-07
D6964 n6965 0 dm2 AREA=4.043e-07
D6965 n6966 0 dm2 AREA=5.735e-07
D6966 n1 0 dm2 AREA=9.947e-07
D6967 n6968 0 dm2 AREA=1.144e-06
D6968 n6969 0 dm2 AREA=7.537e-07
D6969 n6970 0 dm2 AREA=4.644e-07
D6970 n6971 0 dm2 AREA=1.353e-06
D6971 n6972 0 dm2 AREA=8.013e-07
D6972 n6973 0 dm2 AREA=1.212e-06
D6973 n6974 0 dm2 AREA=1.491e-06
D6974 n6975 0 dm2 AREA=1.386e-06
D6975 n6976 0 dm2 AREA=1.459e-06
D6976 n6977 0 dm2 AREA=1.784e-06
D6977 n6978 0 dm2 AREA=9.489e-07
D6978 n6979 0 dm2 AREA=3.092e-06
D6979 n6980 0 dm2 AREA=1.211e-06
D6980 n6981 0 dm2 AREA=1.158e-06
D6981 n6982 0 dm2 AREA=1.968e-07
D6982 n6983 0 dm2 AREA=1.517e-06
D6983 n6984 0 dm2 AREA=8.104e-07
D6984 n6985 0 dm2 AREA=1.540e-06
D6985 n6986 0 dm2 AREA=1.185e-06
D6986 n6987 0 dm2 AREA=1.243e-06
D6987 n6988 0 dm2 AREA=9.465e-07
D6988 n6989 0 dm2 AREA=2.917e-07
D6989 n6990 0 dm2 AREA=9.217e-07
D6990 n6991 0 dm2 AREA=8.959e-07
D6991 n6992 0 dm2 AREA=5.382e-07
D6992 n6993 0 dm2 AREA=7.519e-07
D6993 n6994 0 dm2 AREA=5.570e-07
D6994 n6995 0 dm2 AREA=1.343e-06
D6995 n6996 0 dm2 AREA=2.363e-06
D6996 n6997 0 dm2 AREA=4.763e-07
D6997 n6998 0 dm2 AREA=9.587e-07
D6998 n6999 0 dm2 AREA=1.291e-06
D6999 n7000 0 dm2 AREA=8.534e-07
D7000 n7001 0 dm2 AREA=1.430e-06
D7001 n7002 0 dm2 AREA=1.094e-06
D7002 n7003 0 dm2 AREA=1.465e-06
D7003 n7004 0 dm2 AREA=3.908e-07
D7004 n7005 0 dm2 AREA=1.113e-06
D7005 n7006 0 dm2 AREA=4.659e-07
D7006 n7007 0 dm2 AREA=3.397e-07
D7007 n7008 0 dm2 AREA=1.049e-06
D7008 n7009 0 dm2 AREA=1.610e-06
D7009 n7010 0 dm2 AREA=2.779e-07
D7010 n7011 0 dm2 AREA=2.283e-06
D7011 n7012 0 dm2 AREA=7.668e-07
D7012 n7013 0 dm2 AREA=1.465e-06
D7013 n7014 0 dm2 AREA=5.483e-07
D7014 n7015 0 dm2 AREA=1.041e-06
D7015 n7016 0 dm2 AREA=5.779e-07
D7016 n7017 0 dm2 AREA=1.601e-06
D7017 n7018 0 dm2 AREA=9.453e-07
D7018 n7019 0 dm2 AREA=3.403e-07
D7019 n7020 0 dm2 AREA=1.302e-06
D7020 n7021 0 dm2 AREA=1.596e-06
D7021 n7022 0 dm2 AREA=1.274e-06
D7022 n7023 0 dm2 AREA=8.337e-07
D7023 n7024 0 dm2 AREA=2.032e-06
D7024 n7025 0 dm2 AREA=2.562e-06
D7025 n7026 0 dm2 AREA=5.656e-07
D7026 n7027 0 dm2 AREA=1.071e-06
D7027 n7028 0 dm2 AREA=2.336e-07
D7028 n7029 0 dm2 AREA=6.749e-07
D7029 n7030 0 dm2 AREA=9.179e-07
D7030 n7031 0 dm2 AREA=8.291e-07
D7031 n7032 0 dm2 AREA=1.646e-06
D7032 n7033 0 dm2 AREA=5.224e-07
D7033 n7034 0 dm2 AREA=1.550e-06
D7034 n7035 0 dm2 AREA=1.647e-06
D7035 n7036 0 dm2 AREA=9.247e-07
D7036 n7037 0 dm2 AREA=2.030e-06
D7037 n7038 0 dm2 AREA=4.414e-07
D7038 n7039 0 dm2 AREA=7.460e-07
D7039 n7040 0 dm2 AREA=9.684e-07
D7040 n7041 0 dm2 AREA=5.859e-07
D7041 n7042 0 dm2 AREA=7.725e-07
D7042 n7043 0 dm2 AREA=1.294e-06
D7043 n7044 0 dm2 AREA=1.473e-06
D7044 n7045 0 dm2 AREA=1.040e-06
D7045 n7046 0 dm2 AREA=8.834e-07
D7046 n7047 0 dm2 AREA=5.770e-07
D7047 n7048 0 dm2 AREA=2.158e-06
D7048 n7049 0 dm2 AREA=1.331e-06
D7049 n7050 0 dm2 AREA=7.726e-07
D7050 n7051 0 dm2 AREA=6.000e-07
D7051 n7052 0 dm2 AREA=6.619e-07
D7052 n7053 0 dm2 AREA=1.062e-06
D7053 n7054 0 dm2 AREA=1.015e-06
D7054 n7055 0 dm2 AREA=6.597e-07
D7055 n7056 0 dm2 AREA=1.480e-06
D7056 n7057 0 dm2 AREA=3.103e-07
D7057 n7058 0 dm2 AREA=1.006e-06
D7058 n7059 0 dm2 AREA=7.023e-07
D7059 n7060 0 dm2 AREA=1.959e-06
D7060 n7061 0 dm2 AREA=5.816e-07
D7061 n7062 0 dm2 AREA=5.212e-07
D7062 n7063 0 dm2 AREA=4.260e-07
D7063 n7064 0 dm2 AREA=1.826e-07
D7064 n7065 0 dm2 AREA=1.394e-06
D7065 n7066 0 dm2 AREA=6.308e-07
D7066 n7067 0 dm2 AREA=5.022e-07
D7067 n7068 0 dm2 AREA=1.884e-06
D7068 n7069 0 dm2 AREA=2.279e-07
D7069 n7070 0 dm2 AREA=2.187e-06
D7070 n7071 0 dm2 AREA=1.931e-06
D7071 n7072 0 dm2 AREA=2.472e-06
D7072 n7073 0 dm2 AREA=6.439e-07
D7073 n7074 0 dm2 AREA=3.844e-07
D7074 n7075 0 dm2 AREA=6.873e-07
D7075 n7076 0 dm2 AREA=1.470e-07
D7076 n7077 0 dm2 AREA=1.304e-06
D7077 n7078 0 dm2 AREA=4.348e-07
D7078 n7079 0 dm2 AREA=7.727e-07
D7079 n7080 0 dm2 AREA=9.182e-07
D7080 n7081 0 dm2 AREA=2.813e-07
D7081 n7082 0 dm2 AREA=3.319e-07
D7082 n7083 0 dm2 AREA=1.566e-06
D7083 n7084 0 dm2 AREA=1.473e-06
D7084 n7085 0 dm2 AREA=9.273e-07
D7085 n7086 0 dm2 AREA=8.056e-07
D7086 n7087 0 dm2 AREA=1.654e-06
D7087 n7088 0 dm2 AREA=1.189e-06
D7088 n7089 0 dm2 AREA=1.665e-06
D7089 n7090 0 dm2 AREA=7.547e-07
D7090 n7091 0 dm2 AREA=6.267e-07
D7091 n7092 0 dm2 AREA=1.049e-06
D7092 n7093 0 dm2 AREA=2.965e-07
D7093 n7094 0 dm2 AREA=9.268e-07
D7094 n7095 0 dm2 AREA=1.708e-06
D7095 n7096 0 dm2 AREA=1.572e-06
D7096 n7097 0 dm2 AREA=6.366e-07
D7097 n7098 0 dm2 AREA=5.886e-07
D7098 n7099 0 dm2 AREA=9.092e-07
D7099 n7100 0 dm2 AREA=7.124e-07
D7100 n7101 0 dm2 AREA=3.977e-07
D7101 n7102 0 dm2 AREA=8.346e-07
D7102 n7103 0 dm2 AREA=7.280e-07
D7103 n7104 0 dm2 AREA=1.731e-06
D7104 n7105 0 dm2 AREA=1.202e-06
D7105 n7106 0 dm2 AREA=8.896e-07
D7106 n7107 0 dm2 AREA=1.003e-06
D7107 n7108 0 dm2 AREA=1.038e-06
D7108 n7109 0 dm2 AREA=1.710e-06
D7109 n7110 0 dm2 AREA=1.376e-06
D7110 n7111 0 dm2 AREA=9.394e-07
D7111 n7112 0 dm2 AREA=4.070e-07
D7112 n7113 0 dm2 AREA=7.383e-07
D7113 n7114 0 dm2 AREA=1.750e-06
D7114 n7115 0 dm2 AREA=5.983e-07
D7115 n7116 0 dm2 AREA=7.256e-07
D7116 n7117 0 dm2 AREA=4.086e-07
D7117 n7118 0 dm2 AREA=1.071e-06
D7118 n7119 0 dm2 AREA=9.850e-07
D7119 n7120 0 dm2 AREA=8.707e-07
D7120 n7121 0 dm2 AREA=5.258e-07
D7121 n7122 0 dm2 AREA=1.946e-06
D7122 n7123 0 dm2 AREA=1.501e-06
D7123 n7124 0 dm2 AREA=9.663e-07
D7124 n7125 0 dm2 AREA=1.201e-06
D7125 n7126 0 dm2 AREA=5.408e-07
D7126 n7127 0 dm2 AREA=5.228e-07
D7127 n7128 0 dm2 AREA=5.673e-07
D7128 n7129 0 dm2 AREA=1.450e-06
D7129 n7130 0 dm2 AREA=2.014e-06
D7130 n7131 0 dm2 AREA=4.032e-07
D7131 n7132 0 dm2 AREA=1.277e-06
D7132 n7133 0 dm2 AREA=3.672e-07
D7133 n7134 0 dm2 AREA=6.914e-07
D7134 n7135 0 dm2 AREA=6.702e-07
D7135 n7136 0 dm2 AREA=7.833e-07
D7136 n7137 0 dm2 AREA=8.382e-07
D7137 n7138 0 dm2 AREA=9.768e-07
D7138 n7139 0 dm2 AREA=6.094e-07
D7139 n7140 0 dm2 AREA=1.566e-06
D7140 n7141 0 dm2 AREA=1.420e-06
D7141 n7142 0 dm2 AREA=1.510e-06
D7142 n7143 0 dm2 AREA=1.999e-06
D7143 n7144 0 dm2 AREA=9.565e-07
D7144 n7145 0 dm2 AREA=2.887e-06
D7145 n7146 0 dm2 AREA=2.899e-06
D7146 n7147 0 dm2 AREA=7.631e-07
D7147 n7148 0 dm2 AREA=8.377e-07
D7148 n7149 0 dm2 AREA=7.269e-07
D7149 n7150 0 dm2 AREA=7.925e-08
D7150 n7151 0 dm2 AREA=1.055e-06
D7151 n7152 0 dm2 AREA=2.811e-07
D7152 n7153 0 dm2 AREA=1.554e-06
D7153 n7154 0 dm2 AREA=4.659e-07
D7154 n7155 0 dm2 AREA=8.588e-07
D7155 n7156 0 dm2 AREA=6.181e-07
D7156 n7157 0 dm2 AREA=1.700e-06
D7157 n7158 0 dm2 AREA=1.163e-06
D7158 n7159 0 dm2 AREA=1.043e-06
D7159 n7160 0 dm2 AREA=1.388e-06
D7160 n7161 0 dm2 AREA=1.229e-06
D7161 n7162 0 dm2 AREA=1.402e-06
D7162 n7163 0 dm2 AREA=5.519e-07
D7163 n7164 0 dm2 AREA=5.390e-07
D7164 n7165 0 dm2 AREA=9.722e-07
D7165 n7166 0 dm2 AREA=1.028e-06
D7166 n7167 0 dm2 AREA=7.649e-07
D7167 n7168 0 dm2 AREA=1.025e-06
D7168 n1 0 dm2 AREA=2.157e-07
D7169 n7170 0 dm2 AREA=6.130e-07
D7170 n7171 0 dm2 AREA=4.804e-07
D7171 n7172 0 dm2 AREA=4.851e-07
D7172 n7173 0 dm2 AREA=9.342e-07
D7173 n7174 0 dm2 AREA=6.431e-07
D7174 n7175 0 dm2 AREA=1.863e-06
D7175 n7176 0 dm2 AREA=1.040e-06
D7176 n7177 0 dm2 AREA=2.819e-07
D7177 n7178 0 dm2 AREA=2.412e-07
D7178 n7179 0 dm2 AREA=1.141e-06
D7179 n7180 0 dm2 AREA=2.357e-06
D7180 n7181 0 dm2 AREA=7.857e-07
D7181 n7182 0 dm2 AREA=6.407e-07
D7182 n7183 0 dm2 AREA=1.955e-06
D7183 n7184 0 dm2 AREA=6.504e-07
D7184 n7185 0 dm2 AREA=3.403e-07
D7185 n7186 0 dm2 AREA=7.053e-07
D7186 n7187 0 dm2 AREA=7.651e-07
D7187 n7188 0 dm2 AREA=1.448e-06
D7188 n7189 0 dm2 AREA=1.513e-06
D7189 n7190 0 dm2 AREA=1.313e-06
D7190 n7191 0 dm2 AREA=1.129e-06
D7191 n7192 0 dm2 AREA=1.855e-06
D7192 n7193 0 dm2 AREA=4.948e-07
D7193 n7194 0 dm2 AREA=9.615e-07
D7194 n7195 0 dm2 AREA=1.969e-06
D7195 n7196 0 dm2 AREA=1.127e-06
D7196 n7197 0 dm2 AREA=1.328e-06
D7197 n7198 0 dm2 AREA=1.405e-06
D7198 n7199 0 dm2 AREA=3.735e-07
D7199 n7200 0 dm2 AREA=1.830e-06
D7200 n7201 0 dm2 AREA=4.236e-07
D7201 n7202 0 dm2 AREA=6.751e-07
D7202 n7203 0 dm2 AREA=4.161e-07
D7203 n7204 0 dm2 AREA=1.953e-07
D7204 n7205 0 dm2 AREA=1.256e-06
D7205 n7206 0 dm2 AREA=7.722e-07
D7206 n7207 0 dm2 AREA=9.701e-07
D7207 n7208 0 dm2 AREA=1.554e-06
D7208 n7209 0 dm2 AREA=8.120e-07
D7209 n7210 0 dm2 AREA=1.195e-06
D7210 n7211 0 dm2 AREA=4.135e-07
D7211 n7212 0 dm2 AREA=1.245e-06
D7212 n7213 0 dm2 AREA=5.599e-07
D7213 n7214 0 dm2 AREA=2.744e-06
D7214 n7215 0 dm2 AREA=2.750e-07
D7215 n7216 0 dm2 AREA=1.457e-06
D7216 n7217 0 dm2 AREA=1.643e-06
D7217 n7218 0 dm2 AREA=7.085e-07
D7218 n7219 0 dm2 AREA=1.601e-07
D7219 n7220 0 dm2 AREA=4.437e-07
D7220 n7221 0 dm2 AREA=1.671e-06
D7221 n7222 0 dm2 AREA=6.532e-07
D7222 n7223 0 dm2 AREA=1.304e-06
D7223 n7224 0 dm2 AREA=8.250e-07
D7224 n7225 0 dm2 AREA=9.751e-07
D7225 n7226 0 dm2 AREA=2.748e-07
D7226 n7227 0 dm2 AREA=1.723e-07
D7227 n7228 0 dm2 AREA=5.698e-07
D7228 n7229 0 dm2 AREA=3.792e-07
D7229 n7230 0 dm2 AREA=1.195e-06
D7230 n7231 0 dm2 AREA=1.618e-06
D7231 n7232 0 dm2 AREA=4.217e-07
D7232 n7233 0 dm2 AREA=1.027e-06
D7233 n7234 0 dm2 AREA=1.191e-06
D7234 n7235 0 dm2 AREA=7.241e-07
D7235 n7236 0 dm2 AREA=8.282e-07
D7236 n7237 0 dm2 AREA=1.365e-07
D7237 n7238 0 dm2 AREA=1.038e-06
D7238 n7239 0 dm2 AREA=7.584e-07
D7239 n7240 0 dm2 AREA=5.862e-07
D7240 n7241 0 dm2 AREA=3.322e-07
D7241 n7242 0 dm2 AREA=7.144e-07
D7242 n7243 0 dm2 AREA=1.668e-06
D7243 n7244 0 dm2 AREA=1.887e-06
D7244 n7245 0 dm2 AREA=5.332e-07
D7245 n7246 0 dm2 AREA=1.044e-06
D7246 n7247 0 dm2 AREA=8.767e-07
D7247 n7248 0 dm2 AREA=7.168e-07
D7248 n7249 0 dm2 AREA=9.362e-07
D7249 n7250 0 dm2 AREA=1.955e-07
D7250 n7251 0 dm2 AREA=7.274e-07
D7251 n7252 0 dm2 AREA=1.132e-06
D7252 n7253 0 dm2 AREA=4.233e-07
D7253 n7254 0 dm2 AREA=7.261e-07
D7254 n7255 0 dm2 AREA=3.955e-07
D7255 n7256 0 dm2 AREA=1.073e-06
D7256 n7257 0 dm2 AREA=1.116e-06
D7257 n7258 0 dm2 AREA=2.573e-06
D7258 n7259 0 dm2 AREA=5.721e-07
D7259 n7260 0 dm2 AREA=4.995e-07
D7260 n7261 0 dm2 AREA=1.318e-06
D7261 n7262 0 dm2 AREA=4.409e-07
D7262 n7263 0 dm2 AREA=2.338e-06
D7263 n7264 0 dm2 AREA=2.512e-07
D7264 n7265 0 dm2 AREA=9.688e-07
D7265 n7266 0 dm2 AREA=2.193e-06
D7266 n7267 0 dm2 AREA=1.596e-06
D7267 n7268 0 dm2 AREA=1.262e-06
D7268 n7269 0 dm2 AREA=5.034e-07
D7269 n7270 0 dm2 AREA=7.614e-07
D7270 n7271 0 dm2 AREA=1.059e-06
D7271 n7272 0 dm2 AREA=7.370e-07
D7272 n7273 0 dm2 AREA=6.558e-07
D7273 n7274 0 dm2 AREA=6.700e-07
D7274 n7275 0 dm2 AREA=1.008e-06
D7275 n7276 0 dm2 AREA=7.501e-07
D7276 n7277 0 dm2 AREA=7.231e-07
D7277 n7278 0 dm2 AREA=1.271e-06
D7278 n7279 0 dm2 AREA=7.572e-07
D7279 n7280 0 dm2 AREA=3.924e-07
D7280 n7281 0 dm2 AREA=1.288e-06
D7281 n7282 0 dm2 AREA=2.309e-06
D7282 n7283 0 dm2 AREA=1.534e-07
D7283 n7284 0 dm2 AREA=7.591e-07
D7284 n7285 0 dm2 AREA=2.274e-06
D7285 n7286 0 dm2 AREA=4.608e-07
D7286 n7287 0 dm2 AREA=2.044e-06
D7287 n7288 0 dm2 AREA=8.991e-07
D7288 n7289 0 dm2 AREA=1.070e-06
D7289 n7290 0 dm2 AREA=7.958e-07
D7290 n7291 0 dm2 AREA=8.421e-07
D7291 n7292 0 dm2 AREA=8.275e-07
D7292 n7293 0 dm2 AREA=1.405e-06
D7293 n7294 0 dm2 AREA=1.352e-06
D7294 n7295 0 dm2 AREA=8.157e-07
D7295 n7296 0 dm2 AREA=1.919e-07
D7296 n7297 0 dm2 AREA=2.770e-07
D7297 n7298 0 dm2 AREA=8.808e-07
D7298 n7299 0 dm2 AREA=4.074e-07
D7299 n7300 0 dm2 AREA=8.466e-07
D7300 n7301 0 dm2 AREA=9.741e-07
D7301 n7302 0 dm2 AREA=7.697e-07
D7302 n1 0 dm2 AREA=5.582e-07
D7303 n7304 0 dm2 AREA=1.827e-06
D7304 n7305 0 dm2 AREA=3.252e-07
D7305 n7306 0 dm2 AREA=9.146e-07
D7306 n7307 0 dm2 AREA=1.002e-06
D7307 n7308 0 dm2 AREA=1.369e-06
D7308 n7309 0 dm2 AREA=3.427e-07
D7309 n7310 0 dm2 AREA=1.134e-06
D7310 n7311 0 dm2 AREA=1.193e-06
D7311 n7312 0 dm2 AREA=1.098e-06
D7312 n7313 0 dm2 AREA=3.291e-07
D7313 n7314 0 dm2 AREA=7.687e-07
D7314 n7315 0 dm2 AREA=1.167e-06
D7315 n7316 0 dm2 AREA=3.866e-07
D7316 n7317 0 dm2 AREA=6.600e-07
D7317 n7318 0 dm2 AREA=5.777e-07
D7318 n7319 0 dm2 AREA=1.285e-06
D7319 n7320 0 dm2 AREA=4.769e-07
D7320 n7321 0 dm2 AREA=8.444e-07
D7321 n7322 0 dm2 AREA=9.524e-07
D7322 n7323 0 dm2 AREA=5.435e-07
D7323 n7324 0 dm2 AREA=5.643e-07
D7324 n7325 0 dm2 AREA=6.546e-07
D7325 n7326 0 dm2 AREA=5.614e-07
D7326 n7327 0 dm2 AREA=1.215e-06
D7327 n7328 0 dm2 AREA=6.938e-07
D7328 n7329 0 dm2 AREA=8.416e-07
D7329 n7330 0 dm2 AREA=1.878e-06
D7330 n7331 0 dm2 AREA=9.678e-07
D7331 n7332 0 dm2 AREA=1.241e-06
D7332 n7333 0 dm2 AREA=9.197e-07
D7333 n7334 0 dm2 AREA=1.408e-06
D7334 n7335 0 dm2 AREA=2.494e-07
D7335 n7336 0 dm2 AREA=2.633e-07
D7336 n7337 0 dm2 AREA=4.856e-07
D7337 n7338 0 dm2 AREA=2.840e-06
D7338 n7339 0 dm2 AREA=1.495e-06
D7339 n7340 0 dm2 AREA=1.350e-06
D7340 n7341 0 dm2 AREA=8.138e-07
D7341 n7342 0 dm2 AREA=2.322e-07
D7342 n7343 0 dm2 AREA=7.464e-07
D7343 n7344 0 dm2 AREA=5.700e-07
D7344 n7345 0 dm2 AREA=3.381e-07
D7345 n7346 0 dm2 AREA=3.973e-07
D7346 n7347 0 dm2 AREA=1.028e-06
D7347 n7348 0 dm2 AREA=1.256e-06
D7348 n7349 0 dm2 AREA=6.274e-07
D7349 n7350 0 dm2 AREA=1.378e-06
D7350 n7351 0 dm2 AREA=8.366e-07
D7351 n7352 0 dm2 AREA=2.198e-06
D7352 n7353 0 dm2 AREA=5.838e-07
D7353 n7354 0 dm2 AREA=1.244e-06
D7354 n7355 0 dm2 AREA=5.011e-07
D7355 n7356 0 dm2 AREA=4.776e-07
D7356 n7357 0 dm2 AREA=9.031e-07
D7357 n7358 0 dm2 AREA=3.016e-07
D7358 n1 0 dm2 AREA=1.692e-06
D7359 n7360 0 dm2 AREA=3.038e-07
D7360 n7361 0 dm2 AREA=1.520e-06
D7361 n7362 0 dm2 AREA=5.084e-07
D7362 n7363 0 dm2 AREA=1.454e-06
D7363 n7364 0 dm2 AREA=1.436e-06
D7364 n7365 0 dm2 AREA=1.165e-06
D7365 n7366 0 dm2 AREA=4.343e-07
D7366 n7367 0 dm2 AREA=8.132e-07
D7367 n7368 0 dm2 AREA=6.955e-07
D7368 n7369 0 dm2 AREA=9.732e-07
D7369 n7370 0 dm2 AREA=1.566e-06
D7370 n7371 0 dm2 AREA=1.732e-06
D7371 n7372 0 dm2 AREA=7.832e-07
D7372 n7373 0 dm2 AREA=2.188e-07
D7373 n7374 0 dm2 AREA=1.016e-06
D7374 n7375 0 dm2 AREA=8.235e-07
D7375 n7376 0 dm2 AREA=5.771e-07
D7376 n7377 0 dm2 AREA=6.190e-07
D7377 n7378 0 dm2 AREA=1.513e-06
D7378 n7379 0 dm2 AREA=8.198e-07
D7379 n7380 0 dm2 AREA=1.421e-06
D7380 n7381 0 dm2 AREA=1.052e-06
D7381 n7382 0 dm2 AREA=1.065e-06
D7382 n7383 0 dm2 AREA=1.871e-06
D7383 n7384 0 dm2 AREA=8.737e-07
D7384 n7385 0 dm2 AREA=8.845e-07
D7385 n7386 0 dm2 AREA=5.056e-07
D7386 n7387 0 dm2 AREA=1.211e-06
D7387 n7388 0 dm2 AREA=4.795e-07
D7388 n7389 0 dm2 AREA=5.676e-07
D7389 n7390 0 dm2 AREA=2.304e-06
D7390 n7391 0 dm2 AREA=1.222e-06
D7391 n7392 0 dm2 AREA=1.118e-06
D7392 n7393 0 dm2 AREA=2.474e-07
D7393 n7394 0 dm2 AREA=3.583e-07
D7394 n7395 0 dm2 AREA=1.240e-06
D7395 n7396 0 dm2 AREA=7.290e-07
D7396 n7397 0 dm2 AREA=1.382e-06
D7397 n7398 0 dm2 AREA=1.176e-06
D7398 n7399 0 dm2 AREA=6.219e-07
D7399 n7400 0 dm2 AREA=1.348e-06
D7400 n7401 0 dm2 AREA=1.185e-06
D7401 n7402 0 dm2 AREA=9.452e-07
D7402 n7403 0 dm2 AREA=1.178e-06
D7403 n7404 0 dm2 AREA=2.067e-06
D7404 n7405 0 dm2 AREA=8.935e-07
D7405 n7406 0 dm2 AREA=1.506e-06
D7406 n7407 0 dm2 AREA=9.980e-07
D7407 n7408 0 dm2 AREA=4.620e-07
D7408 n7409 0 dm2 AREA=1.189e-06
D7409 n7410 0 dm2 AREA=5.474e-07
D7410 n7411 0 dm2 AREA=5.839e-07
D7411 n7412 0 dm2 AREA=4.622e-07
D7412 n7413 0 dm2 AREA=7.976e-07
D7413 n7414 0 dm2 AREA=9.684e-07
D7414 n7415 0 dm2 AREA=8.500e-07
D7415 n7416 0 dm2 AREA=1.001e-06
D7416 n7417 0 dm2 AREA=1.287e-06
D7417 n7418 0 dm2 AREA=7.768e-07
D7418 n7419 0 dm2 AREA=1.273e-06
D7419 n7420 0 dm2 AREA=9.609e-07
D7420 n7421 0 dm2 AREA=3.158e-07
D7421 n7422 0 dm2 AREA=3.483e-07
D7422 n7423 0 dm2 AREA=4.498e-07
D7423 n7424 0 dm2 AREA=1.500e-06
D7424 n7425 0 dm2 AREA=1.452e-06
D7425 n7426 0 dm2 AREA=1.680e-06
D7426 n7427 0 dm2 AREA=2.822e-07
D7427 n7428 0 dm2 AREA=6.494e-07
D7428 n7429 0 dm2 AREA=3.633e-07
D7429 n7430 0 dm2 AREA=2.643e-06
D7430 n7431 0 dm2 AREA=9.018e-07
D7431 n7432 0 dm2 AREA=7.036e-07
D7432 n7433 0 dm2 AREA=1.018e-06
D7433 n7434 0 dm2 AREA=6.292e-07
D7434 n7435 0 dm2 AREA=7.245e-07
D7435 n7436 0 dm2 AREA=1.430e-06
D7436 n7437 0 dm2 AREA=7.339e-07
D7437 n7438 0 dm2 AREA=6.708e-07
D7438 n7439 0 dm2 AREA=4.812e-07
D7439 n7440 0 dm2 AREA=1.634e-06
D7440 n7441 0 dm2 AREA=1.640e-06
D7441 n7442 0 dm2 AREA=6.083e-07
D7442 n7443 0 dm2 AREA=4.836e-07
D7443 n7444 0 dm2 AREA=5.349e-07
D7444 n7445 0 dm2 AREA=9.998e-07
D7445 n7446 0 dm2 AREA=2.013e-06
D7446 n7447 0 dm2 AREA=8.874e-07
D7447 n7448 0 dm2 AREA=2.197e-06
D7448 n7449 0 dm2 AREA=2.239e-06
D7449 n7450 0 dm2 AREA=9.020e-07
D7450 n7451 0 dm2 AREA=8.751e-07
D7451 n7452 0 dm2 AREA=1.687e-06
D7452 n7453 0 dm2 AREA=4.882e-07
D7453 n7454 0 dm2 AREA=1.472e-06
D7454 n7455 0 dm2 AREA=7.809e-07
D7455 n7456 0 dm2 AREA=1.658e-06
D7456 n7457 0 dm2 AREA=5.311e-07
D7457 n7458 0 dm2 AREA=8.339e-07
D7458 n7459 0 dm2 AREA=7.621e-07
D7459 n7460 0 dm2 AREA=7.168e-07
D7460 n7461 0 dm2 AREA=4.730e-07
D7461 n7462 0 dm2 AREA=1.337e-06
D7462 n7463 0 dm2 AREA=1.249e-06
D7463 n7464 0 dm2 AREA=1.161e-06
D7464 n7465 0 dm2 AREA=2.178e-06
D7465 n7466 0 dm2 AREA=7.020e-07
D7466 n7467 0 dm2 AREA=7.818e-07
D7467 n7468 0 dm2 AREA=1.127e-06
D7468 n7469 0 dm2 AREA=1.060e-06
D7469 n7470 0 dm2 AREA=5.639e-07
D7470 n7471 0 dm2 AREA=7.437e-07
D7471 n7472 0 dm2 AREA=8.445e-07
D7472 n7473 0 dm2 AREA=1.233e-06
D7473 n7474 0 dm2 AREA=1.093e-06
D7474 n7475 0 dm2 AREA=6.380e-07
D7475 n7476 0 dm2 AREA=5.688e-07
D7476 n7477 0 dm2 AREA=7.709e-07
D7477 n7478 0 dm2 AREA=1.573e-06
D7478 n7479 0 dm2 AREA=1.461e-06
D7479 n7480 0 dm2 AREA=8.074e-07
D7480 n7481 0 dm2 AREA=9.682e-07
D7481 n7482 0 dm2 AREA=8.159e-07
D7482 n7483 0 dm2 AREA=9.980e-07
D7483 n7484 0 dm2 AREA=1.150e-06
D7484 n7485 0 dm2 AREA=5.322e-07
D7485 n7486 0 dm2 AREA=8.742e-07
D7486 n7487 0 dm2 AREA=8.402e-07
D7487 n7488 0 dm2 AREA=1.196e-06
D7488 n7489 0 dm2 AREA=8.114e-07
D7489 n7490 0 dm2 AREA=1.231e-06
D7490 n7491 0 dm2 AREA=5.834e-07
D7491 n7492 0 dm2 AREA=3.995e-07
D7492 n7493 0 dm2 AREA=1.013e-06
D7493 n7494 0 dm2 AREA=1.430e-06
D7494 n7495 0 dm2 AREA=8.803e-07
D7495 n7496 0 dm2 AREA=1.011e-06
D7496 n7497 0 dm2 AREA=9.533e-07
D7497 n7498 0 dm2 AREA=1.042e-06
D7498 n7499 0 dm2 AREA=1.331e-06
D7499 n7500 0 dm2 AREA=5.227e-07
D7500 n7501 0 dm2 AREA=1.380e-06
D7501 n7502 0 dm2 AREA=4.645e-07
D7502 n7503 0 dm2 AREA=1.558e-06
D7503 n7504 0 dm2 AREA=4.918e-07
D7504 n7505 0 dm2 AREA=1.587e-06
D7505 n7506 0 dm2 AREA=1.501e-06
D7506 n7507 0 dm2 AREA=4.070e-07
D7507 n7508 0 dm2 AREA=1.098e-06
D7508 n7509 0 dm2 AREA=7.549e-07
D7509 n7510 0 dm2 AREA=1.974e-06
D7510 n7511 0 dm2 AREA=1.581e-06
D7511 n7512 0 dm2 AREA=7.516e-07
D7512 n7513 0 dm2 AREA=1.538e-07
D7513 n7514 0 dm2 AREA=1.302e-06
D7514 n1 0 dm2 AREA=5.050e-07
D7515 n7516 0 dm2 AREA=8.181e-07
D7516 n7517 0 dm2 AREA=4.546e-07
D7517 n7518 0 dm2 AREA=1.881e-06
D7518 n7519 0 dm2 AREA=4.569e-07
D7519 n7520 0 dm2 AREA=1.151e-06
D7520 n7521 0 dm2 AREA=3.993e-07
D7521 n7522 0 dm2 AREA=1.542e-06
D7522 n7523 0 dm2 AREA=8.970e-07
D7523 n7524 0 dm2 AREA=1.708e-06
D7524 n7525 0 dm2 AREA=9.065e-07
D7525 n7526 0 dm2 AREA=6.486e-07
D7526 n7527 0 dm2 AREA=1.114e-06
D7527 n7528 0 dm2 AREA=8.716e-07
D7528 n7529 0 dm2 AREA=9.988e-07
D7529 n7530 0 dm2 AREA=4.090e-07
D7530 n7531 0 dm2 AREA=1.074e-06
D7531 n7532 0 dm2 AREA=5.143e-07
D7532 n7533 0 dm2 AREA=7.824e-07
D7533 n7534 0 dm2 AREA=8.239e-07
D7534 n7535 0 dm2 AREA=1.250e-06
D7535 n7536 0 dm2 AREA=8.255e-07
D7536 n7537 0 dm2 AREA=1.160e-06
D7537 n7538 0 dm2 AREA=8.257e-07
D7538 n7539 0 dm2 AREA=1.288e-06
D7539 n7540 0 dm2 AREA=4.684e-07
D7540 n7541 0 dm2 AREA=9.200e-07
D7541 n7542 0 dm2 AREA=1.405e-06
D7542 n7543 0 dm2 AREA=9.789e-07
D7543 n7544 0 dm2 AREA=1.065e-06
D7544 n7545 0 dm2 AREA=7.058e-07
D7545 n7546 0 dm2 AREA=4.744e-07
D7546 n7547 0 dm2 AREA=4.388e-07
D7547 n7548 0 dm2 AREA=1.015e-06
D7548 n7549 0 dm2 AREA=4.453e-07
D7549 n7550 0 dm2 AREA=1.055e-06
D7550 n7551 0 dm2 AREA=1.123e-06
D7551 n7552 0 dm2 AREA=1.034e-06
D7552 n7553 0 dm2 AREA=9.519e-07
D7553 n7554 0 dm2 AREA=5.281e-07
D7554 n7555 0 dm2 AREA=6.285e-07
D7555 n7556 0 dm2 AREA=7.180e-07
D7556 n7557 0 dm2 AREA=4.330e-07
D7557 n7558 0 dm2 AREA=7.274e-07
D7558 n7559 0 dm2 AREA=9.633e-07
D7559 n7560 0 dm2 AREA=8.713e-07
D7560 n7561 0 dm2 AREA=5.816e-07
D7561 n7562 0 dm2 AREA=6.193e-07
D7562 n7563 0 dm2 AREA=8.196e-07
D7563 n7564 0 dm2 AREA=6.384e-07
D7564 n7565 0 dm2 AREA=9.597e-07
D7565 n7566 0 dm2 AREA=1.050e-06
D7566 n7567 0 dm2 AREA=5.685e-07
D7567 n7568 0 dm2 AREA=6.428e-07
D7568 n7569 0 dm2 AREA=4.103e-07
D7569 n7570 0 dm2 AREA=2.550e-07
D7570 n7571 0 dm2 AREA=8.835e-07
D7571 n7572 0 dm2 AREA=3.101e-07
D7572 n7573 0 dm2 AREA=2.855e-06
D7573 n7574 0 dm2 AREA=7.585e-07
D7574 n7575 0 dm2 AREA=8.891e-07
D7575 n7576 0 dm2 AREA=9.909e-07
D7576 n7577 0 dm2 AREA=7.193e-07
D7577 n7578 0 dm2 AREA=1.138e-06
D7578 n7579 0 dm2 AREA=1.218e-06
D7579 n7580 0 dm2 AREA=1.008e-06
D7580 n7581 0 dm2 AREA=1.334e-06
D7581 n7582 0 dm2 AREA=9.243e-07
D7582 n7583 0 dm2 AREA=3.699e-07
D7583 n7584 0 dm2 AREA=1.244e-06
D7584 n7585 0 dm2 AREA=1.415e-06
D7585 n7586 0 dm2 AREA=3.853e-07
D7586 n7587 0 dm2 AREA=1.441e-07
D7587 n7588 0 dm2 AREA=3.244e-07
D7588 n7589 0 dm2 AREA=5.230e-07
D7589 n7590 0 dm2 AREA=1.142e-06
D7590 n7591 0 dm2 AREA=5.125e-07
D7591 n7592 0 dm2 AREA=4.832e-07
D7592 n7593 0 dm2 AREA=9.224e-07
D7593 n7594 0 dm2 AREA=1.149e-06
D7594 n7595 0 dm2 AREA=5.284e-07
D7595 n7596 0 dm2 AREA=9.653e-07
D7596 n7597 0 dm2 AREA=1.588e-06
D7597 n7598 0 dm2 AREA=1.690e-06
D7598 n7599 0 dm2 AREA=2.368e-06
D7599 n7600 0 dm2 AREA=2.529e-06
D7600 n7601 0 dm2 AREA=3.046e-07
D7601 n7602 0 dm2 AREA=1.235e-06
D7602 n7603 0 dm2 AREA=1.116e-06
D7603 n7604 0 dm2 AREA=4.206e-07
D7604 n7605 0 dm2 AREA=2.353e-06
D7605 n7606 0 dm2 AREA=7.541e-07
D7606 n7607 0 dm2 AREA=1.275e-06
D7607 n7608 0 dm2 AREA=3.515e-07
D7608 n7609 0 dm2 AREA=7.981e-07
D7609 n7610 0 dm2 AREA=9.713e-07
D7610 n7611 0 dm2 AREA=5.022e-07
D7611 n7612 0 dm2 AREA=1.307e-06
D7612 n7613 0 dm2 AREA=1.086e-06
D7613 n7614 0 dm2 AREA=6.084e-07
D7614 n7615 0 dm2 AREA=9.227e-07
D7615 n7616 0 dm2 AREA=1.991e-06
D7616 n7617 0 dm2 AREA=1.260e-06
D7617 n7618 0 dm2 AREA=1.329e-06
D7618 n7619 0 dm2 AREA=8.535e-07
D7619 n7620 0 dm2 AREA=6.375e-07
D7620 n7621 0 dm2 AREA=2.284e-06
D7621 n7622 0 dm2 AREA=9.747e-07
D7622 n7623 0 dm2 AREA=3.618e-07
D7623 n7624 0 dm2 AREA=8.435e-07
D7624 n7625 0 dm2 AREA=1.628e-06
D7625 n7626 0 dm2 AREA=1.243e-06
D7626 n7627 0 dm2 AREA=1.376e-06
D7627 n7628 0 dm2 AREA=5.981e-07
D7628 n7629 0 dm2 AREA=1.293e-06
D7629 n7630 0 dm2 AREA=5.411e-07
D7630 n7631 0 dm2 AREA=1.370e-06
D7631 n7632 0 dm2 AREA=1.120e-06
D7632 n7633 0 dm2 AREA=2.084e-06
D7633 n7634 0 dm2 AREA=1.301e-06
D7634 n7635 0 dm2 AREA=1.825e-06
D7635 n7636 0 dm2 AREA=5.383e-07
D7636 n7637 0 dm2 AREA=5.546e-07
D7637 n7638 0 dm2 AREA=8.041e-07
D7638 n7639 0 dm2 AREA=1.294e-06
D7639 n7640 0 dm2 AREA=1.198e-06
D7640 n7641 0 dm2 AREA=8.128e-07
D7641 n7642 0 dm2 AREA=6.032e-07
D7642 n7643 0 dm2 AREA=5.510e-07
D7643 n7644 0 dm2 AREA=8.744e-07
D7644 n7645 0 dm2 AREA=4.911e-07
D7645 n7646 0 dm2 AREA=1.027e-06
D7646 n7647 0 dm2 AREA=5.796e-07
D7647 n7648 0 dm2 AREA=1.100e-06
D7648 n7649 0 dm2 AREA=6.398e-07
D7649 n7650 0 dm2 AREA=8.292e-07
D7650 n7651 0 dm2 AREA=1.153e-06
D7651 n7652 0 dm2 AREA=1.152e-06
D7652 n7653 0 dm2 AREA=5.723e-07
D7653 n7654 0 dm2 AREA=2.241e-06
D7654 n7655 0 dm2 AREA=1.248e-06
D7655 n7656 0 dm2 AREA=3.017e-07
D7656 n1 0 dm2 AREA=6.673e-07
D7657 n7658 0 dm2 AREA=1.191e-07
D7658 n7659 0 dm2 AREA=1.161e-06
D7659 n7660 0 dm2 AREA=1.148e-06
D7660 n7661 0 dm2 AREA=2.136e-06
D7661 n7662 0 dm2 AREA=1.077e-06
D7662 n1 0 dm2 AREA=5.576e-07
D7663 n7664 0 dm2 AREA=6.536e-07
D7664 n7665 0 dm2 AREA=8.484e-07
D7665 n1 0 dm2 AREA=9.278e-07
D7666 n7667 0 dm2 AREA=1.564e-06
D7667 n7668 0 dm2 AREA=1.658e-06
D7668 n7669 0 dm2 AREA=4.194e-07
D7669 n7670 0 dm2 AREA=3.392e-07
D7670 n7671 0 dm2 AREA=1.062e-06
D7671 n1 0 dm2 AREA=3.988e-07
D7672 n7673 0 dm2 AREA=3.969e-07
D7673 n7674 0 dm2 AREA=1.123e-06
D7674 n7675 0 dm2 AREA=7.594e-07
D7675 n7676 0 dm2 AREA=5.601e-07
D7676 n7677 0 dm2 AREA=5.698e-07
D7677 n7678 0 dm2 AREA=6.344e-07
D7678 n7679 0 dm2 AREA=4.000e-07
D7679 n7680 0 dm2 AREA=5.852e-07
D7680 n7681 0 dm2 AREA=1.139e-06
D7681 n7682 0 dm2 AREA=8.674e-07
D7682 n7683 0 dm2 AREA=9.235e-07
D7683 n7684 0 dm2 AREA=7.192e-07
D7684 n7685 0 dm2 AREA=9.047e-07
D7685 n7686 0 dm2 AREA=1.986e-06
D7686 n7687 0 dm2 AREA=1.550e-06
D7687 n7688 0 dm2 AREA=1.161e-06
D7688 n7689 0 dm2 AREA=2.423e-07
D7689 n7690 0 dm2 AREA=1.869e-07
D7690 n7691 0 dm2 AREA=3.734e-07
D7691 n7692 0 dm2 AREA=9.912e-07
D7692 n7693 0 dm2 AREA=8.905e-07
D7693 n7694 0 dm2 AREA=3.963e-07
D7694 n7695 0 dm2 AREA=7.328e-07
D7695 n7696 0 dm2 AREA=6.905e-07
D7696 n7697 0 dm2 AREA=2.717e-07
D7697 n7698 0 dm2 AREA=2.036e-06
D7698 n7699 0 dm2 AREA=1.102e-06
D7699 n7700 0 dm2 AREA=8.297e-07
D7700 n7701 0 dm2 AREA=1.173e-06
D7701 n7702 0 dm2 AREA=8.486e-07
D7702 n7703 0 dm2 AREA=5.647e-07
D7703 n7704 0 dm2 AREA=9.189e-07
D7704 n7705 0 dm2 AREA=1.018e-06
D7705 n7706 0 dm2 AREA=7.757e-07
D7706 n7707 0 dm2 AREA=1.190e-06
D7707 n7708 0 dm2 AREA=9.113e-07
D7708 n7709 0 dm2 AREA=1.876e-06
D7709 n7710 0 dm2 AREA=9.122e-07
D7710 n7711 0 dm2 AREA=1.709e-06
D7711 n7712 0 dm2 AREA=6.687e-07
D7712 n7713 0 dm2 AREA=1.410e-06
D7713 n7714 0 dm2 AREA=9.542e-07
D7714 n7715 0 dm2 AREA=9.616e-07
D7715 n7716 0 dm2 AREA=1.284e-06
D7716 n7717 0 dm2 AREA=1.608e-06
D7717 n7718 0 dm2 AREA=4.990e-07
D7718 n7719 0 dm2 AREA=7.244e-07
D7719 n7720 0 dm2 AREA=4.080e-07
D7720 n7721 0 dm2 AREA=5.511e-07
D7721 n7722 0 dm2 AREA=1.248e-06
D7722 n7723 0 dm2 AREA=3.098e-06
D7723 n7724 0 dm2 AREA=1.420e-06
D7724 n7725 0 dm2 AREA=1.398e-06
D7725 n7726 0 dm2 AREA=1.102e-06
D7726 n7727 0 dm2 AREA=5.744e-07
D7727 n7728 0 dm2 AREA=6.643e-07
D7728 n7729 0 dm2 AREA=5.972e-07
D7729 n7730 0 dm2 AREA=6.957e-08
D7730 n7731 0 dm2 AREA=3.259e-07
D7731 n7732 0 dm2 AREA=7.692e-07
D7732 n7733 0 dm2 AREA=8.632e-07
D7733 n7734 0 dm2 AREA=5.618e-07
D7734 n7735 0 dm2 AREA=2.131e-06
D7735 n7736 0 dm2 AREA=1.578e-06
D7736 n7737 0 dm2 AREA=2.757e-06
D7737 n7738 0 dm2 AREA=1.321e-06
D7738 n7739 0 dm2 AREA=4.567e-07
D7739 n7740 0 dm2 AREA=1.119e-06
D7740 n7741 0 dm2 AREA=8.131e-07
D7741 n7742 0 dm2 AREA=9.904e-07
D7742 n7743 0 dm2 AREA=7.914e-07
D7743 n7744 0 dm2 AREA=1.510e-06
D7744 n7745 0 dm2 AREA=2.207e-06
D7745 n7746 0 dm2 AREA=1.075e-06
D7746 n7747 0 dm2 AREA=4.896e-07
D7747 n7748 0 dm2 AREA=6.865e-07
D7748 n7749 0 dm2 AREA=1.022e-06
D7749 n7750 0 dm2 AREA=1.056e-06
D7750 n7751 0 dm2 AREA=9.825e-07
D7751 n7752 0 dm2 AREA=7.903e-07
D7752 n7753 0 dm2 AREA=1.655e-06
D7753 n7754 0 dm2 AREA=6.858e-07
D7754 n7755 0 dm2 AREA=1.032e-06
D7755 n7756 0 dm2 AREA=1.168e-06
D7756 n7757 0 dm2 AREA=1.116e-06
D7757 n7758 0 dm2 AREA=1.233e-06
D7758 n7759 0 dm2 AREA=9.662e-07
D7759 n7760 0 dm2 AREA=1.747e-06
D7760 n7761 0 dm2 AREA=4.529e-07
D7761 n7762 0 dm2 AREA=5.438e-07
D7762 n7763 0 dm2 AREA=1.332e-06
D7763 n7764 0 dm2 AREA=1.677e-06
D7764 n7765 0 dm2 AREA=1.824e-06
D7765 n7766 0 dm2 AREA=9.977e-07
D7766 n7767 0 dm2 AREA=5.362e-07
D7767 n7768 0 dm2 AREA=2.457e-07
D7768 n7769 0 dm2 AREA=1.338e-06
D7769 n7770 0 dm2 AREA=3.461e-07
D7770 n7771 0 dm2 AREA=1.604e-06
D7771 n7772 0 dm2 AREA=7.745e-07
D7772 n7773 0 dm2 AREA=2.735e-07
D7773 n7774 0 dm2 AREA=4.038e-07
D7774 n7775 0 dm2 AREA=1.496e-06
D7775 n7776 0 dm2 AREA=1.007e-06
D7776 n7777 0 dm2 AREA=2.166e-06
D7777 n7778 0 dm2 AREA=1.465e-06
D7778 n7779 0 dm2 AREA=4.061e-07
D7779 n7780 0 dm2 AREA=9.804e-07
D7780 n7781 0 dm2 AREA=5.059e-07
D7781 n7782 0 dm2 AREA=6.154e-07
D7782 n7783 0 dm2 AREA=1.198e-06
D7783 n7784 0 dm2 AREA=4.736e-07
D7784 n7785 0 dm2 AREA=1.245e-06
D7785 n7786 0 dm2 AREA=1.445e-06
D7786 n7787 0 dm2 AREA=1.805e-06
D7787 n7788 0 dm2 AREA=8.905e-07
D7788 n7789 0 dm2 AREA=2.219e-06
D7789 n7790 0 dm2 AREA=3.115e-07
D7790 n7791 0 dm2 AREA=1.522e-07
D7791 n7792 0 dm2 AREA=5.349e-07
D7792 n7793 0 dm2 AREA=1.264e-06
D7793 n7794 0 dm2 AREA=2.118e-07
D7794 n7795 0 dm2 AREA=5.231e-07
D7795 n7796 0 dm2 AREA=1.114e-06
D7796 n7797 0 dm2 AREA=1.902e-06
D7797 n7798 0 dm2 AREA=1.775e-06
D7798 n7799 0 dm2 AREA=1.234e-06
D7799 n7800 0 dm2 AREA=3.007e-07
D7800 n7801 0 dm2 AREA=1.255e-06
D7801 n7802 0 dm2 AREA=1.212e-06
D7802 n7803 0 dm2 AREA=5.286e-07
D7803 n7804 0 dm2 AREA=8.566e-07
D7804 n7805 0 dm2 AREA=9.838e-07
D7805 n7806 0 dm2 AREA=1.911e-06
D7806 n1 0 dm2 AREA=3.627e-07
D7807 n7808 0 dm2 AREA=2.222e-06
D7808 n7809 0 dm2 AREA=4.761e-07
D7809 n7810 0 dm2 AREA=1.605e-06
D7810 n7811 0 dm2 AREA=1.464e-06
D7811 n7812 0 dm2 AREA=7.727e-07
D7812 n7813 0 dm2 AREA=9.829e-07
D7813 n7814 0 dm2 AREA=9.861e-07
D7814 n7815 0 dm2 AREA=3.563e-07
D7815 n7816 0 dm2 AREA=4.682e-07
D7816 n7817 0 dm2 AREA=8.995e-07
D7817 n7818 0 dm2 AREA=2.375e-07
D7818 n7819 0 dm2 AREA=6.766e-07
D7819 n7820 0 dm2 AREA=1.255e-06
D7820 n7821 0 dm2 AREA=4.247e-07
D7821 n7822 0 dm2 AREA=8.593e-07
D7822 n7823 0 dm2 AREA=6.122e-07
D7823 n7824 0 dm2 AREA=4.446e-07
D7824 n7825 0 dm2 AREA=1.516e-06
D7825 n1 0 dm2 AREA=5.610e-07
D7826 n7827 0 dm2 AREA=6.663e-07
D7827 n7828 0 dm2 AREA=1.358e-06
D7828 n7829 0 dm2 AREA=9.265e-07
D7829 n7830 0 dm2 AREA=7.171e-07
D7830 n7831 0 dm2 AREA=1.474e-06
D7831 n7832 0 dm2 AREA=2.003e-06
D7832 n7833 0 dm2 AREA=1.158e-06
D7833 n7834 0 dm2 AREA=2.626e-07
D7834 n7835 0 dm2 AREA=4.736e-07
D7835 n7836 0 dm2 AREA=1.689e-06
D7836 n7837 0 dm2 AREA=2.022e-06
D7837 n7838 0 dm2 AREA=9.069e-07
D7838 n7839 0 dm2 AREA=6.343e-07
D7839 n7840 0 dm2 AREA=2.009e-06
D7840 n7841 0 dm2 AREA=4.397e-07
D7841 n7842 0 dm2 AREA=7.559e-07
D7842 n7843 0 dm2 AREA=1.029e-06
D7843 n7844 0 dm2 AREA=6.381e-07
D7844 n7845 0 dm2 AREA=9.299e-07
D7845 n7846 0 dm2 AREA=6.607e-07
D7846 n7847 0 dm2 AREA=4.663e-07
D7847 n7848 0 dm2 AREA=5.681e-07
D7848 n7849 0 dm2 AREA=2.536e-06
D7849 n7850 0 dm2 AREA=2.269e-06
D7850 n7851 0 dm2 AREA=8.052e-07
D7851 n7852 0 dm2 AREA=1.546e-06
D7852 n7853 0 dm2 AREA=1.190e-06
D7853 n7854 0 dm2 AREA=2.317e-06
D7854 n7855 0 dm2 AREA=1.431e-06
D7855 n7856 0 dm2 AREA=1.500e-06
D7856 n7857 0 dm2 AREA=4.210e-07
D7857 n7858 0 dm2 AREA=1.009e-06
D7858 n7859 0 dm2 AREA=7.930e-07
D7859 n7860 0 dm2 AREA=1.154e-06
D7860 n7861 0 dm2 AREA=6.969e-07
D7861 n7862 0 dm2 AREA=6.672e-07
D7862 n7863 0 dm2 AREA=6.432e-07
D7863 n7864 0 dm2 AREA=4.478e-07
D7864 n7865 0 dm2 AREA=9.490e-07
D7865 n7866 0 dm2 AREA=5.386e-07
D7866 n7867 0 dm2 AREA=6.077e-07
D7867 n7868 0 dm2 AREA=9.515e-07
D7868 n7869 0 dm2 AREA=1.336e-06
D7869 n7870 0 dm2 AREA=1.447e-06
D7870 n7871 0 dm2 AREA=1.179e-06
D7871 n7872 0 dm2 AREA=8.869e-07
D7872 n7873 0 dm2 AREA=1.165e-06
D7873 n7874 0 dm2 AREA=1.028e-06
D7874 n7875 0 dm2 AREA=4.669e-07
D7875 n7876 0 dm2 AREA=1.438e-06
D7876 n7877 0 dm2 AREA=1.075e-06
D7877 n7878 0 dm2 AREA=1.470e-06
D7878 n7879 0 dm2 AREA=8.046e-07
D7879 n7880 0 dm2 AREA=1.155e-06
D7880 n7881 0 dm2 AREA=3.630e-07
D7881 n7882 0 dm2 AREA=1.861e-06
D7882 n7883 0 dm2 AREA=9.297e-07
D7883 n7884 0 dm2 AREA=7.089e-07
D7884 n7885 0 dm2 AREA=9.986e-07
D7885 n7886 0 dm2 AREA=1.108e-06
D7886 n7887 0 dm2 AREA=5.536e-07
D7887 n7888 0 dm2 AREA=1.441e-06
D7888 n7889 0 dm2 AREA=5.300e-07
D7889 n7890 0 dm2 AREA=1.002e-06
D7890 n7891 0 dm2 AREA=9.058e-07
D7891 n7892 0 dm2 AREA=3.691e-07
D7892 n7893 0 dm2 AREA=5.531e-07
D7893 n7894 0 dm2 AREA=1.222e-06
D7894 n7895 0 dm2 AREA=8.421e-07
D7895 n7896 0 dm2 AREA=9.613e-07
D7896 n7897 0 dm2 AREA=1.683e-06
D7897 n7898 0 dm2 AREA=1.370e-06
D7898 n7899 0 dm2 AREA=6.829e-07
D7899 n7900 0 dm2 AREA=4.567e-07
D7900 n7901 0 dm2 AREA=1.348e-06
D7901 n7902 0 dm2 AREA=4.237e-07
D7902 n7903 0 dm2 AREA=1.029e-06
D7903 n7904 0 dm2 AREA=1.522e-06
D7904 n7905 0 dm2 AREA=7.412e-07
D7905 n7906 0 dm2 AREA=1.180e-06
D7906 n7907 0 dm2 AREA=4.152e-07
D7907 n7908 0 dm2 AREA=1.478e-06
D7908 n7909 0 dm2 AREA=1.183e-06
D7909 n7910 0 dm2 AREA=1.408e-06
D7910 n7911 0 dm2 AREA=6.143e-07
D7911 n7912 0 dm2 AREA=9.944e-07
D7912 n7913 0 dm2 AREA=1.053e-06
D7913 n7914 0 dm2 AREA=9.484e-07
D7914 n7915 0 dm2 AREA=1.206e-06
D7915 n7916 0 dm2 AREA=2.851e-08
D7916 n7917 0 dm2 AREA=8.234e-07
D7917 n7918 0 dm2 AREA=1.207e-06
D7918 n7919 0 dm2 AREA=3.484e-07
D7919 n7920 0 dm2 AREA=6.511e-07
D7920 n7921 0 dm2 AREA=7.537e-07
D7921 n7922 0 dm2 AREA=1.576e-06
D7922 n7923 0 dm2 AREA=5.858e-07
D7923 n7924 0 dm2 AREA=2.099e-06
D7924 n7925 0 dm2 AREA=1.148e-06
D7925 n7926 0 dm2 AREA=3.292e-07
D7926 n7927 0 dm2 AREA=9.641e-07
D7927 n7928 0 dm2 AREA=8.302e-07
D7928 n7929 0 dm2 AREA=5.178e-07
D7929 n7930 0 dm2 AREA=1.034e-06
D7930 n7931 0 dm2 AREA=1.041e-06
D7931 n7932 0 dm2 AREA=5.863e-07
D7932 n7933 0 dm2 AREA=1.168e-06
D7933 n7934 0 dm2 AREA=1.028e-06
D7934 n7935 0 dm2 AREA=1.119e-06
D7935 n7936 0 dm2 AREA=9.933e-07
D7936 n7937 0 dm2 AREA=1.291e-06
D7937 n7938 0 dm2 AREA=1.902e-06
D7938 n1 0 dm2 AREA=8.455e-07
D7939 n7940 0 dm2 AREA=4.854e-07
D7940 n7941 0 dm2 AREA=7.771e-07
D7941 n7942 0 dm2 AREA=1.853e-07
D7942 n7943 0 dm2 AREA=4.712e-07
D7943 n7944 0 dm2 AREA=4.998e-07
D7944 n7945 0 dm2 AREA=1.876e-07
D7945 n7946 0 dm2 AREA=6.624e-07
D7946 n7947 0 dm2 AREA=1.038e-06
D7947 n7948 0 dm2 AREA=1.052e-06
D7948 n7949 0 dm2 AREA=1.082e-06
D7949 n7950 0 dm2 AREA=8.409e-07
D7950 n7951 0 dm2 AREA=1.255e-06
D7951 n7952 0 dm2 AREA=6.414e-07
D7952 n7953 0 dm2 AREA=5.953e-07
D7953 n7954 0 dm2 AREA=1.434e-06
D7954 n7955 0 dm2 AREA=4.020e-07
D7955 n7956 0 dm2 AREA=8.956e-07
D7956 n7957 0 dm2 AREA=8.795e-07
D7957 n7958 0 dm2 AREA=6.071e-07
D7958 n7959 0 dm2 AREA=1.215e-06
D7959 n7960 0 dm2 AREA=9.190e-07
D7960 n7961 0 dm2 AREA=8.318e-07
D7961 n7962 0 dm2 AREA=6.217e-07
D7962 n7963 0 dm2 AREA=8.332e-07
D7963 n7964 0 dm2 AREA=6.619e-07
D7964 n7965 0 dm2 AREA=3.967e-07
D7965 n7966 0 dm2 AREA=1.776e-06
D7966 n7967 0 dm2 AREA=5.473e-07
D7967 n7968 0 dm2 AREA=1.459e-06
D7968 n7969 0 dm2 AREA=1.249e-06
D7969 n7970 0 dm2 AREA=7.431e-07
D7970 n7971 0 dm2 AREA=4.115e-07
D7971 n7972 0 dm2 AREA=3.317e-07
D7972 n7973 0 dm2 AREA=1.122e-06
D7973 n7974 0 dm2 AREA=1.035e-06
D7974 n7975 0 dm2 AREA=6.196e-07
D7975 n7976 0 dm2 AREA=1.062e-06
D7976 n7977 0 dm2 AREA=1.007e-06
D7977 n7978 0 dm2 AREA=6.824e-07
D7978 n7979 0 dm2 AREA=4.080e-07
D7979 n7980 0 dm2 AREA=4.399e-07
D7980 n7981 0 dm2 AREA=1.112e-06
D7981 n7982 0 dm2 AREA=6.414e-07
D7982 n7983 0 dm2 AREA=1.472e-06
D7983 n7984 0 dm2 AREA=4.651e-07
D7984 n7985 0 dm2 AREA=5.185e-07
D7985 n7986 0 dm2 AREA=2.676e-07
D7986 n7987 0 dm2 AREA=3.398e-07
D7987 n7988 0 dm2 AREA=8.779e-07
D7988 n7989 0 dm2 AREA=7.090e-07
D7989 n7990 0 dm2 AREA=1.219e-06
D7990 n7991 0 dm2 AREA=1.244e-06
D7991 n7992 0 dm2 AREA=6.295e-07
D7992 n7993 0 dm2 AREA=8.855e-07
D7993 n7994 0 dm2 AREA=1.120e-06
D7994 n7995 0 dm2 AREA=5.021e-07
D7995 n7996 0 dm2 AREA=6.254e-07
D7996 n7997 0 dm2 AREA=1.191e-06
D7997 n7998 0 dm2 AREA=5.113e-07
D7998 n7999 0 dm2 AREA=1.622e-06
D7999 n8000 0 dm2 AREA=7.915e-07
D8000 n8001 0 dm2 AREA=4.627e-07
D8001 n8002 0 dm2 AREA=1.489e-06
D8002 n8003 0 dm2 AREA=1.173e-06
D8003 n8004 0 dm2 AREA=1.410e-06
D8004 n8005 0 dm2 AREA=6.948e-07
D8005 n8006 0 dm2 AREA=1.344e-06
D8006 n8007 0 dm2 AREA=3.262e-07
D8007 n8008 0 dm2 AREA=1.383e-06
D8008 n8009 0 dm2 AREA=1.623e-06
D8009 n8010 0 dm2 AREA=1.485e-06
D8010 n8011 0 dm2 AREA=5.388e-07
D8011 n8012 0 dm2 AREA=1.351e-06
D8012 n8013 0 dm2 AREA=1.350e-06
D8013 n8014 0 dm2 AREA=7.921e-07
D8014 n8015 0 dm2 AREA=4.867e-07
D8015 n8016 0 dm2 AREA=3.358e-07
D8016 n8017 0 dm2 AREA=1.300e-06
D8017 n8018 0 dm2 AREA=1.254e-06
D8018 n8019 0 dm2 AREA=7.777e-07
D8019 n8020 0 dm2 AREA=9.437e-07
D8020 n8021 0 dm2 AREA=6.240e-07
D8021 n8022 0 dm2 AREA=7.386e-07
D8022 n8023 0 dm2 AREA=1.213e-06
D8023 n8024 0 dm2 AREA=3.256e-07
D8024 n8025 0 dm2 AREA=1.201e-06
D8025 n8026 0 dm2 AREA=7.565e-07
D8026 n8027 0 dm2 AREA=2.179e-06
D8027 n8028 0 dm2 AREA=1.486e-06
D8028 n8029 0 dm2 AREA=2.182e-06
D8029 n8030 0 dm2 AREA=3.756e-07
D8030 n8031 0 dm2 AREA=1.009e-06
D8031 n8032 0 dm2 AREA=1.223e-06
D8032 n8033 0 dm2 AREA=4.855e-07
D8033 n8034 0 dm2 AREA=1.871e-06
D8034 n8035 0 dm2 AREA=1.497e-06
D8035 n8036 0 dm2 AREA=9.460e-07
D8036 n8037 0 dm2 AREA=1.566e-06
D8037 n8038 0 dm2 AREA=1.242e-06
D8038 n8039 0 dm2 AREA=3.360e-07
D8039 n8040 0 dm2 AREA=1.614e-06
D8040 n8041 0 dm2 AREA=8.769e-07
D8041 n8042 0 dm2 AREA=6.633e-07
D8042 n8043 0 dm2 AREA=7.020e-07
D8043 n8044 0 dm2 AREA=5.206e-07
D8044 n8045 0 dm2 AREA=1.167e-06
D8045 n8046 0 dm2 AREA=1.883e-06
D8046 n8047 0 dm2 AREA=4.481e-07
D8047 n8048 0 dm2 AREA=1.423e-06
D8048 n8049 0 dm2 AREA=9.216e-07
D8049 n8050 0 dm2 AREA=3.392e-07
D8050 n8051 0 dm2 AREA=1.533e-06
D8051 n8052 0 dm2 AREA=9.892e-07
D8052 n8053 0 dm2 AREA=1.238e-06
D8053 n8054 0 dm2 AREA=2.761e-07
D8054 n8055 0 dm2 AREA=9.362e-08
D8055 n8056 0 dm2 AREA=7.718e-07
D8056 n8057 0 dm2 AREA=1.331e-06
D8057 n8058 0 dm2 AREA=1.058e-06
D8058 n8059 0 dm2 AREA=1.064e-06
D8059 n8060 0 dm2 AREA=7.125e-07
D8060 n8061 0 dm2 AREA=8.303e-07
D8061 n8062 0 dm2 AREA=1.606e-06
D8062 n8063 0 dm2 AREA=5.895e-07
D8063 n8064 0 dm2 AREA=2.873e-07
D8064 n8065 0 dm2 AREA=4.793e-07
D8065 n8066 0 dm2 AREA=1.860e-06
D8066 n8067 0 dm2 AREA=9.930e-07
D8067 n8068 0 dm2 AREA=1.104e-06
D8068 n8069 0 dm2 AREA=7.210e-07
D8069 n8070 0 dm2 AREA=3.556e-07
D8070 n8071 0 dm2 AREA=2.005e-07
D8071 n8072 0 dm2 AREA=1.023e-06
D8072 n8073 0 dm2 AREA=4.102e-07
D8073 n8074 0 dm2 AREA=8.362e-07
D8074 n8075 0 dm2 AREA=8.057e-07
D8075 n8076 0 dm2 AREA=1.030e-06
D8076 n8077 0 dm2 AREA=8.188e-07
D8077 n8078 0 dm2 AREA=1.053e-06
D8078 n8079 0 dm2 AREA=1.648e-06
D8079 n8080 0 dm2 AREA=1.209e-06
D8080 n8081 0 dm2 AREA=1.597e-06
D8081 n8082 0 dm2 AREA=6.713e-07
D8082 n8083 0 dm2 AREA=1.366e-06
D8083 n8084 0 dm2 AREA=9.593e-07
D8084 n8085 0 dm2 AREA=7.823e-07
D8085 n8086 0 dm2 AREA=6.863e-07
D8086 n8087 0 dm2 AREA=1.430e-06
D8087 n8088 0 dm2 AREA=5.645e-07
D8088 n8089 0 dm2 AREA=2.105e-06
D8089 n8090 0 dm2 AREA=1.359e-06
D8090 n8091 0 dm2 AREA=1.475e-06
D8091 n8092 0 dm2 AREA=7.592e-07
D8092 n8093 0 dm2 AREA=8.607e-07
D8093 n8094 0 dm2 AREA=6.221e-07
D8094 n8095 0 dm2 AREA=1.683e-06
D8095 n8096 0 dm2 AREA=9.482e-07
D8096 n8097 0 dm2 AREA=1.499e-07
D8097 n8098 0 dm2 AREA=5.174e-07
D8098 n8099 0 dm2 AREA=3.083e-07
D8099 n8100 0 dm2 AREA=8.234e-07
D8100 n8101 0 dm2 AREA=1.549e-06
D8101 n8102 0 dm2 AREA=1.190e-06
D8102 n8103 0 dm2 AREA=7.780e-07
D8103 n8104 0 dm2 AREA=7.054e-07
D8104 n8105 0 dm2 AREA=7.703e-07
D8105 n8106 0 dm2 AREA=9.988e-07
D8106 n8107 0 dm2 AREA=5.761e-07
D8107 n8108 0 dm2 AREA=1.921e-06
D8108 n8109 0 dm2 AREA=9.327e-07
D8109 n8110 0 dm2 AREA=1.493e-06
D8110 n8111 0 dm2 AREA=9.993e-07
D8111 n8112 0 dm2 AREA=6.825e-07
D8112 n8113 0 dm2 AREA=6.481e-07
D8113 n8114 0 dm2 AREA=3.010e-07
D8114 n8115 0 dm2 AREA=1.539e-06
D8115 n8116 0 dm2 AREA=4.940e-07
D8116 n8117 0 dm2 AREA=1.732e-06
D8117 n8118 0 dm2 AREA=1.652e-06
D8118 n8119 0 dm2 AREA=1.002e-06
D8119 n8120 0 dm2 AREA=1.376e-06
D8120 n8121 0 dm2 AREA=1.812e-06
D8121 n8122 0 dm2 AREA=1.012e-06
D8122 n8123 0 dm2 AREA=4.968e-07
D8123 n8124 0 dm2 AREA=9.051e-07
D8124 n8125 0 dm2 AREA=6.042e-07
D8125 n8126 0 dm2 AREA=1.319e-06
D8126 n8127 0 dm2 AREA=1.109e-06
D8127 n8128 0 dm2 AREA=1.366e-06
D8128 n8129 0 dm2 AREA=1.278e-06
D8129 n8130 0 dm2 AREA=1.646e-06
D8130 n8131 0 dm2 AREA=3.926e-07
D8131 n8132 0 dm2 AREA=1.849e-07
D8132 n8133 0 dm2 AREA=5.811e-07
D8133 n8134 0 dm2 AREA=7.916e-07
D8134 n8135 0 dm2 AREA=7.805e-07
D8135 n8136 0 dm2 AREA=1.022e-06
D8136 n8137 0 dm2 AREA=3.020e-07
D8137 n8138 0 dm2 AREA=1.423e-06
D8138 n8139 0 dm2 AREA=7.098e-07
D8139 n8140 0 dm2 AREA=1.232e-06
D8140 n8141 0 dm2 AREA=9.960e-07
D8141 n8142 0 dm2 AREA=2.998e-07
D8142 n8143 0 dm2 AREA=1.152e-06
D8143 n8144 0 dm2 AREA=9.159e-07
D8144 n8145 0 dm2 AREA=5.629e-07
D8145 n8146 0 dm2 AREA=2.398e-07
D8146 n8147 0 dm2 AREA=1.397e-06
D8147 n8148 0 dm2 AREA=6.326e-07
D8148 n8149 0 dm2 AREA=8.175e-07
D8149 n8150 0 dm2 AREA=8.541e-07
D8150 n8151 0 dm2 AREA=9.879e-07
D8151 n8152 0 dm2 AREA=1.232e-06
D8152 n8153 0 dm2 AREA=2.055e-06
D8153 n8154 0 dm2 AREA=1.192e-06
D8154 n8155 0 dm2 AREA=1.217e-06
D8155 n8156 0 dm2 AREA=5.826e-07
D8156 n8157 0 dm2 AREA=1.226e-06
D8157 n8158 0 dm2 AREA=9.656e-07
D8158 n8159 0 dm2 AREA=1.122e-06
D8159 n8160 0 dm2 AREA=5.119e-07
D8160 n8161 0 dm2 AREA=8.551e-07
D8161 n8162 0 dm2 AREA=1.261e-06
D8162 n8163 0 dm2 AREA=3.068e-07
D8163 n8164 0 dm2 AREA=6.763e-07
D8164 n8165 0 dm2 AREA=6.280e-07
D8165 n8166 0 dm2 AREA=6.969e-07
D8166 n8167 0 dm2 AREA=1.924e-06
D8167 n8168 0 dm2 AREA=1.109e-07
D8168 n8169 0 dm2 AREA=1.057e-06
D8169 n8170 0 dm2 AREA=1.138e-06
D8170 n8171 0 dm2 AREA=1.380e-06
D8171 n8172 0 dm2 AREA=2.041e-07
D8172 n8173 0 dm2 AREA=8.880e-07
D8173 n8174 0 dm2 AREA=1.316e-06
D8174 n8175 0 dm2 AREA=9.538e-07
D8175 n8176 0 dm2 AREA=1.061e-06
D8176 n8177 0 dm2 AREA=1.092e-06
D8177 n8178 0 dm2 AREA=1.308e-06
D8178 n8179 0 dm2 AREA=5.974e-07
D8179 n8180 0 dm2 AREA=8.163e-07
D8180 n8181 0 dm2 AREA=5.807e-07
D8181 n8182 0 dm2 AREA=9.041e-07
D8182 n8183 0 dm2 AREA=1.577e-06
D8183 n8184 0 dm2 AREA=1.774e-06
D8184 n8185 0 dm2 AREA=4.401e-07
D8185 n8186 0 dm2 AREA=5.740e-07
D8186 n8187 0 dm2 AREA=1.697e-06
D8187 n8188 0 dm2 AREA=1.428e-06
D8188 n8189 0 dm2 AREA=9.402e-07
D8189 n8190 0 dm2 AREA=8.040e-07
D8190 n8191 0 dm2 AREA=3.503e-07
D8191 n8192 0 dm2 AREA=8.223e-07
D8192 n8193 0 dm2 AREA=5.379e-07
D8193 n8194 0 dm2 AREA=2.291e-06
D8194 n8195 0 dm2 AREA=3.980e-07
D8195 n8196 0 dm2 AREA=2.072e-06
D8196 n8197 0 dm2 AREA=4.762e-07
D8197 n8198 0 dm2 AREA=6.692e-07
D8198 n8199 0 dm2 AREA=1.039e-06
D8199 n8200 0 dm2 AREA=9.675e-07
D8200 n8201 0 dm2 AREA=4.992e-07
D8201 n8202 0 dm2 AREA=1.396e-06
D8202 n8203 0 dm2 AREA=2.398e-06
D8203 n8204 0 dm2 AREA=1.077e-06
D8204 n8205 0 dm2 AREA=6.006e-07
D8205 n8206 0 dm2 AREA=1.047e-06
D8206 n8207 0 dm2 AREA=1.601e-06
D8207 n8208 0 dm2 AREA=6.009e-07
D8208 n8209 0 dm2 AREA=2.195e-06
D8209 n8210 0 dm2 AREA=7.265e-07
D8210 n8211 0 dm2 AREA=2.782e-06
D8211 n8212 0 dm2 AREA=1.275e-06
D8212 n8213 0 dm2 AREA=4.230e-07
D8213 n8214 0 dm2 AREA=1.691e-06
D8214 n8215 0 dm2 AREA=7.046e-07
D8215 n8216 0 dm2 AREA=1.608e-06
D8216 n8217 0 dm2 AREA=1.866e-07
D8217 n8218 0 dm2 AREA=4.917e-08
D8218 n8219 0 dm2 AREA=5.441e-07
D8219 n8220 0 dm2 AREA=1.230e-06
D8220 n8221 0 dm2 AREA=2.032e-06
D8221 n8222 0 dm2 AREA=1.357e-06
D8222 n8223 0 dm2 AREA=7.357e-07
D8223 n8224 0 dm2 AREA=8.597e-07
D8224 n8225 0 dm2 AREA=8.222e-07
D8225 n8226 0 dm2 AREA=6.762e-07
D8226 n8227 0 dm2 AREA=6.390e-07
D8227 n8228 0 dm2 AREA=4.982e-07
D8228 n8229 0 dm2 AREA=4.149e-07
D8229 n8230 0 dm2 AREA=4.051e-07
D8230 n8231 0 dm2 AREA=1.072e-06
D8231 n8232 0 dm2 AREA=1.004e-06
D8232 n8233 0 dm2 AREA=2.312e-07
D8233 n8234 0 dm2 AREA=1.426e-06
D8234 n8235 0 dm2 AREA=8.799e-07
D8235 n8236 0 dm2 AREA=1.027e-06
D8236 n8237 0 dm2 AREA=1.091e-06
D8237 n8238 0 dm2 AREA=2.104e-06
D8238 n8239 0 dm2 AREA=9.711e-07
D8239 n8240 0 dm2 AREA=1.332e-06
D8240 n8241 0 dm2 AREA=5.763e-07
D8241 n8242 0 dm2 AREA=1.637e-06
D8242 n8243 0 dm2 AREA=9.211e-07
D8243 n8244 0 dm2 AREA=5.966e-07
D8244 n8245 0 dm2 AREA=1.446e-06
D8245 n8246 0 dm2 AREA=7.274e-07
D8246 n8247 0 dm2 AREA=5.752e-07
D8247 n8248 0 dm2 AREA=5.628e-07
D8248 n8249 0 dm2 AREA=1.776e-06
D8249 n8250 0 dm2 AREA=6.455e-07
D8250 n8251 0 dm2 AREA=2.080e-06
D8251 n8252 0 dm2 AREA=6.941e-07
D8252 n8253 0 dm2 AREA=6.554e-07
D8253 n8254 0 dm2 AREA=8.357e-07
D8254 n8255 0 dm2 AREA=7.659e-07
D8255 n8256 0 dm2 AREA=7.018e-07
D8256 n8257 0 dm2 AREA=1.717e-06
D8257 n8258 0 dm2 AREA=5.295e-07
D8258 n8259 0 dm2 AREA=2.127e-07
D8259 n8260 0 dm2 AREA=1.462e-06
D8260 n8261 0 dm2 AREA=1.221e-06
D8261 n8262 0 dm2 AREA=1.404e-07
D8262 n8263 0 dm2 AREA=1.779e-06
D8263 n8264 0 dm2 AREA=9.885e-07
D8264 n8265 0 dm2 AREA=5.906e-07
D8265 n8266 0 dm2 AREA=1.097e-06
D8266 n8267 0 dm2 AREA=2.135e-06
D8267 n8268 0 dm2 AREA=7.794e-07
D8268 n8269 0 dm2 AREA=2.273e-07
D8269 n8270 0 dm2 AREA=7.562e-07
D8270 n8271 0 dm2 AREA=1.009e-06
D8271 n8272 0 dm2 AREA=1.077e-06
D8272 n8273 0 dm2 AREA=1.897e-06
D8273 n8274 0 dm2 AREA=4.341e-07
D8274 n8275 0 dm2 AREA=1.435e-06
D8275 n8276 0 dm2 AREA=1.296e-06
D8276 n8277 0 dm2 AREA=8.529e-07
D8277 n8278 0 dm2 AREA=1.005e-06
D8278 n8279 0 dm2 AREA=1.847e-07
D8279 n8280 0 dm2 AREA=3.579e-07
D8280 n8281 0 dm2 AREA=8.749e-07
D8281 n8282 0 dm2 AREA=9.731e-07
D8282 n8283 0 dm2 AREA=1.260e-06
D8283 n8284 0 dm2 AREA=1.347e-06
D8284 n8285 0 dm2 AREA=6.752e-07
D8285 n8286 0 dm2 AREA=5.426e-07
D8286 n8287 0 dm2 AREA=9.413e-07
D8287 n8288 0 dm2 AREA=8.981e-07
D8288 n8289 0 dm2 AREA=5.531e-07
D8289 n8290 0 dm2 AREA=6.316e-07
D8290 n8291 0 dm2 AREA=9.583e-07
D8291 n8292 0 dm2 AREA=1.059e-06
D8292 n8293 0 dm2 AREA=1.306e-06
D8293 n8294 0 dm2 AREA=4.084e-07
D8294 n8295 0 dm2 AREA=7.025e-07
D8295 n8296 0 dm2 AREA=2.998e-06
D8296 n8297 0 dm2 AREA=9.305e-07
D8297 n8298 0 dm2 AREA=2.316e-07
D8298 n8299 0 dm2 AREA=1.640e-06
D8299 n8300 0 dm2 AREA=5.490e-07
D8300 n8301 0 dm2 AREA=1.508e-06
D8301 n8302 0 dm2 AREA=5.213e-07
D8302 n8303 0 dm2 AREA=5.682e-07
D8303 n8304 0 dm2 AREA=5.614e-07
D8304 n8305 0 dm2 AREA=1.520e-06
D8305 n8306 0 dm2 AREA=3.270e-07
D8306 n8307 0 dm2 AREA=1.247e-06
D8307 n8308 0 dm2 AREA=7.401e-07
D8308 n8309 0 dm2 AREA=8.496e-07
D8309 n8310 0 dm2 AREA=6.512e-07
D8310 n8311 0 dm2 AREA=4.617e-07
D8311 n8312 0 dm2 AREA=2.019e-06
D8312 n8313 0 dm2 AREA=7.104e-07
D8313 n8314 0 dm2 AREA=1.328e-06
D8314 n8315 0 dm2 AREA=4.541e-07
D8315 n8316 0 dm2 AREA=1.714e-06
D8316 n8317 0 dm2 AREA=8.444e-07
D8317 n8318 0 dm2 AREA=7.923e-07
D8318 n8319 0 dm2 AREA=7.954e-07
D8319 n8320 0 dm2 AREA=8.273e-07
D8320 n8321 0 dm2 AREA=1.487e-06
D8321 n8322 0 dm2 AREA=6.010e-07
D8322 n8323 0 dm2 AREA=1.705e-06
D8323 n8324 0 dm2 AREA=1.100e-06
D8324 n8325 0 dm2 AREA=6.657e-07
D8325 n8326 0 dm2 AREA=2.807e-06
D8326 n8327 0 dm2 AREA=8.329e-07
D8327 n8328 0 dm2 AREA=1.310e-06
D8328 n8329 0 dm2 AREA=8.375e-07
D8329 n8330 0 dm2 AREA=8.945e-07
D8330 n8331 0 dm2 AREA=9.520e-07
D8331 n8332 0 dm2 AREA=4.570e-07
D8332 n8333 0 dm2 AREA=1.328e-06
D8333 n8334 0 dm2 AREA=2.020e-06
D8334 n8335 0 dm2 AREA=1.295e-06
D8335 n1 0 dm2 AREA=7.580e-07
D8336 n8337 0 dm2 AREA=7.282e-07
D8337 n8338 0 dm2 AREA=5.484e-07
D8338 n8339 0 dm2 AREA=1.571e-06
D8339 n8340 0 dm2 AREA=3.353e-07
D8340 n8341 0 dm2 AREA=7.773e-07
D8341 n8342 0 dm2 AREA=2.163e-06
D8342 n8343 0 dm2 AREA=1.448e-06
D8343 n8344 0 dm2 AREA=1.218e-06
D8344 n8345 0 dm2 AREA=1.365e-06
D8345 n8346 0 dm2 AREA=7.695e-07
D8346 n8347 0 dm2 AREA=6.941e-07
D8347 n8348 0 dm2 AREA=1.470e-06
D8348 n8349 0 dm2 AREA=1.879e-06
D8349 n8350 0 dm2 AREA=4.187e-07
D8350 n8351 0 dm2 AREA=1.778e-06
D8351 n8352 0 dm2 AREA=1.124e-06
D8352 n8353 0 dm2 AREA=7.452e-07
D8353 n8354 0 dm2 AREA=1.626e-06
D8354 n8355 0 dm2 AREA=5.695e-07
D8355 n8356 0 dm2 AREA=1.031e-06
D8356 n8357 0 dm2 AREA=1.286e-06
D8357 n8358 0 dm2 AREA=5.097e-07
D8358 n8359 0 dm2 AREA=1.813e-06
D8359 n8360 0 dm2 AREA=8.388e-07
D8360 n8361 0 dm2 AREA=1.250e-06
D8361 n8362 0 dm2 AREA=1.158e-06
D8362 n8363 0 dm2 AREA=1.468e-06
D8363 n8364 0 dm2 AREA=9.459e-07
D8364 n8365 0 dm2 AREA=1.751e-06
D8365 n8366 0 dm2 AREA=1.636e-06
D8366 n8367 0 dm2 AREA=8.188e-07
D8367 n8368 0 dm2 AREA=1.044e-06
D8368 n8369 0 dm2 AREA=4.239e-07
D8369 n8370 0 dm2 AREA=1.953e-06
D8370 n8371 0 dm2 AREA=1.440e-06
D8371 n8372 0 dm2 AREA=8.623e-07
D8372 n8373 0 dm2 AREA=1.128e-06
D8373 n8374 0 dm2 AREA=1.608e-06
D8374 n8375 0 dm2 AREA=3.257e-07
D8375 n8376 0 dm2 AREA=8.712e-07
D8376 n8377 0 dm2 AREA=1.156e-07
D8377 n8378 0 dm2 AREA=1.106e-06
D8378 n8379 0 dm2 AREA=1.911e-06
D8379 n8380 0 dm2 AREA=4.154e-07
D8380 n8381 0 dm2 AREA=1.275e-06
D8381 n8382 0 dm2 AREA=1.122e-06
D8382 n8383 0 dm2 AREA=1.047e-06
D8383 n8384 0 dm2 AREA=8.114e-07
D8384 n8385 0 dm2 AREA=6.747e-07
D8385 n8386 0 dm2 AREA=7.907e-07
D8386 n8387 0 dm2 AREA=6.636e-07
D8387 n8388 0 dm2 AREA=1.306e-06
D8388 n8389 0 dm2 AREA=7.447e-07
D8389 n8390 0 dm2 AREA=8.345e-07
D8390 n8391 0 dm2 AREA=1.287e-06
D8391 n8392 0 dm2 AREA=1.421e-06
D8392 n8393 0 dm2 AREA=4.537e-07
D8393 n8394 0 dm2 AREA=8.069e-07
D8394 n8395 0 dm2 AREA=1.358e-06
D8395 n8396 0 dm2 AREA=9.198e-07
D8396 n8397 0 dm2 AREA=1.044e-06
D8397 n8398 0 dm2 AREA=1.494e-06
D8398 n8399 0 dm2 AREA=4.679e-07
D8399 n8400 0 dm2 AREA=8.088e-07
D8400 n8401 0 dm2 AREA=3.056e-07
D8401 n8402 0 dm2 AREA=1.137e-06
D8402 n8403 0 dm2 AREA=4.072e-07
D8403 n8404 0 dm2 AREA=7.339e-07
D8404 n8405 0 dm2 AREA=1.346e-06
D8405 n8406 0 dm2 AREA=8.335e-07
D8406 n8407 0 dm2 AREA=8.332e-07
D8407 n8408 0 dm2 AREA=6.860e-07
D8408 n8409 0 dm2 AREA=5.952e-07
D8409 n8410 0 dm2 AREA=2.278e-06
D8410 n8411 0 dm2 AREA=1.034e-06
D8411 n8412 0 dm2 AREA=1.137e-06
D8412 n8413 0 dm2 AREA=1.856e-06
D8413 n8414 0 dm2 AREA=4.483e-07
D8414 n8415 0 dm2 AREA=1.558e-06
D8415 n8416 0 dm2 AREA=7.434e-07
D8416 n8417 0 dm2 AREA=7.654e-07
D8417 n8418 0 dm2 AREA=2.803e-07
D8418 n8419 0 dm2 AREA=1.737e-06
D8419 n8420 0 dm2 AREA=8.571e-07
D8420 n8421 0 dm2 AREA=3.650e-07
D8421 n8422 0 dm2 AREA=4.245e-07
D8422 n8423 0 dm2 AREA=1.011e-06
D8423 n8424 0 dm2 AREA=5.437e-07
D8424 n8425 0 dm2 AREA=1.135e-06
D8425 n8426 0 dm2 AREA=2.922e-07
D8426 n8427 0 dm2 AREA=6.819e-07
D8427 n8428 0 dm2 AREA=1.568e-06
D8428 n8429 0 dm2 AREA=1.724e-06
D8429 n8430 0 dm2 AREA=1.275e-06
D8430 n8431 0 dm2 AREA=5.141e-07
D8431 n8432 0 dm2 AREA=1.077e-06
D8432 n8433 0 dm2 AREA=8.707e-07
D8433 n8434 0 dm2 AREA=7.797e-07
D8434 n8435 0 dm2 AREA=1.357e-06
D8435 n8436 0 dm2 AREA=1.161e-06
D8436 n8437 0 dm2 AREA=9.856e-07
D8437 n8438 0 dm2 AREA=1.045e-06
D8438 n8439 0 dm2 AREA=9.230e-07
D8439 n8440 0 dm2 AREA=3.564e-07
D8440 n8441 0 dm2 AREA=6.268e-07
D8441 n8442 0 dm2 AREA=6.613e-07
D8442 n8443 0 dm2 AREA=8.356e-07
D8443 n8444 0 dm2 AREA=3.703e-06
D8444 n8445 0 dm2 AREA=1.127e-06
D8445 n8446 0 dm2 AREA=1.193e-06
D8446 n8447 0 dm2 AREA=9.124e-07
D8447 n8448 0 dm2 AREA=1.041e-06
D8448 n8449 0 dm2 AREA=6.359e-07
D8449 n8450 0 dm2 AREA=1.411e-06
D8450 n8451 0 dm2 AREA=1.223e-06
D8451 n8452 0 dm2 AREA=1.476e-06
D8452 n8453 0 dm2 AREA=7.388e-07
D8453 n8454 0 dm2 AREA=6.355e-07
D8454 n8455 0 dm2 AREA=9.496e-07
D8455 n8456 0 dm2 AREA=9.936e-07
D8456 n8457 0 dm2 AREA=7.761e-07
D8457 n8458 0 dm2 AREA=1.167e-06
D8458 n8459 0 dm2 AREA=7.232e-07
D8459 n8460 0 dm2 AREA=7.545e-07
D8460 n8461 0 dm2 AREA=1.426e-06
D8461 n8462 0 dm2 AREA=5.643e-07
D8462 n8463 0 dm2 AREA=2.067e-06
D8463 n8464 0 dm2 AREA=1.126e-06
D8464 n8465 0 dm2 AREA=1.473e-06
D8465 n8466 0 dm2 AREA=9.068e-07
D8466 n8467 0 dm2 AREA=5.198e-07
D8467 n8468 0 dm2 AREA=7.193e-07
D8468 n8469 0 dm2 AREA=3.674e-07
D8469 n8470 0 dm2 AREA=1.526e-06
D8470 n8471 0 dm2 AREA=6.629e-07
D8471 n8472 0 dm2 AREA=1.048e-06
D8472 n8473 0 dm2 AREA=4.785e-07
D8473 n8474 0 dm2 AREA=1.118e-06
D8474 n8475 0 dm2 AREA=2.012e-06
D8475 n8476 0 dm2 AREA=1.196e-06
D8476 n8477 0 dm2 AREA=1.139e-06
D8477 n8478 0 dm2 AREA=9.284e-07
D8478 n8479 0 dm2 AREA=1.380e-06
D8479 n8480 0 dm2 AREA=8.864e-07
D8480 n8481 0 dm2 AREA=9.299e-07
D8481 n8482 0 dm2 AREA=1.135e-06
D8482 n8483 0 dm2 AREA=1.545e-06
D8483 n8484 0 dm2 AREA=1.427e-06
D8484 n8485 0 dm2 AREA=5.715e-07
D8485 n8486 0 dm2 AREA=6.800e-07
D8486 n8487 0 dm2 AREA=1.236e-06
D8487 n8488 0 dm2 AREA=8.403e-07
D8488 n8489 0 dm2 AREA=1.085e-06
D8489 n8490 0 dm2 AREA=1.489e-06
D8490 n8491 0 dm2 AREA=1.724e-06
D8491 n8492 0 dm2 AREA=1.421e-06
D8492 n8493 0 dm2 AREA=1.669e-06
D8493 n8494 0 dm2 AREA=1.138e-06
D8494 n8495 0 dm2 AREA=1.116e-06
D8495 n8496 0 dm2 AREA=5.361e-07
D8496 n8497 0 dm2 AREA=6.079e-07
D8497 n8498 0 dm2 AREA=1.326e-06
D8498 n8499 0 dm2 AREA=6.128e-07
D8499 n1 0 dm2 AREA=3.641e-07
D8500 n8501 0 dm2 AREA=6.395e-07
D8501 n8502 0 dm2 AREA=1.210e-06
D8502 n8503 0 dm2 AREA=1.207e-06
D8503 n8504 0 dm2 AREA=5.439e-07
D8504 n8505 0 dm2 AREA=1.924e-06
D8505 n8506 0 dm2 AREA=1.474e-06
D8506 n8507 0 dm2 AREA=1.262e-06
D8507 n8508 0 dm2 AREA=4.675e-07
D8508 n8509 0 dm2 AREA=1.409e-06
D8509 n8510 0 dm2 AREA=7.203e-07
D8510 n8511 0 dm2 AREA=4.354e-07
D8511 n8512 0 dm2 AREA=1.179e-06
D8512 n8513 0 dm2 AREA=3.753e-07
D8513 n8514 0 dm2 AREA=8.431e-07
D8514 n8515 0 dm2 AREA=7.982e-07
D8515 n8516 0 dm2 AREA=2.148e-07
D8516 n8517 0 dm2 AREA=7.741e-07
D8517 n8518 0 dm2 AREA=5.689e-07
D8518 n8519 0 dm2 AREA=4.964e-07
D8519 n8520 0 dm2 AREA=7.436e-07
D8520 n8521 0 dm2 AREA=1.890e-06
D8521 n8522 0 dm2 AREA=1.400e-06
D8522 n8523 0 dm2 AREA=5.859e-07
D8523 n8524 0 dm2 AREA=1.062e-06
D8524 n8525 0 dm2 AREA=1.300e-06
D8525 n8526 0 dm2 AREA=1.558e-06
D8526 n8527 0 dm2 AREA=1.355e-06
D8527 n8528 0 dm2 AREA=1.621e-06
D8528 n8529 0 dm2 AREA=1.741e-06
D8529 n8530 0 dm2 AREA=7.159e-07
D8530 n8531 0 dm2 AREA=6.573e-07
D8531 n8532 0 dm2 AREA=9.314e-07
D8532 n8533 0 dm2 AREA=6.240e-07
D8533 n8534 0 dm2 AREA=1.377e-06
D8534 n8535 0 dm2 AREA=1.628e-06
D8535 n8536 0 dm2 AREA=9.093e-07
D8536 n8537 0 dm2 AREA=2.763e-06
D8537 n8538 0 dm2 AREA=9.538e-07
D8538 n8539 0 dm2 AREA=1.412e-06
D8539 n8540 0 dm2 AREA=3.315e-07
D8540 n8541 0 dm2 AREA=5.841e-07
D8541 n8542 0 dm2 AREA=1.327e-06
D8542 n8543 0 dm2 AREA=1.243e-06
D8543 n8544 0 dm2 AREA=1.109e-06
D8544 n8545 0 dm2 AREA=1.447e-06
D8545 n8546 0 dm2 AREA=3.683e-07
D8546 n8547 0 dm2 AREA=2.888e-07
D8547 n8548 0 dm2 AREA=8.267e-07
D8548 n8549 0 dm2 AREA=4.284e-07
D8549 n8550 0 dm2 AREA=2.490e-06
D8550 n8551 0 dm2 AREA=6.979e-07
D8551 n8552 0 dm2 AREA=4.526e-07
D8552 n8553 0 dm2 AREA=1.427e-06
D8553 n8554 0 dm2 AREA=6.424e-07
D8554 n1 0 dm2 AREA=7.927e-07
D8555 n8556 0 dm2 AREA=9.533e-07
D8556 n8557 0 dm2 AREA=7.741e-07
D8557 n8558 0 dm2 AREA=1.224e-06
D8558 n8559 0 dm2 AREA=2.445e-06
D8559 n8560 0 dm2 AREA=7.838e-07
D8560 n8561 0 dm2 AREA=1.003e-06
D8561 n8562 0 dm2 AREA=1.295e-06
D8562 n8563 0 dm2 AREA=9.073e-07
D8563 n8564 0 dm2 AREA=2.132e-06
D8564 n8565 0 dm2 AREA=9.938e-07
D8565 n8566 0 dm2 AREA=7.318e-07
D8566 n8567 0 dm2 AREA=1.371e-06
D8567 n8568 0 dm2 AREA=1.118e-06
D8568 n8569 0 dm2 AREA=1.597e-06
D8569 n8570 0 dm2 AREA=7.243e-07
D8570 n8571 0 dm2 AREA=5.995e-07
D8571 n8572 0 dm2 AREA=1.154e-06
D8572 n8573 0 dm2 AREA=6.540e-07
D8573 n8574 0 dm2 AREA=1.812e-06
D8574 n8575 0 dm2 AREA=6.273e-07
D8575 n8576 0 dm2 AREA=8.487e-07
D8576 n8577 0 dm2 AREA=6.084e-07
D8577 n8578 0 dm2 AREA=1.972e-06
D8578 n8579 0 dm2 AREA=5.680e-07
D8579 n8580 0 dm2 AREA=7.897e-07
D8580 n8581 0 dm2 AREA=6.079e-07
D8581 n8582 0 dm2 AREA=7.741e-07
D8582 n8583 0 dm2 AREA=1.343e-06
D8583 n8584 0 dm2 AREA=6.097e-07
D8584 n8585 0 dm2 AREA=8.297e-07
D8585 n8586 0 dm2 AREA=5.502e-07
D8586 n8587 0 dm2 AREA=9.626e-07
D8587 n8588 0 dm2 AREA=1.600e-06
D8588 n8589 0 dm2 AREA=4.946e-07
D8589 n8590 0 dm2 AREA=2.626e-07
D8590 n8591 0 dm2 AREA=6.820e-07
D8591 n8592 0 dm2 AREA=1.949e-06
D8592 n8593 0 dm2 AREA=3.029e-07
D8593 n8594 0 dm2 AREA=1.966e-06
D8594 n8595 0 dm2 AREA=4.270e-07
D8595 n8596 0 dm2 AREA=1.104e-06
D8596 n8597 0 dm2 AREA=2.187e-07
D8597 n8598 0 dm2 AREA=3.899e-07
D8598 n8599 0 dm2 AREA=2.384e-06
D8599 n8600 0 dm2 AREA=7.257e-07
D8600 n8601 0 dm2 AREA=4.163e-07
D8601 n8602 0 dm2 AREA=4.046e-07
D8602 n1 0 dm2 AREA=1.378e-06
D8603 n8604 0 dm2 AREA=7.068e-07
D8604 n8605 0 dm2 AREA=8.184e-07
D8605 n8606 0 dm2 AREA=1.381e-06
D8606 n8607 0 dm2 AREA=1.388e-06
D8607 n8608 0 dm2 AREA=6.637e-07
D8608 n8609 0 dm2 AREA=2.686e-07
D8609 n8610 0 dm2 AREA=1.634e-06
D8610 n8611 0 dm2 AREA=1.245e-06
D8611 n8612 0 dm2 AREA=6.811e-07
D8612 n8613 0 dm2 AREA=9.537e-07
D8613 n8614 0 dm2 AREA=3.403e-07
D8614 n8615 0 dm2 AREA=9.037e-07
D8615 n8616 0 dm2 AREA=8.665e-07
D8616 n8617 0 dm2 AREA=7.988e-07
D8617 n8618 0 dm2 AREA=5.663e-07
D8618 n8619 0 dm2 AREA=1.240e-06
D8619 n8620 0 dm2 AREA=2.017e-06
D8620 n8621 0 dm2 AREA=1.224e-06
D8621 n8622 0 dm2 AREA=1.047e-06
D8622 n8623 0 dm2 AREA=8.764e-07
D8623 n8624 0 dm2 AREA=1.901e-06
D8624 n8625 0 dm2 AREA=1.940e-07
D8625 n8626 0 dm2 AREA=4.094e-07
D8626 n8627 0 dm2 AREA=9.609e-07
D8627 n8628 0 dm2 AREA=1.360e-06
D8628 n8629 0 dm2 AREA=1.043e-06
D8629 n8630 0 dm2 AREA=1.561e-06
D8630 n8631 0 dm2 AREA=8.270e-07
D8631 n8632 0 dm2 AREA=1.492e-06
D8632 n8633 0 dm2 AREA=9.758e-07
D8633 n8634 0 dm2 AREA=5.700e-07
D8634 n8635 0 dm2 AREA=7.943e-07
D8635 n8636 0 dm2 AREA=7.884e-08
D8636 n8637 0 dm2 AREA=8.708e-07
D8637 n8638 0 dm2 AREA=1.231e-06
D8638 n8639 0 dm2 AREA=5.934e-07
D8639 n8640 0 dm2 AREA=8.490e-07
D8640 n8641 0 dm2 AREA=5.933e-07
D8641 n8642 0 dm2 AREA=1.299e-06
D8642 n8643 0 dm2 AREA=4.241e-07
D8643 n8644 0 dm2 AREA=7.564e-07
D8644 n8645 0 dm2 AREA=1.169e-06
D8645 n8646 0 dm2 AREA=1.258e-06
D8646 n8647 0 dm2 AREA=1.027e-06
D8647 n8648 0 dm2 AREA=6.677e-07
D8648 n8649 0 dm2 AREA=2.551e-06
D8649 n8650 0 dm2 AREA=1.090e-06
D8650 n8651 0 dm2 AREA=7.045e-07
D8651 n8652 0 dm2 AREA=1.018e-06
D8652 n8653 0 dm2 AREA=1.529e-06
D8653 n8654 0 dm2 AREA=9.381e-07
D8654 n8655 0 dm2 AREA=2.773e-06
D8655 n8656 0 dm2 AREA=1.484e-06
D8656 n8657 0 dm2 AREA=1.414e-06
D8657 n8658 0 dm2 AREA=8.773e-07
D8658 n8659 0 dm2 AREA=4.288e-07
D8659 n8660 0 dm2 AREA=2.052e-06
D8660 n8661 0 dm2 AREA=1.040e-06
D8661 n8662 0 dm2 AREA=2.408e-06
D8662 n8663 0 dm2 AREA=1.295e-06
D8663 n8664 0 dm2 AREA=7.860e-07
D8664 n8665 0 dm2 AREA=1.703e-06
D8665 n8666 0 dm2 AREA=9.438e-07
D8666 n8667 0 dm2 AREA=2.915e-07
D8667 n8668 0 dm2 AREA=2.466e-07
D8668 n8669 0 dm2 AREA=8.897e-07
D8669 n8670 0 dm2 AREA=1.644e-06
D8670 n8671 0 dm2 AREA=1.426e-06
D8671 n8672 0 dm2 AREA=9.967e-07
D8672 n8673 0 dm2 AREA=1.155e-06
D8673 n8674 0 dm2 AREA=1.001e-06
D8674 n8675 0 dm2 AREA=1.053e-06
D8675 n8676 0 dm2 AREA=8.792e-07
D8676 n8677 0 dm2 AREA=6.576e-07
D8677 n8678 0 dm2 AREA=9.566e-07
D8678 n8679 0 dm2 AREA=1.663e-06
D8679 n1 0 dm2 AREA=2.254e-06
D8680 n8681 0 dm2 AREA=8.748e-07
D8681 n8682 0 dm2 AREA=8.824e-07
D8682 n8683 0 dm2 AREA=7.074e-07
D8683 n8684 0 dm2 AREA=7.425e-07
D8684 n8685 0 dm2 AREA=5.064e-07
D8685 n8686 0 dm2 AREA=1.142e-06
D8686 n8687 0 dm2 AREA=1.146e-06
D8687 n8688 0 dm2 AREA=1.314e-06
D8688 n8689 0 dm2 AREA=1.044e-06
D8689 n8690 0 dm2 AREA=1.066e-06
D8690 n8691 0 dm2 AREA=1.749e-06
D8691 n8692 0 dm2 AREA=1.113e-06
D8692 n8693 0 dm2 AREA=1.107e-06
D8693 n8694 0 dm2 AREA=1.530e-06
D8694 n8695 0 dm2 AREA=1.775e-07
D8695 n8696 0 dm2 AREA=2.835e-06
D8696 n8697 0 dm2 AREA=8.172e-07
D8697 n8698 0 dm2 AREA=1.166e-06
D8698 n8699 0 dm2 AREA=2.946e-06
D8699 n8700 0 dm2 AREA=7.459e-07
D8700 n8701 0 dm2 AREA=1.400e-06
D8701 n8702 0 dm2 AREA=6.136e-07
D8702 n8703 0 dm2 AREA=7.112e-07
D8703 n8704 0 dm2 AREA=6.242e-07
D8704 n8705 0 dm2 AREA=7.956e-07
D8705 n8706 0 dm2 AREA=9.065e-07
D8706 n8707 0 dm2 AREA=4.139e-07
D8707 n8708 0 dm2 AREA=5.939e-07
D8708 n8709 0 dm2 AREA=8.796e-07
D8709 n8710 0 dm2 AREA=1.204e-06
D8710 n8711 0 dm2 AREA=9.914e-07
D8711 n8712 0 dm2 AREA=2.595e-06
D8712 n8713 0 dm2 AREA=1.097e-06
D8713 n8714 0 dm2 AREA=3.618e-07
D8714 n8715 0 dm2 AREA=1.793e-06
D8715 n8716 0 dm2 AREA=6.386e-07
D8716 n8717 0 dm2 AREA=7.106e-07
D8717 n8718 0 dm2 AREA=8.367e-07
D8718 n8719 0 dm2 AREA=1.308e-06
D8719 n8720 0 dm2 AREA=1.298e-06
D8720 n8721 0 dm2 AREA=5.374e-07
D8721 n8722 0 dm2 AREA=1.865e-06
D8722 n8723 0 dm2 AREA=1.905e-06
D8723 n8724 0 dm2 AREA=3.030e-06
D8724 n8725 0 dm2 AREA=2.144e-06
D8725 n8726 0 dm2 AREA=1.296e-06
D8726 n8727 0 dm2 AREA=1.058e-06
D8727 n8728 0 dm2 AREA=1.029e-06
D8728 n8729 0 dm2 AREA=9.098e-07
D8729 n8730 0 dm2 AREA=1.297e-06
D8730 n8731 0 dm2 AREA=1.393e-06
D8731 n8732 0 dm2 AREA=1.123e-06
D8732 n8733 0 dm2 AREA=1.685e-07
D8733 n8734 0 dm2 AREA=1.893e-06
D8734 n8735 0 dm2 AREA=2.523e-07
D8735 n8736 0 dm2 AREA=1.577e-06
D8736 n8737 0 dm2 AREA=7.469e-07
D8737 n8738 0 dm2 AREA=1.050e-06
D8738 n8739 0 dm2 AREA=8.956e-07
D8739 n8740 0 dm2 AREA=3.008e-07
D8740 n8741 0 dm2 AREA=5.832e-07
D8741 n8742 0 dm2 AREA=1.272e-06
D8742 n8743 0 dm2 AREA=6.180e-07
D8743 n8744 0 dm2 AREA=1.147e-06
D8744 n8745 0 dm2 AREA=9.276e-07
D8745 n8746 0 dm2 AREA=4.592e-07
D8746 n8747 0 dm2 AREA=1.356e-06
D8747 n8748 0 dm2 AREA=7.304e-07
D8748 n8749 0 dm2 AREA=1.742e-06
D8749 n8750 0 dm2 AREA=2.045e-06
D8750 n8751 0 dm2 AREA=1.287e-06
D8751 n8752 0 dm2 AREA=7.048e-07
D8752 n8753 0 dm2 AREA=7.723e-07
D8753 n8754 0 dm2 AREA=7.600e-07
D8754 n8755 0 dm2 AREA=8.372e-07
D8755 n8756 0 dm2 AREA=8.985e-07
D8756 n8757 0 dm2 AREA=1.078e-06
D8757 n8758 0 dm2 AREA=1.126e-06
D8758 n8759 0 dm2 AREA=1.260e-06
D8759 n8760 0 dm2 AREA=1.015e-06
D8760 n8761 0 dm2 AREA=3.491e-07
D8761 n8762 0 dm2 AREA=1.001e-06
D8762 n8763 0 dm2 AREA=4.964e-07
D8763 n8764 0 dm2 AREA=8.046e-07
D8764 n8765 0 dm2 AREA=6.222e-07
D8765 n8766 0 dm2 AREA=1.321e-06
D8766 n8767 0 dm2 AREA=6.594e-07
D8767 n8768 0 dm2 AREA=1.457e-06
D8768 n8769 0 dm2 AREA=7.518e-07
D8769 n8770 0 dm2 AREA=2.084e-07
D8770 n8771 0 dm2 AREA=4.180e-07
D8771 n8772 0 dm2 AREA=6.294e-07
D8772 n8773 0 dm2 AREA=1.768e-06
D8773 n8774 0 dm2 AREA=3.343e-07
D8774 n8775 0 dm2 AREA=1.187e-06
D8775 n8776 0 dm2 AREA=9.757e-07
D8776 n8777 0 dm2 AREA=4.021e-07
D8777 n8778 0 dm2 AREA=1.347e-06
D8778 n8779 0 dm2 AREA=8.157e-07
D8779 n8780 0 dm2 AREA=1.726e-06
D8780 n8781 0 dm2 AREA=1.729e-06
D8781 n8782 0 dm2 AREA=8.279e-07
D8782 n8783 0 dm2 AREA=1.303e-06
D8783 n8784 0 dm2 AREA=8.220e-07
D8784 n8785 0 dm2 AREA=5.080e-07
D8785 n8786 0 dm2 AREA=8.189e-07
D8786 n8787 0 dm2 AREA=6.051e-07
D8787 n8788 0 dm2 AREA=1.453e-06
D8788 n8789 0 dm2 AREA=3.933e-07
D8789 n8790 0 dm2 AREA=1.373e-06
D8790 n8791 0 dm2 AREA=8.576e-07
D8791 n8792 0 dm2 AREA=9.655e-07
D8792 n8793 0 dm2 AREA=1.121e-06
D8793 n8794 0 dm2 AREA=3.740e-07
D8794 n8795 0 dm2 AREA=1.114e-06
D8795 n8796 0 dm2 AREA=5.100e-07
D8796 n8797 0 dm2 AREA=1.358e-06
D8797 n8798 0 dm2 AREA=1.571e-06
D8798 n8799 0 dm2 AREA=1.028e-06
D8799 n8800 0 dm2 AREA=7.581e-07
D8800 n8801 0 dm2 AREA=2.774e-06
D8801 n8802 0 dm2 AREA=7.150e-07
D8802 n8803 0 dm2 AREA=1.169e-06
D8803 n8804 0 dm2 AREA=7.196e-07
D8804 n8805 0 dm2 AREA=1.451e-06
D8805 n8806 0 dm2 AREA=8.751e-07
D8806 n8807 0 dm2 AREA=5.427e-07
D8807 n8808 0 dm2 AREA=2.700e-07
D8808 n8809 0 dm2 AREA=9.725e-07
D8809 n8810 0 dm2 AREA=5.221e-07
D8810 n8811 0 dm2 AREA=8.544e-07
D8811 n8812 0 dm2 AREA=1.059e-06
D8812 n8813 0 dm2 AREA=3.483e-07
D8813 n8814 0 dm2 AREA=1.912e-06
D8814 n8815 0 dm2 AREA=1.176e-06
D8815 n8816 0 dm2 AREA=1.467e-06
D8816 n8817 0 dm2 AREA=4.763e-07
D8817 n8818 0 dm2 AREA=8.863e-07
D8818 n8819 0 dm2 AREA=4.045e-07
D8819 n8820 0 dm2 AREA=8.199e-07
D8820 n8821 0 dm2 AREA=1.361e-06
D8821 n8822 0 dm2 AREA=8.228e-07
D8822 n8823 0 dm2 AREA=3.655e-07
D8823 n8824 0 dm2 AREA=1.777e-06
D8824 n8825 0 dm2 AREA=3.124e-07
D8825 n8826 0 dm2 AREA=8.386e-07
D8826 n8827 0 dm2 AREA=5.746e-07
D8827 n8828 0 dm2 AREA=8.156e-07
D8828 n8829 0 dm2 AREA=9.755e-07
D8829 n8830 0 dm2 AREA=6.554e-07
D8830 n8831 0 dm2 AREA=5.330e-07
D8831 n8832 0 dm2 AREA=1.615e-06
D8832 n8833 0 dm2 AREA=1.087e-06
D8833 n8834 0 dm2 AREA=3.380e-07
D8834 n8835 0 dm2 AREA=8.059e-07
D8835 n8836 0 dm2 AREA=7.331e-07
D8836 n8837 0 dm2 AREA=9.147e-07
D8837 n8838 0 dm2 AREA=1.473e-06
D8838 n8839 0 dm2 AREA=1.223e-06
D8839 n8840 0 dm2 AREA=1.774e-06
D8840 n8841 0 dm2 AREA=5.318e-07
D8841 n8842 0 dm2 AREA=9.419e-07
D8842 n1 0 dm2 AREA=1.409e-06
D8843 n8844 0 dm2 AREA=1.585e-06
D8844 n8845 0 dm2 AREA=9.685e-07
D8845 n8846 0 dm2 AREA=9.943e-07
D8846 n8847 0 dm2 AREA=9.164e-07
D8847 n8848 0 dm2 AREA=5.550e-07
D8848 n8849 0 dm2 AREA=1.298e-06
D8849 n8850 0 dm2 AREA=1.351e-06
D8850 n8851 0 dm2 AREA=7.609e-07
D8851 n8852 0 dm2 AREA=1.249e-06
D8852 n8853 0 dm2 AREA=1.083e-06
D8853 n8854 0 dm2 AREA=1.021e-06
D8854 n8855 0 dm2 AREA=1.521e-06
D8855 n8856 0 dm2 AREA=7.684e-07
D8856 n8857 0 dm2 AREA=8.424e-07
D8857 n8858 0 dm2 AREA=1.623e-06
D8858 n8859 0 dm2 AREA=1.616e-06
D8859 n8860 0 dm2 AREA=9.313e-07
D8860 n8861 0 dm2 AREA=5.559e-07
D8861 n8862 0 dm2 AREA=9.609e-07
D8862 n8863 0 dm2 AREA=1.257e-06
D8863 n8864 0 dm2 AREA=2.931e-07
D8864 n8865 0 dm2 AREA=1.501e-06
D8865 n8866 0 dm2 AREA=8.047e-07
D8866 n8867 0 dm2 AREA=1.412e-06
D8867 n8868 0 dm2 AREA=1.268e-06
D8868 n8869 0 dm2 AREA=1.230e-06
D8869 n8870 0 dm2 AREA=1.241e-06
D8870 n8871 0 dm2 AREA=6.378e-07
D8871 n8872 0 dm2 AREA=1.112e-06
D8872 n8873 0 dm2 AREA=1.221e-07
D8873 n8874 0 dm2 AREA=1.165e-07
D8874 n8875 0 dm2 AREA=7.613e-07
D8875 n8876 0 dm2 AREA=8.237e-07
D8876 n8877 0 dm2 AREA=8.698e-07
D8877 n8878 0 dm2 AREA=9.569e-07
D8878 n8879 0 dm2 AREA=4.140e-07
D8879 n8880 0 dm2 AREA=8.338e-07
D8880 n8881 0 dm2 AREA=1.003e-06
D8881 n8882 0 dm2 AREA=1.025e-06
D8882 n8883 0 dm2 AREA=8.868e-07
D8883 n8884 0 dm2 AREA=2.821e-06
D8884 n8885 0 dm2 AREA=3.296e-07
D8885 n8886 0 dm2 AREA=1.504e-06
D8886 n8887 0 dm2 AREA=5.538e-07
D8887 n8888 0 dm2 AREA=6.406e-07
D8888 n8889 0 dm2 AREA=5.921e-07
D8889 n8890 0 dm2 AREA=2.608e-07
D8890 n8891 0 dm2 AREA=1.761e-06
D8891 n8892 0 dm2 AREA=6.937e-07
D8892 n8893 0 dm2 AREA=8.129e-07
D8893 n8894 0 dm2 AREA=7.372e-07
D8894 n8895 0 dm2 AREA=5.805e-07
D8895 n8896 0 dm2 AREA=1.670e-06
D8896 n8897 0 dm2 AREA=6.345e-07
D8897 n8898 0 dm2 AREA=2.142e-06
D8898 n8899 0 dm2 AREA=9.214e-07
D8899 n8900 0 dm2 AREA=1.203e-06
D8900 n8901 0 dm2 AREA=1.260e-06
D8901 n8902 0 dm2 AREA=9.908e-07
D8902 n8903 0 dm2 AREA=2.469e-06
D8903 n8904 0 dm2 AREA=9.955e-07
D8904 n8905 0 dm2 AREA=6.653e-07
D8905 n8906 0 dm2 AREA=6.382e-07
D8906 n8907 0 dm2 AREA=8.489e-07
D8907 n8908 0 dm2 AREA=1.120e-06
D8908 n8909 0 dm2 AREA=1.202e-06
D8909 n8910 0 dm2 AREA=1.033e-06
D8910 n8911 0 dm2 AREA=9.804e-07
D8911 n8912 0 dm2 AREA=1.646e-06
D8912 n8913 0 dm2 AREA=2.431e-06
D8913 n8914 0 dm2 AREA=1.145e-06
D8914 n8915 0 dm2 AREA=1.019e-06
D8915 n8916 0 dm2 AREA=4.440e-07
D8916 n8917 0 dm2 AREA=9.123e-07
D8917 n8918 0 dm2 AREA=4.410e-07
D8918 n8919 0 dm2 AREA=1.759e-06
D8919 n8920 0 dm2 AREA=6.015e-07
D8920 n8921 0 dm2 AREA=1.571e-06
D8921 n8922 0 dm2 AREA=8.554e-07
D8922 n8923 0 dm2 AREA=7.187e-07
D8923 n8924 0 dm2 AREA=8.595e-07
D8924 n8925 0 dm2 AREA=6.887e-07
D8925 n1 0 dm2 AREA=1.243e-06
D8926 n8927 0 dm2 AREA=8.942e-07
D8927 n8928 0 dm2 AREA=1.125e-06
D8928 n8929 0 dm2 AREA=1.430e-06
D8929 n8930 0 dm2 AREA=1.490e-06
D8930 n8931 0 dm2 AREA=2.069e-06
D8931 n8932 0 dm2 AREA=2.034e-06
D8932 n8933 0 dm2 AREA=9.720e-07
D8933 n8934 0 dm2 AREA=1.112e-06
D8934 n8935 0 dm2 AREA=6.576e-07
D8935 n8936 0 dm2 AREA=4.585e-07
D8936 n8937 0 dm2 AREA=9.042e-07
D8937 n8938 0 dm2 AREA=1.346e-06
D8938 n8939 0 dm2 AREA=1.410e-06
D8939 n8940 0 dm2 AREA=9.564e-07
D8940 n8941 0 dm2 AREA=1.448e-06
D8941 n8942 0 dm2 AREA=3.437e-07
D8942 n8943 0 dm2 AREA=2.215e-06
D8943 n8944 0 dm2 AREA=5.784e-07
D8944 n8945 0 dm2 AREA=1.235e-06
D8945 n8946 0 dm2 AREA=1.954e-06
D8946 n8947 0 dm2 AREA=9.974e-07
D8947 n8948 0 dm2 AREA=1.268e-06
D8948 n8949 0 dm2 AREA=9.905e-07
D8949 n8950 0 dm2 AREA=7.282e-07
D8950 n8951 0 dm2 AREA=1.223e-06
D8951 n8952 0 dm2 AREA=5.635e-07
D8952 n8953 0 dm2 AREA=7.921e-07
D8953 n8954 0 dm2 AREA=4.451e-07
D8954 n8955 0 dm2 AREA=1.970e-06
D8955 n8956 0 dm2 AREA=4.373e-07
D8956 n8957 0 dm2 AREA=2.754e-07
D8957 n8958 0 dm2 AREA=9.027e-07
D8958 n8959 0 dm2 AREA=2.252e-07
D8959 n8960 0 dm2 AREA=3.282e-06
D8960 n8961 0 dm2 AREA=1.438e-06
D8961 n8962 0 dm2 AREA=5.836e-07
D8962 n8963 0 dm2 AREA=1.643e-06
D8963 n8964 0 dm2 AREA=2.665e-06
D8964 n8965 0 dm2 AREA=3.931e-07
D8965 n8966 0 dm2 AREA=5.072e-07
D8966 n8967 0 dm2 AREA=1.463e-06
D8967 n8968 0 dm2 AREA=1.781e-06
D8968 n8969 0 dm2 AREA=2.032e-06
D8969 n8970 0 dm2 AREA=5.819e-07
D8970 n8971 0 dm2 AREA=6.728e-07
D8971 n8972 0 dm2 AREA=7.511e-07
D8972 n8973 0 dm2 AREA=4.492e-07
D8973 n8974 0 dm2 AREA=1.374e-06
D8974 n8975 0 dm2 AREA=8.079e-07
D8975 n8976 0 dm2 AREA=5.310e-07
D8976 n8977 0 dm2 AREA=7.747e-07
D8977 n8978 0 dm2 AREA=9.098e-07
D8978 n8979 0 dm2 AREA=1.647e-06
D8979 n8980 0 dm2 AREA=6.084e-07
D8980 n8981 0 dm2 AREA=1.896e-06
D8981 n8982 0 dm2 AREA=5.815e-07
D8982 n8983 0 dm2 AREA=5.442e-07
D8983 n8984 0 dm2 AREA=1.176e-06
D8984 n8985 0 dm2 AREA=6.935e-07
D8985 n8986 0 dm2 AREA=1.065e-06
D8986 n8987 0 dm2 AREA=9.514e-07
D8987 n8988 0 dm2 AREA=1.381e-06
D8988 n8989 0 dm2 AREA=3.901e-07
D8989 n8990 0 dm2 AREA=9.942e-07
D8990 n8991 0 dm2 AREA=9.665e-07
D8991 n8992 0 dm2 AREA=1.258e-06
D8992 n8993 0 dm2 AREA=7.123e-07
D8993 n8994 0 dm2 AREA=5.796e-07
D8994 n8995 0 dm2 AREA=1.145e-06
D8995 n8996 0 dm2 AREA=6.296e-07
D8996 n8997 0 dm2 AREA=1.764e-06
D8997 n8998 0 dm2 AREA=1.057e-06
D8998 n8999 0 dm2 AREA=6.413e-07
D8999 n9000 0 dm2 AREA=6.026e-07
D9000 n9001 0 dm2 AREA=8.239e-07
D9001 n9002 0 dm2 AREA=1.866e-06
D9002 n9003 0 dm2 AREA=7.406e-07
D9003 n9004 0 dm2 AREA=1.187e-06
D9004 n9005 0 dm2 AREA=1.085e-06
D9005 n9006 0 dm2 AREA=7.505e-07
D9006 n9007 0 dm2 AREA=1.995e-06
D9007 n9008 0 dm2 AREA=9.828e-07
D9008 n9009 0 dm2 AREA=9.845e-07
D9009 n9010 0 dm2 AREA=7.399e-07
D9010 n9011 0 dm2 AREA=8.087e-07
D9011 n9012 0 dm2 AREA=1.320e-06
D9012 n9013 0 dm2 AREA=2.064e-06
D9013 n9014 0 dm2 AREA=1.222e-06
D9014 n9015 0 dm2 AREA=2.237e-07
D9015 n9016 0 dm2 AREA=7.645e-07
D9016 n9017 0 dm2 AREA=7.945e-07
D9017 n9018 0 dm2 AREA=2.052e-06
D9018 n9019 0 dm2 AREA=1.054e-06
D9019 n9020 0 dm2 AREA=7.870e-07
D9020 n9021 0 dm2 AREA=1.008e-06
D9021 n9022 0 dm2 AREA=6.151e-07
D9022 n9023 0 dm2 AREA=1.905e-06
D9023 n9024 0 dm2 AREA=4.870e-07
D9024 n9025 0 dm2 AREA=4.918e-07
D9025 n9026 0 dm2 AREA=1.302e-06
D9026 n9027 0 dm2 AREA=6.473e-07
D9027 n9028 0 dm2 AREA=5.801e-07
D9028 n9029 0 dm2 AREA=1.006e-06
D9029 n9030 0 dm2 AREA=1.042e-06
D9030 n9031 0 dm2 AREA=1.081e-06
D9031 n9032 0 dm2 AREA=1.764e-06
D9032 n9033 0 dm2 AREA=2.372e-06
D9033 n9034 0 dm2 AREA=2.778e-06
D9034 n9035 0 dm2 AREA=1.824e-06
D9035 n9036 0 dm2 AREA=1.092e-06
D9036 n9037 0 dm2 AREA=1.497e-06
D9037 n9038 0 dm2 AREA=5.802e-07
D9038 n9039 0 dm2 AREA=8.344e-07
D9039 n9040 0 dm2 AREA=1.086e-06
D9040 n9041 0 dm2 AREA=4.746e-07
D9041 n9042 0 dm2 AREA=1.090e-06
D9042 n9043 0 dm2 AREA=1.050e-06
D9043 n9044 0 dm2 AREA=1.191e-06
D9044 n9045 0 dm2 AREA=1.840e-06
D9045 n9046 0 dm2 AREA=1.210e-06
D9046 n9047 0 dm2 AREA=7.141e-07
D9047 n9048 0 dm2 AREA=3.731e-07
D9048 n9049 0 dm2 AREA=1.156e-06
D9049 n9050 0 dm2 AREA=6.473e-07
D9050 n9051 0 dm2 AREA=1.389e-06
D9051 n9052 0 dm2 AREA=8.005e-07
D9052 n9053 0 dm2 AREA=6.064e-07
D9053 n9054 0 dm2 AREA=9.150e-07
D9054 n9055 0 dm2 AREA=9.920e-07
D9055 n9056 0 dm2 AREA=2.222e-06
D9056 n9057 0 dm2 AREA=1.598e-06
D9057 n9058 0 dm2 AREA=2.153e-06
D9058 n9059 0 dm2 AREA=1.173e-06
D9059 n9060 0 dm2 AREA=1.144e-06
D9060 n9061 0 dm2 AREA=8.236e-07
D9061 n9062 0 dm2 AREA=9.046e-07
D9062 n9063 0 dm2 AREA=1.055e-06
D9063 n9064 0 dm2 AREA=9.348e-07
D9064 n9065 0 dm2 AREA=1.640e-06
D9065 n9066 0 dm2 AREA=5.204e-07
D9066 n9067 0 dm2 AREA=1.033e-06
D9067 n9068 0 dm2 AREA=1.016e-06
D9068 n9069 0 dm2 AREA=4.885e-07
D9069 n9070 0 dm2 AREA=9.719e-07
D9070 n9071 0 dm2 AREA=9.486e-07
D9071 n9072 0 dm2 AREA=1.875e-07
D9072 n9073 0 dm2 AREA=7.134e-07
D9073 n9074 0 dm2 AREA=8.170e-07
D9074 n9075 0 dm2 AREA=6.665e-07
D9075 n9076 0 dm2 AREA=5.630e-07
D9076 n9077 0 dm2 AREA=9.007e-07
D9077 n9078 0 dm2 AREA=7.448e-07
D9078 n9079 0 dm2 AREA=1.035e-06
D9079 n9080 0 dm2 AREA=1.763e-06
D9080 n9081 0 dm2 AREA=1.173e-06
D9081 n1 0 dm2 AREA=9.370e-07
D9082 n9083 0 dm2 AREA=6.217e-07
D9083 n9084 0 dm2 AREA=4.770e-07
D9084 n9085 0 dm2 AREA=1.312e-06
D9085 n9086 0 dm2 AREA=7.326e-07
D9086 n9087 0 dm2 AREA=7.066e-07
D9087 n9088 0 dm2 AREA=1.615e-06
D9088 n9089 0 dm2 AREA=1.514e-06
D9089 n9090 0 dm2 AREA=9.708e-07
D9090 n9091 0 dm2 AREA=5.126e-07
D9091 n9092 0 dm2 AREA=4.423e-07
D9092 n9093 0 dm2 AREA=7.587e-07
D9093 n9094 0 dm2 AREA=1.859e-06
D9094 n9095 0 dm2 AREA=1.779e-07
D9095 n9096 0 dm2 AREA=7.933e-07
D9096 n9097 0 dm2 AREA=8.364e-07
D9097 n9098 0 dm2 AREA=9.857e-07
D9098 n9099 0 dm2 AREA=1.232e-06
D9099 n9100 0 dm2 AREA=1.204e-06
D9100 n9101 0 dm2 AREA=2.840e-06
D9101 n9102 0 dm2 AREA=5.841e-07
D9102 n9103 0 dm2 AREA=2.478e-06
D9103 n9104 0 dm2 AREA=4.680e-07
D9104 n9105 0 dm2 AREA=2.315e-06
D9105 n9106 0 dm2 AREA=1.483e-06
D9106 n9107 0 dm2 AREA=1.380e-06
D9107 n9108 0 dm2 AREA=1.184e-06
D9108 n9109 0 dm2 AREA=1.093e-06
D9109 n9110 0 dm2 AREA=1.111e-06
D9110 n9111 0 dm2 AREA=6.597e-07
D9111 n9112 0 dm2 AREA=2.559e-07
D9112 n9113 0 dm2 AREA=5.110e-07
D9113 n9114 0 dm2 AREA=1.655e-06
D9114 n9115 0 dm2 AREA=1.036e-06
D9115 n9116 0 dm2 AREA=6.803e-07
D9116 n9117 0 dm2 AREA=4.589e-07
D9117 n9118 0 dm2 AREA=3.260e-06
D9118 n9119 0 dm2 AREA=6.220e-07
D9119 n9120 0 dm2 AREA=1.499e-06
D9120 n9121 0 dm2 AREA=6.944e-07
D9121 n9122 0 dm2 AREA=1.475e-06
D9122 n9123 0 dm2 AREA=5.548e-07
D9123 n9124 0 dm2 AREA=1.175e-06
D9124 n9125 0 dm2 AREA=3.769e-07
D9125 n9126 0 dm2 AREA=2.746e-06
D9126 n9127 0 dm2 AREA=1.436e-06
D9127 n9128 0 dm2 AREA=9.416e-07
D9128 n9129 0 dm2 AREA=6.171e-07
D9129 n9130 0 dm2 AREA=7.856e-07
D9130 n9131 0 dm2 AREA=1.264e-06
D9131 n9132 0 dm2 AREA=9.014e-07
D9132 n9133 0 dm2 AREA=1.325e-06
D9133 n9134 0 dm2 AREA=5.441e-07
D9134 n9135 0 dm2 AREA=4.225e-07
D9135 n9136 0 dm2 AREA=1.005e-06
D9136 n9137 0 dm2 AREA=6.365e-07
D9137 n1 0 dm2 AREA=1.855e-06
D9138 n9139 0 dm2 AREA=1.633e-06
D9139 n9140 0 dm2 AREA=9.594e-07
D9140 n9141 0 dm2 AREA=9.904e-07
D9141 n9142 0 dm2 AREA=8.540e-07
D9142 n9143 0 dm2 AREA=7.636e-07
D9143 n9144 0 dm2 AREA=3.969e-07
D9144 n9145 0 dm2 AREA=8.321e-07
D9145 n9146 0 dm2 AREA=8.587e-07
D9146 n9147 0 dm2 AREA=9.099e-07
D9147 n9148 0 dm2 AREA=7.646e-07
D9148 n9149 0 dm2 AREA=1.185e-06
D9149 n9150 0 dm2 AREA=1.739e-06
D9150 n9151 0 dm2 AREA=6.121e-07
D9151 n9152 0 dm2 AREA=5.068e-07
D9152 n9153 0 dm2 AREA=3.735e-07
D9153 n9154 0 dm2 AREA=2.117e-06
D9154 n9155 0 dm2 AREA=6.947e-07
D9155 n9156 0 dm2 AREA=1.116e-06
D9156 n9157 0 dm2 AREA=9.158e-07
D9157 n9158 0 dm2 AREA=1.597e-06
D9158 n9159 0 dm2 AREA=3.499e-07
D9159 n9160 0 dm2 AREA=8.128e-07
D9160 n9161 0 dm2 AREA=4.126e-07
D9161 n9162 0 dm2 AREA=5.300e-07
D9162 n9163 0 dm2 AREA=1.212e-06
D9163 n9164 0 dm2 AREA=4.911e-07
D9164 n9165 0 dm2 AREA=3.226e-07
D9165 n9166 0 dm2 AREA=8.434e-07
D9166 n9167 0 dm2 AREA=1.844e-06
D9167 n9168 0 dm2 AREA=1.994e-06
D9168 n9169 0 dm2 AREA=1.664e-06
D9169 n9170 0 dm2 AREA=1.693e-07
D9170 n9171 0 dm2 AREA=5.608e-07
D9171 n9172 0 dm2 AREA=1.186e-06
D9172 n9173 0 dm2 AREA=4.959e-07
D9173 n9174 0 dm2 AREA=6.902e-07
D9174 n9175 0 dm2 AREA=6.850e-07
D9175 n9176 0 dm2 AREA=5.440e-07
D9176 n9177 0 dm2 AREA=1.456e-06
D9177 n9178 0 dm2 AREA=1.354e-06
D9178 n9179 0 dm2 AREA=6.425e-07
D9179 n9180 0 dm2 AREA=9.429e-07
D9180 n9181 0 dm2 AREA=8.092e-07
D9181 n9182 0 dm2 AREA=8.470e-07
D9182 n9183 0 dm2 AREA=2.738e-07
D9183 n9184 0 dm2 AREA=2.340e-07
D9184 n9185 0 dm2 AREA=5.094e-07
D9185 n9186 0 dm2 AREA=1.107e-06
D9186 n9187 0 dm2 AREA=5.820e-07
D9187 n9188 0 dm2 AREA=7.728e-07
D9188 n9189 0 dm2 AREA=1.347e-06
D9189 n9190 0 dm2 AREA=5.425e-07
D9190 n9191 0 dm2 AREA=1.077e-06
D9191 n9192 0 dm2 AREA=5.925e-07
D9192 n9193 0 dm2 AREA=3.080e-07
D9193 n9194 0 dm2 AREA=8.663e-07
D9194 n9195 0 dm2 AREA=1.242e-07
D9195 n9196 0 dm2 AREA=1.748e-07
D9196 n9197 0 dm2 AREA=3.020e-07
D9197 n9198 0 dm2 AREA=1.269e-06
D9198 n9199 0 dm2 AREA=7.740e-07
D9199 n9200 0 dm2 AREA=1.074e-06
D9200 n9201 0 dm2 AREA=5.049e-07
D9201 n9202 0 dm2 AREA=1.825e-06
D9202 n9203 0 dm2 AREA=1.271e-06
D9203 n9204 0 dm2 AREA=1.557e-06
D9204 n9205 0 dm2 AREA=2.537e-06
D9205 n9206 0 dm2 AREA=1.177e-06
D9206 n9207 0 dm2 AREA=1.151e-06
D9207 n9208 0 dm2 AREA=8.917e-07
D9208 n9209 0 dm2 AREA=9.338e-07
D9209 n9210 0 dm2 AREA=1.934e-06
D9210 n9211 0 dm2 AREA=7.611e-07
D9211 n9212 0 dm2 AREA=2.270e-06
D9212 n9213 0 dm2 AREA=1.177e-06
D9213 n9214 0 dm2 AREA=9.970e-07
D9214 n9215 0 dm2 AREA=3.758e-07
D9215 n9216 0 dm2 AREA=1.271e-06
D9216 n9217 0 dm2 AREA=9.860e-07
D9217 n9218 0 dm2 AREA=7.411e-07
D9218 n9219 0 dm2 AREA=4.153e-07
D9219 n9220 0 dm2 AREA=1.100e-06
D9220 n9221 0 dm2 AREA=1.376e-06
D9221 n9222 0 dm2 AREA=1.106e-06
D9222 n9223 0 dm2 AREA=6.913e-07
D9223 n9224 0 dm2 AREA=7.855e-07
D9224 n9225 0 dm2 AREA=9.579e-07
D9225 n9226 0 dm2 AREA=1.427e-07
D9226 n9227 0 dm2 AREA=5.797e-07
D9227 n9228 0 dm2 AREA=1.162e-06
D9228 n9229 0 dm2 AREA=1.303e-06
D9229 n9230 0 dm2 AREA=1.014e-06
D9230 n9231 0 dm2 AREA=1.837e-06
D9231 n9232 0 dm2 AREA=4.486e-07
D9232 n9233 0 dm2 AREA=8.420e-07
D9233 n9234 0 dm2 AREA=1.223e-06
D9234 n9235 0 dm2 AREA=1.072e-06
D9235 n9236 0 dm2 AREA=6.895e-07
D9236 n9237 0 dm2 AREA=1.488e-06
D9237 n9238 0 dm2 AREA=4.379e-07
D9238 n9239 0 dm2 AREA=7.838e-07
D9239 n9240 0 dm2 AREA=1.094e-06
D9240 n9241 0 dm2 AREA=9.197e-07
D9241 n9242 0 dm2 AREA=2.238e-07
D9242 n9243 0 dm2 AREA=8.006e-07
D9243 n9244 0 dm2 AREA=1.000e-06
D9244 n9245 0 dm2 AREA=7.979e-07
D9245 n9246 0 dm2 AREA=5.401e-07
D9246 n9247 0 dm2 AREA=7.731e-07
D9247 n9248 0 dm2 AREA=8.708e-07
D9248 n9249 0 dm2 AREA=1.458e-06
D9249 n9250 0 dm2 AREA=8.660e-07
D9250 n9251 0 dm2 AREA=7.692e-07
D9251 n9252 0 dm2 AREA=1.181e-06
D9252 n9253 0 dm2 AREA=1.160e-06
D9253 n9254 0 dm2 AREA=1.507e-06
D9254 n9255 0 dm2 AREA=7.987e-07
D9255 n9256 0 dm2 AREA=9.246e-07
D9256 n9257 0 dm2 AREA=1.928e-06
D9257 n9258 0 dm2 AREA=1.170e-06
D9258 n9259 0 dm2 AREA=5.751e-07
D9259 n9260 0 dm2 AREA=3.619e-07
D9260 n9261 0 dm2 AREA=6.095e-07
D9261 n9262 0 dm2 AREA=2.847e-07
D9262 n9263 0 dm2 AREA=1.003e-06
D9263 n9264 0 dm2 AREA=1.065e-06
D9264 n9265 0 dm2 AREA=4.645e-07
D9265 n9266 0 dm2 AREA=1.106e-06
D9266 n9267 0 dm2 AREA=4.273e-07
D9267 n9268 0 dm2 AREA=8.742e-07
D9268 n9269 0 dm2 AREA=4.871e-07
D9269 n9270 0 dm2 AREA=7.915e-07
D9270 n9271 0 dm2 AREA=1.443e-06
D9271 n9272 0 dm2 AREA=2.170e-06
D9272 n9273 0 dm2 AREA=4.834e-07
D9273 n9274 0 dm2 AREA=4.411e-07
D9274 n9275 0 dm2 AREA=1.416e-06
D9275 n9276 0 dm2 AREA=1.547e-06
D9276 n9277 0 dm2 AREA=8.223e-07
D9277 n9278 0 dm2 AREA=1.893e-07
D9278 n9279 0 dm2 AREA=8.586e-07
D9279 n9280 0 dm2 AREA=7.546e-07
D9280 n9281 0 dm2 AREA=3.663e-07
D9281 n9282 0 dm2 AREA=1.730e-06
D9282 n9283 0 dm2 AREA=9.320e-07
D9283 n9284 0 dm2 AREA=1.109e-06
D9284 n9285 0 dm2 AREA=9.532e-07
D9285 n9286 0 dm2 AREA=1.414e-06
D9286 n9287 0 dm2 AREA=7.385e-07
D9287 n9288 0 dm2 AREA=1.432e-06
D9288 n9289 0 dm2 AREA=1.943e-06
D9289 n9290 0 dm2 AREA=1.584e-06
D9290 n9291 0 dm2 AREA=4.575e-07
D9291 n9292 0 dm2 AREA=1.620e-06
D9292 n9293 0 dm2 AREA=1.076e-06
D9293 n9294 0 dm2 AREA=5.032e-07
D9294 n9295 0 dm2 AREA=1.326e-06
D9295 n9296 0 dm2 AREA=9.752e-07
D9296 n9297 0 dm2 AREA=3.649e-07
D9297 n9298 0 dm2 AREA=2.807e-06
D9298 n9299 0 dm2 AREA=1.604e-06
D9299 n9300 0 dm2 AREA=2.830e-07
D9300 n9301 0 dm2 AREA=6.572e-07
D9301 n9302 0 dm2 AREA=5.747e-07
D9302 n9303 0 dm2 AREA=1.681e-06
D9303 n9304 0 dm2 AREA=1.004e-06
D9304 n9305 0 dm2 AREA=3.317e-07
D9305 n9306 0 dm2 AREA=1.716e-06
D9306 n9307 0 dm2 AREA=1.914e-06
D9307 n9308 0 dm2 AREA=8.640e-07
D9308 n9309 0 dm2 AREA=1.657e-06
D9309 n9310 0 dm2 AREA=7.621e-07
D9310 n9311 0 dm2 AREA=9.867e-07
D9311 n9312 0 dm2 AREA=4.117e-07
D9312 n9313 0 dm2 AREA=1.366e-06
D9313 n9314 0 dm2 AREA=3.528e-07
D9314 n9315 0 dm2 AREA=1.322e-06
D9315 n9316 0 dm2 AREA=8.340e-07
D9316 n9317 0 dm2 AREA=6.045e-07
D9317 n9318 0 dm2 AREA=8.800e-07
D9318 n9319 0 dm2 AREA=7.363e-07
D9319 n9320 0 dm2 AREA=1.266e-06
D9320 n9321 0 dm2 AREA=1.445e-06
D9321 n9322 0 dm2 AREA=1.959e-06
D9322 n9323 0 dm2 AREA=1.407e-06
D9323 n9324 0 dm2 AREA=7.654e-07
D9324 n1 0 dm2 AREA=9.194e-07
D9325 n9326 0 dm2 AREA=5.794e-07
D9326 n9327 0 dm2 AREA=1.413e-06
D9327 n9328 0 dm2 AREA=5.108e-07
D9328 n9329 0 dm2 AREA=4.352e-07
D9329 n9330 0 dm2 AREA=2.216e-07
D9330 n9331 0 dm2 AREA=5.426e-07
D9331 n9332 0 dm2 AREA=1.917e-06
D9332 n9333 0 dm2 AREA=1.038e-06
D9333 n9334 0 dm2 AREA=6.376e-07
D9334 n9335 0 dm2 AREA=3.560e-07
D9335 n9336 0 dm2 AREA=1.352e-07
D9336 n9337 0 dm2 AREA=4.764e-07
D9337 n9338 0 dm2 AREA=1.040e-06
D9338 n9339 0 dm2 AREA=1.784e-06
D9339 n9340 0 dm2 AREA=3.271e-07
D9340 n9341 0 dm2 AREA=3.134e-07
D9341 n9342 0 dm2 AREA=2.185e-06
D9342 n9343 0 dm2 AREA=2.946e-07
D9343 n9344 0 dm2 AREA=1.260e-06
D9344 n9345 0 dm2 AREA=1.001e-06
D9345 n9346 0 dm2 AREA=1.429e-06
D9346 n9347 0 dm2 AREA=1.361e-06
D9347 n9348 0 dm2 AREA=4.281e-07
D9348 n9349 0 dm2 AREA=1.296e-06
D9349 n9350 0 dm2 AREA=6.922e-07
D9350 n9351 0 dm2 AREA=6.154e-07
D9351 n9352 0 dm2 AREA=6.006e-07
D9352 n9353 0 dm2 AREA=8.781e-07
D9353 n9354 0 dm2 AREA=1.306e-06
D9354 n9355 0 dm2 AREA=1.285e-06
D9355 n9356 0 dm2 AREA=6.447e-07
D9356 n9357 0 dm2 AREA=2.246e-07
D9357 n9358 0 dm2 AREA=7.244e-07
D9358 n9359 0 dm2 AREA=7.382e-07
D9359 n9360 0 dm2 AREA=5.200e-07
D9360 n9361 0 dm2 AREA=8.816e-07
D9361 n9362 0 dm2 AREA=4.203e-07
D9362 n9363 0 dm2 AREA=6.849e-07
D9363 n9364 0 dm2 AREA=9.534e-07
D9364 n9365 0 dm2 AREA=1.670e-06
D9365 n9366 0 dm2 AREA=1.254e-06
D9366 n9367 0 dm2 AREA=5.298e-07
D9367 n9368 0 dm2 AREA=9.960e-07
D9368 n9369 0 dm2 AREA=1.227e-06
D9369 n9370 0 dm2 AREA=1.460e-06
D9370 n9371 0 dm2 AREA=4.797e-07
D9371 n9372 0 dm2 AREA=4.509e-07
D9372 n9373 0 dm2 AREA=1.497e-06
D9373 n9374 0 dm2 AREA=5.381e-07
D9374 n9375 0 dm2 AREA=1.034e-06
D9375 n9376 0 dm2 AREA=4.288e-07
D9376 n9377 0 dm2 AREA=8.231e-07
D9377 n9378 0 dm2 AREA=1.783e-06
D9378 n9379 0 dm2 AREA=1.662e-06
D9379 n9380 0 dm2 AREA=1.190e-06
D9380 n9381 0 dm2 AREA=7.706e-07
D9381 n9382 0 dm2 AREA=2.200e-07
D9382 n9383 0 dm2 AREA=8.227e-07
D9383 n9384 0 dm2 AREA=6.616e-07
D9384 n9385 0 dm2 AREA=5.589e-07
D9385 n9386 0 dm2 AREA=1.075e-06
D9386 n9387 0 dm2 AREA=1.821e-06
D9387 n9388 0 dm2 AREA=2.202e-06
D9388 n9389 0 dm2 AREA=6.938e-07
D9389 n9390 0 dm2 AREA=5.198e-07
D9390 n9391 0 dm2 AREA=7.991e-07
D9391 n9392 0 dm2 AREA=5.208e-07
D9392 n9393 0 dm2 AREA=1.003e-06
D9393 n9394 0 dm2 AREA=7.983e-07
D9394 n9395 0 dm2 AREA=5.863e-07
D9395 n9396 0 dm2 AREA=2.169e-07
D9396 n9397 0 dm2 AREA=2.355e-07
D9397 n9398 0 dm2 AREA=2.596e-07
D9398 n9399 0 dm2 AREA=3.143e-07
D9399 n9400 0 dm2 AREA=1.151e-06
D9400 n9401 0 dm2 AREA=7.042e-07
D9401 n9402 0 dm2 AREA=7.218e-07
D9402 n9403 0 dm2 AREA=7.292e-07
D9403 n9404 0 dm2 AREA=5.938e-07
D9404 n9405 0 dm2 AREA=1.936e-06
D9405 n9406 0 dm2 AREA=7.133e-07
D9406 n9407 0 dm2 AREA=9.208e-07
D9407 n9408 0 dm2 AREA=1.420e-06
D9408 n9409 0 dm2 AREA=1.093e-06
D9409 n9410 0 dm2 AREA=4.933e-07
D9410 n9411 0 dm2 AREA=7.933e-07
D9411 n9412 0 dm2 AREA=1.038e-06
D9412 n9413 0 dm2 AREA=1.623e-06
D9413 n9414 0 dm2 AREA=3.005e-07
D9414 n9415 0 dm2 AREA=6.112e-07
D9415 n9416 0 dm2 AREA=1.242e-06
D9416 n9417 0 dm2 AREA=1.571e-06
D9417 n9418 0 dm2 AREA=2.266e-06
D9418 n9419 0 dm2 AREA=1.034e-06
D9419 n9420 0 dm2 AREA=7.575e-07
D9420 n9421 0 dm2 AREA=6.052e-07
D9421 n9422 0 dm2 AREA=8.355e-07
D9422 n9423 0 dm2 AREA=9.919e-07
D9423 n9424 0 dm2 AREA=7.359e-07
D9424 n9425 0 dm2 AREA=1.493e-06
D9425 n9426 0 dm2 AREA=2.462e-07
D9426 n9427 0 dm2 AREA=5.893e-07
D9427 n9428 0 dm2 AREA=4.235e-07
D9428 n9429 0 dm2 AREA=7.408e-07
D9429 n9430 0 dm2 AREA=5.185e-07
D9430 n9431 0 dm2 AREA=6.979e-07
D9431 n9432 0 dm2 AREA=8.173e-07
D9432 n9433 0 dm2 AREA=1.193e-06
D9433 n9434 0 dm2 AREA=8.609e-07
D9434 n9435 0 dm2 AREA=1.429e-06
D9435 n9436 0 dm2 AREA=3.458e-06
D9436 n9437 0 dm2 AREA=1.120e-06
D9437 n9438 0 dm2 AREA=1.146e-07
D9438 n9439 0 dm2 AREA=8.051e-07
D9439 n9440 0 dm2 AREA=1.068e-06
D9440 n9441 0 dm2 AREA=7.821e-07
D9441 n9442 0 dm2 AREA=3.458e-07
D9442 n9443 0 dm2 AREA=1.338e-06
D9443 n9444 0 dm2 AREA=1.536e-06
D9444 n9445 0 dm2 AREA=2.610e-06
D9445 n9446 0 dm2 AREA=1.369e-06
D9446 n9447 0 dm2 AREA=6.551e-07
D9447 n9448 0 dm2 AREA=9.482e-07
D9448 n9449 0 dm2 AREA=1.038e-06
D9449 n9450 0 dm2 AREA=1.521e-06
D9450 n9451 0 dm2 AREA=2.089e-06
D9451 n9452 0 dm2 AREA=1.398e-06
D9452 n9453 0 dm2 AREA=1.007e-06
D9453 n9454 0 dm2 AREA=6.556e-07
D9454 n9455 0 dm2 AREA=1.641e-07
D9455 n9456 0 dm2 AREA=1.272e-06
D9456 n9457 0 dm2 AREA=4.481e-07
D9457 n9458 0 dm2 AREA=9.561e-07
D9458 n9459 0 dm2 AREA=3.976e-07
D9459 n9460 0 dm2 AREA=5.475e-07
D9460 n9461 0 dm2 AREA=1.143e-06
D9461 n9462 0 dm2 AREA=1.515e-06
D9462 n9463 0 dm2 AREA=7.430e-07
D9463 n9464 0 dm2 AREA=1.416e-06
D9464 n9465 0 dm2 AREA=1.050e-06
D9465 n9466 0 dm2 AREA=4.960e-07
D9466 n9467 0 dm2 AREA=4.925e-07
D9467 n9468 0 dm2 AREA=7.081e-07
D9468 n9469 0 dm2 AREA=1.526e-06
D9469 n9470 0 dm2 AREA=8.594e-07
D9470 n9471 0 dm2 AREA=1.062e-06
D9471 n9472 0 dm2 AREA=1.281e-06
D9472 n9473 0 dm2 AREA=7.555e-07
D9473 n9474 0 dm2 AREA=7.517e-07
D9474 n9475 0 dm2 AREA=9.537e-07
D9475 n9476 0 dm2 AREA=5.160e-07
D9476 n9477 0 dm2 AREA=6.872e-07
D9477 n9478 0 dm2 AREA=3.708e-07
D9478 n9479 0 dm2 AREA=1.022e-06
D9479 n9480 0 dm2 AREA=1.646e-06
D9480 n9481 0 dm2 AREA=1.643e-06
D9481 n9482 0 dm2 AREA=6.375e-07
D9482 n9483 0 dm2 AREA=9.534e-07
D9483 n9484 0 dm2 AREA=2.337e-07
D9484 n9485 0 dm2 AREA=9.238e-07
D9485 n9486 0 dm2 AREA=6.732e-07
D9486 n9487 0 dm2 AREA=1.816e-06
D9487 n9488 0 dm2 AREA=7.160e-07
D9488 n9489 0 dm2 AREA=6.668e-07
D9489 n9490 0 dm2 AREA=1.067e-06
D9490 n9491 0 dm2 AREA=1.108e-06
D9491 n9492 0 dm2 AREA=4.998e-07
D9492 n9493 0 dm2 AREA=1.928e-06
D9493 n9494 0 dm2 AREA=1.155e-06
D9494 n9495 0 dm2 AREA=1.040e-06
D9495 n9496 0 dm2 AREA=6.379e-07
D9496 n9497 0 dm2 AREA=6.973e-07
D9497 n9498 0 dm2 AREA=3.038e-07
D9498 n9499 0 dm2 AREA=7.334e-07
D9499 n9500 0 dm2 AREA=1.474e-07
D9500 n9501 0 dm2 AREA=3.476e-07
D9501 n9502 0 dm2 AREA=6.793e-07
D9502 n9503 0 dm2 AREA=1.510e-06
D9503 n9504 0 dm2 AREA=3.998e-07
D9504 n9505 0 dm2 AREA=8.567e-07
D9505 n9506 0 dm2 AREA=1.991e-06
D9506 n9507 0 dm2 AREA=1.582e-06
D9507 n9508 0 dm2 AREA=6.213e-07
D9508 n9509 0 dm2 AREA=5.476e-07
D9509 n9510 0 dm2 AREA=4.532e-06
D9510 n1 0 dm2 AREA=7.783e-07
D9511 n9512 0 dm2 AREA=1.631e-06
D9512 n9513 0 dm2 AREA=6.741e-07
D9513 n9514 0 dm2 AREA=6.873e-07
D9514 n9515 0 dm2 AREA=2.652e-06
D9515 n9516 0 dm2 AREA=7.689e-07
D9516 n9517 0 dm2 AREA=1.182e-06
D9517 n9518 0 dm2 AREA=5.291e-07
D9518 n9519 0 dm2 AREA=9.869e-07
D9519 n9520 0 dm2 AREA=9.682e-07
D9520 n9521 0 dm2 AREA=8.429e-07
D9521 n9522 0 dm2 AREA=1.521e-06
D9522 n9523 0 dm2 AREA=8.640e-07
D9523 n9524 0 dm2 AREA=5.145e-07
D9524 n9525 0 dm2 AREA=3.031e-06
D9525 n9526 0 dm2 AREA=9.136e-07
D9526 n9527 0 dm2 AREA=6.582e-07
D9527 n9528 0 dm2 AREA=9.429e-07
D9528 n9529 0 dm2 AREA=1.863e-06
D9529 n9530 0 dm2 AREA=6.212e-07
D9530 n9531 0 dm2 AREA=3.090e-07
D9531 n9532 0 dm2 AREA=6.298e-07
D9532 n9533 0 dm2 AREA=5.710e-07
D9533 n9534 0 dm2 AREA=8.921e-07
D9534 n9535 0 dm2 AREA=1.170e-06
D9535 n9536 0 dm2 AREA=1.010e-06
D9536 n9537 0 dm2 AREA=7.272e-07
D9537 n9538 0 dm2 AREA=7.079e-07
D9538 n9539 0 dm2 AREA=2.616e-07
D9539 n9540 0 dm2 AREA=4.876e-07
D9540 n9541 0 dm2 AREA=6.972e-07
D9541 n9542 0 dm2 AREA=8.982e-07
D9542 n9543 0 dm2 AREA=8.724e-07
D9543 n9544 0 dm2 AREA=3.367e-07
D9544 n9545 0 dm2 AREA=6.689e-07
D9545 n9546 0 dm2 AREA=2.181e-06
D9546 n9547 0 dm2 AREA=1.097e-06
D9547 n9548 0 dm2 AREA=1.864e-06
D9548 n9549 0 dm2 AREA=9.513e-07
D9549 n9550 0 dm2 AREA=1.146e-06
D9550 n9551 0 dm2 AREA=1.317e-06
D9551 n9552 0 dm2 AREA=5.920e-07
D9552 n9553 0 dm2 AREA=5.551e-07
D9553 n9554 0 dm2 AREA=5.016e-07
D9554 n9555 0 dm2 AREA=6.088e-07
D9555 n9556 0 dm2 AREA=3.976e-07
D9556 n9557 0 dm2 AREA=3.396e-07
D9557 n9558 0 dm2 AREA=9.007e-07
D9558 n9559 0 dm2 AREA=1.675e-06
D9559 n9560 0 dm2 AREA=1.837e-06
D9560 n9561 0 dm2 AREA=1.150e-06
D9561 n9562 0 dm2 AREA=1.023e-06
D9562 n9563 0 dm2 AREA=1.431e-06
D9563 n9564 0 dm2 AREA=9.924e-07
D9564 n9565 0 dm2 AREA=1.052e-06
D9565 n9566 0 dm2 AREA=2.047e-06
D9566 n9567 0 dm2 AREA=1.060e-06
D9567 n9568 0 dm2 AREA=2.610e-06
D9568 n9569 0 dm2 AREA=7.388e-07
D9569 n9570 0 dm2 AREA=1.067e-06
D9570 n9571 0 dm2 AREA=8.288e-07
D9571 n9572 0 dm2 AREA=4.478e-07
D9572 n9573 0 dm2 AREA=1.655e-06
D9573 n9574 0 dm2 AREA=6.132e-07
D9574 n9575 0 dm2 AREA=4.920e-07
D9575 n9576 0 dm2 AREA=5.715e-07
D9576 n9577 0 dm2 AREA=7.866e-07
D9577 n9578 0 dm2 AREA=1.138e-06
D9578 n9579 0 dm2 AREA=1.030e-06
D9579 n9580 0 dm2 AREA=1.506e-06
D9580 n9581 0 dm2 AREA=1.267e-06
D9581 n9582 0 dm2 AREA=7.889e-07
D9582 n9583 0 dm2 AREA=8.314e-07
D9583 n9584 0 dm2 AREA=1.004e-06
D9584 n9585 0 dm2 AREA=8.009e-07
D9585 n9586 0 dm2 AREA=7.611e-07
D9586 n9587 0 dm2 AREA=4.170e-07
D9587 n9588 0 dm2 AREA=1.871e-06
D9588 n9589 0 dm2 AREA=9.054e-07
D9589 n9590 0 dm2 AREA=1.432e-06
D9590 n9591 0 dm2 AREA=1.533e-06
D9591 n9592 0 dm2 AREA=5.691e-07
D9592 n9593 0 dm2 AREA=8.998e-07
D9593 n9594 0 dm2 AREA=7.398e-07
D9594 n9595 0 dm2 AREA=1.034e-06
D9595 n9596 0 dm2 AREA=7.818e-07
D9596 n9597 0 dm2 AREA=5.203e-07
D9597 n9598 0 dm2 AREA=8.172e-07
D9598 n9599 0 dm2 AREA=8.415e-07
D9599 n9600 0 dm2 AREA=5.248e-07
D9600 n9601 0 dm2 AREA=1.139e-06
D9601 n9602 0 dm2 AREA=1.373e-06
D9602 n9603 0 dm2 AREA=9.635e-07
D9603 n9604 0 dm2 AREA=7.291e-07
D9604 n9605 0 dm2 AREA=9.277e-07
D9605 n9606 0 dm2 AREA=1.231e-06
D9606 n9607 0 dm2 AREA=8.469e-07
D9607 n9608 0 dm2 AREA=1.300e-06
D9608 n9609 0 dm2 AREA=6.015e-07
D9609 n9610 0 dm2 AREA=5.326e-07
D9610 n9611 0 dm2 AREA=9.348e-07
D9611 n9612 0 dm2 AREA=7.769e-07
D9612 n9613 0 dm2 AREA=9.402e-07
D9613 n9614 0 dm2 AREA=8.846e-07
D9614 n9615 0 dm2 AREA=8.852e-07
D9615 n9616 0 dm2 AREA=6.610e-07
D9616 n9617 0 dm2 AREA=1.097e-06
D9617 n9618 0 dm2 AREA=3.541e-07
D9618 n9619 0 dm2 AREA=1.657e-06
D9619 n9620 0 dm2 AREA=1.480e-06
D9620 n9621 0 dm2 AREA=8.351e-07
D9621 n9622 0 dm2 AREA=1.346e-06
D9622 n9623 0 dm2 AREA=6.994e-07
D9623 n9624 0 dm2 AREA=1.522e-06
D9624 n9625 0 dm2 AREA=9.017e-07
D9625 n9626 0 dm2 AREA=1.305e-06
D9626 n9627 0 dm2 AREA=1.050e-06
D9627 n9628 0 dm2 AREA=7.879e-07
D9628 n9629 0 dm2 AREA=4.125e-07
D9629 n9630 0 dm2 AREA=9.480e-07
D9630 n9631 0 dm2 AREA=8.513e-07
D9631 n9632 0 dm2 AREA=1.032e-06
D9632 n9633 0 dm2 AREA=1.223e-06
D9633 n9634 0 dm2 AREA=4.641e-07
D9634 n9635 0 dm2 AREA=1.153e-06
D9635 n9636 0 dm2 AREA=1.725e-06
D9636 n9637 0 dm2 AREA=4.619e-07
D9637 n9638 0 dm2 AREA=6.284e-07
D9638 n9639 0 dm2 AREA=1.666e-07
D9639 n9640 0 dm2 AREA=6.907e-07
D9640 n9641 0 dm2 AREA=8.435e-07
D9641 n9642 0 dm2 AREA=1.141e-06
D9642 n9643 0 dm2 AREA=4.235e-07
D9643 n9644 0 dm2 AREA=6.501e-07
D9644 n9645 0 dm2 AREA=8.644e-07
D9645 n9646 0 dm2 AREA=8.490e-07
D9646 n9647 0 dm2 AREA=3.355e-07
D9647 n9648 0 dm2 AREA=2.073e-07
D9648 n9649 0 dm2 AREA=1.876e-06
D9649 n9650 0 dm2 AREA=7.931e-07
D9650 n9651 0 dm2 AREA=1.499e-06
D9651 n9652 0 dm2 AREA=5.959e-07
D9652 n9653 0 dm2 AREA=1.234e-06
D9653 n9654 0 dm2 AREA=1.266e-07
D9654 n9655 0 dm2 AREA=7.865e-07
D9655 n9656 0 dm2 AREA=1.410e-06
D9656 n9657 0 dm2 AREA=8.365e-07
D9657 n9658 0 dm2 AREA=2.736e-07
D9658 n9659 0 dm2 AREA=5.500e-07
D9659 n9660 0 dm2 AREA=5.077e-07
D9660 n9661 0 dm2 AREA=2.851e-06
D9661 n9662 0 dm2 AREA=3.874e-07
D9662 n9663 0 dm2 AREA=1.899e-07
D9663 n9664 0 dm2 AREA=1.124e-06
D9664 n9665 0 dm2 AREA=9.594e-07
D9665 n9666 0 dm2 AREA=1.198e-06
D9666 n9667 0 dm2 AREA=3.388e-07
D9667 n9668 0 dm2 AREA=7.647e-07
D9668 n9669 0 dm2 AREA=1.153e-06
D9669 n9670 0 dm2 AREA=1.519e-06
D9670 n9671 0 dm2 AREA=9.150e-07
D9671 n9672 0 dm2 AREA=2.656e-07
D9672 n9673 0 dm2 AREA=5.401e-07
D9673 n9674 0 dm2 AREA=1.041e-06
D9674 n9675 0 dm2 AREA=6.627e-07
D9675 n9676 0 dm2 AREA=1.828e-06
D9676 n9677 0 dm2 AREA=1.393e-06
D9677 n9678 0 dm2 AREA=7.512e-07
D9678 n9679 0 dm2 AREA=1.307e-06
D9679 n9680 0 dm2 AREA=1.295e-06
D9680 n9681 0 dm2 AREA=1.027e-06
D9681 n9682 0 dm2 AREA=1.021e-06
D9682 n9683 0 dm2 AREA=1.589e-06
D9683 n9684 0 dm2 AREA=1.120e-06
D9684 n9685 0 dm2 AREA=6.454e-07
D9685 n9686 0 dm2 AREA=7.855e-07
D9686 n9687 0 dm2 AREA=3.530e-07
D9687 n9688 0 dm2 AREA=6.499e-07
D9688 n9689 0 dm2 AREA=9.164e-07
D9689 n9690 0 dm2 AREA=8.907e-07
D9690 n9691 0 dm2 AREA=6.591e-07
D9691 n9692 0 dm2 AREA=3.735e-07
D9692 n9693 0 dm2 AREA=7.748e-07
D9693 n9694 0 dm14 AREA=3.488e-07

*** current source definition
I2 0 n3 3.361e-02A M=4.190e-07
I3 0 n4 3.361e-02A M=3.064e-07
I4 0 n5 3.361e-02A M=5.062e-07
I5 0 n6 3.361e-02A M=2.541e-07
I6 0 n7 3.361e-02A M=4.298e-07
I7 0 n8 3.361e-02A M=8.625e-07
I8 0 n9 3.361e-02A M=9.339e-07
I9 0 n10 3.361e-02A M=5.878e-07
I10 0 n11 3.361e-02A M=1.559e-06
I11 0 n12 3.361e-02A M=1.225e-06
I12 0 n13 3.361e-02A M=1.127e-06
I13 0 n14 3.361e-02A M=6.810e-07
I14 0 n15 3.361e-02A M=9.285e-07
I15 0 n16 3.361e-02A M=1.314e-06
I16 0 n17 3.361e-02A M=6.018e-07
I17 0 n18 3.361e-02A M=1.235e-06
I18 0 n19 3.361e-02A M=2.556e-07
I19 0 n20 3.361e-02A M=4.861e-07
I20 0 n21 3.361e-02A M=1.103e-06
I21 0 n22 3.361e-02A M=5.660e-07
I22 0 n23 3.361e-02A M=4.605e-07
I23 0 n24 3.361e-02A M=6.236e-07
I24 0 n25 3.361e-02A M=6.088e-07
I25 0 n26 3.361e-02A M=1.298e-06
I26 0 n27 3.361e-02A M=7.569e-07
I27 0 n28 3.361e-02A M=3.530e-07
I28 0 n29 3.361e-02A M=4.491e-07
I29 0 n30 3.361e-02A M=6.631e-07
I30 0 n31 3.361e-02A M=1.128e-06
I31 0 n32 3.361e-02A M=8.167e-07
I32 0 n33 3.361e-02A M=7.455e-07
I33 0 n34 3.361e-02A M=7.323e-07
I34 0 n35 3.361e-02A M=9.119e-07
I35 0 n36 3.361e-02A M=4.246e-07
I36 0 n37 3.361e-02A M=7.176e-07
I37 0 n38 3.361e-02A M=1.426e-06
I38 0 n39 3.361e-02A M=1.314e-06
I39 0 n40 3.361e-02A M=1.214e-06
I40 0 n41 3.361e-02A M=1.936e-06
I41 0 n42 3.361e-02A M=6.377e-07
I42 0 n43 3.361e-02A M=9.413e-07
I43 0 n44 3.361e-02A M=7.136e-07
I44 0 n45 3.361e-02A M=1.331e-06
I45 0 n46 3.361e-02A M=7.655e-07
I46 0 n47 3.361e-02A M=7.247e-07
I47 0 n48 3.361e-02A M=2.307e-07
I48 0 n49 3.361e-02A M=1.277e-06
I49 0 n50 3.361e-02A M=2.119e-06
I50 0 n51 3.361e-02A M=7.286e-07
I51 0 n52 3.361e-02A M=4.096e-07
I52 0 n53 3.361e-02A M=4.957e-07
I53 0 n54 3.361e-02A M=6.202e-07
I54 0 n55 3.361e-02A M=8.884e-07
I55 0 n56 3.361e-02A M=1.846e-06
I56 0 n57 3.361e-02A M=5.088e-07
I57 0 n58 3.361e-02A M=1.370e-06
I58 0 n59 3.361e-02A M=9.885e-07
I59 0 n60 3.361e-02A M=7.307e-07
I60 0 n61 3.361e-02A M=1.574e-06
I61 0 n62 3.361e-02A M=4.701e-07
I62 0 n63 3.361e-02A M=3.521e-07
I63 0 n64 3.361e-02A M=1.134e-06
I64 0 n65 3.361e-02A M=6.607e-07
I65 0 n66 3.361e-02A M=6.719e-07
I66 0 n67 3.361e-02A M=2.565e-06
I67 0 n68 3.361e-02A M=3.700e-07
I68 0 n69 3.361e-02A M=1.314e-06
I69 0 n70 3.361e-02A M=1.633e-06
I70 0 n71 3.361e-02A M=1.193e-06
I71 0 n72 3.361e-02A M=8.711e-07
I72 0 n73 3.361e-02A M=6.286e-07
I73 0 n74 3.361e-02A M=3.611e-07
I74 0 n75 3.361e-02A M=1.399e-06
I75 0 n76 3.361e-02A M=1.387e-06
I76 0 n77 3.361e-02A M=1.630e-06
I77 0 n78 3.361e-02A M=6.776e-07
I78 0 n79 3.361e-02A M=1.236e-06
I79 0 n80 3.361e-02A M=6.540e-07
I80 0 n81 3.361e-02A M=9.424e-07
I81 0 n82 3.361e-02A M=1.068e-06
I82 0 n83 3.361e-02A M=8.713e-07
I83 0 n84 3.361e-02A M=1.235e-06
I84 0 n85 3.361e-02A M=1.127e-06
I85 0 n86 3.361e-02A M=9.646e-07
I86 0 n87 3.361e-02A M=5.929e-07
I87 0 n88 3.361e-02A M=8.341e-07
I88 0 n89 3.361e-02A M=4.546e-07
I89 0 n90 3.361e-02A M=1.055e-06
I90 0 n91 3.361e-02A M=8.806e-07
I91 0 n92 3.361e-02A M=7.549e-07
I92 0 n93 3.361e-02A M=6.124e-07
I93 0 n94 3.361e-02A M=1.046e-06
I94 0 n95 3.361e-02A M=7.094e-07
I95 0 n96 3.361e-02A M=7.010e-07
I96 0 n97 3.361e-02A M=9.498e-07
I97 0 n98 3.361e-02A M=6.611e-07
I98 0 n99 3.361e-02A M=1.736e-06
I99 0 n100 3.361e-02A M=1.062e-06
I100 0 n101 3.361e-02A M=5.478e-07
I101 0 n102 3.361e-02A M=1.304e-06
I102 0 n103 3.361e-02A M=1.498e-06
I103 0 n104 3.361e-02A M=9.375e-07
I104 0 n105 3.361e-02A M=1.111e-06
I105 0 n106 3.361e-02A M=6.419e-07
I106 0 n107 3.361e-02A M=7.029e-07
I107 0 n108 3.361e-02A M=1.010e-06
I108 0 n109 3.361e-02A M=2.309e-06
I109 0 n110 3.361e-02A M=1.723e-06
I110 0 n111 3.361e-02A M=1.128e-06
I111 0 n112 3.361e-02A M=8.483e-07
I112 0 n113 3.361e-02A M=1.161e-06
I113 0 n114 3.361e-02A M=9.833e-07
I114 0 n115 3.361e-02A M=7.142e-07
I115 0 n116 3.361e-02A M=1.951e-06
I116 0 n117 3.361e-02A M=9.904e-07
I117 0 n118 3.361e-02A M=1.572e-06
I118 0 n119 3.361e-02A M=9.237e-07
I119 0 n120 3.361e-02A M=9.627e-07
I120 0 n121 3.361e-02A M=7.365e-07
I121 0 n122 3.361e-02A M=1.908e-06
I122 0 n123 3.361e-02A M=1.114e-06
I123 0 n124 3.361e-02A M=5.429e-07
I124 0 n125 3.361e-02A M=8.227e-07
I125 0 n126 3.361e-02A M=5.163e-07
I126 0 n127 3.361e-02A M=9.082e-07
I127 0 n128 3.361e-02A M=1.799e-06
I128 0 n129 3.361e-02A M=7.372e-07
I129 0 n130 3.361e-02A M=1.142e-06
I130 0 n131 3.361e-02A M=2.547e-07
I131 0 n132 3.361e-02A M=2.459e-06
I132 0 n133 3.361e-02A M=1.634e-06
I133 0 n134 3.361e-02A M=6.828e-07
I134 0 n135 3.361e-02A M=1.258e-06
I135 0 n136 3.361e-02A M=9.633e-07
I136 0 n137 3.361e-02A M=1.437e-06
I137 0 n138 3.361e-02A M=9.349e-07
I138 0 n139 3.361e-02A M=1.189e-06
I139 0 n140 3.361e-02A M=6.119e-07
I140 0 n141 3.361e-02A M=6.820e-07
I141 0 n142 3.361e-02A M=3.288e-07
I142 0 n143 3.361e-02A M=7.578e-07
I143 0 n144 3.361e-02A M=1.446e-06
I144 0 n145 3.361e-02A M=9.524e-07
I145 0 n146 3.361e-02A M=7.706e-07
I146 0 n147 3.361e-02A M=7.518e-07
I147 0 n148 3.361e-02A M=1.021e-06
I148 0 n149 3.361e-02A M=2.872e-07
I149 0 n150 3.361e-02A M=1.280e-06
I150 0 n151 3.361e-02A M=7.318e-07
I151 0 n152 3.361e-02A M=6.110e-07
I152 0 n153 3.361e-02A M=3.461e-07
I153 0 n154 3.361e-02A M=1.031e-06
I154 0 n155 3.361e-02A M=1.276e-06
I155 0 n156 3.361e-02A M=1.061e-06
I156 0 n157 3.361e-02A M=1.520e-06
I157 0 n158 3.361e-02A M=2.784e-07
I158 0 n159 3.361e-02A M=8.815e-07
I159 0 n160 3.361e-02A M=1.736e-06
I160 0 n161 3.361e-02A M=7.552e-07
I161 0 n162 3.361e-02A M=1.031e-06
I162 0 n163 3.361e-02A M=9.168e-07
I163 0 n164 3.361e-02A M=1.022e-06
I164 0 n165 3.361e-02A M=1.863e-06
I165 0 n166 3.361e-02A M=1.403e-07
I166 0 n167 3.361e-02A M=7.623e-07
I167 0 n168 3.361e-02A M=1.116e-06
I168 0 n169 3.361e-02A M=6.604e-07
I169 0 n170 3.361e-02A M=7.253e-07
I170 0 n171 3.361e-02A M=8.543e-07
I171 0 n172 3.361e-02A M=8.213e-07
I172 0 n173 3.361e-02A M=1.388e-06
I173 0 n174 3.361e-02A M=7.550e-07
I174 0 n1 3.361e-02A M=3.116e-07
I175 0 n176 3.361e-02A M=1.088e-06
I176 0 n177 3.361e-02A M=6.280e-07
I177 0 n178 3.361e-02A M=8.084e-07
I178 0 n179 3.361e-02A M=2.384e-06
I179 0 n180 3.361e-02A M=6.449e-07
I180 0 n181 3.361e-02A M=6.942e-07
I181 0 n182 3.361e-02A M=1.509e-06
I182 0 n183 3.361e-02A M=9.229e-07
I183 0 n184 3.361e-02A M=1.682e-06
I184 0 n185 3.361e-02A M=1.518e-06
I185 0 n186 3.361e-02A M=4.404e-07
I186 0 n187 3.361e-02A M=6.991e-07
I187 0 n188 3.361e-02A M=5.162e-07
I188 0 n189 3.361e-02A M=5.656e-07
I189 0 n190 3.361e-02A M=8.403e-07
I190 0 n191 3.361e-02A M=8.540e-07
I191 0 n192 3.361e-02A M=9.868e-07
I192 0 n193 3.361e-02A M=8.153e-07
I193 0 n194 3.361e-02A M=9.817e-07
I194 0 n195 3.361e-02A M=1.354e-06
I195 0 n196 3.361e-02A M=7.490e-07
I196 0 n197 3.361e-02A M=1.812e-06
I197 0 n198 3.361e-02A M=6.654e-07
I198 0 n199 3.361e-02A M=7.075e-07
I199 0 n200 3.361e-02A M=4.573e-07
I200 0 n201 3.361e-02A M=5.507e-07
I201 0 n202 3.361e-02A M=8.823e-07
I202 0 n203 3.361e-02A M=6.509e-07
I203 0 n204 3.361e-02A M=1.134e-06
I204 0 n205 3.361e-02A M=9.513e-07
I205 0 n206 3.361e-02A M=9.713e-07
I206 0 n207 3.361e-02A M=2.493e-07
I207 0 n208 3.361e-02A M=6.778e-07
I208 0 n209 3.361e-02A M=4.802e-07
I209 0 n210 3.361e-02A M=1.116e-06
I210 0 n211 3.361e-02A M=6.809e-07
I211 0 n212 3.361e-02A M=1.257e-06
I212 0 n213 3.361e-02A M=4.486e-07
I213 0 n214 3.361e-02A M=6.301e-07
I214 0 n215 3.361e-02A M=6.827e-07
I215 0 n216 3.361e-02A M=1.134e-06
I216 0 n217 3.361e-02A M=5.581e-07
I217 0 n218 3.361e-02A M=9.403e-07
I218 0 n219 3.361e-02A M=2.426e-06
I219 0 n220 3.361e-02A M=1.740e-06
I220 0 n221 3.361e-02A M=7.440e-07
I221 0 n222 3.361e-02A M=6.907e-07
I222 0 n223 3.361e-02A M=7.625e-07
I223 0 n224 3.361e-02A M=1.246e-06
I224 0 n225 3.361e-02A M=8.199e-07
I225 0 n226 3.361e-02A M=2.846e-07
I226 0 n227 3.361e-02A M=1.329e-06
I227 0 n228 3.361e-02A M=8.607e-07
I228 0 n229 3.361e-02A M=4.208e-07
I229 0 n230 3.361e-02A M=1.091e-06
I230 0 n231 3.361e-02A M=7.345e-07
I231 0 n1 3.361e-02A M=5.216e-07
I232 0 n233 3.361e-02A M=8.843e-07
I233 0 n234 3.361e-02A M=9.722e-07
I234 0 n235 3.361e-02A M=5.683e-07
I235 0 n236 3.361e-02A M=1.589e-06
I236 0 n237 3.361e-02A M=1.701e-06
I237 0 n238 3.361e-02A M=6.146e-07
I238 0 n239 3.361e-02A M=4.949e-07
I239 0 n240 3.361e-02A M=8.789e-07
I240 0 n241 3.361e-02A M=5.355e-07
I241 0 n242 3.361e-02A M=8.667e-07
I242 0 n243 3.361e-02A M=1.357e-06
I243 0 n244 3.361e-02A M=1.330e-06
I244 0 n245 3.361e-02A M=2.681e-06
I245 0 n246 3.361e-02A M=3.731e-07
I246 0 n247 3.361e-02A M=4.759e-07
I247 0 n248 3.361e-02A M=5.027e-07
I248 0 n249 3.361e-02A M=6.673e-07
I249 0 n250 3.361e-02A M=6.688e-07
I250 0 n251 3.361e-02A M=3.095e-07
I251 0 n252 3.361e-02A M=5.354e-07
I252 0 n253 3.361e-02A M=1.169e-06
I253 0 n254 3.361e-02A M=7.403e-07
I254 0 n255 3.361e-02A M=1.281e-06
I255 0 n256 3.361e-02A M=1.042e-06
I256 0 n257 3.361e-02A M=8.482e-07
I257 0 n258 3.361e-02A M=8.679e-07
I258 0 n259 3.361e-02A M=8.126e-07
I259 0 n260 3.361e-02A M=3.252e-07
I260 0 n261 3.361e-02A M=9.272e-07
I261 0 n262 3.361e-02A M=1.268e-06
I262 0 n263 3.361e-02A M=9.098e-07
I263 0 n264 3.361e-02A M=1.573e-06
I264 0 n265 3.361e-02A M=7.835e-07
I265 0 n266 3.361e-02A M=7.864e-07
I266 0 n267 3.361e-02A M=9.937e-07
I267 0 n268 3.361e-02A M=7.115e-07
I268 0 n269 3.361e-02A M=1.178e-06
I269 0 n270 3.361e-02A M=1.136e-06
I270 0 n271 3.361e-02A M=6.752e-07
I271 0 n272 3.361e-02A M=1.939e-06
I272 0 n273 3.361e-02A M=1.347e-06
I273 0 n274 3.361e-02A M=3.438e-07
I274 0 n275 3.361e-02A M=1.341e-06
I275 0 n276 3.361e-02A M=1.514e-06
I276 0 n277 3.361e-02A M=2.482e-07
I277 0 n278 3.361e-02A M=1.151e-06
I278 0 n1 3.361e-02A M=9.026e-07
I279 0 n280 3.361e-02A M=1.337e-06
I280 0 n281 3.361e-02A M=7.364e-07
I281 0 n282 3.361e-02A M=9.972e-07
I282 0 n283 3.361e-02A M=1.071e-06
I283 0 n284 3.361e-02A M=7.243e-07
I284 0 n285 3.361e-02A M=7.236e-07
I285 0 n286 3.361e-02A M=1.355e-06
I286 0 n287 3.361e-02A M=2.349e-07
I287 0 n288 3.361e-02A M=1.070e-06
I288 0 n289 3.361e-02A M=8.990e-07
I289 0 n290 3.361e-02A M=2.352e-07
I290 0 n291 3.361e-02A M=9.428e-07
I291 0 n292 3.361e-02A M=6.823e-07
I292 0 n293 3.361e-02A M=1.057e-06
I293 0 n294 3.361e-02A M=7.779e-07
I294 0 n295 3.361e-02A M=6.273e-07
I295 0 n296 3.361e-02A M=4.362e-07
I296 0 n297 3.361e-02A M=9.841e-07
I297 0 n298 3.361e-02A M=1.390e-06
I298 0 n299 3.361e-02A M=6.086e-07
I299 0 n300 3.361e-02A M=4.720e-07
I300 0 n301 3.361e-02A M=4.765e-07
I301 0 n302 3.361e-02A M=6.769e-07
I302 0 n303 3.361e-02A M=1.955e-06
I303 0 n304 3.361e-02A M=4.579e-07
I304 0 n305 3.361e-02A M=5.280e-07
I305 0 n306 3.361e-02A M=1.382e-06
I306 0 n307 3.361e-02A M=5.889e-07
I307 0 n308 3.361e-02A M=2.202e-07
I308 0 n309 3.361e-02A M=6.689e-07
I309 0 n310 3.361e-02A M=9.813e-07
I310 0 n311 3.361e-02A M=1.336e-06
I311 0 n312 3.361e-02A M=8.846e-07
I312 0 n313 3.361e-02A M=7.759e-07
I313 0 n314 3.361e-02A M=1.305e-06
I314 0 n315 3.361e-02A M=4.139e-07
I315 0 n1 3.361e-02A M=7.449e-07
I316 0 n317 3.361e-02A M=4.299e-07
I317 0 n318 3.361e-02A M=1.609e-06
I318 0 n319 3.361e-02A M=7.397e-07
I319 0 n320 3.361e-02A M=1.098e-06
I320 0 n321 3.361e-02A M=3.681e-07
I321 0 n322 3.361e-02A M=6.883e-07
I322 0 n323 3.361e-02A M=7.436e-07
I323 0 n324 3.361e-02A M=7.772e-07
I324 0 n325 3.361e-02A M=1.470e-06
I325 0 n326 3.361e-02A M=1.354e-06
I326 0 n327 3.361e-02A M=5.480e-07
I327 0 n328 3.361e-02A M=2.118e-06
I328 0 n329 3.361e-02A M=1.825e-06
I329 0 n330 3.361e-02A M=9.061e-07
I330 0 n331 3.361e-02A M=1.019e-06
I331 0 n332 3.361e-02A M=2.233e-06
I332 0 n333 3.361e-02A M=2.277e-06
I333 0 n334 3.361e-02A M=1.181e-06
I334 0 n335 3.361e-02A M=1.263e-06
I335 0 n336 3.361e-02A M=4.404e-07
I336 0 n337 3.361e-02A M=1.720e-06
I337 0 n338 3.361e-02A M=1.274e-06
I338 0 n339 3.361e-02A M=1.582e-06
I339 0 n340 3.361e-02A M=1.324e-06
I340 0 n341 3.361e-02A M=4.545e-07
I341 0 n342 3.361e-02A M=1.200e-06
I342 0 n343 3.361e-02A M=1.324e-06
I343 0 n344 3.361e-02A M=6.992e-07
I344 0 n345 3.361e-02A M=2.438e-07
I345 0 n346 3.361e-02A M=4.069e-07
I346 0 n347 3.361e-02A M=5.276e-07
I347 0 n348 3.361e-02A M=1.262e-06
I348 0 n349 3.361e-02A M=1.625e-06
I349 0 n350 3.361e-02A M=1.254e-06
I350 0 n351 3.361e-02A M=8.401e-07
I351 0 n352 3.361e-02A M=1.061e-06
I352 0 n353 3.361e-02A M=1.533e-06
I353 0 n354 3.361e-02A M=6.102e-07
I354 0 n355 3.361e-02A M=1.656e-06
I355 0 n356 3.361e-02A M=3.360e-07
I356 0 n357 3.361e-02A M=5.933e-07
I357 0 n358 3.361e-02A M=3.864e-07
I358 0 n359 3.361e-02A M=1.766e-06
I359 0 n360 3.361e-02A M=1.469e-06
I360 0 n361 3.361e-02A M=7.867e-07
I361 0 n362 3.361e-02A M=1.945e-06
I362 0 n363 3.361e-02A M=1.010e-06
I363 0 n364 3.361e-02A M=8.332e-07
I364 0 n365 3.361e-02A M=5.336e-07
I365 0 n366 3.361e-02A M=1.826e-06
I366 0 n367 3.361e-02A M=2.866e-06
I367 0 n368 3.361e-02A M=2.610e-06
I368 0 n369 3.361e-02A M=1.125e-06
I369 0 n370 3.361e-02A M=1.360e-06
I370 0 n371 3.361e-02A M=7.868e-07
I371 0 n372 3.361e-02A M=2.445e-06
I372 0 n373 3.361e-02A M=9.505e-07
I373 0 n374 3.361e-02A M=2.399e-06
I374 0 n375 3.361e-02A M=4.883e-07
I375 0 n376 3.361e-02A M=1.763e-06
I376 0 n377 3.361e-02A M=3.044e-07
I377 0 n378 3.361e-02A M=8.654e-07
I378 0 n379 3.361e-02A M=6.796e-07
I379 0 n380 3.361e-02A M=6.514e-07
I380 0 n381 3.361e-02A M=7.339e-07
I381 0 n382 3.361e-02A M=2.187e-06
I382 0 n383 3.361e-02A M=1.229e-06
I383 0 n384 3.361e-02A M=1.327e-06
I384 0 n385 3.361e-02A M=3.797e-07
I385 0 n386 3.361e-02A M=7.583e-07
I386 0 n387 3.361e-02A M=9.801e-07
I387 0 n388 3.361e-02A M=3.110e-07
I388 0 n389 3.361e-02A M=5.515e-07
I389 0 n390 3.361e-02A M=9.278e-07
I390 0 n391 3.361e-02A M=9.598e-07
I391 0 n392 3.361e-02A M=6.058e-07
I392 0 n393 3.361e-02A M=1.298e-06
I393 0 n394 3.361e-02A M=1.708e-06
I394 0 n395 3.361e-02A M=7.262e-07
I395 0 n396 3.361e-02A M=7.621e-07
I396 0 n397 3.361e-02A M=7.406e-07
I397 0 n398 3.361e-02A M=3.543e-07
I398 0 n1 3.361e-02A M=2.022e-06
I399 0 n400 3.361e-02A M=9.956e-07
I400 0 n401 3.361e-02A M=6.255e-07
I401 0 n402 3.361e-02A M=2.440e-06
I402 0 n403 3.361e-02A M=1.041e-06
I403 0 n404 3.361e-02A M=1.239e-06
I404 0 n405 3.361e-02A M=1.294e-06
I405 0 n406 3.361e-02A M=5.010e-07
I406 0 n407 3.361e-02A M=6.876e-07
I407 0 n408 3.361e-02A M=5.898e-07
I408 0 n409 3.361e-02A M=7.510e-07
I409 0 n410 3.361e-02A M=1.159e-06
I410 0 n411 3.361e-02A M=5.910e-07
I411 0 n412 3.361e-02A M=9.142e-07
I412 0 n413 3.361e-02A M=1.595e-06
I413 0 n414 3.361e-02A M=1.823e-07
I414 0 n415 3.361e-02A M=1.948e-06
I415 0 n416 3.361e-02A M=4.165e-07
I416 0 n417 3.361e-02A M=5.817e-07
I417 0 n418 3.361e-02A M=8.565e-07
I418 0 n419 3.361e-02A M=4.761e-07
I419 0 n420 3.361e-02A M=4.035e-07
I420 0 n421 3.361e-02A M=1.128e-06
I421 0 n422 3.361e-02A M=1.595e-07
I422 0 n423 3.361e-02A M=2.733e-06
I423 0 n424 3.361e-02A M=2.891e-06
I424 0 n425 3.361e-02A M=1.096e-06
I425 0 n426 3.361e-02A M=1.094e-06
I426 0 n427 3.361e-02A M=7.784e-07
I427 0 n428 3.361e-02A M=1.669e-06
I428 0 n429 3.361e-02A M=1.020e-06
I429 0 n430 3.361e-02A M=1.547e-06
I430 0 n431 3.361e-02A M=8.184e-07
I431 0 n432 3.361e-02A M=6.470e-07
I432 0 n433 3.361e-02A M=6.844e-07
I433 0 n434 3.361e-02A M=1.030e-06
I434 0 n435 3.361e-02A M=9.088e-07
I435 0 n436 3.361e-02A M=1.017e-06
I436 0 n437 3.361e-02A M=8.821e-07
I437 0 n438 3.361e-02A M=1.395e-06
I438 0 n439 3.361e-02A M=5.393e-07
I439 0 n440 3.361e-02A M=7.949e-07
I440 0 n441 3.361e-02A M=1.985e-06
I441 0 n442 3.361e-02A M=1.463e-07
I442 0 n443 3.361e-02A M=1.672e-06
I443 0 n444 3.361e-02A M=1.318e-06
I444 0 n445 3.361e-02A M=1.108e-06
I445 0 n446 3.361e-02A M=5.204e-07
I446 0 n447 3.361e-02A M=1.397e-06
I447 0 n448 3.361e-02A M=1.727e-06
I448 0 n449 3.361e-02A M=4.613e-07
I449 0 n450 3.361e-02A M=5.923e-07
I450 0 n451 3.361e-02A M=1.643e-06
I451 0 n452 3.361e-02A M=4.584e-07
I452 0 n453 3.361e-02A M=1.333e-06
I453 0 n454 3.361e-02A M=9.004e-07
I454 0 n455 3.361e-02A M=3.383e-07
I455 0 n456 3.361e-02A M=8.690e-07
I456 0 n457 3.361e-02A M=1.395e-06
I457 0 n458 3.361e-02A M=1.516e-06
I458 0 n459 3.361e-02A M=3.992e-07
I459 0 n460 3.361e-02A M=1.329e-06
I460 0 n461 3.361e-02A M=9.907e-07
I461 0 n462 3.361e-02A M=1.011e-06
I462 0 n463 3.361e-02A M=2.384e-07
I463 0 n464 3.361e-02A M=1.321e-06
I464 0 n465 3.361e-02A M=2.070e-07
I465 0 n466 3.361e-02A M=8.158e-07
I466 0 n467 3.361e-02A M=9.289e-07
I467 0 n468 3.361e-02A M=9.012e-07
I468 0 n469 3.361e-02A M=8.395e-07
I469 0 n470 3.361e-02A M=1.493e-06
I470 0 n471 3.361e-02A M=1.527e-06
I471 0 n472 3.361e-02A M=1.243e-06
I472 0 n473 3.361e-02A M=1.916e-06
I473 0 n474 3.361e-02A M=4.917e-07
I474 0 n475 3.361e-02A M=5.112e-07
I475 0 n476 3.361e-02A M=4.157e-07
I476 0 n477 3.361e-02A M=2.187e-06
I477 0 n478 3.361e-02A M=8.166e-07
I478 0 n479 3.361e-02A M=1.621e-06
I479 0 n480 3.361e-02A M=7.468e-07
I480 0 n481 3.361e-02A M=4.014e-07
I481 0 n482 3.361e-02A M=1.442e-06
I482 0 n483 3.361e-02A M=3.818e-07
I483 0 n1 3.361e-02A M=1.741e-06
I484 0 n485 3.361e-02A M=1.495e-06
I485 0 n486 3.361e-02A M=2.334e-06
I486 0 n487 3.361e-02A M=6.252e-07
I487 0 n488 3.361e-02A M=9.676e-07
I488 0 n489 3.361e-02A M=1.114e-06
I489 0 n490 3.361e-02A M=1.564e-07
I490 0 n491 3.361e-02A M=2.065e-07
I491 0 n492 3.361e-02A M=5.031e-07
I492 0 n493 3.361e-02A M=2.327e-07
I493 0 n494 3.361e-02A M=9.968e-07
I494 0 n495 3.361e-02A M=7.256e-07
I495 0 n496 3.361e-02A M=8.804e-07
I496 0 n497 3.361e-02A M=6.504e-07
I497 0 n498 3.361e-02A M=7.260e-07
I498 0 n499 3.361e-02A M=5.206e-07
I499 0 n500 3.361e-02A M=7.546e-07
I500 0 n501 3.361e-02A M=1.110e-06
I501 0 n502 3.361e-02A M=5.420e-07
I502 0 n503 3.361e-02A M=5.765e-07
I503 0 n504 3.361e-02A M=1.127e-06
I504 0 n505 3.361e-02A M=1.644e-06
I505 0 n506 3.361e-02A M=6.800e-07
I506 0 n507 3.361e-02A M=1.084e-06
I507 0 n508 3.361e-02A M=8.842e-07
I508 0 n509 3.361e-02A M=1.732e-06
I509 0 n510 3.361e-02A M=6.401e-07
I510 0 n511 3.361e-02A M=1.119e-06
I511 0 n512 3.361e-02A M=6.554e-07
I512 0 n513 3.361e-02A M=1.146e-06
I513 0 n514 3.361e-02A M=5.660e-07
I514 0 n515 3.361e-02A M=7.115e-07
I515 0 n516 3.361e-02A M=3.132e-07
I516 0 n517 3.361e-02A M=7.536e-07
I517 0 n518 3.361e-02A M=4.545e-07
I518 0 n519 3.361e-02A M=6.963e-07
I519 0 n520 3.361e-02A M=1.551e-06
I520 0 n521 3.361e-02A M=6.956e-07
I521 0 n522 3.361e-02A M=4.249e-07
I522 0 n523 3.361e-02A M=2.653e-06
I523 0 n524 3.361e-02A M=4.144e-07
I524 0 n525 3.361e-02A M=1.132e-06
I525 0 n526 3.361e-02A M=4.858e-07
I526 0 n527 3.361e-02A M=1.065e-06
I527 0 n528 3.361e-02A M=5.348e-07
I528 0 n529 3.361e-02A M=1.303e-06
I529 0 n530 3.361e-02A M=9.905e-07
I530 0 n531 3.361e-02A M=2.518e-06
I531 0 n532 3.361e-02A M=3.039e-07
I532 0 n533 3.361e-02A M=2.148e-06
I533 0 n534 3.361e-02A M=1.418e-06
I534 0 n535 3.361e-02A M=3.358e-07
I535 0 n536 3.361e-02A M=1.002e-06
I536 0 n537 3.361e-02A M=2.771e-06
I537 0 n538 3.361e-02A M=1.420e-06
I538 0 n539 3.361e-02A M=8.497e-07
I539 0 n540 3.361e-02A M=6.195e-07
I540 0 n541 3.361e-02A M=7.575e-07
I541 0 n542 3.361e-02A M=5.202e-07
I542 0 n543 3.361e-02A M=1.725e-06
I543 0 n544 3.361e-02A M=1.543e-06
I544 0 n545 3.361e-02A M=1.047e-06
I545 0 n546 3.361e-02A M=1.214e-06
I546 0 n547 3.361e-02A M=7.092e-07
I547 0 n548 3.361e-02A M=1.039e-06
I548 0 n549 3.361e-02A M=8.370e-07
I549 0 n550 3.361e-02A M=1.026e-06
I550 0 n551 3.361e-02A M=1.716e-06
I551 0 n552 3.361e-02A M=1.060e-06
I552 0 n553 3.361e-02A M=1.036e-06
I553 0 n554 3.361e-02A M=8.584e-07
I554 0 n555 3.361e-02A M=1.142e-06
I555 0 n556 3.361e-02A M=2.729e-07
I556 0 n557 3.361e-02A M=1.723e-06
I557 0 n558 3.361e-02A M=1.134e-06
I558 0 n559 3.361e-02A M=8.916e-07
I559 0 n560 3.361e-02A M=1.157e-06
I560 0 n561 3.361e-02A M=1.700e-06
I561 0 n562 3.361e-02A M=5.669e-07
I562 0 n563 3.361e-02A M=1.389e-06
I563 0 n564 3.361e-02A M=8.302e-07
I564 0 n565 3.361e-02A M=3.631e-07
I565 0 n566 3.361e-02A M=1.395e-06
I566 0 n567 3.361e-02A M=8.817e-07
I567 0 n568 3.361e-02A M=1.328e-06
I568 0 n569 3.361e-02A M=1.430e-07
I569 0 n570 3.361e-02A M=1.166e-06
I570 0 n571 3.361e-02A M=3.760e-07
I571 0 n572 3.361e-02A M=3.458e-07
I572 0 n573 3.361e-02A M=1.021e-06
I573 0 n574 3.361e-02A M=1.208e-06
I574 0 n575 3.361e-02A M=6.848e-07
I575 0 n576 3.361e-02A M=1.041e-06
I576 0 n577 3.361e-02A M=1.532e-06
I577 0 n578 3.361e-02A M=2.659e-07
I578 0 n579 3.361e-02A M=1.078e-06
I579 0 n580 3.361e-02A M=1.701e-06
I580 0 n581 3.361e-02A M=2.596e-06
I581 0 n582 3.361e-02A M=6.833e-07
I582 0 n583 3.361e-02A M=1.255e-06
I583 0 n584 3.361e-02A M=1.144e-06
I584 0 n585 3.361e-02A M=1.042e-06
I585 0 n586 3.361e-02A M=9.609e-07
I586 0 n587 3.361e-02A M=1.201e-06
I587 0 n588 3.361e-02A M=7.061e-07
I588 0 n589 3.361e-02A M=4.006e-07
I589 0 n590 3.361e-02A M=7.860e-07
I590 0 n591 3.361e-02A M=1.772e-06
I591 0 n592 3.361e-02A M=2.688e-07
I592 0 n593 3.361e-02A M=1.070e-06
I593 0 n594 3.361e-02A M=1.358e-06
I594 0 n595 3.361e-02A M=1.045e-06
I595 0 n596 3.361e-02A M=1.221e-06
I596 0 n597 3.361e-02A M=9.846e-07
I597 0 n598 3.361e-02A M=8.173e-07
I598 0 n599 3.361e-02A M=5.454e-07
I599 0 n600 3.361e-02A M=5.407e-07
I600 0 n601 3.361e-02A M=7.823e-07
I601 0 n602 3.361e-02A M=1.302e-06
I602 0 n603 3.361e-02A M=9.015e-07
I603 0 n604 3.361e-02A M=3.196e-07
I604 0 n605 3.361e-02A M=1.333e-06
I605 0 n606 3.361e-02A M=1.468e-06
I606 0 n607 3.361e-02A M=1.006e-06
I607 0 n608 3.361e-02A M=7.249e-07
I608 0 n609 3.361e-02A M=1.080e-06
I609 0 n610 3.361e-02A M=5.515e-07
I610 0 n611 3.361e-02A M=1.474e-07
I611 0 n612 3.361e-02A M=1.182e-06
I612 0 n613 3.361e-02A M=8.533e-07
I613 0 n614 3.361e-02A M=1.245e-06
I614 0 n615 3.361e-02A M=9.486e-07
I615 0 n616 3.361e-02A M=4.132e-07
I616 0 n617 3.361e-02A M=2.537e-06
I617 0 n618 3.361e-02A M=1.319e-06
I618 0 n619 3.361e-02A M=1.278e-06
I619 0 n620 3.361e-02A M=7.625e-07
I620 0 n621 3.361e-02A M=6.512e-07
I621 0 n622 3.361e-02A M=4.605e-07
I622 0 n623 3.361e-02A M=1.017e-06
I623 0 n624 3.361e-02A M=7.482e-07
I624 0 n625 3.361e-02A M=6.140e-07
I625 0 n626 3.361e-02A M=9.329e-07
I626 0 n627 3.361e-02A M=2.441e-07
I627 0 n628 3.361e-02A M=6.617e-07
I628 0 n629 3.361e-02A M=5.607e-07
I629 0 n630 3.361e-02A M=1.689e-06
I630 0 n631 3.361e-02A M=4.120e-07
I631 0 n632 3.361e-02A M=1.529e-06
I632 0 n633 3.361e-02A M=4.789e-07
I633 0 n634 3.361e-02A M=6.100e-07
I634 0 n635 3.361e-02A M=2.032e-06
I635 0 n636 3.361e-02A M=8.097e-07
I636 0 n637 3.361e-02A M=4.979e-07
I637 0 n638 3.361e-02A M=6.579e-07
I638 0 n639 3.361e-02A M=2.312e-06
I639 0 n640 3.361e-02A M=8.503e-07
I640 0 n641 3.361e-02A M=8.522e-07
I641 0 n642 3.361e-02A M=1.832e-06
I642 0 n643 3.361e-02A M=6.469e-07
I643 0 n644 3.361e-02A M=1.411e-06
I644 0 n645 3.361e-02A M=4.632e-07
I645 0 n646 3.361e-02A M=4.822e-07
I646 0 n647 3.361e-02A M=2.553e-06
I647 0 n648 3.361e-02A M=1.207e-06
I648 0 n649 3.361e-02A M=1.278e-06
I649 0 n650 3.361e-02A M=2.471e-06
I650 0 n651 3.361e-02A M=8.734e-07
I651 0 n652 3.361e-02A M=8.160e-07
I652 0 n653 3.361e-02A M=6.939e-07
I653 0 n654 3.361e-02A M=1.272e-06
I654 0 n655 3.361e-02A M=8.753e-07
I655 0 n656 3.361e-02A M=4.091e-07
I656 0 n657 3.361e-02A M=8.357e-07
I657 0 n658 3.361e-02A M=4.424e-07
I658 0 n659 3.361e-02A M=6.915e-07
I659 0 n660 3.361e-02A M=1.832e-06
I660 0 n661 3.361e-02A M=1.621e-06
I661 0 n662 3.361e-02A M=5.807e-07
I662 0 n663 3.361e-02A M=7.805e-07
I663 0 n664 3.361e-02A M=5.706e-07
I664 0 n665 3.361e-02A M=7.901e-07
I665 0 n666 3.361e-02A M=3.967e-07
I666 0 n667 3.361e-02A M=1.208e-06
I667 0 n668 3.361e-02A M=6.328e-07
I668 0 n669 3.361e-02A M=9.679e-07
I669 0 n670 3.361e-02A M=1.012e-06
I670 0 n671 3.361e-02A M=6.815e-07
I671 0 n672 3.361e-02A M=2.757e-06
I672 0 n673 3.361e-02A M=1.220e-06
I673 0 n674 3.361e-02A M=7.116e-07
I674 0 n675 3.361e-02A M=5.721e-07
I675 0 n676 3.361e-02A M=7.830e-07
I676 0 n677 3.361e-02A M=1.020e-06
I677 0 n678 3.361e-02A M=8.388e-07
I678 0 n679 3.361e-02A M=6.864e-07
I679 0 n680 3.361e-02A M=4.344e-07
I680 0 n681 3.361e-02A M=1.602e-06
I681 0 n682 3.361e-02A M=7.698e-07
I682 0 n683 3.361e-02A M=9.344e-07
I683 0 n684 3.361e-02A M=7.830e-07
I684 0 n685 3.361e-02A M=2.538e-07
I685 0 n686 3.361e-02A M=1.614e-06
I686 0 n687 3.361e-02A M=7.077e-07
I687 0 n688 3.361e-02A M=2.719e-06
I688 0 n689 3.361e-02A M=1.071e-06
I689 0 n690 3.361e-02A M=1.302e-06
I690 0 n691 3.361e-02A M=9.688e-07
I691 0 n692 3.361e-02A M=1.310e-06
I692 0 n1 3.361e-02A M=9.627e-07
I693 0 n694 3.361e-02A M=8.444e-07
I694 0 n695 3.361e-02A M=1.319e-06
I695 0 n696 3.361e-02A M=9.658e-07
I696 0 n697 3.361e-02A M=5.479e-07
I697 0 n698 3.361e-02A M=8.982e-07
I698 0 n699 3.361e-02A M=2.068e-06
I699 0 n700 3.361e-02A M=1.241e-07
I700 0 n701 3.361e-02A M=4.449e-07
I701 0 n702 3.361e-02A M=6.839e-07
I702 0 n703 3.361e-02A M=8.093e-07
I703 0 n704 3.361e-02A M=8.449e-07
I704 0 n705 3.361e-02A M=4.703e-07
I705 0 n706 3.361e-02A M=1.589e-06
I706 0 n707 3.361e-02A M=1.006e-06
I707 0 n708 3.361e-02A M=4.137e-07
I708 0 n709 3.361e-02A M=2.921e-06
I709 0 n710 3.361e-02A M=7.562e-07
I710 0 n711 3.361e-02A M=1.619e-06
I711 0 n712 3.361e-02A M=1.436e-06
I712 0 n713 3.361e-02A M=4.636e-07
I713 0 n714 3.361e-02A M=9.167e-07
I714 0 n715 3.361e-02A M=1.103e-06
I715 0 n716 3.361e-02A M=7.594e-07
I716 0 n717 3.361e-02A M=7.290e-07
I717 0 n718 3.361e-02A M=5.351e-07
I718 0 n719 3.361e-02A M=1.626e-06
I719 0 n720 3.361e-02A M=7.818e-07
I720 0 n721 3.361e-02A M=9.533e-07
I721 0 n722 3.361e-02A M=1.174e-06
I722 0 n723 3.361e-02A M=2.427e-07
I723 0 n724 3.361e-02A M=3.644e-07
I724 0 n725 3.361e-02A M=1.509e-06
I725 0 n726 3.361e-02A M=1.380e-06
I726 0 n727 3.361e-02A M=1.082e-06
I727 0 n728 3.361e-02A M=1.043e-06
I728 0 n729 3.361e-02A M=7.722e-07
I729 0 n730 3.361e-02A M=1.048e-06
I730 0 n731 3.361e-02A M=6.595e-07
I731 0 n732 3.361e-02A M=1.301e-06
I732 0 n733 3.361e-02A M=4.704e-07
I733 0 n734 3.361e-02A M=3.492e-07
I734 0 n735 3.361e-02A M=1.642e-06
I735 0 n736 3.361e-02A M=9.426e-07
I736 0 n737 3.361e-02A M=1.462e-06
I737 0 n738 3.361e-02A M=2.224e-06
I738 0 n739 3.361e-02A M=1.663e-06
I739 0 n740 3.361e-02A M=4.546e-07
I740 0 n741 3.361e-02A M=1.365e-06
I741 0 n742 3.361e-02A M=8.754e-07
I742 0 n743 3.361e-02A M=4.151e-07
I743 0 n744 3.361e-02A M=9.681e-07
I744 0 n745 3.361e-02A M=7.806e-07
I745 0 n746 3.361e-02A M=7.657e-07
I746 0 n747 3.361e-02A M=1.069e-06
I747 0 n748 3.361e-02A M=8.348e-07
I748 0 n749 3.361e-02A M=8.844e-07
I749 0 n750 3.361e-02A M=4.445e-07
I750 0 n751 3.361e-02A M=1.017e-06
I751 0 n752 3.361e-02A M=8.947e-07
I752 0 n753 3.361e-02A M=2.024e-06
I753 0 n754 3.361e-02A M=1.145e-06
I754 0 n755 3.361e-02A M=2.592e-06
I755 0 n756 3.361e-02A M=4.768e-07
I756 0 n757 3.361e-02A M=5.990e-07
I757 0 n758 3.361e-02A M=2.135e-06
I758 0 n759 3.361e-02A M=1.491e-06
I759 0 n760 3.361e-02A M=6.513e-07
I760 0 n761 3.361e-02A M=7.460e-07
I761 0 n762 3.361e-02A M=1.779e-06
I762 0 n763 3.361e-02A M=2.858e-07
I763 0 n764 3.361e-02A M=6.881e-07
I764 0 n765 3.361e-02A M=1.110e-06
I765 0 n766 3.361e-02A M=8.967e-07
I766 0 n767 3.361e-02A M=1.082e-06
I767 0 n768 3.361e-02A M=1.366e-06
I768 0 n769 3.361e-02A M=1.290e-06
I769 0 n770 3.361e-02A M=5.053e-07
I770 0 n771 3.361e-02A M=8.371e-07
I771 0 n772 3.361e-02A M=3.644e-06
I772 0 n773 3.361e-02A M=4.643e-07
I773 0 n774 3.361e-02A M=7.137e-07
I774 0 n775 3.361e-02A M=8.266e-07
I775 0 n776 3.361e-02A M=7.646e-07
I776 0 n777 3.361e-02A M=4.175e-07
I777 0 n778 3.361e-02A M=8.160e-07
I778 0 n779 3.361e-02A M=1.271e-06
I779 0 n780 3.361e-02A M=9.448e-07
I780 0 n781 3.361e-02A M=1.181e-06
I781 0 n782 3.361e-02A M=8.394e-07
I782 0 n783 3.361e-02A M=1.034e-06
I783 0 n784 3.361e-02A M=1.016e-06
I784 0 n785 3.361e-02A M=1.579e-06
I785 0 n786 3.361e-02A M=2.905e-07
I786 0 n787 3.361e-02A M=8.890e-07
I787 0 n788 3.361e-02A M=1.613e-06
I788 0 n789 3.361e-02A M=1.568e-06
I789 0 n790 3.361e-02A M=6.790e-07
I790 0 n791 3.361e-02A M=5.599e-07
I791 0 n792 3.361e-02A M=4.254e-07
I792 0 n793 3.361e-02A M=1.426e-06
I793 0 n794 3.361e-02A M=1.074e-06
I794 0 n795 3.361e-02A M=1.205e-06
I795 0 n796 3.361e-02A M=2.887e-07
I796 0 n797 3.361e-02A M=1.008e-06
I797 0 n798 3.361e-02A M=8.800e-07
I798 0 n799 3.361e-02A M=1.179e-06
I799 0 n800 3.361e-02A M=8.074e-07
I800 0 n801 3.361e-02A M=1.492e-06
I801 0 n802 3.361e-02A M=2.088e-07
I802 0 n803 3.361e-02A M=5.726e-07
I803 0 n804 3.361e-02A M=5.478e-07
I804 0 n805 3.361e-02A M=4.491e-07
I805 0 n806 3.361e-02A M=1.179e-06
I806 0 n807 3.361e-02A M=1.456e-06
I807 0 n808 3.361e-02A M=1.467e-06
I808 0 n809 3.361e-02A M=1.305e-06
I809 0 n810 3.361e-02A M=9.733e-07
I810 0 n811 3.361e-02A M=6.564e-07
I811 0 n812 3.361e-02A M=1.036e-06
I812 0 n813 3.361e-02A M=1.277e-06
I813 0 n814 3.361e-02A M=1.457e-06
I814 0 n815 3.361e-02A M=1.073e-06
I815 0 n816 3.361e-02A M=9.696e-07
I816 0 n817 3.361e-02A M=1.324e-06
I817 0 n818 3.361e-02A M=7.199e-07
I818 0 n819 3.361e-02A M=1.143e-06
I819 0 n820 3.361e-02A M=5.278e-07
I820 0 n821 3.361e-02A M=1.282e-06
I821 0 n822 3.361e-02A M=3.693e-07
I822 0 n823 3.361e-02A M=1.002e-06
I823 0 n824 3.361e-02A M=9.389e-07
I824 0 n825 3.361e-02A M=9.990e-07
I825 0 n826 3.361e-02A M=8.635e-07
I826 0 n827 3.361e-02A M=2.124e-06
I827 0 n828 3.361e-02A M=3.769e-07
I828 0 n829 3.361e-02A M=1.358e-06
I829 0 n830 3.361e-02A M=1.949e-06
I830 0 n831 3.361e-02A M=8.666e-07
I831 0 n832 3.361e-02A M=1.415e-06
I832 0 n833 3.361e-02A M=1.190e-06
I833 0 n834 3.361e-02A M=7.378e-07
I834 0 n835 3.361e-02A M=1.567e-06
I835 0 n836 3.361e-02A M=3.189e-06
I836 0 n837 3.361e-02A M=4.309e-07
I837 0 n838 3.361e-02A M=1.753e-06
I838 0 n839 3.361e-02A M=5.664e-07
I839 0 n840 3.361e-02A M=6.919e-07
I840 0 n841 3.361e-02A M=1.223e-06
I841 0 n842 3.361e-02A M=1.605e-06
I842 0 n843 3.361e-02A M=2.555e-07
I843 0 n844 3.361e-02A M=1.040e-06
I844 0 n845 3.361e-02A M=5.596e-07
I845 0 n846 3.361e-02A M=1.171e-06
I846 0 n847 3.361e-02A M=6.538e-07
I847 0 n848 3.361e-02A M=1.390e-06
I848 0 n849 3.361e-02A M=7.676e-07
I849 0 n850 3.361e-02A M=7.106e-07
I850 0 n851 3.361e-02A M=1.389e-06
I851 0 n852 3.361e-02A M=7.680e-07
I852 0 n853 3.361e-02A M=1.879e-06
I853 0 n854 3.361e-02A M=6.843e-07
I854 0 n855 3.361e-02A M=1.364e-06
I855 0 n856 3.361e-02A M=9.267e-07
I856 0 n857 3.361e-02A M=7.744e-07
I857 0 n858 3.361e-02A M=1.019e-06
I858 0 n859 3.361e-02A M=3.636e-07
I859 0 n860 3.361e-02A M=1.017e-06
I860 0 n861 3.361e-02A M=2.092e-06
I861 0 n862 3.361e-02A M=2.075e-06
I862 0 n863 3.361e-02A M=6.749e-07
I863 0 n864 3.361e-02A M=1.304e-06
I864 0 n865 3.361e-02A M=8.745e-07
I865 0 n866 3.361e-02A M=1.672e-06
I866 0 n867 3.361e-02A M=1.071e-06
I867 0 n868 3.361e-02A M=2.817e-07
I868 0 n869 3.361e-02A M=7.103e-07
I869 0 n870 3.361e-02A M=1.391e-06
I870 0 n871 3.361e-02A M=1.427e-06
I871 0 n872 3.361e-02A M=6.206e-07
I872 0 n873 3.361e-02A M=6.815e-07
I873 0 n874 3.361e-02A M=1.925e-06
I874 0 n875 3.361e-02A M=1.044e-06
I875 0 n876 3.361e-02A M=1.427e-06
I876 0 n877 3.361e-02A M=5.266e-07
I877 0 n878 3.361e-02A M=9.314e-07
I878 0 n879 3.361e-02A M=1.726e-06
I879 0 n880 3.361e-02A M=6.483e-07
I880 0 n881 3.361e-02A M=4.396e-07
I881 0 n882 3.361e-02A M=1.986e-06
I882 0 n883 3.361e-02A M=5.710e-07
I883 0 n884 3.361e-02A M=9.865e-07
I884 0 n885 3.361e-02A M=1.026e-06
I885 0 n886 3.361e-02A M=1.249e-06
I886 0 n887 3.361e-02A M=7.298e-07
I887 0 n888 3.361e-02A M=4.309e-07
I888 0 n889 3.361e-02A M=2.308e-06
I889 0 n890 3.361e-02A M=5.330e-07
I890 0 n891 3.361e-02A M=8.695e-07
I891 0 n892 3.361e-02A M=7.167e-07
I892 0 n893 3.361e-02A M=1.016e-06
I893 0 n894 3.361e-02A M=8.941e-07
I894 0 n895 3.361e-02A M=7.573e-07
I895 0 n896 3.361e-02A M=4.494e-07
I896 0 n897 3.361e-02A M=8.369e-07
I897 0 n1 3.361e-02A M=3.474e-07
I898 0 n899 3.361e-02A M=4.221e-07
I899 0 n900 3.361e-02A M=8.044e-07
I900 0 n901 3.361e-02A M=2.745e-06
I901 0 n902 3.361e-02A M=6.682e-07
I902 0 n903 3.361e-02A M=5.532e-07
I903 0 n904 3.361e-02A M=1.791e-06
I904 0 n905 3.361e-02A M=2.092e-06
I905 0 n906 3.361e-02A M=8.343e-07
I906 0 n907 3.361e-02A M=1.247e-06
I907 0 n908 3.361e-02A M=1.603e-06
I908 0 n909 3.361e-02A M=4.201e-07
I909 0 n910 3.361e-02A M=6.467e-07
I910 0 n911 3.361e-02A M=1.276e-06
I911 0 n912 3.361e-02A M=2.583e-07
I912 0 n913 3.361e-02A M=5.773e-07
I913 0 n914 3.361e-02A M=8.539e-07
I914 0 n915 3.361e-02A M=1.703e-06
I915 0 n916 3.361e-02A M=4.126e-07
I916 0 n917 3.361e-02A M=6.244e-07
I917 0 n918 3.361e-02A M=1.805e-06
I918 0 n919 3.361e-02A M=6.465e-07
I919 0 n920 3.361e-02A M=8.689e-07
I920 0 n921 3.361e-02A M=1.794e-06
I921 0 n922 3.361e-02A M=1.821e-06
I922 0 n923 3.361e-02A M=5.181e-07
I923 0 n924 3.361e-02A M=7.770e-07
I924 0 n925 3.361e-02A M=5.572e-07
I925 0 n926 3.361e-02A M=1.186e-06
I926 0 n927 3.361e-02A M=4.811e-07
I927 0 n928 3.361e-02A M=5.656e-07
I928 0 n929 3.361e-02A M=2.113e-07
I929 0 n930 3.361e-02A M=1.283e-06
I930 0 n931 3.361e-02A M=7.515e-07
I931 0 n932 3.361e-02A M=1.894e-06
I932 0 n933 3.361e-02A M=3.893e-07
I933 0 n934 3.361e-02A M=1.885e-06
I934 0 n935 3.361e-02A M=1.004e-06
I935 0 n936 3.361e-02A M=1.174e-07
I936 0 n937 3.361e-02A M=8.418e-07
I937 0 n938 3.361e-02A M=1.972e-06
I938 0 n939 3.361e-02A M=1.454e-06
I939 0 n940 3.361e-02A M=6.385e-07
I940 0 n941 3.361e-02A M=4.262e-07
I941 0 n942 3.361e-02A M=2.533e-07
I942 0 n943 3.361e-02A M=3.632e-07
I943 0 n944 3.361e-02A M=3.034e-06
I944 0 n945 3.361e-02A M=5.936e-07
I945 0 n946 3.361e-02A M=1.266e-06
I946 0 n947 3.361e-02A M=5.694e-07
I947 0 n948 3.361e-02A M=6.230e-07
I948 0 n949 3.361e-02A M=9.865e-07
I949 0 n950 3.361e-02A M=6.750e-07
I950 0 n951 3.361e-02A M=1.849e-06
I951 0 n952 3.361e-02A M=4.723e-07
I952 0 n953 3.361e-02A M=4.261e-07
I953 0 n954 3.361e-02A M=7.252e-07
I954 0 n955 3.361e-02A M=6.333e-07
I955 0 n956 3.361e-02A M=7.875e-07
I956 0 n957 3.361e-02A M=1.393e-06
I957 0 n958 3.361e-02A M=1.471e-06
I958 0 n959 3.361e-02A M=4.816e-07
I959 0 n960 3.361e-02A M=9.772e-07
I960 0 n961 3.361e-02A M=9.283e-07
I961 0 n962 3.361e-02A M=1.130e-06
I962 0 n963 3.361e-02A M=7.910e-07
I963 0 n964 3.361e-02A M=1.520e-06
I964 0 n965 3.361e-02A M=7.043e-07
I965 0 n966 3.361e-02A M=1.570e-06
I966 0 n967 3.361e-02A M=4.621e-07
I967 0 n968 3.361e-02A M=1.207e-06
I968 0 n969 3.361e-02A M=9.323e-07
I969 0 n970 3.361e-02A M=3.421e-06
I970 0 n971 3.361e-02A M=7.537e-07
I971 0 n972 3.361e-02A M=8.525e-07
I972 0 n973 3.361e-02A M=1.162e-06
I973 0 n974 3.361e-02A M=1.139e-06
I974 0 n975 3.361e-02A M=1.602e-06
I975 0 n976 3.361e-02A M=4.875e-07
I976 0 n977 3.361e-02A M=9.979e-07
I977 0 n978 3.361e-02A M=2.139e-06
I978 0 n979 3.361e-02A M=5.706e-07
I979 0 n980 3.361e-02A M=4.605e-07
I980 0 n981 3.361e-02A M=3.420e-07
I981 0 n982 3.361e-02A M=1.517e-06
I982 0 n983 3.361e-02A M=2.095e-06
I983 0 n984 3.361e-02A M=6.055e-07
I984 0 n985 3.361e-02A M=9.141e-07
I985 0 n986 3.361e-02A M=1.347e-06
I986 0 n987 3.361e-02A M=1.205e-07
I987 0 n988 3.361e-02A M=1.856e-06
I988 0 n989 3.361e-02A M=3.983e-07
I989 0 n990 3.361e-02A M=4.008e-07
I990 0 n991 3.361e-02A M=1.597e-06
I991 0 n992 3.361e-02A M=1.200e-06
I992 0 n993 3.361e-02A M=8.942e-07
I993 0 n994 3.361e-02A M=9.340e-07
I994 0 n995 3.361e-02A M=7.421e-07
I995 0 n996 3.361e-02A M=8.892e-07
I996 0 n997 3.361e-02A M=7.726e-07
I997 0 n998 3.361e-02A M=1.198e-06
I998 0 n999 3.361e-02A M=1.302e-06
I999 0 n1000 3.361e-02A M=1.729e-06
I1000 0 n1001 3.361e-02A M=1.284e-06
I1001 0 n1002 3.361e-02A M=5.222e-07
I1002 0 n1003 3.361e-02A M=4.123e-07
I1003 0 n1004 3.361e-02A M=8.629e-07
I1004 0 n1005 3.361e-02A M=7.233e-07
I1005 0 n1006 3.361e-02A M=1.454e-06
I1006 0 n1007 3.361e-02A M=4.087e-07
I1007 0 n1008 3.361e-02A M=5.867e-07
I1008 0 n1009 3.361e-02A M=1.072e-06
I1009 0 n1010 3.361e-02A M=1.232e-06
I1010 0 n1011 3.361e-02A M=7.836e-07
I1011 0 n1012 3.361e-02A M=2.219e-07
I1012 0 n1013 3.361e-02A M=1.337e-06
I1013 0 n1014 3.361e-02A M=6.436e-07
I1014 0 n1015 3.361e-02A M=1.038e-06
I1015 0 n1016 3.361e-02A M=5.271e-07
I1016 0 n1017 3.361e-02A M=8.883e-07
I1017 0 n1018 3.361e-02A M=6.726e-07
I1018 0 n1019 3.361e-02A M=4.937e-07
I1019 0 n1020 3.361e-02A M=9.001e-07
I1020 0 n1021 3.361e-02A M=2.020e-06
I1021 0 n1022 3.361e-02A M=5.327e-07
I1022 0 n1023 3.361e-02A M=4.563e-07
I1023 0 n1024 3.361e-02A M=1.484e-06
I1024 0 n1025 3.361e-02A M=8.412e-07
I1025 0 n1026 3.361e-02A M=1.425e-06
I1026 0 n1027 3.361e-02A M=9.694e-07
I1027 0 n1028 3.361e-02A M=4.368e-07
I1028 0 n1029 3.361e-02A M=4.314e-07
I1029 0 n1030 3.361e-02A M=5.495e-07
I1030 0 n1031 3.361e-02A M=1.402e-06
I1031 0 n1032 3.361e-02A M=3.140e-07
I1032 0 n1033 3.361e-02A M=6.079e-07
I1033 0 n1034 3.361e-02A M=3.358e-07
I1034 0 n1035 3.361e-02A M=9.251e-07
I1035 0 n1036 3.361e-02A M=9.467e-07
I1036 0 n1037 3.361e-02A M=9.816e-07
I1037 0 n1038 3.361e-02A M=2.402e-07
I1038 0 n1039 3.361e-02A M=9.594e-07
I1039 0 n1040 3.361e-02A M=8.810e-07
I1040 0 n1041 3.361e-02A M=1.001e-06
I1041 0 n1042 3.361e-02A M=1.579e-06
I1042 0 n1043 3.361e-02A M=4.856e-07
I1043 0 n1044 3.361e-02A M=1.007e-06
I1044 0 n1045 3.361e-02A M=7.230e-07
I1045 0 n1046 3.361e-02A M=6.866e-07
I1046 0 n1047 3.361e-02A M=1.012e-06
I1047 0 n1048 3.361e-02A M=1.467e-06
I1048 0 n1049 3.361e-02A M=5.830e-07
I1049 0 n1050 3.361e-02A M=7.527e-07
I1050 0 n1051 3.361e-02A M=6.642e-07
I1051 0 n1052 3.361e-02A M=5.666e-07
I1052 0 n1053 3.361e-02A M=9.839e-07
I1053 0 n1054 3.361e-02A M=1.556e-06
I1054 0 n1055 3.361e-02A M=5.277e-07
I1055 0 n1056 3.361e-02A M=1.248e-06
I1056 0 n1057 3.361e-02A M=1.159e-06
I1057 0 n1058 3.361e-02A M=2.892e-07
I1058 0 n1059 3.361e-02A M=3.389e-07
I1059 0 n1060 3.361e-02A M=4.291e-07
I1060 0 n1061 3.361e-02A M=5.826e-07
I1061 0 n1062 3.361e-02A M=1.196e-06
I1062 0 n1063 3.361e-02A M=3.238e-07
I1063 0 n1064 3.361e-02A M=1.000e-06
I1064 0 n1065 3.361e-02A M=1.679e-07
I1065 0 n1066 3.361e-02A M=1.662e-06
I1066 0 n1067 3.361e-02A M=1.260e-06
I1067 0 n1068 3.361e-02A M=2.223e-06
I1068 0 n1069 3.361e-02A M=4.112e-07
I1069 0 n1070 3.361e-02A M=2.479e-07
I1070 0 n1071 3.361e-02A M=1.118e-06
I1071 0 n1072 3.361e-02A M=6.374e-07
I1072 0 n1073 3.361e-02A M=8.490e-07
I1073 0 n1074 3.361e-02A M=1.363e-06
I1074 0 n1075 3.361e-02A M=8.383e-07
I1075 0 n1076 3.361e-02A M=1.312e-06
I1076 0 n1077 3.361e-02A M=8.454e-07
I1077 0 n1078 3.361e-02A M=9.880e-07
I1078 0 n1079 3.361e-02A M=6.704e-07
I1079 0 n1080 3.361e-02A M=1.256e-06
I1080 0 n1081 3.361e-02A M=5.184e-07
I1081 0 n1082 3.361e-02A M=7.780e-07
I1082 0 n1083 3.361e-02A M=1.457e-06
I1083 0 n1084 3.361e-02A M=9.524e-07
I1084 0 n1085 3.361e-02A M=1.620e-06
I1085 0 n1086 3.361e-02A M=4.643e-07
I1086 0 n1087 3.361e-02A M=3.534e-07
I1087 0 n1088 3.361e-02A M=2.927e-06
I1088 0 n1089 3.361e-02A M=9.416e-07
I1089 0 n1090 3.361e-02A M=7.030e-07
I1090 0 n1091 3.361e-02A M=1.343e-06
I1091 0 n1092 3.361e-02A M=5.547e-07
I1092 0 n1093 3.361e-02A M=1.104e-06
I1093 0 n1094 3.361e-02A M=4.889e-07
I1094 0 n1095 3.361e-02A M=1.405e-06
I1095 0 n1096 3.361e-02A M=1.881e-06
I1096 0 n1097 3.361e-02A M=1.346e-06
I1097 0 n1098 3.361e-02A M=4.977e-07
I1098 0 n1099 3.361e-02A M=1.340e-06
I1099 0 n1100 3.361e-02A M=9.670e-07
I1100 0 n1101 3.361e-02A M=5.549e-07
I1101 0 n1102 3.361e-02A M=1.047e-06
I1102 0 n1103 3.361e-02A M=3.417e-07
I1103 0 n1104 3.361e-02A M=2.496e-07
I1104 0 n1105 3.361e-02A M=9.603e-07
I1105 0 n1106 3.361e-02A M=8.420e-07
I1106 0 n1107 3.361e-02A M=7.632e-07
I1107 0 n1108 3.361e-02A M=6.593e-07
I1108 0 n1109 3.361e-02A M=1.149e-06
I1109 0 n1110 3.361e-02A M=9.321e-07
I1110 0 n1111 3.361e-02A M=9.308e-07
I1111 0 n1112 3.361e-02A M=5.469e-07
I1112 0 n1113 3.361e-02A M=4.603e-07
I1113 0 n1114 3.361e-02A M=1.602e-06
I1114 0 n1115 3.361e-02A M=7.956e-07
I1115 0 n1116 3.361e-02A M=1.039e-06
I1116 0 n1117 3.361e-02A M=6.046e-07
I1117 0 n1118 3.361e-02A M=6.844e-07
I1118 0 n1119 3.361e-02A M=1.054e-06
I1119 0 n1120 3.361e-02A M=1.216e-06
I1120 0 n1121 3.361e-02A M=1.002e-06
I1121 0 n1122 3.361e-02A M=1.671e-06
I1122 0 n1123 3.361e-02A M=1.216e-06
I1123 0 n1124 3.361e-02A M=1.888e-06
I1124 0 n1125 3.361e-02A M=5.609e-07
I1125 0 n1126 3.361e-02A M=6.535e-07
I1126 0 n1127 3.361e-02A M=8.262e-07
I1127 0 n1128 3.361e-02A M=7.725e-07
I1128 0 n1129 3.361e-02A M=1.012e-06
I1129 0 n1130 3.361e-02A M=1.503e-07
I1130 0 n1131 3.361e-02A M=1.233e-06
I1131 0 n1132 3.361e-02A M=6.558e-07
I1132 0 n1133 3.361e-02A M=4.904e-07
I1133 0 n1134 3.361e-02A M=1.348e-07
I1134 0 n1135 3.361e-02A M=5.693e-07
I1135 0 n1136 3.361e-02A M=1.921e-06
I1136 0 n1137 3.361e-02A M=6.643e-07
I1137 0 n1138 3.361e-02A M=1.544e-06
I1138 0 n1139 3.361e-02A M=2.000e-06
I1139 0 n1140 3.361e-02A M=9.005e-07
I1140 0 n1141 3.361e-02A M=1.078e-06
I1141 0 n1142 3.361e-02A M=5.338e-07
I1142 0 n1143 3.361e-02A M=1.645e-06
I1143 0 n1144 3.361e-02A M=5.375e-07
I1144 0 n1145 3.361e-02A M=1.101e-06
I1145 0 n1146 3.361e-02A M=5.534e-07
I1146 0 n1147 3.361e-02A M=9.812e-07
I1147 0 n1148 3.361e-02A M=5.272e-07
I1148 0 n1149 3.361e-02A M=1.079e-06
I1149 0 n1150 3.361e-02A M=1.069e-06
I1150 0 n1151 3.361e-02A M=1.024e-06
I1151 0 n1152 3.361e-02A M=1.674e-06
I1152 0 n1153 3.361e-02A M=6.382e-07
I1153 0 n1154 3.361e-02A M=1.262e-06
I1154 0 n1 3.361e-02A M=1.467e-07
I1155 0 n1156 3.361e-02A M=3.325e-07
I1156 0 n1157 3.361e-02A M=2.280e-06
I1157 0 n1158 3.361e-02A M=3.235e-07
I1158 0 n1159 3.361e-02A M=6.261e-07
I1159 0 n1160 3.361e-02A M=4.874e-07
I1160 0 n1161 3.361e-02A M=1.195e-06
I1161 0 n1162 3.361e-02A M=2.748e-07
I1162 0 n1163 3.361e-02A M=1.147e-06
I1163 0 n1164 3.361e-02A M=9.839e-07
I1164 0 n1165 3.361e-02A M=8.702e-07
I1165 0 n1166 3.361e-02A M=1.089e-06
I1166 0 n1167 3.361e-02A M=1.753e-06
I1167 0 n1168 3.361e-02A M=1.059e-06
I1168 0 n1169 3.361e-02A M=5.824e-07
I1169 0 n1170 3.361e-02A M=5.200e-07
I1170 0 n1171 3.361e-02A M=4.780e-07
I1171 0 n1172 3.361e-02A M=6.333e-07
I1172 0 n1173 3.361e-02A M=6.107e-07
I1173 0 n1174 3.361e-02A M=1.589e-06
I1174 0 n1175 3.361e-02A M=3.762e-07
I1175 0 n1176 3.361e-02A M=6.843e-07
I1176 0 n1177 3.361e-02A M=1.946e-06
I1177 0 n1178 3.361e-02A M=1.198e-06
I1178 0 n1179 3.361e-02A M=1.049e-06
I1179 0 n1 3.361e-02A M=1.754e-07
I1180 0 n1181 3.361e-02A M=1.066e-06
I1181 0 n1182 3.361e-02A M=2.980e-06
I1182 0 n1183 3.361e-02A M=6.420e-07
I1183 0 n1184 3.361e-02A M=1.789e-06
I1184 0 n1185 3.361e-02A M=6.495e-07
I1185 0 n1186 3.361e-02A M=1.157e-06
I1186 0 n1187 3.361e-02A M=3.745e-06
I1187 0 n1188 3.361e-02A M=1.505e-06
I1188 0 n1189 3.361e-02A M=7.910e-07
I1189 0 n1190 3.361e-02A M=3.087e-07
I1190 0 n1191 3.361e-02A M=9.167e-07
I1191 0 n1192 3.361e-02A M=1.443e-06
I1192 0 n1193 3.361e-02A M=9.274e-07
I1193 0 n1194 3.361e-02A M=8.541e-07
I1194 0 n1195 3.361e-02A M=1.803e-06
I1195 0 n1196 3.361e-02A M=9.266e-07
I1196 0 n1197 3.361e-02A M=9.330e-07
I1197 0 n1198 3.361e-02A M=7.810e-07
I1198 0 n1199 3.361e-02A M=1.517e-06
I1199 0 n1200 3.361e-02A M=6.532e-07
I1200 0 n1201 3.361e-02A M=9.095e-07
I1201 0 n1 3.361e-02A M=7.429e-07
I1202 0 n1203 3.361e-02A M=1.222e-06
I1203 0 n1204 3.361e-02A M=3.085e-07
I1204 0 n1205 3.361e-02A M=6.816e-07
I1205 0 n1206 3.361e-02A M=1.046e-06
I1206 0 n1207 3.361e-02A M=1.549e-06
I1207 0 n1208 3.361e-02A M=4.001e-07
I1208 0 n1209 3.361e-02A M=3.081e-07
I1209 0 n1210 3.361e-02A M=1.452e-06
I1210 0 n1211 3.361e-02A M=4.018e-07
I1211 0 n1212 3.361e-02A M=8.383e-07
I1212 0 n1213 3.361e-02A M=1.097e-06
I1213 0 n1214 3.361e-02A M=5.261e-07
I1214 0 n1215 3.361e-02A M=1.340e-06
I1215 0 n1216 3.361e-02A M=8.519e-07
I1216 0 n1217 3.361e-02A M=5.907e-07
I1217 0 n1218 3.361e-02A M=4.965e-07
I1218 0 n1219 3.361e-02A M=1.076e-06
I1219 0 n1220 3.361e-02A M=9.905e-07
I1220 0 n1221 3.361e-02A M=1.373e-06
I1221 0 n1222 3.361e-02A M=9.037e-07
I1222 0 n1223 3.361e-02A M=1.445e-06
I1223 0 n1224 3.361e-02A M=1.089e-06
I1224 0 n1225 3.361e-02A M=2.026e-06
I1225 0 n1226 3.361e-02A M=6.371e-07
I1226 0 n1227 3.361e-02A M=1.102e-06
I1227 0 n1228 3.361e-02A M=1.423e-06
I1228 0 n1229 3.361e-02A M=6.930e-07
I1229 0 n1230 3.361e-02A M=5.410e-07
I1230 0 n1231 3.361e-02A M=1.181e-06
I1231 0 n1232 3.361e-02A M=7.902e-07
I1232 0 n1233 3.361e-02A M=1.906e-06
I1233 0 n1234 3.361e-02A M=1.627e-06
I1234 0 n1235 3.361e-02A M=9.834e-07
I1235 0 n1236 3.361e-02A M=7.134e-07
I1236 0 n1237 3.361e-02A M=5.238e-07
I1237 0 n1238 3.361e-02A M=1.039e-06
I1238 0 n1239 3.361e-02A M=4.796e-07
I1239 0 n1240 3.361e-02A M=1.231e-06
I1240 0 n1241 3.361e-02A M=2.033e-06
I1241 0 n1242 3.361e-02A M=1.468e-06
I1242 0 n1243 3.361e-02A M=1.187e-06
I1243 0 n1244 3.361e-02A M=8.674e-07
I1244 0 n1245 3.361e-02A M=1.402e-06
I1245 0 n1246 3.361e-02A M=4.845e-07
I1246 0 n1247 3.361e-02A M=2.072e-06
I1247 0 n1248 3.361e-02A M=1.837e-06
I1248 0 n1249 3.361e-02A M=1.429e-06
I1249 0 n1250 3.361e-02A M=1.072e-06
I1250 0 n1251 3.361e-02A M=2.997e-06
I1251 0 n1252 3.361e-02A M=9.704e-07
I1252 0 n1253 3.361e-02A M=2.445e-06
I1253 0 n1254 3.361e-02A M=5.237e-07
I1254 0 n1255 3.361e-02A M=5.501e-07
I1255 0 n1256 3.361e-02A M=7.598e-07
I1256 0 n1257 3.361e-02A M=3.154e-07
I1257 0 n1258 3.361e-02A M=1.677e-06
I1258 0 n1259 3.361e-02A M=5.373e-07
I1259 0 n1260 3.361e-02A M=2.585e-06
I1260 0 n1261 3.361e-02A M=9.400e-07
I1261 0 n1262 3.361e-02A M=1.394e-06
I1262 0 n1263 3.361e-02A M=6.791e-07
I1263 0 n1264 3.361e-02A M=1.149e-06
I1264 0 n1265 3.361e-02A M=1.494e-06
I1265 0 n1266 3.361e-02A M=1.845e-06
I1266 0 n1267 3.361e-02A M=4.265e-07
I1267 0 n1268 3.361e-02A M=5.703e-07
I1268 0 n1269 3.361e-02A M=6.306e-07
I1269 0 n1270 3.361e-02A M=1.273e-06
I1270 0 n1271 3.361e-02A M=9.577e-07
I1271 0 n1 3.361e-02A M=1.202e-06
I1272 0 n1273 3.361e-02A M=7.172e-07
I1273 0 n1 3.361e-02A M=1.467e-06
I1274 0 n1275 3.361e-02A M=6.894e-07
I1275 0 n1276 3.361e-02A M=5.128e-07
I1276 0 n1277 3.361e-02A M=6.178e-07
I1277 0 n1278 3.361e-02A M=1.030e-06
I1278 0 n1279 3.361e-02A M=1.459e-06
I1279 0 n1280 3.361e-02A M=1.112e-06
I1280 0 n1281 3.361e-02A M=5.704e-07
I1281 0 n1282 3.361e-02A M=9.410e-07
I1282 0 n1283 3.361e-02A M=5.494e-07
I1283 0 n1284 3.361e-02A M=3.777e-07
I1284 0 n1285 3.361e-02A M=8.725e-07
I1285 0 n1286 3.361e-02A M=8.546e-07
I1286 0 n1287 3.361e-02A M=9.583e-07
I1287 0 n1288 3.361e-02A M=8.806e-07
I1288 0 n1289 3.361e-02A M=1.037e-06
I1289 0 n1290 3.361e-02A M=1.736e-06
I1290 0 n1291 3.361e-02A M=8.460e-07
I1291 0 n1292 3.361e-02A M=1.094e-06
I1292 0 n1293 3.361e-02A M=2.990e-07
I1293 0 n1294 3.361e-02A M=3.277e-06
I1294 0 n1295 3.361e-02A M=8.789e-07
I1295 0 n1296 3.361e-02A M=7.119e-07
I1296 0 n1297 3.361e-02A M=2.204e-07
I1297 0 n1298 3.361e-02A M=5.487e-07
I1298 0 n1299 3.361e-02A M=2.187e-06
I1299 0 n1300 3.361e-02A M=8.579e-07
I1300 0 n1301 3.361e-02A M=4.424e-07
I1301 0 n1302 3.361e-02A M=1.099e-06
I1302 0 n1303 3.361e-02A M=1.027e-06
I1303 0 n1304 3.361e-02A M=9.992e-07
I1304 0 n1305 3.361e-02A M=3.724e-07
I1305 0 n1306 3.361e-02A M=6.971e-07
I1306 0 n1307 3.361e-02A M=6.495e-07
I1307 0 n1308 3.361e-02A M=1.654e-06
I1308 0 n1309 3.361e-02A M=7.685e-07
I1309 0 n1310 3.361e-02A M=2.753e-07
I1310 0 n1311 3.361e-02A M=6.639e-07
I1311 0 n1312 3.361e-02A M=1.112e-06
I1312 0 n1313 3.361e-02A M=9.638e-07
I1313 0 n1314 3.361e-02A M=1.336e-06
I1314 0 n1315 3.361e-02A M=9.499e-07
I1315 0 n1316 3.361e-02A M=7.674e-07
I1316 0 n1317 3.361e-02A M=1.118e-06
I1317 0 n1318 3.361e-02A M=6.136e-07
I1318 0 n1319 3.361e-02A M=8.260e-07
I1319 0 n1320 3.361e-02A M=5.301e-07
I1320 0 n1321 3.361e-02A M=1.634e-06
I1321 0 n1322 3.361e-02A M=1.078e-06
I1322 0 n1 3.361e-02A M=8.366e-07
I1323 0 n1324 3.361e-02A M=9.161e-07
I1324 0 n1325 3.361e-02A M=5.830e-07
I1325 0 n1326 3.361e-02A M=7.678e-07
I1326 0 n1327 3.361e-02A M=1.152e-06
I1327 0 n1328 3.361e-02A M=5.169e-07
I1328 0 n1329 3.361e-02A M=1.268e-06
I1329 0 n1330 3.361e-02A M=1.589e-06
I1330 0 n1331 3.361e-02A M=5.159e-07
I1331 0 n1332 3.361e-02A M=1.541e-06
I1332 0 n1333 3.361e-02A M=5.760e-07
I1333 0 n1334 3.361e-02A M=1.636e-06
I1334 0 n1335 3.361e-02A M=6.405e-07
I1335 0 n1336 3.361e-02A M=1.263e-06
I1336 0 n1337 3.361e-02A M=3.747e-07
I1337 0 n1338 3.361e-02A M=1.078e-06
I1338 0 n1339 3.361e-02A M=4.879e-07
I1339 0 n1340 3.361e-02A M=5.668e-07
I1340 0 n1341 3.361e-02A M=6.375e-07
I1341 0 n1342 3.361e-02A M=1.525e-06
I1342 0 n1343 3.361e-02A M=5.264e-07
I1343 0 n1344 3.361e-02A M=1.118e-06
I1344 0 n1345 3.361e-02A M=1.133e-06
I1345 0 n1346 3.361e-02A M=1.223e-06
I1346 0 n1347 3.361e-02A M=9.810e-07
I1347 0 n1348 3.361e-02A M=2.095e-07
I1348 0 n1349 3.361e-02A M=1.405e-06
I1349 0 n1350 3.361e-02A M=1.018e-06
I1350 0 n1351 3.361e-02A M=8.551e-07
I1351 0 n1352 3.361e-02A M=7.011e-07
I1352 0 n1353 3.361e-02A M=1.951e-07
I1353 0 n1354 3.361e-02A M=2.472e-06
I1354 0 n1355 3.361e-02A M=1.340e-06
I1355 0 n1356 3.361e-02A M=5.189e-07
I1356 0 n1357 3.361e-02A M=1.393e-06
I1357 0 n1358 3.361e-02A M=4.310e-07
I1358 0 n1359 3.361e-02A M=6.278e-07
I1359 0 n1360 3.361e-02A M=1.474e-06
I1360 0 n1361 3.361e-02A M=1.389e-06
I1361 0 n1362 3.361e-02A M=1.314e-06
I1362 0 n1363 3.361e-02A M=2.150e-07
I1363 0 n1364 3.361e-02A M=9.767e-07
I1364 0 n1365 3.361e-02A M=1.025e-06
I1365 0 n1366 3.361e-02A M=1.153e-06
I1366 0 n1367 3.361e-02A M=9.387e-07
I1367 0 n1368 3.361e-02A M=1.071e-06
I1368 0 n1369 3.361e-02A M=6.779e-07
I1369 0 n1370 3.361e-02A M=4.364e-07
I1370 0 n1371 3.361e-02A M=2.038e-06
I1371 0 n1372 3.361e-02A M=5.232e-07
I1372 0 n1373 3.361e-02A M=9.390e-07
I1373 0 n1374 3.361e-02A M=1.048e-06
I1374 0 n1375 3.361e-02A M=1.848e-06
I1375 0 n1376 3.361e-02A M=9.124e-07
I1376 0 n1377 3.361e-02A M=3.800e-07
I1377 0 n1378 3.361e-02A M=5.474e-07
I1378 0 n1379 3.361e-02A M=6.509e-07
I1379 0 n1380 3.361e-02A M=6.121e-07
I1380 0 n1381 3.361e-02A M=1.382e-06
I1381 0 n1382 3.361e-02A M=1.841e-06
I1382 0 n1383 3.361e-02A M=1.845e-06
I1383 0 n1384 3.361e-02A M=1.273e-06
I1384 0 n1385 3.361e-02A M=1.008e-06
I1385 0 n1386 3.361e-02A M=8.960e-07
I1386 0 n1387 3.361e-02A M=6.383e-07
I1387 0 n1388 3.361e-02A M=8.634e-07
I1388 0 n1389 3.361e-02A M=6.428e-07
I1389 0 n1390 3.361e-02A M=1.337e-06
I1390 0 n1391 3.361e-02A M=1.438e-06
I1391 0 n1392 3.361e-02A M=1.274e-06
I1392 0 n1393 3.361e-02A M=1.400e-06
I1393 0 n1394 3.361e-02A M=2.447e-06
I1394 0 n1395 3.361e-02A M=3.376e-07
I1395 0 n1396 3.361e-02A M=1.658e-06
I1396 0 n1397 3.361e-02A M=4.320e-07
I1397 0 n1398 3.361e-02A M=2.145e-07
I1398 0 n1399 3.361e-02A M=3.584e-07
I1399 0 n1400 3.361e-02A M=3.593e-07
I1400 0 n1401 3.361e-02A M=1.448e-06
I1401 0 n1402 3.361e-02A M=1.679e-07
I1402 0 n1403 3.361e-02A M=9.943e-07
I1403 0 n1404 3.361e-02A M=6.620e-07
I1404 0 n1405 3.361e-02A M=1.620e-06
I1405 0 n1406 3.361e-02A M=8.143e-07
I1406 0 n1407 3.361e-02A M=1.284e-06
I1407 0 n1408 3.361e-02A M=8.231e-07
I1408 0 n1409 3.361e-02A M=1.554e-06
I1409 0 n1410 3.361e-02A M=2.068e-06
I1410 0 n1411 3.361e-02A M=6.382e-07
I1411 0 n1412 3.361e-02A M=4.692e-07
I1412 0 n1413 3.361e-02A M=1.344e-06
I1413 0 n1414 3.361e-02A M=8.122e-07
I1414 0 n1415 3.361e-02A M=7.427e-07
I1415 0 n1416 3.361e-02A M=1.848e-06
I1416 0 n1417 3.361e-02A M=1.176e-06
I1417 0 n1418 3.361e-02A M=1.085e-06
I1418 0 n1419 3.361e-02A M=5.629e-07
I1419 0 n1420 3.361e-02A M=2.393e-07
I1420 0 n1421 3.361e-02A M=1.366e-06
I1421 0 n1422 3.361e-02A M=1.650e-06
I1422 0 n1423 3.361e-02A M=5.174e-07
I1423 0 n1424 3.361e-02A M=1.771e-06
I1424 0 n1425 3.361e-02A M=5.781e-07
I1425 0 n1426 3.361e-02A M=2.063e-07
I1426 0 n1427 3.361e-02A M=4.956e-07
I1427 0 n1428 3.361e-02A M=1.519e-06
I1428 0 n1429 3.361e-02A M=4.957e-07
I1429 0 n1430 3.361e-02A M=4.583e-07
I1430 0 n1431 3.361e-02A M=1.300e-06
I1431 0 n1432 3.361e-02A M=4.333e-07
I1432 0 n1433 3.361e-02A M=5.188e-07
I1433 0 n1434 3.361e-02A M=2.466e-06
I1434 0 n1435 3.361e-02A M=8.620e-07
I1435 0 n1436 3.361e-02A M=9.649e-07
I1436 0 n1437 3.361e-02A M=5.923e-07
I1437 0 n1438 3.361e-02A M=1.521e-06
I1438 0 n1439 3.361e-02A M=5.792e-07
I1439 0 n1440 3.361e-02A M=1.517e-06
I1440 0 n1441 3.361e-02A M=9.445e-07
I1441 0 n1442 3.361e-02A M=4.794e-07
I1442 0 n1443 3.361e-02A M=1.693e-06
I1443 0 n1444 3.361e-02A M=2.112e-06
I1444 0 n1445 3.361e-02A M=2.636e-06
I1445 0 n1446 3.361e-02A M=6.804e-07
I1446 0 n1447 3.361e-02A M=7.208e-07
I1447 0 n1448 3.361e-02A M=7.877e-07
I1448 0 n1449 3.361e-02A M=8.382e-07
I1449 0 n1450 3.361e-02A M=1.134e-06
I1450 0 n1451 3.361e-02A M=1.611e-06
I1451 0 n1452 3.361e-02A M=1.241e-06
I1452 0 n1453 3.361e-02A M=4.432e-07
I1453 0 n1454 3.361e-02A M=1.787e-07
I1454 0 n1455 3.361e-02A M=1.588e-06
I1455 0 n1456 3.361e-02A M=7.620e-07
I1456 0 n1457 3.361e-02A M=9.841e-07
I1457 0 n1458 3.361e-02A M=1.817e-06
I1458 0 n1459 3.361e-02A M=1.642e-06
I1459 0 n1460 3.361e-02A M=9.306e-07
I1460 0 n1461 3.361e-02A M=3.214e-07
I1461 0 n1462 3.361e-02A M=1.567e-06
I1462 0 n1463 3.361e-02A M=5.108e-07
I1463 0 n1464 3.361e-02A M=6.833e-07
I1464 0 n1465 3.361e-02A M=5.559e-07
I1465 0 n1466 3.361e-02A M=1.508e-06
I1466 0 n1467 3.361e-02A M=2.585e-06
I1467 0 n1468 3.361e-02A M=1.476e-06
I1468 0 n1469 3.361e-02A M=2.525e-07
I1469 0 n1470 3.361e-02A M=7.834e-07
I1470 0 n1471 3.361e-02A M=1.247e-06
I1471 0 n1472 3.361e-02A M=8.702e-07
I1472 0 n1473 3.361e-02A M=6.867e-07
I1473 0 n1474 3.361e-02A M=4.001e-07
I1474 0 n1475 3.361e-02A M=2.025e-06
I1475 0 n1476 3.361e-02A M=1.834e-06
I1476 0 n1477 3.361e-02A M=1.915e-06
I1477 0 n1478 3.361e-02A M=2.319e-06
I1478 0 n1479 3.361e-02A M=6.918e-07
I1479 0 n1480 3.361e-02A M=5.841e-07
I1480 0 n1481 3.361e-02A M=7.324e-07
I1481 0 n1482 3.361e-02A M=4.942e-07
I1482 0 n1483 3.361e-02A M=4.433e-07
I1483 0 n1484 3.361e-02A M=8.009e-07
I1484 0 n1 3.361e-02A M=2.441e-06
I1485 0 n1486 3.361e-02A M=1.522e-06
I1486 0 n1487 3.361e-02A M=1.151e-06
I1487 0 n1488 3.361e-02A M=1.370e-06
I1488 0 n1489 3.361e-02A M=6.660e-07
I1489 0 n1490 3.361e-02A M=7.215e-07
I1490 0 n1491 3.361e-02A M=9.714e-07
I1491 0 n1492 3.361e-02A M=7.258e-08
I1492 0 n1493 3.361e-02A M=1.252e-06
I1493 0 n1494 3.361e-02A M=6.670e-07
I1494 0 n1495 3.361e-02A M=1.106e-06
I1495 0 n1496 3.361e-02A M=3.938e-07
I1496 0 n1497 3.361e-02A M=8.470e-07
I1497 0 n1498 3.361e-02A M=6.571e-07
I1498 0 n1499 3.361e-02A M=1.482e-07
I1499 0 n1500 3.361e-02A M=3.626e-07
I1500 0 n1501 3.361e-02A M=1.443e-06
I1501 0 n1502 3.361e-02A M=2.580e-07
I1502 0 n1503 3.361e-02A M=1.633e-06
I1503 0 n1504 3.361e-02A M=4.322e-07
I1504 0 n1505 3.361e-02A M=3.472e-07
I1505 0 n1506 3.361e-02A M=1.051e-06
I1506 0 n1507 3.361e-02A M=8.320e-07
I1507 0 n1508 3.361e-02A M=1.092e-06
I1508 0 n1509 3.361e-02A M=1.177e-06
I1509 0 n1510 3.361e-02A M=1.280e-06
I1510 0 n1511 3.361e-02A M=2.356e-06
I1511 0 n1512 3.361e-02A M=7.682e-07
I1512 0 n1513 3.361e-02A M=1.136e-06
I1513 0 n1514 3.361e-02A M=7.346e-07
I1514 0 n1515 3.361e-02A M=1.323e-06
I1515 0 n1516 3.361e-02A M=8.245e-07
I1516 0 n1517 3.361e-02A M=1.191e-06
I1517 0 n1518 3.361e-02A M=1.186e-06
I1518 0 n1519 3.361e-02A M=1.377e-06
I1519 0 n1520 3.361e-02A M=1.207e-06
I1520 0 n1521 3.361e-02A M=9.599e-07
I1521 0 n1522 3.361e-02A M=8.889e-07
I1522 0 n1523 3.361e-02A M=4.371e-07
I1523 0 n1524 3.361e-02A M=5.879e-07
I1524 0 n1525 3.361e-02A M=2.363e-07
I1525 0 n1526 3.361e-02A M=7.867e-07
I1526 0 n1527 3.361e-02A M=1.772e-06
I1527 0 n1528 3.361e-02A M=3.266e-07
I1528 0 n1529 3.361e-02A M=3.685e-07
I1529 0 n1530 3.361e-02A M=1.592e-06
I1530 0 n1531 3.361e-02A M=5.660e-07
I1531 0 n1532 3.361e-02A M=9.475e-07
I1532 0 n1533 3.361e-02A M=5.495e-07
I1533 0 n1534 3.361e-02A M=1.688e-06
I1534 0 n1535 3.361e-02A M=5.259e-07
I1535 0 n1536 3.361e-02A M=2.000e-06
I1536 0 n1537 3.361e-02A M=6.422e-07
I1537 0 n1538 3.361e-02A M=3.411e-07
I1538 0 n1539 3.361e-02A M=1.046e-06
I1539 0 n1540 3.361e-02A M=8.563e-07
I1540 0 n1541 3.361e-02A M=1.542e-06
I1541 0 n1542 3.361e-02A M=1.511e-06
I1542 0 n1543 3.361e-02A M=1.311e-06
I1543 0 n1544 3.361e-02A M=1.150e-06
I1544 0 n1545 3.361e-02A M=2.770e-07
I1545 0 n1546 3.361e-02A M=2.137e-06
I1546 0 n1547 3.361e-02A M=4.020e-07
I1547 0 n1548 3.361e-02A M=4.176e-07
I1548 0 n1549 3.361e-02A M=5.471e-07
I1549 0 n1550 3.361e-02A M=1.423e-06
I1550 0 n1551 3.361e-02A M=6.671e-07
I1551 0 n1552 3.361e-02A M=1.348e-06
I1552 0 n1553 3.361e-02A M=1.624e-06
I1553 0 n1554 3.361e-02A M=1.076e-06
I1554 0 n1555 3.361e-02A M=8.792e-07
I1555 0 n1556 3.361e-02A M=1.050e-06
I1556 0 n1557 3.361e-02A M=5.171e-07
I1557 0 n1558 3.361e-02A M=1.216e-06
I1558 0 n1559 3.361e-02A M=7.760e-07
I1559 0 n1560 3.361e-02A M=1.282e-06
I1560 0 n1561 3.361e-02A M=1.700e-07
I1561 0 n1562 3.361e-02A M=4.044e-07
I1562 0 n1563 3.361e-02A M=3.267e-07
I1563 0 n1564 3.361e-02A M=7.686e-07
I1564 0 n1565 3.361e-02A M=5.320e-07
I1565 0 n1566 3.361e-02A M=1.378e-06
I1566 0 n1567 3.361e-02A M=1.707e-06
I1567 0 n1568 3.361e-02A M=1.455e-06
I1568 0 n1569 3.361e-02A M=2.792e-07
I1569 0 n1570 3.361e-02A M=1.724e-06
I1570 0 n1571 3.361e-02A M=5.279e-07
I1571 0 n1572 3.361e-02A M=1.869e-06
I1572 0 n1573 3.361e-02A M=3.975e-07
I1573 0 n1574 3.361e-02A M=8.179e-07
I1574 0 n1575 3.361e-02A M=1.257e-06
I1575 0 n1576 3.361e-02A M=8.441e-07
I1576 0 n1577 3.361e-02A M=8.631e-07
I1577 0 n1578 3.361e-02A M=5.867e-07
I1578 0 n1579 3.361e-02A M=1.396e-06
I1579 0 n1580 3.361e-02A M=1.290e-06
I1580 0 n1581 3.361e-02A M=8.227e-07
I1581 0 n1582 3.361e-02A M=4.127e-07
I1582 0 n1583 3.361e-02A M=1.042e-06
I1583 0 n1584 3.361e-02A M=1.422e-06
I1584 0 n1585 3.361e-02A M=5.237e-07
I1585 0 n1586 3.361e-02A M=3.643e-07
I1586 0 n1587 3.361e-02A M=6.516e-07
I1587 0 n1588 3.361e-02A M=1.373e-06
I1588 0 n1589 3.361e-02A M=1.645e-06
I1589 0 n1590 3.361e-02A M=1.219e-06
I1590 0 n1591 3.361e-02A M=3.071e-07
I1591 0 n1592 3.361e-02A M=9.230e-07
I1592 0 n1593 3.361e-02A M=1.356e-06
I1593 0 n1594 3.361e-02A M=1.701e-06
I1594 0 n1595 3.361e-02A M=2.293e-06
I1595 0 n1596 3.361e-02A M=1.317e-06
I1596 0 n1597 3.361e-02A M=5.399e-07
I1597 0 n1598 3.361e-02A M=1.530e-06
I1598 0 n1599 3.361e-02A M=2.610e-07
I1599 0 n1600 3.361e-02A M=2.750e-07
I1600 0 n1601 3.361e-02A M=6.347e-07
I1601 0 n1602 3.361e-02A M=1.458e-06
I1602 0 n1603 3.361e-02A M=1.151e-06
I1603 0 n1604 3.361e-02A M=6.874e-07
I1604 0 n1605 3.361e-02A M=4.000e-07
I1605 0 n1606 3.361e-02A M=1.063e-06
I1606 0 n1607 3.361e-02A M=5.919e-07
I1607 0 n1608 3.361e-02A M=1.112e-06
I1608 0 n1609 3.361e-02A M=4.463e-07
I1609 0 n1610 3.361e-02A M=7.720e-07
I1610 0 n1611 3.361e-02A M=8.309e-07
I1611 0 n1612 3.361e-02A M=1.308e-06
I1612 0 n1613 3.361e-02A M=1.858e-07
I1613 0 n1614 3.361e-02A M=7.999e-07
I1614 0 n1615 3.361e-02A M=4.644e-07
I1615 0 n1616 3.361e-02A M=1.214e-06
I1616 0 n1617 3.361e-02A M=4.887e-07
I1617 0 n1618 3.361e-02A M=2.029e-06
I1618 0 n1619 3.361e-02A M=7.213e-07
I1619 0 n1620 3.361e-02A M=1.791e-06
I1620 0 n1621 3.361e-02A M=9.214e-07
I1621 0 n1622 3.361e-02A M=1.473e-06
I1622 0 n1623 3.361e-02A M=5.973e-07
I1623 0 n1624 3.361e-02A M=6.955e-07
I1624 0 n1625 3.361e-02A M=1.976e-06
I1625 0 n1626 3.361e-02A M=1.012e-06
I1626 0 n1627 3.361e-02A M=9.802e-07
I1627 0 n1628 3.361e-02A M=1.100e-06
I1628 0 n1629 3.361e-02A M=8.828e-07
I1629 0 n1630 3.361e-02A M=1.344e-06
I1630 0 n1631 3.361e-02A M=1.563e-06
I1631 0 n1632 3.361e-02A M=2.469e-06
I1632 0 n1633 3.361e-02A M=4.903e-07
I1633 0 n1634 3.361e-02A M=1.271e-06
I1634 0 n1635 3.361e-02A M=2.287e-06
I1635 0 n1636 3.361e-02A M=1.674e-06
I1636 0 n1637 3.361e-02A M=6.028e-07
I1637 0 n1638 3.361e-02A M=1.107e-06
I1638 0 n1639 3.361e-02A M=7.926e-07
I1639 0 n1640 3.361e-02A M=4.163e-07
I1640 0 n1641 3.361e-02A M=7.916e-07
I1641 0 n1642 3.361e-02A M=4.510e-07
I1642 0 n1643 3.361e-02A M=9.843e-07
I1643 0 n1644 3.361e-02A M=6.114e-07
I1644 0 n1645 3.361e-02A M=1.208e-06
I1645 0 n1646 3.361e-02A M=9.548e-07
I1646 0 n1647 3.361e-02A M=6.574e-07
I1647 0 n1648 3.361e-02A M=1.075e-06
I1648 0 n1649 3.361e-02A M=1.077e-06
I1649 0 n1650 3.361e-02A M=1.215e-06
I1650 0 n1651 3.361e-02A M=1.056e-06
I1651 0 n1652 3.361e-02A M=1.607e-06
I1652 0 n1653 3.361e-02A M=9.603e-07
I1653 0 n1654 3.361e-02A M=5.439e-07
I1654 0 n1655 3.361e-02A M=9.337e-07
I1655 0 n1656 3.361e-02A M=5.451e-07
I1656 0 n1657 3.361e-02A M=1.646e-06
I1657 0 n1658 3.361e-02A M=4.881e-07
I1658 0 n1659 3.361e-02A M=6.663e-07
I1659 0 n1660 3.361e-02A M=7.476e-07
I1660 0 n1661 3.361e-02A M=1.675e-06
I1661 0 n1662 3.361e-02A M=1.186e-06
I1662 0 n1663 3.361e-02A M=6.357e-07
I1663 0 n1664 3.361e-02A M=6.737e-07
I1664 0 n1665 3.361e-02A M=1.154e-06
I1665 0 n1666 3.361e-02A M=9.069e-07
I1666 0 n1667 3.361e-02A M=3.178e-07
I1667 0 n1668 3.361e-02A M=7.407e-07
I1668 0 n1669 3.361e-02A M=9.807e-07
I1669 0 n1670 3.361e-02A M=7.755e-07
I1670 0 n1671 3.361e-02A M=4.743e-07
I1671 0 n1672 3.361e-02A M=5.850e-07
I1672 0 n1673 3.361e-02A M=1.202e-06
I1673 0 n1674 3.361e-02A M=8.740e-07
I1674 0 n1675 3.361e-02A M=1.185e-06
I1675 0 n1676 3.361e-02A M=8.754e-07
I1676 0 n1677 3.361e-02A M=4.244e-07
I1677 0 n1678 3.361e-02A M=1.017e-06
I1678 0 n1679 3.361e-02A M=4.769e-07
I1679 0 n1680 3.361e-02A M=1.834e-06
I1680 0 n1681 3.361e-02A M=7.844e-07
I1681 0 n1682 3.361e-02A M=1.285e-06
I1682 0 n1683 3.361e-02A M=1.127e-06
I1683 0 n1684 3.361e-02A M=9.389e-07
I1684 0 n1685 3.361e-02A M=1.079e-06
I1685 0 n1686 3.361e-02A M=1.207e-06
I1686 0 n1687 3.361e-02A M=2.989e-07
I1687 0 n1688 3.361e-02A M=7.529e-07
I1688 0 n1689 3.361e-02A M=1.773e-06
I1689 0 n1690 3.361e-02A M=7.151e-07
I1690 0 n1691 3.361e-02A M=1.445e-06
I1691 0 n1692 3.361e-02A M=1.425e-06
I1692 0 n1693 3.361e-02A M=4.119e-07
I1693 0 n1694 3.361e-02A M=1.584e-06
I1694 0 n1695 3.361e-02A M=2.493e-06
I1695 0 n1696 3.361e-02A M=7.896e-07
I1696 0 n1697 3.361e-02A M=6.651e-07
I1697 0 n1698 3.361e-02A M=6.255e-07
I1698 0 n1699 3.361e-02A M=6.275e-07
I1699 0 n1700 3.361e-02A M=1.346e-06
I1700 0 n1701 3.361e-02A M=4.850e-07
I1701 0 n1702 3.361e-02A M=5.788e-07
I1702 0 n1703 3.361e-02A M=1.174e-06
I1703 0 n1704 3.361e-02A M=3.997e-07
I1704 0 n1705 3.361e-02A M=2.494e-07
I1705 0 n1706 3.361e-02A M=1.732e-06
I1706 0 n1707 3.361e-02A M=7.541e-07
I1707 0 n1708 3.361e-02A M=8.102e-07
I1708 0 n1 3.361e-02A M=1.761e-06
I1709 0 n1710 3.361e-02A M=1.113e-06
I1710 0 n1711 3.361e-02A M=8.577e-07
I1711 0 n1712 3.361e-02A M=5.294e-07
I1712 0 n1713 3.361e-02A M=5.657e-07
I1713 0 n1714 3.361e-02A M=5.179e-07
I1714 0 n1715 3.361e-02A M=7.940e-07
I1715 0 n1716 3.361e-02A M=1.025e-06
I1716 0 n1717 3.361e-02A M=7.158e-07
I1717 0 n1718 3.361e-02A M=8.097e-07
I1718 0 n1719 3.361e-02A M=1.363e-06
I1719 0 n1720 3.361e-02A M=5.915e-07
I1720 0 n1721 3.361e-02A M=5.939e-07
I1721 0 n1722 3.361e-02A M=1.247e-06
I1722 0 n1723 3.361e-02A M=9.818e-07
I1723 0 n1724 3.361e-02A M=9.705e-07
I1724 0 n1725 3.361e-02A M=2.419e-07
I1725 0 n1726 3.361e-02A M=1.146e-06
I1726 0 n1727 3.361e-02A M=1.975e-07
I1727 0 n1 3.361e-02A M=1.355e-06
I1728 0 n1729 3.361e-02A M=2.292e-07
I1729 0 n1730 3.361e-02A M=6.168e-07
I1730 0 n1731 3.361e-02A M=6.029e-07
I1731 0 n1732 3.361e-02A M=5.500e-07
I1732 0 n1733 3.361e-02A M=4.763e-07
I1733 0 n1734 3.361e-02A M=4.356e-07
I1734 0 n1735 3.361e-02A M=7.707e-07
I1735 0 n1736 3.361e-02A M=1.029e-06
I1736 0 n1737 3.361e-02A M=5.111e-07
I1737 0 n1738 3.361e-02A M=8.900e-07
I1738 0 n1739 3.361e-02A M=8.738e-07
I1739 0 n1740 3.361e-02A M=1.168e-06
I1740 0 n1741 3.361e-02A M=5.439e-07
I1741 0 n1742 3.361e-02A M=4.817e-07
I1742 0 n1743 3.361e-02A M=1.134e-06
I1743 0 n1744 3.361e-02A M=6.644e-07
I1744 0 n1745 3.361e-02A M=4.353e-07
I1745 0 n1746 3.361e-02A M=1.511e-06
I1746 0 n1747 3.361e-02A M=9.676e-07
I1747 0 n1748 3.361e-02A M=2.045e-07
I1748 0 n1749 3.361e-02A M=1.126e-06
I1749 0 n1750 3.361e-02A M=4.397e-07
I1750 0 n1751 3.361e-02A M=3.881e-07
I1751 0 n1752 3.361e-02A M=6.570e-07
I1752 0 n1753 3.361e-02A M=4.137e-07
I1753 0 n1754 3.361e-02A M=5.638e-07
I1754 0 n1755 3.361e-02A M=8.747e-07
I1755 0 n1756 3.361e-02A M=1.916e-06
I1756 0 n1757 3.361e-02A M=5.311e-07
I1757 0 n1758 3.361e-02A M=7.075e-07
I1758 0 n1759 3.361e-02A M=7.066e-07
I1759 0 n1760 3.361e-02A M=8.914e-07
I1760 0 n1761 3.361e-02A M=2.158e-06
I1761 0 n1762 3.361e-02A M=7.873e-07
I1762 0 n1763 3.361e-02A M=1.685e-06
I1763 0 n1764 3.361e-02A M=8.157e-07
I1764 0 n1765 3.361e-02A M=8.651e-07
I1765 0 n1766 3.361e-02A M=5.382e-07
I1766 0 n1767 3.361e-02A M=7.450e-07
I1767 0 n1768 3.361e-02A M=9.319e-07
I1768 0 n1769 3.361e-02A M=9.541e-07
I1769 0 n1770 3.361e-02A M=1.103e-06
I1770 0 n1771 3.361e-02A M=1.572e-06
I1771 0 n1772 3.361e-02A M=8.179e-07
I1772 0 n1773 3.361e-02A M=6.183e-07
I1773 0 n1774 3.361e-02A M=1.322e-06
I1774 0 n1775 3.361e-02A M=8.398e-07
I1775 0 n1776 3.361e-02A M=1.217e-06
I1776 0 n1777 3.361e-02A M=1.311e-06
I1777 0 n1778 3.361e-02A M=6.064e-07
I1778 0 n1779 3.361e-02A M=8.320e-07
I1779 0 n1 3.361e-02A M=8.696e-07
I1780 0 n1781 3.361e-02A M=1.507e-06
I1781 0 n1782 3.361e-02A M=3.721e-07
I1782 0 n1783 3.361e-02A M=3.797e-07
I1783 0 n1784 3.361e-02A M=5.793e-07
I1784 0 n1785 3.361e-02A M=1.820e-06
I1785 0 n1786 3.361e-02A M=1.533e-06
I1786 0 n1787 3.361e-02A M=1.111e-06
I1787 0 n1788 3.361e-02A M=8.177e-07
I1788 0 n1789 3.361e-02A M=1.631e-06
I1789 0 n1790 3.361e-02A M=2.270e-07
I1790 0 n1791 3.361e-02A M=2.160e-06
I1791 0 n1792 3.361e-02A M=6.184e-07
I1792 0 n1793 3.361e-02A M=7.211e-07
I1793 0 n1794 3.361e-02A M=5.235e-07
I1794 0 n1795 3.361e-02A M=3.409e-07
I1795 0 n1796 3.361e-02A M=8.828e-07
I1796 0 n1797 3.361e-02A M=9.487e-07
I1797 0 n1798 3.361e-02A M=1.057e-06
I1798 0 n1799 3.361e-02A M=9.554e-07
I1799 0 n1800 3.361e-02A M=8.900e-07
I1800 0 n1801 3.361e-02A M=1.936e-06
I1801 0 n1802 3.361e-02A M=7.800e-07
I1802 0 n1803 3.361e-02A M=1.100e-06
I1803 0 n1804 3.361e-02A M=1.349e-06
I1804 0 n1805 3.361e-02A M=4.342e-07
I1805 0 n1806 3.361e-02A M=1.128e-06
I1806 0 n1807 3.361e-02A M=1.009e-06
I1807 0 n1808 3.361e-02A M=1.054e-06
I1808 0 n1809 3.361e-02A M=7.419e-07
I1809 0 n1810 3.361e-02A M=1.314e-06
I1810 0 n1811 3.361e-02A M=4.422e-07
I1811 0 n1812 3.361e-02A M=5.065e-07
I1812 0 n1813 3.361e-02A M=2.391e-06
I1813 0 n1814 3.361e-02A M=1.926e-07
I1814 0 n1815 3.361e-02A M=7.329e-07
I1815 0 n1816 3.361e-02A M=1.278e-06
I1816 0 n1817 3.361e-02A M=5.955e-07
I1817 0 n1818 3.361e-02A M=1.687e-06
I1818 0 n1819 3.361e-02A M=3.173e-07
I1819 0 n1820 3.361e-02A M=1.580e-06
I1820 0 n1821 3.361e-02A M=1.134e-06
I1821 0 n1822 3.361e-02A M=1.168e-06
I1822 0 n1823 3.361e-02A M=5.286e-07
I1823 0 n1824 3.361e-02A M=5.607e-07
I1824 0 n1825 3.361e-02A M=5.255e-07
I1825 0 n1826 3.361e-02A M=9.545e-07
I1826 0 n1827 3.361e-02A M=1.373e-06
I1827 0 n1828 3.361e-02A M=1.903e-06
I1828 0 n1829 3.361e-02A M=1.101e-06
I1829 0 n1830 3.361e-02A M=1.456e-06
I1830 0 n1831 3.361e-02A M=7.024e-07
I1831 0 n1832 3.361e-02A M=7.832e-07
I1832 0 n1833 3.361e-02A M=6.755e-07
I1833 0 n1834 3.361e-02A M=1.466e-06
I1834 0 n1835 3.361e-02A M=1.033e-06
I1835 0 n1836 3.361e-02A M=4.725e-07
I1836 0 n1837 3.361e-02A M=9.210e-07
I1837 0 n1838 3.361e-02A M=8.962e-07
I1838 0 n1839 3.361e-02A M=3.838e-07
I1839 0 n1 3.361e-02A M=9.107e-07
I1840 0 n1841 3.361e-02A M=5.733e-07
I1841 0 n1842 3.361e-02A M=3.929e-07
I1842 0 n1843 3.361e-02A M=5.914e-07
I1843 0 n1844 3.361e-02A M=1.077e-06
I1844 0 n1845 3.361e-02A M=5.239e-07
I1845 0 n1846 3.361e-02A M=1.382e-06
I1846 0 n1847 3.361e-02A M=6.928e-07
I1847 0 n1848 3.361e-02A M=3.247e-07
I1848 0 n1849 3.361e-02A M=1.503e-06
I1849 0 n1850 3.361e-02A M=2.990e-07
I1850 0 n1851 3.361e-02A M=1.144e-06
I1851 0 n1852 3.361e-02A M=1.354e-06
I1852 0 n1853 3.361e-02A M=2.272e-07
I1853 0 n1854 3.361e-02A M=6.682e-07
I1854 0 n1855 3.361e-02A M=9.590e-07
I1855 0 n1856 3.361e-02A M=1.176e-06
I1856 0 n1857 3.361e-02A M=1.351e-06
I1857 0 n1858 3.361e-02A M=2.460e-06
I1858 0 n1859 3.361e-02A M=3.457e-07
I1859 0 n1860 3.361e-02A M=8.739e-07
I1860 0 n1861 3.361e-02A M=5.680e-07
I1861 0 n1862 3.361e-02A M=1.812e-06
I1862 0 n1863 3.361e-02A M=1.108e-06
I1863 0 n1864 3.361e-02A M=2.142e-06
I1864 0 n1865 3.361e-02A M=1.450e-06
I1865 0 n1866 3.361e-02A M=1.452e-06
I1866 0 n1867 3.361e-02A M=4.373e-07
I1867 0 n1868 3.361e-02A M=3.395e-06
I1868 0 n1869 3.361e-02A M=1.463e-06
I1869 0 n1870 3.361e-02A M=6.692e-07
I1870 0 n1871 3.361e-02A M=7.720e-07
I1871 0 n1872 3.361e-02A M=6.258e-07
I1872 0 n1873 3.361e-02A M=1.567e-06
I1873 0 n1874 3.361e-02A M=5.428e-07
I1874 0 n1875 3.361e-02A M=1.265e-06
I1875 0 n1876 3.361e-02A M=9.783e-07
I1876 0 n1877 3.361e-02A M=3.971e-07
I1877 0 n1878 3.361e-02A M=1.812e-07
I1878 0 n1879 3.361e-02A M=5.318e-07
I1879 0 n1880 3.361e-02A M=1.979e-06
I1880 0 n1881 3.361e-02A M=1.549e-06
I1881 0 n1882 3.361e-02A M=8.546e-07
I1882 0 n1883 3.361e-02A M=7.570e-07
I1883 0 n1884 3.361e-02A M=1.481e-06
I1884 0 n1885 3.361e-02A M=1.527e-06
I1885 0 n1886 3.361e-02A M=5.426e-07
I1886 0 n1887 3.361e-02A M=1.632e-06
I1887 0 n1888 3.361e-02A M=9.617e-07
I1888 0 n1889 3.361e-02A M=1.371e-06
I1889 0 n1 3.361e-02A M=1.945e-06
I1890 0 n1891 3.361e-02A M=6.287e-07
I1891 0 n1892 3.361e-02A M=4.215e-07
I1892 0 n1893 3.361e-02A M=1.331e-06
I1893 0 n1894 3.361e-02A M=1.685e-06
I1894 0 n1895 3.361e-02A M=5.664e-07
I1895 0 n1896 3.361e-02A M=1.140e-06
I1896 0 n1897 3.361e-02A M=6.472e-07
I1897 0 n1898 3.361e-02A M=5.483e-07
I1898 0 n1899 3.361e-02A M=2.713e-07
I1899 0 n1900 3.361e-02A M=6.003e-07
I1900 0 n1901 3.361e-02A M=5.354e-07
I1901 0 n1902 3.361e-02A M=1.838e-06
I1902 0 n1903 3.361e-02A M=1.767e-06
I1903 0 n1904 3.361e-02A M=7.617e-07
I1904 0 n1905 3.361e-02A M=1.074e-06
I1905 0 n1906 3.361e-02A M=1.049e-06
I1906 0 n1907 3.361e-02A M=1.433e-06
I1907 0 n1908 3.361e-02A M=9.792e-07
I1908 0 n1909 3.361e-02A M=8.329e-07
I1909 0 n1910 3.361e-02A M=1.620e-06
I1910 0 n1911 3.361e-02A M=9.725e-07
I1911 0 n1912 3.361e-02A M=9.399e-07
I1912 0 n1913 3.361e-02A M=7.100e-07
I1913 0 n1914 3.361e-02A M=8.681e-07
I1914 0 n1915 3.361e-02A M=3.674e-07
I1915 0 n1916 3.361e-02A M=8.930e-07
I1916 0 n1917 3.361e-02A M=1.263e-06
I1917 0 n1918 3.361e-02A M=7.159e-07
I1918 0 n1919 3.361e-02A M=4.992e-07
I1919 0 n1920 3.361e-02A M=2.990e-07
I1920 0 n1921 3.361e-02A M=5.317e-07
I1921 0 n1922 3.361e-02A M=1.403e-06
I1922 0 n1923 3.361e-02A M=1.171e-06
I1923 0 n1924 3.361e-02A M=1.828e-06
I1924 0 n1925 3.361e-02A M=5.098e-07
I1925 0 n1926 3.361e-02A M=8.252e-07
I1926 0 n1927 3.361e-02A M=1.780e-06
I1927 0 n1928 3.361e-02A M=5.749e-07
I1928 0 n1929 3.361e-02A M=1.676e-06
I1929 0 n1930 3.361e-02A M=8.815e-07
I1930 0 n1931 3.361e-02A M=2.486e-06
I1931 0 n1932 3.361e-02A M=7.559e-07
I1932 0 n1933 3.361e-02A M=5.553e-07
I1933 0 n1934 3.361e-02A M=2.311e-07
I1934 0 n1935 3.361e-02A M=1.905e-06
I1935 0 n1936 3.361e-02A M=1.660e-06
I1936 0 n1937 3.361e-02A M=1.035e-06
I1937 0 n1938 3.361e-02A M=1.131e-06
I1938 0 n1939 3.361e-02A M=4.850e-07
I1939 0 n1940 3.361e-02A M=8.489e-07
I1940 0 n1941 3.361e-02A M=5.676e-07
I1941 0 n1942 3.361e-02A M=1.102e-06
I1942 0 n1943 3.361e-02A M=5.554e-07
I1943 0 n1944 3.361e-02A M=1.114e-06
I1944 0 n1945 3.361e-02A M=2.621e-07
I1945 0 n1946 3.361e-02A M=1.251e-06
I1946 0 n1947 3.361e-02A M=1.272e-06
I1947 0 n1948 3.361e-02A M=8.436e-07
I1948 0 n1949 3.361e-02A M=7.420e-07
I1949 0 n1950 3.361e-02A M=2.302e-06
I1950 0 n1951 3.361e-02A M=8.677e-07
I1951 0 n1952 3.361e-02A M=9.340e-07
I1952 0 n1953 3.361e-02A M=7.134e-07
I1953 0 n1954 3.361e-02A M=9.262e-07
I1954 0 n1955 3.361e-02A M=5.572e-07
I1955 0 n1956 3.361e-02A M=5.127e-07
I1956 0 n1957 3.361e-02A M=1.276e-06
I1957 0 n1958 3.361e-02A M=6.688e-07
I1958 0 n1959 3.361e-02A M=1.231e-06
I1959 0 n1960 3.361e-02A M=7.938e-07
I1960 0 n1961 3.361e-02A M=8.031e-07
I1961 0 n1962 3.361e-02A M=8.574e-07
I1962 0 n1963 3.361e-02A M=7.206e-07
I1963 0 n1964 3.361e-02A M=4.988e-07
I1964 0 n1965 3.361e-02A M=3.581e-07
I1965 0 n1966 3.361e-02A M=6.842e-07
I1966 0 n1967 3.361e-02A M=9.246e-07
I1967 0 n1968 3.361e-02A M=4.888e-07
I1968 0 n1969 3.361e-02A M=6.645e-07
I1969 0 n1970 3.361e-02A M=1.438e-06
I1970 0 n1971 3.361e-02A M=6.130e-07
I1971 0 n1972 3.361e-02A M=9.062e-07
I1972 0 n1973 3.361e-02A M=1.131e-06
I1973 0 n1974 3.361e-02A M=9.959e-07
I1974 0 n1975 3.361e-02A M=2.902e-07
I1975 0 n1976 3.361e-02A M=1.210e-06
I1976 0 n1977 3.361e-02A M=6.489e-07
I1977 0 n1978 3.361e-02A M=5.623e-07
I1978 0 n1979 3.361e-02A M=5.890e-07
I1979 0 n1980 3.361e-02A M=9.539e-07
I1980 0 n1981 3.361e-02A M=9.019e-07
I1981 0 n1982 3.361e-02A M=6.243e-07
I1982 0 n1983 3.361e-02A M=2.000e-07
I1983 0 n1984 3.361e-02A M=1.057e-06
I1984 0 n1985 3.361e-02A M=1.035e-06
I1985 0 n1986 3.361e-02A M=2.327e-07
I1986 0 n1987 3.361e-02A M=1.612e-06
I1987 0 n1988 3.361e-02A M=2.959e-07
I1988 0 n1989 3.361e-02A M=9.459e-07
I1989 0 n1990 3.361e-02A M=1.021e-06
I1990 0 n1991 3.361e-02A M=6.459e-07
I1991 0 n1992 3.361e-02A M=1.777e-07
I1992 0 n1993 3.361e-02A M=1.181e-06
I1993 0 n1994 3.361e-02A M=5.034e-07
I1994 0 n1995 3.361e-02A M=3.116e-07
I1995 0 n1996 3.361e-02A M=1.757e-06
I1996 0 n1 3.361e-02A M=2.182e-07
I1997 0 n1998 3.361e-02A M=5.162e-07
I1998 0 n1999 3.361e-02A M=9.234e-08
I1999 0 n2000 3.361e-02A M=7.823e-07
I2000 0 n2001 3.361e-02A M=6.867e-07
I2001 0 n2002 3.361e-02A M=6.581e-07
I2002 0 n2003 3.361e-02A M=5.059e-07
I2003 0 n2004 3.361e-02A M=1.097e-06
I2004 0 n2005 3.361e-02A M=1.000e-06
I2005 0 n2006 3.361e-02A M=2.263e-06
I2006 0 n2007 3.361e-02A M=7.413e-07
I2007 0 n2008 3.361e-02A M=3.027e-07
I2008 0 n2009 3.361e-02A M=1.505e-06
I2009 0 n2010 3.361e-02A M=7.689e-07
I2010 0 n2011 3.361e-02A M=1.843e-06
I2011 0 n2012 3.361e-02A M=6.532e-07
I2012 0 n2013 3.361e-02A M=8.499e-07
I2013 0 n2014 3.361e-02A M=1.216e-06
I2014 0 n2015 3.361e-02A M=9.929e-07
I2015 0 n2016 3.361e-02A M=1.165e-06
I2016 0 n2017 3.361e-02A M=9.895e-07
I2017 0 n2018 3.361e-02A M=1.855e-06
I2018 0 n2019 3.361e-02A M=1.189e-06
I2019 0 n2020 3.361e-02A M=1.426e-06
I2020 0 n2021 3.361e-02A M=2.278e-07
I2021 0 n2022 3.361e-02A M=1.057e-06
I2022 0 n2023 3.361e-02A M=5.373e-07
I2023 0 n2024 3.361e-02A M=1.290e-06
I2024 0 n2025 3.361e-02A M=4.603e-07
I2025 0 n2026 3.361e-02A M=3.859e-07
I2026 0 n2027 3.361e-02A M=7.638e-07
I2027 0 n2028 3.361e-02A M=1.768e-06
I2028 0 n2029 3.361e-02A M=1.986e-06
I2029 0 n2030 3.361e-02A M=6.722e-07
I2030 0 n2031 3.361e-02A M=8.353e-07
I2031 0 n2032 3.361e-02A M=8.105e-07
I2032 0 n2033 3.361e-02A M=9.030e-07
I2033 0 n2034 3.361e-02A M=1.670e-06
I2034 0 n2035 3.361e-02A M=8.652e-07
I2035 0 n2036 3.361e-02A M=9.608e-07
I2036 0 n2037 3.361e-02A M=8.426e-07
I2037 0 n2038 3.361e-02A M=2.499e-07
I2038 0 n2039 3.361e-02A M=8.031e-07
I2039 0 n2040 3.361e-02A M=1.334e-06
I2040 0 n2041 3.361e-02A M=9.767e-07
I2041 0 n2042 3.361e-02A M=1.655e-06
I2042 0 n2043 3.361e-02A M=4.985e-07
I2043 0 n2044 3.361e-02A M=8.287e-07
I2044 0 n2045 3.361e-02A M=5.938e-07
I2045 0 n2046 3.361e-02A M=6.605e-07
I2046 0 n1 3.361e-02A M=1.342e-06
I2047 0 n2048 3.361e-02A M=8.033e-07
I2048 0 n2049 3.361e-02A M=3.635e-07
I2049 0 n2050 3.361e-02A M=7.804e-07
I2050 0 n2051 3.361e-02A M=1.177e-06
I2051 0 n2052 3.361e-02A M=1.547e-06
I2052 0 n2053 3.361e-02A M=1.432e-06
I2053 0 n2054 3.361e-02A M=8.775e-07
I2054 0 n2055 3.361e-02A M=2.473e-06
I2055 0 n2056 3.361e-02A M=7.864e-07
I2056 0 n2057 3.361e-02A M=6.706e-07
I2057 0 n2058 3.361e-02A M=6.701e-07
I2058 0 n2059 3.361e-02A M=1.046e-06
I2059 0 n2060 3.361e-02A M=5.647e-07
I2060 0 n2061 3.361e-02A M=1.498e-06
I2061 0 n2062 3.361e-02A M=7.948e-07
I2062 0 n2063 3.361e-02A M=3.449e-07
I2063 0 n1 3.361e-02A M=1.298e-06
I2064 0 n2065 3.361e-02A M=1.233e-06
I2065 0 n2066 3.361e-02A M=8.322e-07
I2066 0 n2067 3.361e-02A M=9.901e-08
I2067 0 n2068 3.361e-02A M=1.405e-06
I2068 0 n2069 3.361e-02A M=6.567e-07
I2069 0 n2070 3.361e-02A M=6.759e-07
I2070 0 n2071 3.361e-02A M=1.327e-06
I2071 0 n2072 3.361e-02A M=9.444e-07
I2072 0 n2073 3.361e-02A M=7.577e-07
I2073 0 n2074 3.361e-02A M=2.917e-06
I2074 0 n2075 3.361e-02A M=7.127e-07
I2075 0 n2076 3.361e-02A M=8.658e-07
I2076 0 n2077 3.361e-02A M=1.321e-06
I2077 0 n2078 3.361e-02A M=6.208e-07
I2078 0 n2079 3.361e-02A M=1.302e-06
I2079 0 n2080 3.361e-02A M=3.437e-07
I2080 0 n2081 3.361e-02A M=2.784e-06
I2081 0 n2082 3.361e-02A M=9.780e-07
I2082 0 n2083 3.361e-02A M=8.265e-07
I2083 0 n2084 3.361e-02A M=8.540e-07
I2084 0 n2085 3.361e-02A M=7.410e-07
I2085 0 n2086 3.361e-02A M=5.644e-07
I2086 0 n2087 3.361e-02A M=1.194e-06
I2087 0 n2088 3.361e-02A M=1.243e-06
I2088 0 n2089 3.361e-02A M=6.347e-07
I2089 0 n2090 3.361e-02A M=8.021e-07
I2090 0 n2091 3.361e-02A M=6.030e-07
I2091 0 n1 3.361e-02A M=7.243e-07
I2092 0 n2093 3.361e-02A M=5.088e-07
I2093 0 n2094 3.361e-02A M=1.932e-06
I2094 0 n2095 3.361e-02A M=2.083e-06
I2095 0 n2096 3.361e-02A M=1.405e-06
I2096 0 n2097 3.361e-02A M=3.500e-07
I2097 0 n2098 3.361e-02A M=6.614e-07
I2098 0 n2099 3.361e-02A M=1.235e-06
I2099 0 n2100 3.361e-02A M=2.291e-06
I2100 0 n2101 3.361e-02A M=1.549e-06
I2101 0 n2102 3.361e-02A M=9.375e-07
I2102 0 n2103 3.361e-02A M=1.239e-06
I2103 0 n2104 3.361e-02A M=6.257e-07
I2104 0 n2105 3.361e-02A M=7.990e-07
I2105 0 n2106 3.361e-02A M=2.039e-06
I2106 0 n2107 3.361e-02A M=1.122e-06
I2107 0 n2108 3.361e-02A M=1.017e-06
I2108 0 n2109 3.361e-02A M=1.618e-06
I2109 0 n2110 3.361e-02A M=6.361e-07
I2110 0 n2111 3.361e-02A M=1.836e-06
I2111 0 n2112 3.361e-02A M=1.302e-06
I2112 0 n2113 3.361e-02A M=7.981e-07
I2113 0 n2114 3.361e-02A M=7.469e-07
I2114 0 n2115 3.361e-02A M=1.063e-06
I2115 0 n2116 3.361e-02A M=1.786e-06
I2116 0 n2117 3.361e-02A M=9.167e-07
I2117 0 n2118 3.361e-02A M=1.659e-06
I2118 0 n2119 3.361e-02A M=1.126e-06
I2119 0 n2120 3.361e-02A M=1.783e-06
I2120 0 n2121 3.361e-02A M=4.838e-07
I2121 0 n2122 3.361e-02A M=1.865e-07
I2122 0 n2123 3.361e-02A M=4.438e-07
I2123 0 n2124 3.361e-02A M=8.383e-07
I2124 0 n2125 3.361e-02A M=7.571e-07
I2125 0 n2126 3.361e-02A M=8.509e-07
I2126 0 n2127 3.361e-02A M=4.608e-07
I2127 0 n2128 3.361e-02A M=5.149e-07
I2128 0 n2129 3.361e-02A M=1.741e-06
I2129 0 n2130 3.361e-02A M=2.036e-07
I2130 0 n2131 3.361e-02A M=4.481e-07
I2131 0 n2132 3.361e-02A M=6.967e-07
I2132 0 n2133 3.361e-02A M=6.966e-07
I2133 0 n2134 3.361e-02A M=4.792e-07
I2134 0 n2135 3.361e-02A M=1.373e-06
I2135 0 n2136 3.361e-02A M=1.397e-06
I2136 0 n2137 3.361e-02A M=3.190e-07
I2137 0 n2138 3.361e-02A M=1.173e-06
I2138 0 n2139 3.361e-02A M=9.706e-07
I2139 0 n2140 3.361e-02A M=6.463e-07
I2140 0 n2141 3.361e-02A M=1.744e-06
I2141 0 n2142 3.361e-02A M=1.434e-07
I2142 0 n2143 3.361e-02A M=9.602e-07
I2143 0 n2144 3.361e-02A M=9.740e-07
I2144 0 n2145 3.361e-02A M=4.950e-07
I2145 0 n2146 3.361e-02A M=6.387e-07
I2146 0 n2147 3.361e-02A M=7.913e-07
I2147 0 n2148 3.361e-02A M=1.062e-06
I2148 0 n2149 3.361e-02A M=7.029e-07
I2149 0 n2150 3.361e-02A M=8.487e-07
I2150 0 n2151 3.361e-02A M=9.049e-07
I2151 0 n2152 3.361e-02A M=4.044e-07
I2152 0 n2153 3.361e-02A M=9.971e-07
I2153 0 n2154 3.361e-02A M=8.425e-07
I2154 0 n2155 3.361e-02A M=2.906e-06
I2155 0 n2156 3.361e-02A M=8.577e-07
I2156 0 n2157 3.361e-02A M=6.364e-07
I2157 0 n2158 3.361e-02A M=1.213e-06
I2158 0 n2159 3.361e-02A M=1.787e-06
I2159 0 n2160 3.361e-02A M=4.385e-07
I2160 0 n2161 3.361e-02A M=1.577e-06
I2161 0 n2162 3.361e-02A M=1.406e-07
I2162 0 n2163 3.361e-02A M=4.220e-07
I2163 0 n2164 3.361e-02A M=2.298e-06
I2164 0 n2165 3.361e-02A M=2.135e-06
I2165 0 n2166 3.361e-02A M=4.399e-07
I2166 0 n2167 3.361e-02A M=1.004e-06
I2167 0 n2168 3.361e-02A M=6.744e-07
I2168 0 n2169 3.361e-02A M=1.557e-06
I2169 0 n2170 3.361e-02A M=9.895e-07
I2170 0 n2171 3.361e-02A M=4.565e-07
I2171 0 n2172 3.361e-02A M=7.064e-07
I2172 0 n2173 3.361e-02A M=2.167e-06
I2173 0 n2174 3.361e-02A M=8.865e-07
I2174 0 n2175 3.361e-02A M=1.032e-06
I2175 0 n2176 3.361e-02A M=5.922e-07
I2176 0 n2177 3.361e-02A M=1.342e-06
I2177 0 n2178 3.361e-02A M=8.342e-07
I2178 0 n2179 3.361e-02A M=8.205e-07
I2179 0 n2180 3.361e-02A M=6.534e-07
I2180 0 n2181 3.361e-02A M=8.362e-07
I2181 0 n2182 3.361e-02A M=8.987e-07
I2182 0 n2183 3.361e-02A M=4.565e-07
I2183 0 n2184 3.361e-02A M=2.401e-06
I2184 0 n2185 3.361e-02A M=9.465e-07
I2185 0 n2186 3.361e-02A M=6.285e-07
I2186 0 n2187 3.361e-02A M=9.879e-07
I2187 0 n2188 3.361e-02A M=7.897e-07
I2188 0 n2189 3.361e-02A M=1.046e-06
I2189 0 n2190 3.361e-02A M=1.663e-06
I2190 0 n2191 3.361e-02A M=4.882e-07
I2191 0 n2192 3.361e-02A M=1.737e-06
I2192 0 n2193 3.361e-02A M=1.034e-06
I2193 0 n2194 3.361e-02A M=1.200e-06
I2194 0 n2195 3.361e-02A M=1.549e-06
I2195 0 n2196 3.361e-02A M=1.215e-06
I2196 0 n2197 3.361e-02A M=2.714e-07
I2197 0 n2198 3.361e-02A M=3.861e-07
I2198 0 n1 3.361e-02A M=3.887e-07
I2199 0 n2200 3.361e-02A M=3.319e-07
I2200 0 n2201 3.361e-02A M=2.867e-07
I2201 0 n2202 3.361e-02A M=9.656e-07
I2202 0 n2203 3.361e-02A M=6.323e-07
I2203 0 n2204 3.361e-02A M=6.459e-07
I2204 0 n2205 3.361e-02A M=5.207e-07
I2205 0 n2206 3.361e-02A M=1.634e-06
I2206 0 n2207 3.361e-02A M=1.210e-06
I2207 0 n2208 3.361e-02A M=4.689e-07
I2208 0 n2209 3.361e-02A M=4.464e-07
I2209 0 n2210 3.361e-02A M=8.206e-07
I2210 0 n2211 3.361e-02A M=2.393e-07
I2211 0 n2212 3.361e-02A M=2.062e-06
I2212 0 n2213 3.361e-02A M=7.537e-07
I2213 0 n2214 3.361e-02A M=2.761e-06
I2214 0 n2215 3.361e-02A M=6.550e-07
I2215 0 n2216 3.361e-02A M=8.558e-07
I2216 0 n2217 3.361e-02A M=1.511e-06
I2217 0 n2218 3.361e-02A M=7.508e-08
I2218 0 n2219 3.361e-02A M=5.346e-07
I2219 0 n2220 3.361e-02A M=1.361e-06
I2220 0 n2221 3.361e-02A M=2.811e-07
I2221 0 n2222 3.361e-02A M=9.220e-07
I2222 0 n2223 3.361e-02A M=5.009e-07
I2223 0 n2224 3.361e-02A M=5.430e-07
I2224 0 n2225 3.361e-02A M=6.140e-07
I2225 0 n2226 3.361e-02A M=1.192e-06
I2226 0 n2227 3.361e-02A M=9.044e-07
I2227 0 n2228 3.361e-02A M=1.476e-06
I2228 0 n2229 3.361e-02A M=1.875e-06
I2229 0 n2230 3.361e-02A M=9.268e-07
I2230 0 n2231 3.361e-02A M=2.750e-06
I2231 0 n2232 3.361e-02A M=2.554e-06
I2232 0 n2233 3.361e-02A M=8.788e-07
I2233 0 n2234 3.361e-02A M=1.265e-06
I2234 0 n2235 3.361e-02A M=1.327e-06
I2235 0 n2236 3.361e-02A M=4.242e-07
I2236 0 n2237 3.361e-02A M=4.978e-07
I2237 0 n2238 3.361e-02A M=1.125e-06
I2238 0 n2239 3.361e-02A M=6.187e-07
I2239 0 n2240 3.361e-02A M=7.677e-07
I2240 0 n2241 3.361e-02A M=4.882e-07
I2241 0 n2242 3.361e-02A M=5.364e-07
I2242 0 n2243 3.361e-02A M=7.884e-07
I2243 0 n2244 3.361e-02A M=9.529e-07
I2244 0 n2245 3.361e-02A M=1.449e-06
I2245 0 n2246 3.361e-02A M=7.995e-07
I2246 0 n2247 3.361e-02A M=1.856e-07
I2247 0 n2248 3.361e-02A M=1.395e-06
I2248 0 n2249 3.361e-02A M=4.439e-07
I2249 0 n2250 3.361e-02A M=1.138e-06
I2250 0 n2251 3.361e-02A M=1.429e-06
I2251 0 n2252 3.361e-02A M=8.008e-07
I2252 0 n2253 3.361e-02A M=4.394e-07
I2253 0 n2254 3.361e-02A M=5.451e-07
I2254 0 n2255 3.361e-02A M=6.261e-07
I2255 0 n2256 3.361e-02A M=1.005e-06
I2256 0 n2257 3.361e-02A M=1.515e-06
I2257 0 n2258 3.361e-02A M=1.178e-06
I2258 0 n2259 3.361e-02A M=2.041e-06
I2259 0 n2260 3.361e-02A M=2.133e-06
I2260 0 n2261 3.361e-02A M=4.922e-07
I2261 0 n2262 3.361e-02A M=1.363e-06
I2262 0 n2263 3.361e-02A M=3.755e-07
I2263 0 n2264 3.361e-02A M=1.050e-06
I2264 0 n2265 3.361e-02A M=9.658e-07
I2265 0 n2266 3.361e-02A M=8.345e-07
I2266 0 n2267 3.361e-02A M=5.907e-07
I2267 0 n2268 3.361e-02A M=7.686e-07
I2268 0 n2269 3.361e-02A M=8.875e-07
I2269 0 n2270 3.361e-02A M=5.714e-07
I2270 0 n2271 3.361e-02A M=1.160e-06
I2271 0 n2272 3.361e-02A M=2.971e-07
I2272 0 n2273 3.361e-02A M=5.009e-07
I2273 0 n2274 3.361e-02A M=4.281e-07
I2274 0 n2275 3.361e-02A M=8.384e-07
I2275 0 n2276 3.361e-02A M=1.606e-06
I2276 0 n2277 3.361e-02A M=2.624e-06
I2277 0 n2278 3.361e-02A M=1.203e-06
I2278 0 n2279 3.361e-02A M=5.137e-07
I2279 0 n2280 3.361e-02A M=9.832e-07
I2280 0 n2281 3.361e-02A M=2.251e-06
I2281 0 n2282 3.361e-02A M=3.836e-07
I2282 0 n2283 3.361e-02A M=2.938e-07
I2283 0 n2284 3.361e-02A M=7.985e-07
I2284 0 n2285 3.361e-02A M=1.663e-06
I2285 0 n2286 3.361e-02A M=6.374e-07
I2286 0 n2287 3.361e-02A M=8.369e-07
I2287 0 n2288 3.361e-02A M=9.742e-07
I2288 0 n2289 3.361e-02A M=8.272e-07
I2289 0 n2290 3.361e-02A M=7.935e-07
I2290 0 n2291 3.361e-02A M=1.067e-06
I2291 0 n2292 3.361e-02A M=1.255e-06
I2292 0 n2293 3.361e-02A M=6.951e-07
I2293 0 n2294 3.361e-02A M=9.446e-07
I2294 0 n2295 3.361e-02A M=8.201e-07
I2295 0 n2296 3.361e-02A M=1.428e-06
I2296 0 n2297 3.361e-02A M=2.120e-07
I2297 0 n2298 3.361e-02A M=1.543e-06
I2298 0 n2299 3.361e-02A M=1.925e-06
I2299 0 n2300 3.361e-02A M=7.082e-07
I2300 0 n2301 3.361e-02A M=4.028e-07
I2301 0 n2302 3.361e-02A M=9.104e-07
I2302 0 n2303 3.361e-02A M=2.067e-07
I2303 0 n2304 3.361e-02A M=4.619e-07
I2304 0 n2305 3.361e-02A M=1.323e-06
I2305 0 n2306 3.361e-02A M=7.307e-07
I2306 0 n2307 3.361e-02A M=8.662e-07
I2307 0 n2308 3.361e-02A M=6.367e-07
I2308 0 n2309 3.361e-02A M=2.154e-06
I2309 0 n2310 3.361e-02A M=2.136e-07
I2310 0 n2311 3.361e-02A M=1.175e-06
I2311 0 n2312 3.361e-02A M=8.020e-07
I2312 0 n2313 3.361e-02A M=2.294e-06
I2313 0 n2314 3.361e-02A M=1.538e-06
I2314 0 n2315 3.361e-02A M=5.259e-07
I2315 0 n2316 3.361e-02A M=1.132e-06
I2316 0 n2317 3.361e-02A M=4.362e-07
I2317 0 n2318 3.361e-02A M=2.112e-06
I2318 0 n2319 3.361e-02A M=6.480e-07
I2319 0 n2320 3.361e-02A M=9.173e-07
I2320 0 n2321 3.361e-02A M=3.056e-07
I2321 0 n2322 3.361e-02A M=8.414e-07
I2322 0 n2323 3.361e-02A M=7.563e-07
I2323 0 n2324 3.361e-02A M=1.352e-06
I2324 0 n2325 3.361e-02A M=8.671e-07
I2325 0 n2326 3.361e-02A M=1.518e-06
I2326 0 n2327 3.361e-02A M=1.754e-06
I2327 0 n2328 3.361e-02A M=1.782e-06
I2328 0 n2329 3.361e-02A M=1.475e-06
I2329 0 n2330 3.361e-02A M=9.287e-07
I2330 0 n2331 3.361e-02A M=8.393e-07
I2331 0 n2332 3.361e-02A M=1.769e-06
I2332 0 n2333 3.361e-02A M=1.999e-06
I2333 0 n2334 3.361e-02A M=1.345e-06
I2334 0 n2335 3.361e-02A M=7.447e-07
I2335 0 n2336 3.361e-02A M=4.393e-07
I2336 0 n2337 3.361e-02A M=1.258e-06
I2337 0 n2338 3.361e-02A M=1.236e-06
I2338 0 n2339 3.361e-02A M=1.099e-06
I2339 0 n2340 3.361e-02A M=1.862e-06
I2340 0 n2341 3.361e-02A M=9.950e-07
I2341 0 n2342 3.361e-02A M=1.088e-06
I2342 0 n2343 3.361e-02A M=1.170e-06
I2343 0 n2344 3.361e-02A M=1.531e-06
I2344 0 n2345 3.361e-02A M=8.198e-07
I2345 0 n2346 3.361e-02A M=1.329e-06
I2346 0 n2347 3.361e-02A M=1.320e-06
I2347 0 n2348 3.361e-02A M=7.072e-07
I2348 0 n2349 3.361e-02A M=3.952e-07
I2349 0 n2350 3.361e-02A M=1.853e-06
I2350 0 n2351 3.361e-02A M=7.631e-07
I2351 0 n2352 3.361e-02A M=1.628e-06
I2352 0 n2353 3.361e-02A M=9.407e-07
I2353 0 n2354 3.361e-02A M=8.857e-07
I2354 0 n2355 3.361e-02A M=4.743e-07
I2355 0 n2356 3.361e-02A M=1.207e-06
I2356 0 n2357 3.361e-02A M=6.741e-07
I2357 0 n2358 3.361e-02A M=9.194e-07
I2358 0 n2359 3.361e-02A M=7.249e-07
I2359 0 n2360 3.361e-02A M=1.275e-06
I2360 0 n2361 3.361e-02A M=8.858e-07
I2361 0 n2362 3.361e-02A M=2.503e-06
I2362 0 n2363 3.361e-02A M=5.120e-07
I2363 0 n2364 3.361e-02A M=7.487e-07
I2364 0 n2365 3.361e-02A M=2.591e-07
I2365 0 n2366 3.361e-02A M=2.260e-06
I2366 0 n2367 3.361e-02A M=1.291e-06
I2367 0 n2368 3.361e-02A M=1.565e-06
I2368 0 n2369 3.361e-02A M=7.624e-07
I2369 0 n2370 3.361e-02A M=9.977e-07
I2370 0 n2371 3.361e-02A M=1.933e-06
I2371 0 n2372 3.361e-02A M=1.290e-06
I2372 0 n2373 3.361e-02A M=1.131e-06
I2373 0 n2374 3.361e-02A M=2.511e-07
I2374 0 n2375 3.361e-02A M=9.276e-07
I2375 0 n2376 3.361e-02A M=8.498e-07
I2376 0 n2377 3.361e-02A M=4.500e-07
I2377 0 n2378 3.361e-02A M=3.602e-07
I2378 0 n2379 3.361e-02A M=7.984e-07
I2379 0 n2380 3.361e-02A M=1.047e-06
I2380 0 n2381 3.361e-02A M=1.292e-06
I2381 0 n2382 3.361e-02A M=1.629e-06
I2382 0 n2383 3.361e-02A M=1.893e-06
I2383 0 n2384 3.361e-02A M=1.034e-06
I2384 0 n2385 3.361e-02A M=4.862e-07
I2385 0 n2386 3.361e-02A M=1.734e-06
I2386 0 n2387 3.361e-02A M=4.733e-07
I2387 0 n2388 3.361e-02A M=1.608e-06
I2388 0 n2389 3.361e-02A M=6.259e-07
I2389 0 n2390 3.361e-02A M=7.946e-07
I2390 0 n2391 3.361e-02A M=2.454e-06
I2391 0 n2392 3.361e-02A M=1.308e-06
I2392 0 n2393 3.361e-02A M=1.391e-06
I2393 0 n2394 3.361e-02A M=8.803e-07
I2394 0 n2395 3.361e-02A M=8.492e-07
I2395 0 n1 3.361e-02A M=8.314e-07
I2396 0 n2397 3.361e-02A M=1.646e-06
I2397 0 n2398 3.361e-02A M=4.386e-07
I2398 0 n2399 3.361e-02A M=9.774e-07
I2399 0 n2400 3.361e-02A M=7.101e-07
I2400 0 n2401 3.361e-02A M=4.350e-07
I2401 0 n2402 3.361e-02A M=1.627e-06
I2402 0 n2403 3.361e-02A M=1.000e-06
I2403 0 n2404 3.361e-02A M=1.339e-06
I2404 0 n2405 3.361e-02A M=2.530e-06
I2405 0 n2406 3.361e-02A M=1.793e-07
I2406 0 n2407 3.361e-02A M=4.290e-07
I2407 0 n2408 3.361e-02A M=4.382e-07
I2408 0 n2409 3.361e-02A M=5.815e-07
I2409 0 n2410 3.361e-02A M=1.024e-06
I2410 0 n2411 3.361e-02A M=4.443e-07
I2411 0 n2412 3.361e-02A M=7.058e-07
I2412 0 n2413 3.361e-02A M=1.171e-06
I2413 0 n2414 3.361e-02A M=1.187e-06
I2414 0 n2415 3.361e-02A M=1.574e-07
I2415 0 n2416 3.361e-02A M=1.912e-06
I2416 0 n2417 3.361e-02A M=6.171e-07
I2417 0 n2418 3.361e-02A M=7.303e-07
I2418 0 n2419 3.361e-02A M=1.452e-06
I2419 0 n2420 3.361e-02A M=1.282e-06
I2420 0 n2421 3.361e-02A M=1.507e-06
I2421 0 n2422 3.361e-02A M=1.140e-06
I2422 0 n2423 3.361e-02A M=5.262e-07
I2423 0 n2424 3.361e-02A M=1.772e-06
I2424 0 n2425 3.361e-02A M=7.328e-07
I2425 0 n2426 3.361e-02A M=2.723e-07
I2426 0 n2427 3.361e-02A M=5.149e-07
I2427 0 n2428 3.361e-02A M=1.037e-06
I2428 0 n2429 3.361e-02A M=4.073e-07
I2429 0 n2430 3.361e-02A M=6.099e-07
I2430 0 n2431 3.361e-02A M=7.608e-07
I2431 0 n2432 3.361e-02A M=7.523e-07
I2432 0 n2433 3.361e-02A M=2.105e-06
I2433 0 n2434 3.361e-02A M=1.661e-06
I2434 0 n2435 3.361e-02A M=6.407e-07
I2435 0 n2436 3.361e-02A M=1.241e-06
I2436 0 n2437 3.361e-02A M=1.334e-06
I2437 0 n2438 3.361e-02A M=1.908e-06
I2438 0 n2439 3.361e-02A M=9.100e-07
I2439 0 n1 3.361e-02A M=8.140e-07
I2440 0 n2441 3.361e-02A M=7.192e-07
I2441 0 n2442 3.361e-02A M=6.181e-07
I2442 0 n2443 3.361e-02A M=9.606e-07
I2443 0 n2444 3.361e-02A M=8.612e-07
I2444 0 n2445 3.361e-02A M=5.962e-07
I2445 0 n2446 3.361e-02A M=5.992e-07
I2446 0 n1 3.361e-02A M=6.661e-07
I2447 0 n2448 3.361e-02A M=8.987e-07
I2448 0 n2449 3.361e-02A M=7.015e-07
I2449 0 n2450 3.361e-02A M=8.760e-07
I2450 0 n2451 3.361e-02A M=1.185e-06
I2451 0 n2452 3.361e-02A M=3.762e-07
I2452 0 n2453 3.361e-02A M=8.338e-07
I2453 0 n2454 3.361e-02A M=6.166e-07
I2454 0 n2455 3.361e-02A M=1.850e-06
I2455 0 n2456 3.361e-02A M=3.721e-07
I2456 0 n2457 3.361e-02A M=7.840e-07
I2457 0 n2458 3.361e-02A M=6.574e-07
I2458 0 n2459 3.361e-02A M=1.590e-06
I2459 0 n2460 3.361e-02A M=6.168e-07
I2460 0 n2461 3.361e-02A M=2.128e-06
I2461 0 n2462 3.361e-02A M=2.375e-06
I2462 0 n2463 3.361e-02A M=1.184e-06
I2463 0 n2464 3.361e-02A M=8.589e-07
I2464 0 n2465 3.361e-02A M=8.669e-07
I2465 0 n2466 3.361e-02A M=1.448e-06
I2466 0 n2467 3.361e-02A M=1.253e-06
I2467 0 n2468 3.361e-02A M=1.489e-06
I2468 0 n2469 3.361e-02A M=8.677e-07
I2469 0 n2470 3.361e-02A M=1.065e-06
I2470 0 n2471 3.361e-02A M=8.004e-07
I2471 0 n2472 3.361e-02A M=1.796e-06
I2472 0 n2473 3.361e-02A M=7.839e-07
I2473 0 n2474 3.361e-02A M=1.183e-06
I2474 0 n2475 3.361e-02A M=1.400e-06
I2475 0 n2476 3.361e-02A M=1.799e-06
I2476 0 n2477 3.361e-02A M=1.019e-06
I2477 0 n2478 3.361e-02A M=6.991e-07
I2478 0 n2479 3.361e-02A M=3.040e-07
I2479 0 n2480 3.361e-02A M=2.283e-07
I2480 0 n2481 3.361e-02A M=6.262e-07
I2481 0 n2482 3.361e-02A M=7.751e-07
I2482 0 n2483 3.361e-02A M=1.470e-06
I2483 0 n2484 3.361e-02A M=9.797e-07
I2484 0 n2485 3.361e-02A M=1.165e-06
I2485 0 n2486 3.361e-02A M=1.458e-06
I2486 0 n2487 3.361e-02A M=7.819e-07
I2487 0 n2488 3.361e-02A M=2.581e-06
I2488 0 n2489 3.361e-02A M=1.565e-06
I2489 0 n2490 3.361e-02A M=1.010e-06
I2490 0 n2491 3.361e-02A M=1.366e-06
I2491 0 n2492 3.361e-02A M=1.218e-06
I2492 0 n2493 3.361e-02A M=2.969e-07
I2493 0 n2494 3.361e-02A M=1.901e-06
I2494 0 n2495 3.361e-02A M=6.021e-07
I2495 0 n2496 3.361e-02A M=2.527e-06
I2496 0 n2497 3.361e-02A M=3.817e-07
I2497 0 n2498 3.361e-02A M=1.268e-06
I2498 0 n2499 3.361e-02A M=1.553e-06
I2499 0 n2500 3.361e-02A M=1.166e-06
I2500 0 n2501 3.361e-02A M=1.164e-06
I2501 0 n2502 3.361e-02A M=3.794e-07
I2502 0 n2503 3.361e-02A M=2.255e-07
I2503 0 n2504 3.361e-02A M=1.341e-06
I2504 0 n2505 3.361e-02A M=2.153e-06
I2505 0 n2506 3.361e-02A M=8.914e-07
I2506 0 n2507 3.361e-02A M=5.773e-07
I2507 0 n2508 3.361e-02A M=8.529e-07
I2508 0 n2509 3.361e-02A M=2.473e-06
I2509 0 n2510 3.361e-02A M=5.346e-07
I2510 0 n2511 3.361e-02A M=7.277e-07
I2511 0 n2512 3.361e-02A M=6.381e-07
I2512 0 n2513 3.361e-02A M=2.244e-06
I2513 0 n2514 3.361e-02A M=8.029e-07
I2514 0 n2515 3.361e-02A M=1.078e-06
I2515 0 n2516 3.361e-02A M=9.418e-07
I2516 0 n2517 3.361e-02A M=9.086e-07
I2517 0 n2518 3.361e-02A M=2.688e-07
I2518 0 n2519 3.361e-02A M=7.714e-07
I2519 0 n2520 3.361e-02A M=3.710e-07
I2520 0 n2521 3.361e-02A M=8.298e-07
I2521 0 n2522 3.361e-02A M=7.694e-07
I2522 0 n2523 3.361e-02A M=5.372e-07
I2523 0 n2524 3.361e-02A M=1.260e-06
I2524 0 n2525 3.361e-02A M=1.470e-07
I2525 0 n2526 3.361e-02A M=1.162e-06
I2526 0 n2527 3.361e-02A M=3.333e-07
I2527 0 n2528 3.361e-02A M=3.868e-07
I2528 0 n2529 3.361e-02A M=1.221e-06
I2529 0 n2530 3.361e-02A M=5.357e-07
I2530 0 n2531 3.361e-02A M=3.518e-07
I2531 0 n2532 3.361e-02A M=6.841e-07
I2532 0 n2533 3.361e-02A M=9.216e-07
I2533 0 n2534 3.361e-02A M=1.469e-06
I2534 0 n2535 3.361e-02A M=5.862e-07
I2535 0 n2536 3.361e-02A M=8.243e-07
I2536 0 n2537 3.361e-02A M=1.433e-06
I2537 0 n2538 3.361e-02A M=5.693e-07
I2538 0 n2539 3.361e-02A M=8.337e-07
I2539 0 n2540 3.361e-02A M=1.421e-06
I2540 0 n2541 3.361e-02A M=4.370e-07
I2541 0 n2542 3.361e-02A M=5.394e-07
I2542 0 n2543 3.361e-02A M=3.093e-07
I2543 0 n2544 3.361e-02A M=2.746e-07
I2544 0 n2545 3.361e-02A M=2.135e-06
I2545 0 n2546 3.361e-02A M=6.211e-07
I2546 0 n2547 3.361e-02A M=4.799e-07
I2547 0 n2548 3.361e-02A M=6.559e-07
I2548 0 n2549 3.361e-02A M=3.161e-07
I2549 0 n2550 3.361e-02A M=1.393e-06
I2550 0 n2551 3.361e-02A M=1.157e-06
I2551 0 n2552 3.361e-02A M=8.334e-07
I2552 0 n2553 3.361e-02A M=6.920e-07
I2553 0 n2554 3.361e-02A M=5.610e-07
I2554 0 n2555 3.361e-02A M=6.037e-07
I2555 0 n2556 3.361e-02A M=1.416e-06
I2556 0 n2557 3.361e-02A M=1.097e-06
I2557 0 n2558 3.361e-02A M=5.185e-07
I2558 0 n2559 3.361e-02A M=5.197e-07
I2559 0 n2560 3.361e-02A M=5.407e-07
I2560 0 n2561 3.361e-02A M=6.848e-07
I2561 0 n2562 3.361e-02A M=1.812e-06
I2562 0 n2563 3.361e-02A M=1.781e-06
I2563 0 n2564 3.361e-02A M=1.069e-06
I2564 0 n2565 3.361e-02A M=1.635e-06
I2565 0 n2566 3.361e-02A M=1.360e-06
I2566 0 n2567 3.361e-02A M=5.008e-07
I2567 0 n2568 3.361e-02A M=1.106e-06
I2568 0 n2569 3.361e-02A M=1.779e-06
I2569 0 n2570 3.361e-02A M=6.979e-07
I2570 0 n2571 3.361e-02A M=9.677e-07
I2571 0 n1 3.361e-02A M=9.258e-07
I2572 0 n2573 3.361e-02A M=5.622e-07
I2573 0 n2574 3.361e-02A M=2.028e-07
I2574 0 n2575 3.361e-02A M=1.268e-06
I2575 0 n2576 3.361e-02A M=9.871e-07
I2576 0 n2577 3.361e-02A M=1.046e-06
I2577 0 n2578 3.361e-02A M=1.007e-06
I2578 0 n2579 3.361e-02A M=6.481e-07
I2579 0 n2580 3.361e-02A M=7.577e-07
I2580 0 n2581 3.361e-02A M=3.136e-07
I2581 0 n2582 3.361e-02A M=9.670e-07
I2582 0 n2583 3.361e-02A M=5.466e-07
I2583 0 n2584 3.361e-02A M=1.964e-06
I2584 0 n2585 3.361e-02A M=3.953e-07
I2585 0 n2586 3.361e-02A M=1.016e-06
I2586 0 n2587 3.361e-02A M=6.430e-07
I2587 0 n2588 3.361e-02A M=7.140e-07
I2588 0 n2589 3.361e-02A M=9.229e-07
I2589 0 n2590 3.361e-02A M=5.621e-07
I2590 0 n2591 3.361e-02A M=5.487e-07
I2591 0 n2592 3.361e-02A M=1.060e-06
I2592 0 n2593 3.361e-02A M=1.065e-06
I2593 0 n2594 3.361e-02A M=6.890e-07
I2594 0 n2595 3.361e-02A M=8.534e-07
I2595 0 n2596 3.361e-02A M=1.902e-06
I2596 0 n2597 3.361e-02A M=9.030e-07
I2597 0 n2598 3.361e-02A M=4.148e-07
I2598 0 n2599 3.361e-02A M=4.005e-07
I2599 0 n2600 3.361e-02A M=1.358e-06
I2600 0 n2601 3.361e-02A M=2.236e-07
I2601 0 n2602 3.361e-02A M=9.544e-07
I2602 0 n2603 3.361e-02A M=2.660e-07
I2603 0 n2604 3.361e-02A M=7.735e-07
I2604 0 n2605 3.361e-02A M=1.077e-06
I2605 0 n2606 3.361e-02A M=7.866e-07
I2606 0 n2607 3.361e-02A M=8.451e-07
I2607 0 n2608 3.361e-02A M=1.112e-07
I2608 0 n2609 3.361e-02A M=1.086e-06
I2609 0 n2610 3.361e-02A M=2.092e-07
I2610 0 n1 3.361e-02A M=1.060e-06
I2611 0 n2612 3.361e-02A M=1.952e-07
I2612 0 n2613 3.361e-02A M=1.601e-06
I2613 0 n2614 3.361e-02A M=6.157e-07
I2614 0 n2615 3.361e-02A M=9.849e-07
I2615 0 n2616 3.361e-02A M=5.728e-07
I2616 0 n2617 3.361e-02A M=9.350e-07
I2617 0 n2618 3.361e-02A M=2.005e-06
I2618 0 n2619 3.361e-02A M=6.181e-07
I2619 0 n2620 3.361e-02A M=1.636e-06
I2620 0 n2621 3.361e-02A M=6.408e-07
I2621 0 n2622 3.361e-02A M=4.041e-07
I2622 0 n2623 3.361e-02A M=6.394e-07
I2623 0 n2624 3.361e-02A M=6.523e-07
I2624 0 n2625 3.361e-02A M=1.576e-06
I2625 0 n2626 3.361e-02A M=7.881e-07
I2626 0 n2627 3.361e-02A M=1.539e-06
I2627 0 n2628 3.361e-02A M=4.961e-07
I2628 0 n2629 3.361e-02A M=5.368e-07
I2629 0 n2630 3.361e-02A M=6.427e-07
I2630 0 n2631 3.361e-02A M=1.276e-06
I2631 0 n2632 3.361e-02A M=6.877e-07
I2632 0 n2633 3.361e-02A M=5.634e-07
I2633 0 n2634 3.361e-02A M=1.264e-06
I2634 0 n2635 3.361e-02A M=1.887e-06
I2635 0 n2636 3.361e-02A M=2.043e-06
I2636 0 n2637 3.361e-02A M=1.443e-06
I2637 0 n2638 3.361e-02A M=4.173e-07
I2638 0 n2639 3.361e-02A M=6.590e-07
I2639 0 n2640 3.361e-02A M=2.518e-06
I2640 0 n2641 3.361e-02A M=8.809e-07
I2641 0 n2642 3.361e-02A M=1.543e-06
I2642 0 n2643 3.361e-02A M=5.506e-07
I2643 0 n2644 3.361e-02A M=1.446e-06
I2644 0 n2645 3.361e-02A M=1.418e-06
I2645 0 n2646 3.361e-02A M=1.815e-07
I2646 0 n2647 3.361e-02A M=4.567e-07
I2647 0 n2648 3.361e-02A M=9.418e-07
I2648 0 n2649 3.361e-02A M=7.747e-07
I2649 0 n2650 3.361e-02A M=3.421e-07
I2650 0 n2651 3.361e-02A M=9.129e-07
I2651 0 n2652 3.361e-02A M=2.070e-06
I2652 0 n2653 3.361e-02A M=1.154e-06
I2653 0 n2654 3.361e-02A M=3.262e-07
I2654 0 n2655 3.361e-02A M=1.212e-06
I2655 0 n2656 3.361e-02A M=7.641e-07
I2656 0 n2657 3.361e-02A M=6.564e-07
I2657 0 n2658 3.361e-02A M=2.673e-06
I2658 0 n2659 3.361e-02A M=1.233e-06
I2659 0 n2660 3.361e-02A M=7.925e-07
I2660 0 n2661 3.361e-02A M=1.174e-06
I2661 0 n2662 3.361e-02A M=2.343e-06
I2662 0 n2663 3.361e-02A M=3.245e-07
I2663 0 n2664 3.361e-02A M=4.950e-07
I2664 0 n2665 3.361e-02A M=8.129e-07
I2665 0 n2666 3.361e-02A M=1.073e-06
I2666 0 n2667 3.361e-02A M=7.750e-07
I2667 0 n2668 3.361e-02A M=2.695e-06
I2668 0 n2669 3.361e-02A M=1.210e-06
I2669 0 n2670 3.361e-02A M=3.770e-07
I2670 0 n2671 3.361e-02A M=1.155e-06
I2671 0 n2672 3.361e-02A M=6.021e-07
I2672 0 n2673 3.361e-02A M=1.269e-06
I2673 0 n2674 3.361e-02A M=1.171e-06
I2674 0 n2675 3.361e-02A M=7.859e-07
I2675 0 n2676 3.361e-02A M=3.980e-07
I2676 0 n2677 3.361e-02A M=7.305e-07
I2677 0 n2678 3.361e-02A M=7.919e-07
I2678 0 n2679 3.361e-02A M=1.797e-06
I2679 0 n2680 3.361e-02A M=9.168e-07
I2680 0 n2681 3.361e-02A M=9.091e-07
I2681 0 n2682 3.361e-02A M=9.946e-07
I2682 0 n2683 3.361e-02A M=6.996e-07
I2683 0 n2684 3.361e-02A M=1.247e-06
I2684 0 n2685 3.361e-02A M=6.130e-07
I2685 0 n2686 3.361e-02A M=7.127e-07
I2686 0 n2687 3.361e-02A M=1.634e-06
I2687 0 n2688 3.361e-02A M=1.062e-06
I2688 0 n2689 3.361e-02A M=1.684e-06
I2689 0 n2690 3.361e-02A M=6.999e-07
I2690 0 n2691 3.361e-02A M=9.522e-07
I2691 0 n2692 3.361e-02A M=1.317e-06
I2692 0 n2693 3.361e-02A M=9.925e-07
I2693 0 n2694 3.361e-02A M=7.051e-07
I2694 0 n2695 3.361e-02A M=4.137e-07
I2695 0 n2696 3.361e-02A M=2.306e-06
I2696 0 n2697 3.361e-02A M=9.962e-07
I2697 0 n2698 3.361e-02A M=7.819e-07
I2698 0 n2699 3.361e-02A M=4.075e-07
I2699 0 n2700 3.361e-02A M=9.080e-07
I2700 0 n2701 3.361e-02A M=7.656e-07
I2701 0 n2702 3.361e-02A M=1.282e-06
I2702 0 n2703 3.361e-02A M=8.332e-07
I2703 0 n2704 3.361e-02A M=8.778e-07
I2704 0 n2705 3.361e-02A M=4.092e-07
I2705 0 n2706 3.361e-02A M=1.038e-06
I2706 0 n2707 3.361e-02A M=6.395e-07
I2707 0 n2708 3.361e-02A M=1.412e-06
I2708 0 n2709 3.361e-02A M=1.192e-06
I2709 0 n2710 3.361e-02A M=1.638e-06
I2710 0 n2711 3.361e-02A M=5.842e-07
I2711 0 n2712 3.361e-02A M=1.452e-06
I2712 0 n2713 3.361e-02A M=3.241e-07
I2713 0 n2714 3.361e-02A M=1.218e-06
I2714 0 n2715 3.361e-02A M=6.326e-07
I2715 0 n2716 3.361e-02A M=1.707e-06
I2716 0 n2717 3.361e-02A M=2.573e-06
I2717 0 n2718 3.361e-02A M=8.477e-07
I2718 0 n2719 3.361e-02A M=1.034e-06
I2719 0 n2720 3.361e-02A M=1.845e-06
I2720 0 n2721 3.361e-02A M=1.609e-06
I2721 0 n2722 3.361e-02A M=3.801e-07
I2722 0 n2723 3.361e-02A M=1.482e-07
I2723 0 n2724 3.361e-02A M=6.670e-07
I2724 0 n2725 3.361e-02A M=2.078e-06
I2725 0 n2726 3.361e-02A M=7.247e-07
I2726 0 n2727 3.361e-02A M=7.174e-07
I2727 0 n2728 3.361e-02A M=4.640e-07
I2728 0 n2729 3.361e-02A M=6.898e-07
I2729 0 n2730 3.361e-02A M=1.095e-06
I2730 0 n2731 3.361e-02A M=1.210e-06
I2731 0 n2732 3.361e-02A M=1.050e-06
I2732 0 n2733 3.361e-02A M=8.959e-07
I2733 0 n2734 3.361e-02A M=1.628e-06
I2734 0 n2735 3.361e-02A M=1.478e-06
I2735 0 n2736 3.361e-02A M=1.184e-06
I2736 0 n2737 3.361e-02A M=1.030e-06
I2737 0 n2738 3.361e-02A M=1.347e-06
I2738 0 n2739 3.361e-02A M=1.891e-06
I2739 0 n2740 3.361e-02A M=8.545e-07
I2740 0 n2741 3.361e-02A M=1.286e-06
I2741 0 n2742 3.361e-02A M=1.030e-07
I2742 0 n2743 3.361e-02A M=1.137e-06
I2743 0 n2744 3.361e-02A M=1.062e-06
I2744 0 n2745 3.361e-02A M=9.689e-07
I2745 0 n2746 3.361e-02A M=8.505e-07
I2746 0 n2747 3.361e-02A M=1.003e-06
I2747 0 n1 3.361e-02A M=1.052e-06
I2748 0 n2749 3.361e-02A M=1.481e-06
I2749 0 n2750 3.361e-02A M=1.538e-06
I2750 0 n2751 3.361e-02A M=7.363e-07
I2751 0 n2752 3.361e-02A M=1.575e-06
I2752 0 n2753 3.361e-02A M=1.107e-06
I2753 0 n2754 3.361e-02A M=1.266e-06
I2754 0 n2755 3.361e-02A M=1.026e-06
I2755 0 n2756 3.361e-02A M=1.430e-06
I2756 0 n2757 3.361e-02A M=1.048e-06
I2757 0 n2758 3.361e-02A M=1.748e-06
I2758 0 n2759 3.361e-02A M=1.931e-06
I2759 0 n2760 3.361e-02A M=8.461e-07
I2760 0 n2761 3.361e-02A M=7.410e-07
I2761 0 n2762 3.361e-02A M=2.027e-06
I2762 0 n2763 3.361e-02A M=1.547e-06
I2763 0 n2764 3.361e-02A M=1.144e-06
I2764 0 n2765 3.361e-02A M=3.119e-07
I2765 0 n2766 3.361e-02A M=8.726e-07
I2766 0 n2767 3.361e-02A M=1.141e-06
I2767 0 n2768 3.361e-02A M=1.207e-06
I2768 0 n2769 3.361e-02A M=1.103e-06
I2769 0 n2770 3.361e-02A M=1.084e-06
I2770 0 n2771 3.361e-02A M=1.061e-06
I2771 0 n2772 3.361e-02A M=1.300e-06
I2772 0 n2773 3.361e-02A M=8.614e-08
I2773 0 n2774 3.361e-02A M=1.022e-06
I2774 0 n2775 3.361e-02A M=2.185e-07
I2775 0 n2776 3.361e-02A M=1.037e-06
I2776 0 n2777 3.361e-02A M=3.077e-07
I2777 0 n2778 3.361e-02A M=9.192e-07
I2778 0 n2779 3.361e-02A M=1.286e-06
I2779 0 n2780 3.361e-02A M=7.662e-07
I2780 0 n2781 3.361e-02A M=1.831e-06
I2781 0 n2782 3.361e-02A M=1.630e-06
I2782 0 n2783 3.361e-02A M=5.734e-07
I2783 0 n2784 3.361e-02A M=1.090e-06
I2784 0 n2785 3.361e-02A M=1.100e-06
I2785 0 n2786 3.361e-02A M=1.105e-06
I2786 0 n2787 3.361e-02A M=7.726e-07
I2787 0 n2788 3.361e-02A M=1.031e-06
I2788 0 n2789 3.361e-02A M=7.063e-07
I2789 0 n2790 3.361e-02A M=1.642e-06
I2790 0 n2791 3.361e-02A M=1.397e-06
I2791 0 n2792 3.361e-02A M=6.917e-07
I2792 0 n2793 3.361e-02A M=4.373e-07
I2793 0 n2794 3.361e-02A M=5.513e-07
I2794 0 n2795 3.361e-02A M=1.522e-06
I2795 0 n2796 3.361e-02A M=1.663e-06
I2796 0 n2797 3.361e-02A M=1.144e-06
I2797 0 n2798 3.361e-02A M=4.594e-07
I2798 0 n2799 3.361e-02A M=8.332e-07
I2799 0 n2800 3.361e-02A M=4.595e-07
I2800 0 n2801 3.361e-02A M=4.474e-07
I2801 0 n2802 3.361e-02A M=9.438e-07
I2802 0 n2803 3.361e-02A M=8.881e-07
I2803 0 n2804 3.361e-02A M=4.215e-07
I2804 0 n2805 3.361e-02A M=2.336e-07
I2805 0 n2806 3.361e-02A M=1.539e-06
I2806 0 n2807 3.361e-02A M=2.331e-07
I2807 0 n2808 3.361e-02A M=1.814e-06
I2808 0 n2809 3.361e-02A M=8.649e-07
I2809 0 n2810 3.361e-02A M=1.279e-06
I2810 0 n2811 3.361e-02A M=3.409e-07
I2811 0 n2812 3.361e-02A M=1.205e-06
I2812 0 n2813 3.361e-02A M=1.839e-06
I2813 0 n2814 3.361e-02A M=5.285e-07
I2814 0 n2815 3.361e-02A M=5.084e-07
I2815 0 n2816 3.361e-02A M=1.545e-06
I2816 0 n2817 3.361e-02A M=1.845e-06
I2817 0 n2818 3.361e-02A M=4.437e-07
I2818 0 n2819 3.361e-02A M=1.622e-06
I2819 0 n2820 3.361e-02A M=6.849e-07
I2820 0 n2821 3.361e-02A M=4.758e-07
I2821 0 n2822 3.361e-02A M=1.257e-06
I2822 0 n2823 3.361e-02A M=7.162e-07
I2823 0 n2824 3.361e-02A M=8.013e-07
I2824 0 n2825 3.361e-02A M=2.403e-06
I2825 0 n2826 3.361e-02A M=6.093e-07
I2826 0 n2827 3.361e-02A M=6.514e-07
I2827 0 n2828 3.361e-02A M=9.764e-07
I2828 0 n2829 3.361e-02A M=1.580e-06
I2829 0 n2830 3.361e-02A M=7.741e-07
I2830 0 n2831 3.361e-02A M=7.442e-07
I2831 0 n2832 3.361e-02A M=2.872e-06
I2832 0 n2833 3.361e-02A M=1.100e-06
I2833 0 n2834 3.361e-02A M=1.373e-06
I2834 0 n2835 3.361e-02A M=1.425e-06
I2835 0 n2836 3.361e-02A M=4.089e-07
I2836 0 n2837 3.361e-02A M=1.432e-06
I2837 0 n2838 3.361e-02A M=9.954e-07
I2838 0 n2839 3.361e-02A M=1.586e-06
I2839 0 n2840 3.361e-02A M=1.250e-06
I2840 0 n2841 3.361e-02A M=9.772e-07
I2841 0 n2842 3.361e-02A M=5.573e-07
I2842 0 n2843 3.361e-02A M=1.189e-06
I2843 0 n2844 3.361e-02A M=1.699e-06
I2844 0 n2845 3.361e-02A M=1.263e-06
I2845 0 n2846 3.361e-02A M=5.649e-07
I2846 0 n2847 3.361e-02A M=1.424e-06
I2847 0 n2848 3.361e-02A M=1.232e-06
I2848 0 n2849 3.361e-02A M=8.870e-07
I2849 0 n2850 3.361e-02A M=1.305e-06
I2850 0 n1 3.361e-02A M=1.992e-06
I2851 0 n2852 3.361e-02A M=8.638e-07
I2852 0 n2853 3.361e-02A M=6.221e-07
I2853 0 n2854 3.361e-02A M=1.188e-06
I2854 0 n2855 3.361e-02A M=1.505e-06
I2855 0 n2856 3.361e-02A M=1.845e-06
I2856 0 n2857 3.361e-02A M=2.093e-06
I2857 0 n2858 3.361e-02A M=1.880e-06
I2858 0 n2859 3.361e-02A M=1.558e-06
I2859 0 n2860 3.361e-02A M=6.558e-07
I2860 0 n2861 3.361e-02A M=6.821e-07
I2861 0 n2862 3.361e-02A M=7.736e-07
I2862 0 n2863 3.361e-02A M=1.094e-06
I2863 0 n2864 3.361e-02A M=8.240e-07
I2864 0 n2865 3.361e-02A M=1.115e-06
I2865 0 n2866 3.361e-02A M=6.941e-07
I2866 0 n2867 3.361e-02A M=9.778e-07
I2867 0 n2868 3.361e-02A M=1.121e-06
I2868 0 n2869 3.361e-02A M=4.851e-07
I2869 0 n1 3.361e-02A M=3.150e-07
I2870 0 n2871 3.361e-02A M=1.657e-06
I2871 0 n2872 3.361e-02A M=1.210e-06
I2872 0 n2873 3.361e-02A M=6.970e-07
I2873 0 n2874 3.361e-02A M=2.248e-06
I2874 0 n2875 3.361e-02A M=6.349e-07
I2875 0 n2876 3.361e-02A M=8.074e-07
I2876 0 n2877 3.361e-02A M=6.018e-07
I2877 0 n2878 3.361e-02A M=1.024e-06
I2878 0 n2879 3.361e-02A M=6.078e-07
I2879 0 n2880 3.361e-02A M=6.619e-07
I2880 0 n2881 3.361e-02A M=8.128e-07
I2881 0 n2882 3.361e-02A M=6.642e-07
I2882 0 n2883 3.361e-02A M=1.042e-06
I2883 0 n2884 3.361e-02A M=7.542e-07
I2884 0 n2885 3.361e-02A M=1.413e-06
I2885 0 n2886 3.361e-02A M=6.335e-07
I2886 0 n2887 3.361e-02A M=1.152e-06
I2887 0 n2888 3.361e-02A M=3.106e-07
I2888 0 n2889 3.361e-02A M=1.306e-06
I2889 0 n2890 3.361e-02A M=1.311e-06
I2890 0 n2891 3.361e-02A M=7.706e-07
I2891 0 n2892 3.361e-02A M=8.970e-07
I2892 0 n2893 3.361e-02A M=1.658e-06
I2893 0 n2894 3.361e-02A M=7.981e-07
I2894 0 n2895 3.361e-02A M=9.583e-07
I2895 0 n2896 3.361e-02A M=5.051e-07
I2896 0 n2897 3.361e-02A M=9.950e-07
I2897 0 n2898 3.361e-02A M=1.876e-06
I2898 0 n2899 3.361e-02A M=1.258e-06
I2899 0 n2900 3.361e-02A M=1.429e-06
I2900 0 n1 3.361e-02A M=8.099e-07
I2901 0 n2902 3.361e-02A M=1.261e-06
I2902 0 n2903 3.361e-02A M=7.333e-07
I2903 0 n2904 3.361e-02A M=5.524e-07
I2904 0 n2905 3.361e-02A M=1.059e-06
I2905 0 n2906 3.361e-02A M=4.484e-07
I2906 0 n2907 3.361e-02A M=1.928e-06
I2907 0 n2908 3.361e-02A M=8.942e-07
I2908 0 n2909 3.361e-02A M=7.699e-07
I2909 0 n2910 3.361e-02A M=2.160e-06
I2910 0 n2911 3.361e-02A M=1.768e-06
I2911 0 n2912 3.361e-02A M=7.927e-07
I2912 0 n2913 3.361e-02A M=1.526e-06
I2913 0 n2914 3.361e-02A M=1.288e-06
I2914 0 n2915 3.361e-02A M=1.345e-07
I2915 0 n2916 3.361e-02A M=1.103e-06
I2916 0 n2917 3.361e-02A M=1.096e-06
I2917 0 n2918 3.361e-02A M=8.873e-07
I2918 0 n2919 3.361e-02A M=1.102e-06
I2919 0 n2920 3.361e-02A M=8.306e-07
I2920 0 n2921 3.361e-02A M=8.841e-07
I2921 0 n2922 3.361e-02A M=1.040e-06
I2922 0 n2923 3.361e-02A M=1.748e-06
I2923 0 n2924 3.361e-02A M=4.302e-07
I2924 0 n2925 3.361e-02A M=6.497e-07
I2925 0 n2926 3.361e-02A M=2.193e-06
I2926 0 n2927 3.361e-02A M=1.190e-06
I2927 0 n2928 3.361e-02A M=1.074e-06
I2928 0 n2929 3.361e-02A M=1.288e-06
I2929 0 n2930 3.361e-02A M=6.538e-07
I2930 0 n2931 3.361e-02A M=3.487e-07
I2931 0 n2932 3.361e-02A M=7.912e-07
I2932 0 n2933 3.361e-02A M=6.743e-07
I2933 0 n2934 3.361e-02A M=1.114e-06
I2934 0 n2935 3.361e-02A M=1.387e-06
I2935 0 n2936 3.361e-02A M=6.331e-07
I2936 0 n2937 3.361e-02A M=1.018e-06
I2937 0 n2938 3.361e-02A M=1.276e-06
I2938 0 n2939 3.361e-02A M=1.048e-06
I2939 0 n2940 3.361e-02A M=7.280e-07
I2940 0 n2941 3.361e-02A M=3.393e-07
I2941 0 n2942 3.361e-02A M=3.274e-07
I2942 0 n2943 3.361e-02A M=1.059e-06
I2943 0 n1 3.361e-02A M=4.512e-07
I2944 0 n2945 3.361e-02A M=1.567e-06
I2945 0 n2946 3.361e-02A M=1.507e-06
I2946 0 n2947 3.361e-02A M=1.287e-06
I2947 0 n2948 3.361e-02A M=2.124e-06
I2948 0 n2949 3.361e-02A M=8.761e-07
I2949 0 n2950 3.361e-02A M=2.327e-06
I2950 0 n2951 3.361e-02A M=9.287e-07
I2951 0 n2952 3.361e-02A M=1.378e-06
I2952 0 n2953 3.361e-02A M=6.255e-07
I2953 0 n2954 3.361e-02A M=7.248e-07
I2954 0 n2955 3.361e-02A M=8.598e-07
I2955 0 n2956 3.361e-02A M=4.687e-07
I2956 0 n2957 3.361e-02A M=3.026e-07
I2957 0 n2958 3.361e-02A M=8.844e-07
I2958 0 n2959 3.361e-02A M=1.487e-06
I2959 0 n2960 3.361e-02A M=5.238e-07
I2960 0 n2961 3.361e-02A M=1.042e-06
I2961 0 n2962 3.361e-02A M=1.072e-07
I2962 0 n2963 3.361e-02A M=1.044e-06
I2963 0 n2964 3.361e-02A M=1.201e-06
I2964 0 n2965 3.361e-02A M=4.328e-07
I2965 0 n2966 3.361e-02A M=1.173e-06
I2966 0 n2967 3.361e-02A M=1.057e-06
I2967 0 n2968 3.361e-02A M=1.363e-06
I2968 0 n2969 3.361e-02A M=1.354e-06
I2969 0 n2970 3.361e-02A M=4.780e-07
I2970 0 n2971 3.361e-02A M=3.578e-07
I2971 0 n2972 3.361e-02A M=7.403e-07
I2972 0 n2973 3.361e-02A M=7.584e-07
I2973 0 n2974 3.361e-02A M=7.201e-07
I2974 0 n2975 3.361e-02A M=2.446e-07
I2975 0 n2976 3.361e-02A M=1.103e-06
I2976 0 n2977 3.361e-02A M=1.933e-07
I2977 0 n2978 3.361e-02A M=1.871e-06
I2978 0 n2979 3.361e-02A M=8.287e-07
I2979 0 n2980 3.361e-02A M=6.050e-07
I2980 0 n2981 3.361e-02A M=6.873e-07
I2981 0 n2982 3.361e-02A M=6.928e-07
I2982 0 n2983 3.361e-02A M=9.135e-07
I2983 0 n2984 3.361e-02A M=5.239e-07
I2984 0 n2985 3.361e-02A M=8.435e-07
I2985 0 n2986 3.361e-02A M=2.620e-07
I2986 0 n2987 3.361e-02A M=6.226e-07
I2987 0 n2988 3.361e-02A M=5.507e-07
I2988 0 n2989 3.361e-02A M=7.369e-07
I2989 0 n2990 3.361e-02A M=1.231e-06
I2990 0 n2991 3.361e-02A M=2.365e-06
I2991 0 n2992 3.361e-02A M=3.884e-07
I2992 0 n2993 3.361e-02A M=1.951e-07
I2993 0 n2994 3.361e-02A M=5.448e-07
I2994 0 n2995 3.361e-02A M=8.526e-07
I2995 0 n2996 3.361e-02A M=4.551e-07
I2996 0 n2997 3.361e-02A M=1.071e-06
I2997 0 n2998 3.361e-02A M=9.658e-07
I2998 0 n2999 3.361e-02A M=5.638e-07
I2999 0 n3000 3.361e-02A M=4.506e-07
I3000 0 n3001 3.361e-02A M=1.210e-06
I3001 0 n3002 3.361e-02A M=6.687e-07
I3002 0 n3003 3.361e-02A M=6.748e-07
I3003 0 n3004 3.361e-02A M=1.244e-06
I3004 0 n3005 3.361e-02A M=4.963e-07
I3005 0 n3006 3.361e-02A M=1.479e-06
I3006 0 n3007 3.361e-02A M=1.400e-06
I3007 0 n3008 3.361e-02A M=5.122e-07
I3008 0 n3009 3.361e-02A M=7.978e-07
I3009 0 n3010 3.361e-02A M=9.648e-07
I3010 0 n3011 3.361e-02A M=1.890e-07
I3011 0 n3012 3.361e-02A M=1.283e-06
I3012 0 n3013 3.361e-02A M=3.545e-07
I3013 0 n3014 3.361e-02A M=1.704e-06
I3014 0 n3015 3.361e-02A M=6.319e-07
I3015 0 n3016 3.361e-02A M=6.229e-07
I3016 0 n3017 3.361e-02A M=9.590e-07
I3017 0 n3018 3.361e-02A M=6.316e-07
I3018 0 n3019 3.361e-02A M=4.826e-07
I3019 0 n3020 3.361e-02A M=1.352e-06
I3020 0 n3021 3.361e-02A M=5.110e-07
I3021 0 n3022 3.361e-02A M=7.575e-07
I3022 0 n3023 3.361e-02A M=1.141e-06
I3023 0 n3024 3.361e-02A M=6.584e-07
I3024 0 n3025 3.361e-02A M=1.370e-06
I3025 0 n3026 3.361e-02A M=1.519e-06
I3026 0 n3027 3.361e-02A M=6.546e-07
I3027 0 n3028 3.361e-02A M=8.026e-07
I3028 0 n3029 3.361e-02A M=7.483e-07
I3029 0 n3030 3.361e-02A M=1.624e-06
I3030 0 n3031 3.361e-02A M=1.389e-06
I3031 0 n3032 3.361e-02A M=1.423e-06
I3032 0 n3033 3.361e-02A M=1.145e-06
I3033 0 n3034 3.361e-02A M=1.934e-06
I3034 0 n3035 3.361e-02A M=9.968e-07
I3035 0 n3036 3.361e-02A M=5.329e-07
I3036 0 n3037 3.361e-02A M=2.795e-07
I3037 0 n3038 3.361e-02A M=1.496e-06
I3038 0 n3039 3.361e-02A M=2.314e-06
I3039 0 n1 3.361e-02A M=8.598e-07
I3040 0 n3041 3.361e-02A M=1.105e-06
I3041 0 n3042 3.361e-02A M=6.260e-07
I3042 0 n3043 3.361e-02A M=1.045e-06
I3043 0 n3044 3.361e-02A M=1.040e-06
I3044 0 n3045 3.361e-02A M=5.659e-07
I3045 0 n3046 3.361e-02A M=6.913e-07
I3046 0 n3047 3.361e-02A M=3.177e-07
I3047 0 n3048 3.361e-02A M=2.671e-06
I3048 0 n3049 3.361e-02A M=1.763e-07
I3049 0 n3050 3.361e-02A M=1.509e-06
I3050 0 n3051 3.361e-02A M=1.236e-06
I3051 0 n3052 3.361e-02A M=1.944e-06
I3052 0 n3053 3.361e-02A M=7.637e-07
I3053 0 n3054 3.361e-02A M=4.088e-07
I3054 0 n3055 3.361e-02A M=1.767e-06
I3055 0 n3056 3.361e-02A M=9.397e-07
I3056 0 n3057 3.361e-02A M=9.379e-07
I3057 0 n3058 3.361e-02A M=4.370e-07
I3058 0 n3059 3.361e-02A M=2.346e-06
I3059 0 n3060 3.361e-02A M=1.004e-06
I3060 0 n3061 3.361e-02A M=7.516e-07
I3061 0 n3062 3.361e-02A M=1.238e-06
I3062 0 n3063 3.361e-02A M=8.882e-07
I3063 0 n3064 3.361e-02A M=6.832e-07
I3064 0 n3065 3.361e-02A M=1.197e-06
I3065 0 n3066 3.361e-02A M=7.290e-07
I3066 0 n3067 3.361e-02A M=5.046e-07
I3067 0 n3068 3.361e-02A M=6.312e-07
I3068 0 n3069 3.361e-02A M=9.035e-07
I3069 0 n3070 3.361e-02A M=2.501e-07
I3070 0 n3071 3.361e-02A M=1.431e-06
I3071 0 n3072 3.361e-02A M=7.918e-07
I3072 0 n3073 3.361e-02A M=2.383e-07
I3073 0 n3074 3.361e-02A M=8.397e-07
I3074 0 n3075 3.361e-02A M=1.009e-06
I3075 0 n3076 3.361e-02A M=7.869e-07
I3076 0 n3077 3.361e-02A M=3.836e-07
I3077 0 n3078 3.361e-02A M=1.171e-06
I3078 0 n3079 3.361e-02A M=7.467e-07
I3079 0 n3080 3.361e-02A M=5.089e-07
I3080 0 n3081 3.361e-02A M=7.583e-07
I3081 0 n3082 3.361e-02A M=1.043e-06
I3082 0 n3083 3.361e-02A M=9.499e-07
I3083 0 n3084 3.361e-02A M=7.259e-07
I3084 0 n3085 3.361e-02A M=1.292e-06
I3085 0 n3086 3.361e-02A M=3.168e-06
I3086 0 n3087 3.361e-02A M=9.293e-07
I3087 0 n3088 3.361e-02A M=7.963e-07
I3088 0 n3089 3.361e-02A M=6.874e-07
I3089 0 n3090 3.361e-02A M=5.622e-07
I3090 0 n3091 3.361e-02A M=1.168e-06
I3091 0 n3092 3.361e-02A M=3.077e-07
I3092 0 n3093 3.361e-02A M=8.051e-07
I3093 0 n3094 3.361e-02A M=7.781e-07
I3094 0 n3095 3.361e-02A M=1.969e-06
I3095 0 n3096 3.361e-02A M=5.864e-07
I3096 0 n3097 3.361e-02A M=1.170e-06
I3097 0 n1 3.361e-02A M=8.112e-07
I3098 0 n3099 3.361e-02A M=9.582e-07
I3099 0 n3100 3.361e-02A M=7.084e-07
I3100 0 n3101 3.361e-02A M=1.219e-06
I3101 0 n3102 3.361e-02A M=9.306e-07
I3102 0 n3103 3.361e-02A M=1.219e-06
I3103 0 n3104 3.361e-02A M=6.750e-07
I3104 0 n3105 3.361e-02A M=6.249e-07
I3105 0 n3106 3.361e-02A M=9.499e-07
I3106 0 n3107 3.361e-02A M=1.793e-06
I3107 0 n3108 3.361e-02A M=1.068e-06
I3108 0 n3109 3.361e-02A M=1.819e-06
I3109 0 n3110 3.361e-02A M=2.095e-06
I3110 0 n3111 3.361e-02A M=2.091e-07
I3111 0 n1 3.361e-02A M=6.818e-07
I3112 0 n3113 3.361e-02A M=8.972e-07
I3113 0 n3114 3.361e-02A M=9.313e-07
I3114 0 n3115 3.361e-02A M=8.400e-07
I3115 0 n3116 3.361e-02A M=2.551e-06
I3116 0 n3117 3.361e-02A M=9.038e-07
I3117 0 n3118 3.361e-02A M=1.205e-06
I3118 0 n3119 3.361e-02A M=6.252e-07
I3119 0 n3120 3.361e-02A M=1.306e-06
I3120 0 n3121 3.361e-02A M=1.133e-06
I3121 0 n3122 3.361e-02A M=2.951e-07
I3122 0 n3123 3.361e-02A M=1.065e-06
I3123 0 n3124 3.361e-02A M=3.100e-07
I3124 0 n3125 3.361e-02A M=2.477e-06
I3125 0 n3126 3.361e-02A M=9.202e-07
I3126 0 n3127 3.361e-02A M=8.589e-07
I3127 0 n3128 3.361e-02A M=8.086e-07
I3128 0 n3129 3.361e-02A M=1.199e-06
I3129 0 n3130 3.361e-02A M=2.096e-07
I3130 0 n3131 3.361e-02A M=7.131e-07
I3131 0 n3132 3.361e-02A M=5.885e-07
I3132 0 n3133 3.361e-02A M=6.421e-07
I3133 0 n3134 3.361e-02A M=1.557e-06
I3134 0 n3135 3.361e-02A M=1.333e-06
I3135 0 n3136 3.361e-02A M=4.375e-07
I3136 0 n3137 3.361e-02A M=1.842e-06
I3137 0 n3138 3.361e-02A M=7.350e-07
I3138 0 n3139 3.361e-02A M=8.150e-07
I3139 0 n3140 3.361e-02A M=3.884e-07
I3140 0 n3141 3.361e-02A M=1.122e-06
I3141 0 n3142 3.361e-02A M=1.264e-06
I3142 0 n3143 3.361e-02A M=1.698e-06
I3143 0 n3144 3.361e-02A M=9.457e-07
I3144 0 n3145 3.361e-02A M=3.199e-07
I3145 0 n3146 3.361e-02A M=9.039e-07
I3146 0 n3147 3.361e-02A M=5.886e-07
I3147 0 n3148 3.361e-02A M=1.837e-07
I3148 0 n3149 3.361e-02A M=7.564e-07
I3149 0 n3150 3.361e-02A M=1.911e-06
I3150 0 n3151 3.361e-02A M=3.866e-07
I3151 0 n3152 3.361e-02A M=5.437e-07
I3152 0 n3153 3.361e-02A M=2.471e-06
I3153 0 n3154 3.361e-02A M=1.527e-06
I3154 0 n3155 3.361e-02A M=9.242e-07
I3155 0 n3156 3.361e-02A M=2.815e-07
I3156 0 n3157 3.361e-02A M=4.096e-07
I3157 0 n3158 3.361e-02A M=1.195e-06
I3158 0 n3159 3.361e-02A M=3.585e-07
I3159 0 n3160 3.361e-02A M=1.427e-06
I3160 0 n3161 3.361e-02A M=6.595e-07
I3161 0 n3162 3.361e-02A M=3.674e-07
I3162 0 n3163 3.361e-02A M=5.909e-07
I3163 0 n3164 3.361e-02A M=1.406e-06
I3164 0 n3165 3.361e-02A M=8.995e-07
I3165 0 n3166 3.361e-02A M=1.434e-06
I3166 0 n3167 3.361e-02A M=9.021e-07
I3167 0 n3168 3.361e-02A M=4.819e-07
I3168 0 n1 3.361e-02A M=5.590e-07
I3169 0 n3170 3.361e-02A M=6.624e-07
I3170 0 n3171 3.361e-02A M=1.604e-06
I3171 0 n3172 3.361e-02A M=7.385e-07
I3172 0 n3173 3.361e-02A M=1.737e-06
I3173 0 n3174 3.361e-02A M=4.944e-07
I3174 0 n3175 3.361e-02A M=1.518e-06
I3175 0 n3176 3.361e-02A M=1.206e-06
I3176 0 n3177 3.361e-02A M=9.571e-07
I3177 0 n3178 3.361e-02A M=5.500e-07
I3178 0 n3179 3.361e-02A M=2.243e-06
I3179 0 n3180 3.361e-02A M=2.543e-06
I3180 0 n3181 3.361e-02A M=1.555e-06
I3181 0 n3182 3.361e-02A M=1.292e-06
I3182 0 n3183 3.361e-02A M=7.488e-07
I3183 0 n3184 3.361e-02A M=9.221e-07
I3184 0 n3185 3.361e-02A M=1.035e-06
I3185 0 n3186 3.361e-02A M=8.766e-07
I3186 0 n3187 3.361e-02A M=7.471e-07
I3187 0 n3188 3.361e-02A M=7.138e-07
I3188 0 n3189 3.361e-02A M=1.063e-06
I3189 0 n3190 3.361e-02A M=1.673e-06
I3190 0 n3191 3.361e-02A M=2.002e-06
I3191 0 n3192 3.361e-02A M=1.573e-06
I3192 0 n3193 3.361e-02A M=5.667e-07
I3193 0 n3194 3.361e-02A M=9.128e-07
I3194 0 n3195 3.361e-02A M=1.175e-06
I3195 0 n3196 3.361e-02A M=4.331e-07
I3196 0 n3197 3.361e-02A M=4.904e-07
I3197 0 n3198 3.361e-02A M=1.337e-06
I3198 0 n3199 3.361e-02A M=5.878e-07
I3199 0 n3200 3.361e-02A M=6.193e-07
I3200 0 n3201 3.361e-02A M=9.687e-07
I3201 0 n3202 3.361e-02A M=5.935e-07
I3202 0 n3203 3.361e-02A M=1.650e-06
I3203 0 n3204 3.361e-02A M=8.513e-07
I3204 0 n3205 3.361e-02A M=3.276e-06
I3205 0 n3206 3.361e-02A M=9.200e-07
I3206 0 n3207 3.361e-02A M=2.237e-07
I3207 0 n3208 3.361e-02A M=1.623e-06
I3208 0 n3209 3.361e-02A M=2.144e-06
I3209 0 n3210 3.361e-02A M=7.932e-07
I3210 0 n3211 3.361e-02A M=5.045e-07
I3211 0 n3212 3.361e-02A M=1.642e-06
I3212 0 n3213 3.361e-02A M=1.706e-06
I3213 0 n3214 3.361e-02A M=1.646e-06
I3214 0 n3215 3.361e-02A M=7.743e-07
I3215 0 n3216 3.361e-02A M=1.050e-06
I3216 0 n3217 3.361e-02A M=6.950e-07
I3217 0 n3218 3.361e-02A M=1.650e-06
I3218 0 n3219 3.361e-02A M=9.950e-07
I3219 0 n3220 3.361e-02A M=7.357e-07
I3220 0 n3221 3.361e-02A M=9.130e-07
I3221 0 n3222 3.361e-02A M=1.256e-06
I3222 0 n3223 3.361e-02A M=9.531e-07
I3223 0 n1 3.361e-02A M=1.541e-06
I3224 0 n3225 3.361e-02A M=1.068e-06
I3225 0 n3226 3.361e-02A M=1.586e-06
I3226 0 n3227 3.361e-02A M=3.361e-07
I3227 0 n3228 3.361e-02A M=1.186e-06
I3228 0 n3229 3.361e-02A M=4.805e-07
I3229 0 n3230 3.361e-02A M=1.298e-06
I3230 0 n3231 3.361e-02A M=1.017e-06
I3231 0 n3232 3.361e-02A M=3.678e-07
I3232 0 n3233 3.361e-02A M=1.294e-06
I3233 0 n3234 3.361e-02A M=6.979e-07
I3234 0 n3235 3.361e-02A M=5.370e-07
I3235 0 n3236 3.361e-02A M=2.337e-06
I3236 0 n3237 3.361e-02A M=9.499e-07
I3237 0 n3238 3.361e-02A M=1.205e-06
I3238 0 n3239 3.361e-02A M=3.072e-07
I3239 0 n3240 3.361e-02A M=1.185e-06
I3240 0 n3241 3.361e-02A M=5.544e-07
I3241 0 n3242 3.361e-02A M=1.182e-06
I3242 0 n3243 3.361e-02A M=1.484e-06
I3243 0 n3244 3.361e-02A M=4.547e-07
I3244 0 n3245 3.361e-02A M=1.330e-06
I3245 0 n3246 3.361e-02A M=1.250e-06
I3246 0 n3247 3.361e-02A M=6.190e-07
I3247 0 n3248 3.361e-02A M=1.735e-06
I3248 0 n3249 3.361e-02A M=8.484e-07
I3249 0 n3250 3.361e-02A M=8.984e-07
I3250 0 n3251 3.361e-02A M=1.075e-06
I3251 0 n3252 3.361e-02A M=1.981e-06
I3252 0 n3253 3.361e-02A M=2.834e-07
I3253 0 n3254 3.361e-02A M=7.942e-07
I3254 0 n3255 3.361e-02A M=1.821e-06
I3255 0 n3256 3.361e-02A M=1.178e-06
I3256 0 n3257 3.361e-02A M=1.245e-06
I3257 0 n3258 3.361e-02A M=1.262e-06
I3258 0 n3259 3.361e-02A M=6.216e-07
I3259 0 n3260 3.361e-02A M=1.317e-06
I3260 0 n3261 3.361e-02A M=1.943e-06
I3261 0 n3262 3.361e-02A M=1.014e-06
I3262 0 n3263 3.361e-02A M=7.745e-07
I3263 0 n3264 3.361e-02A M=8.424e-07
I3264 0 n3265 3.361e-02A M=1.671e-06
I3265 0 n3266 3.361e-02A M=9.595e-07
I3266 0 n3267 3.361e-02A M=1.811e-06
I3267 0 n3268 3.361e-02A M=3.827e-07
I3268 0 n3269 3.361e-02A M=9.709e-07
I3269 0 n3270 3.361e-02A M=8.924e-07
I3270 0 n3271 3.361e-02A M=1.354e-06
I3271 0 n3272 3.361e-02A M=1.102e-06
I3272 0 n3273 3.361e-02A M=4.783e-07
I3273 0 n3274 3.361e-02A M=1.675e-06
I3274 0 n3275 3.361e-02A M=3.001e-07
I3275 0 n3276 3.361e-02A M=1.166e-06
I3276 0 n3277 3.361e-02A M=1.204e-06
I3277 0 n3278 3.361e-02A M=1.913e-06
I3278 0 n3279 3.361e-02A M=1.475e-06
I3279 0 n3280 3.361e-02A M=5.593e-07
I3280 0 n3281 3.361e-02A M=3.517e-07
I3281 0 n3282 3.361e-02A M=4.707e-07
I3282 0 n3283 3.361e-02A M=1.963e-06
I3283 0 n3284 3.361e-02A M=8.975e-07
I3284 0 n3285 3.361e-02A M=1.219e-06
I3285 0 n3286 3.361e-02A M=8.695e-07
I3286 0 n3287 3.361e-02A M=1.220e-06
I3287 0 n3288 3.361e-02A M=1.005e-06
I3288 0 n3289 3.361e-02A M=1.195e-06
I3289 0 n3290 3.361e-02A M=1.116e-06
I3290 0 n3291 3.361e-02A M=3.205e-07
I3291 0 n3292 3.361e-02A M=3.278e-07
I3292 0 n3293 3.361e-02A M=4.874e-07
I3293 0 n3294 3.361e-02A M=8.093e-07
I3294 0 n3295 3.361e-02A M=6.401e-07
I3295 0 n3296 3.361e-02A M=1.014e-06
I3296 0 n3297 3.361e-02A M=4.697e-07
I3297 0 n3298 3.361e-02A M=9.805e-07
I3298 0 n3299 3.361e-02A M=2.225e-07
I3299 0 n3300 3.361e-02A M=1.319e-06
I3300 0 n3301 3.361e-02A M=1.168e-06
I3301 0 n3302 3.361e-02A M=1.077e-06
I3302 0 n3303 3.361e-02A M=8.574e-07
I3303 0 n3304 3.361e-02A M=1.037e-06
I3304 0 n3305 3.361e-02A M=9.708e-07
I3305 0 n3306 3.361e-02A M=8.413e-07
I3306 0 n3307 3.361e-02A M=6.561e-07
I3307 0 n3308 3.361e-02A M=1.410e-06
I3308 0 n1 3.361e-02A M=4.512e-07
I3309 0 n3310 3.361e-02A M=3.962e-07
I3310 0 n3311 3.361e-02A M=1.168e-06
I3311 0 n3312 3.361e-02A M=1.559e-06
I3312 0 n3313 3.361e-02A M=1.205e-06
I3313 0 n3314 3.361e-02A M=6.442e-07
I3314 0 n3315 3.361e-02A M=9.995e-07
I3315 0 n3316 3.361e-02A M=7.204e-07
I3316 0 n3317 3.361e-02A M=1.118e-06
I3317 0 n3318 3.361e-02A M=8.018e-07
I3318 0 n3319 3.361e-02A M=1.487e-06
I3319 0 n3320 3.361e-02A M=1.948e-07
I3320 0 n3321 3.361e-02A M=1.329e-06
I3321 0 n3322 3.361e-02A M=1.658e-06
I3322 0 n3323 3.361e-02A M=3.894e-07
I3323 0 n3324 3.361e-02A M=1.165e-06
I3324 0 n3325 3.361e-02A M=7.764e-07
I3325 0 n3326 3.361e-02A M=2.292e-06
I3326 0 n3327 3.361e-02A M=1.103e-06
I3327 0 n3328 3.361e-02A M=6.603e-07
I3328 0 n3329 3.361e-02A M=3.853e-07
I3329 0 n3330 3.361e-02A M=5.541e-07
I3330 0 n3331 3.361e-02A M=7.181e-07
I3331 0 n3332 3.361e-02A M=1.374e-06
I3332 0 n3333 3.361e-02A M=6.538e-07
I3333 0 n3334 3.361e-02A M=1.214e-06
I3334 0 n3335 3.361e-02A M=1.400e-06
I3335 0 n3336 3.361e-02A M=1.720e-07
I3336 0 n3337 3.361e-02A M=7.276e-07
I3337 0 n3338 3.361e-02A M=6.675e-07
I3338 0 n3339 3.361e-02A M=1.317e-06
I3339 0 n3340 3.361e-02A M=4.944e-07
I3340 0 n3341 3.361e-02A M=2.774e-07
I3341 0 n3342 3.361e-02A M=1.085e-06
I3342 0 n3343 3.361e-02A M=5.248e-07
I3343 0 n3344 3.361e-02A M=1.442e-06
I3344 0 n3345 3.361e-02A M=7.903e-07
I3345 0 n3346 3.361e-02A M=8.975e-07
I3346 0 n3347 3.361e-02A M=3.263e-07
I3347 0 n3348 3.361e-02A M=8.164e-07
I3348 0 n3349 3.361e-02A M=1.577e-06
I3349 0 n3350 3.361e-02A M=1.438e-06
I3350 0 n3351 3.361e-02A M=1.158e-06
I3351 0 n3352 3.361e-02A M=1.738e-06
I3352 0 n3353 3.361e-02A M=2.105e-06
I3353 0 n3354 3.361e-02A M=1.195e-06
I3354 0 n3355 3.361e-02A M=8.934e-07
I3355 0 n3356 3.361e-02A M=6.286e-07
I3356 0 n3357 3.361e-02A M=1.577e-06
I3357 0 n3358 3.361e-02A M=1.255e-06
I3358 0 n3359 3.361e-02A M=1.531e-06
I3359 0 n3360 3.361e-02A M=1.168e-06
I3360 0 n3361 3.361e-02A M=6.232e-07
I3361 0 n3362 3.361e-02A M=6.038e-07
I3362 0 n3363 3.361e-02A M=2.118e-07
I3363 0 n3364 3.361e-02A M=4.762e-07
I3364 0 n3365 3.361e-02A M=3.399e-06
I3365 0 n3366 3.361e-02A M=7.991e-07
I3366 0 n3367 3.361e-02A M=7.441e-07
I3367 0 n3368 3.361e-02A M=1.105e-06
I3368 0 n3369 3.361e-02A M=6.136e-07
I3369 0 n3370 3.361e-02A M=9.790e-07
I3370 0 n3371 3.361e-02A M=1.709e-06
I3371 0 n3372 3.361e-02A M=1.329e-06
I3372 0 n3373 3.361e-02A M=5.898e-07
I3373 0 n3374 3.361e-02A M=6.460e-07
I3374 0 n3375 3.361e-02A M=9.353e-07
I3375 0 n3376 3.361e-02A M=4.603e-07
I3376 0 n3377 3.361e-02A M=4.813e-07
I3377 0 n3378 3.361e-02A M=1.112e-06
I3378 0 n3379 3.361e-02A M=5.421e-07
I3379 0 n3380 3.361e-02A M=9.532e-07
I3380 0 n3381 3.361e-02A M=9.892e-07
I3381 0 n3382 3.361e-02A M=1.011e-06
I3382 0 n3383 3.361e-02A M=5.068e-07
I3383 0 n3384 3.361e-02A M=8.408e-07
I3384 0 n3385 3.361e-02A M=1.070e-06
I3385 0 n3386 3.361e-02A M=2.150e-06
I3386 0 n3387 3.361e-02A M=2.400e-06
I3387 0 n3388 3.361e-02A M=1.893e-06
I3388 0 n3389 3.361e-02A M=2.107e-07
I3389 0 n1 3.361e-02A M=1.303e-06
I3390 0 n3391 3.361e-02A M=8.001e-07
I3391 0 n3392 3.361e-02A M=8.373e-07
I3392 0 n3393 3.361e-02A M=4.289e-07
I3393 0 n3394 3.361e-02A M=8.073e-07
I3394 0 n3395 3.361e-02A M=5.557e-07
I3395 0 n3396 3.361e-02A M=4.272e-07
I3396 0 n3397 3.361e-02A M=9.078e-07
I3397 0 n3398 3.361e-02A M=1.197e-06
I3398 0 n3399 3.361e-02A M=1.134e-06
I3399 0 n3400 3.361e-02A M=9.934e-07
I3400 0 n3401 3.361e-02A M=7.343e-07
I3401 0 n3402 3.361e-02A M=6.339e-07
I3402 0 n3403 3.361e-02A M=1.073e-06
I3403 0 n3404 3.361e-02A M=5.057e-07
I3404 0 n3405 3.361e-02A M=4.601e-07
I3405 0 n3406 3.361e-02A M=4.014e-07
I3406 0 n3407 3.361e-02A M=1.278e-06
I3407 0 n3408 3.361e-02A M=6.991e-07
I3408 0 n3409 3.361e-02A M=5.256e-07
I3409 0 n3410 3.361e-02A M=4.602e-07
I3410 0 n3411 3.361e-02A M=6.855e-07
I3411 0 n3412 3.361e-02A M=8.425e-07
I3412 0 n3413 3.361e-02A M=1.047e-06
I3413 0 n3414 3.361e-02A M=6.204e-07
I3414 0 n3415 3.361e-02A M=5.029e-07
I3415 0 n3416 3.361e-02A M=9.759e-07
I3416 0 n3417 3.361e-02A M=2.203e-06
I3417 0 n3418 3.361e-02A M=2.839e-06
I3418 0 n3419 3.361e-02A M=9.128e-07
I3419 0 n3420 3.361e-02A M=6.342e-07
I3420 0 n3421 3.361e-02A M=9.046e-07
I3421 0 n3422 3.361e-02A M=1.046e-06
I3422 0 n3423 3.361e-02A M=1.956e-06
I3423 0 n3424 3.361e-02A M=5.614e-07
I3424 0 n3425 3.361e-02A M=8.055e-07
I3425 0 n3426 3.361e-02A M=6.947e-07
I3426 0 n3427 3.361e-02A M=8.997e-07
I3427 0 n3428 3.361e-02A M=8.377e-07
I3428 0 n3429 3.361e-02A M=6.291e-07
I3429 0 n3430 3.361e-02A M=9.511e-07
I3430 0 n3431 3.361e-02A M=6.853e-07
I3431 0 n3432 3.361e-02A M=4.940e-07
I3432 0 n3433 3.361e-02A M=9.948e-07
I3433 0 n3434 3.361e-02A M=1.039e-06
I3434 0 n3435 3.361e-02A M=6.267e-07
I3435 0 n3436 3.361e-02A M=9.085e-07
I3436 0 n3437 3.361e-02A M=1.018e-06
I3437 0 n3438 3.361e-02A M=1.868e-06
I3438 0 n3439 3.361e-02A M=1.389e-06
I3439 0 n3440 3.361e-02A M=1.234e-06
I3440 0 n3441 3.361e-02A M=1.280e-06
I3441 0 n3442 3.361e-02A M=5.854e-07
I3442 0 n3443 3.361e-02A M=3.899e-07
I3443 0 n3444 3.361e-02A M=8.201e-07
I3444 0 n3445 3.361e-02A M=2.094e-06
I3445 0 n3446 3.361e-02A M=1.419e-06
I3446 0 n3447 3.361e-02A M=1.547e-06
I3447 0 n3448 3.361e-02A M=6.824e-07
I3448 0 n3449 3.361e-02A M=1.199e-06
I3449 0 n3450 3.361e-02A M=1.235e-06
I3450 0 n3451 3.361e-02A M=1.154e-06
I3451 0 n3452 3.361e-02A M=1.001e-06
I3452 0 n3453 3.361e-02A M=1.270e-06
I3453 0 n3454 3.361e-02A M=1.179e-06
I3454 0 n3455 3.361e-02A M=1.038e-06
I3455 0 n3456 3.361e-02A M=8.039e-07
I3456 0 n3457 3.361e-02A M=1.072e-06
I3457 0 n3458 3.361e-02A M=1.196e-06
I3458 0 n3459 3.361e-02A M=6.508e-07
I3459 0 n3460 3.361e-02A M=1.262e-06
I3460 0 n3461 3.361e-02A M=1.130e-06
I3461 0 n3462 3.361e-02A M=1.067e-06
I3462 0 n3463 3.361e-02A M=2.235e-07
I3463 0 n3464 3.361e-02A M=9.599e-07
I3464 0 n3465 3.361e-02A M=1.863e-06
I3465 0 n3466 3.361e-02A M=1.197e-06
I3466 0 n3467 3.361e-02A M=5.227e-07
I3467 0 n3468 3.361e-02A M=1.373e-06
I3468 0 n3469 3.361e-02A M=1.440e-06
I3469 0 n3470 3.361e-02A M=1.922e-06
I3470 0 n3471 3.361e-02A M=1.047e-06
I3471 0 n3472 3.361e-02A M=9.311e-07
I3472 0 n3473 3.361e-02A M=5.262e-07
I3473 0 n3474 3.361e-02A M=5.634e-07
I3474 0 n3475 3.361e-02A M=4.553e-07
I3475 0 n3476 3.361e-02A M=6.511e-07
I3476 0 n3477 3.361e-02A M=8.479e-07
I3477 0 n3478 3.361e-02A M=4.146e-07
I3478 0 n3479 3.361e-02A M=3.726e-07
I3479 0 n3480 3.361e-02A M=1.159e-06
I3480 0 n3481 3.361e-02A M=4.782e-07
I3481 0 n3482 3.361e-02A M=2.054e-06
I3482 0 n3483 3.361e-02A M=1.548e-06
I3483 0 n3484 3.361e-02A M=1.712e-07
I3484 0 n3485 3.361e-02A M=1.472e-07
I3485 0 n3486 3.361e-02A M=7.066e-07
I3486 0 n3487 3.361e-02A M=1.656e-06
I3487 0 n3488 3.361e-02A M=1.123e-06
I3488 0 n3489 3.361e-02A M=6.639e-07
I3489 0 n3490 3.361e-02A M=1.095e-06
I3490 0 n3491 3.361e-02A M=1.486e-06
I3491 0 n3492 3.361e-02A M=1.221e-06
I3492 0 n1 3.361e-02A M=8.609e-07
I3493 0 n3494 3.361e-02A M=1.991e-06
I3494 0 n3495 3.361e-02A M=3.499e-07
I3495 0 n3496 3.361e-02A M=6.659e-07
I3496 0 n3497 3.361e-02A M=1.197e-06
I3497 0 n3498 3.361e-02A M=7.153e-07
I3498 0 n3499 3.361e-02A M=4.466e-07
I3499 0 n3500 3.361e-02A M=9.738e-07
I3500 0 n3501 3.361e-02A M=1.068e-06
I3501 0 n3502 3.361e-02A M=6.088e-07
I3502 0 n3503 3.361e-02A M=1.255e-06
I3503 0 n3504 3.361e-02A M=1.329e-06
I3504 0 n3505 3.361e-02A M=1.168e-06
I3505 0 n3506 3.361e-02A M=4.340e-07
I3506 0 n3507 3.361e-02A M=5.992e-07
I3507 0 n3508 3.361e-02A M=1.200e-06
I3508 0 n3509 3.361e-02A M=1.564e-06
I3509 0 n3510 3.361e-02A M=7.002e-07
I3510 0 n3511 3.361e-02A M=1.360e-06
I3511 0 n3512 3.361e-02A M=1.663e-07
I3512 0 n3513 3.361e-02A M=8.436e-07
I3513 0 n3514 3.361e-02A M=1.075e-06
I3514 0 n3515 3.361e-02A M=1.701e-06
I3515 0 n3516 3.361e-02A M=1.102e-06
I3516 0 n3517 3.361e-02A M=1.729e-06
I3517 0 n3518 3.361e-02A M=1.079e-06
I3518 0 n3519 3.361e-02A M=8.206e-07
I3519 0 n3520 3.361e-02A M=4.018e-07
I3520 0 n3521 3.361e-02A M=4.024e-07
I3521 0 n3522 3.361e-02A M=9.371e-07
I3522 0 n3523 3.361e-02A M=1.169e-06
I3523 0 n3524 3.361e-02A M=5.914e-07
I3524 0 n3525 3.361e-02A M=8.012e-07
I3525 0 n3526 3.361e-02A M=6.652e-07
I3526 0 n3527 3.361e-02A M=6.790e-07
I3527 0 n3528 3.361e-02A M=1.091e-06
I3528 0 n3529 3.361e-02A M=1.311e-06
I3529 0 n3530 3.361e-02A M=1.367e-06
I3530 0 n3531 3.361e-02A M=1.117e-06
I3531 0 n3532 3.361e-02A M=6.338e-07
I3532 0 n3533 3.361e-02A M=4.755e-07
I3533 0 n3534 3.361e-02A M=1.025e-06
I3534 0 n3535 3.361e-02A M=1.193e-06
I3535 0 n3536 3.361e-02A M=1.101e-06
I3536 0 n3537 3.361e-02A M=1.503e-06
I3537 0 n3538 3.361e-02A M=5.089e-07
I3538 0 n3539 3.361e-02A M=1.694e-06
I3539 0 n3540 3.361e-02A M=5.611e-07
I3540 0 n3541 3.361e-02A M=9.565e-07
I3541 0 n3542 3.361e-02A M=3.052e-07
I3542 0 n3543 3.361e-02A M=1.661e-06
I3543 0 n3544 3.361e-02A M=4.717e-07
I3544 0 n3545 3.361e-02A M=5.777e-07
I3545 0 n3546 3.361e-02A M=1.097e-06
I3546 0 n3547 3.361e-02A M=1.057e-06
I3547 0 n3548 3.361e-02A M=1.149e-06
I3548 0 n3549 3.361e-02A M=8.004e-07
I3549 0 n3550 3.361e-02A M=3.880e-07
I3550 0 n3551 3.361e-02A M=8.372e-07
I3551 0 n3552 3.361e-02A M=1.303e-06
I3552 0 n3553 3.361e-02A M=9.362e-07
I3553 0 n3554 3.361e-02A M=1.474e-06
I3554 0 n3555 3.361e-02A M=9.057e-07
I3555 0 n3556 3.361e-02A M=1.265e-06
I3556 0 n3557 3.361e-02A M=1.295e-06
I3557 0 n3558 3.361e-02A M=1.297e-06
I3558 0 n3559 3.361e-02A M=8.131e-07
I3559 0 n3560 3.361e-02A M=5.561e-07
I3560 0 n3561 3.361e-02A M=9.633e-07
I3561 0 n3562 3.361e-02A M=1.347e-06
I3562 0 n3563 3.361e-02A M=3.811e-07
I3563 0 n3564 3.361e-02A M=1.004e-06
I3564 0 n3565 3.361e-02A M=1.225e-06
I3565 0 n3566 3.361e-02A M=6.895e-07
I3566 0 n3567 3.361e-02A M=9.378e-07
I3567 0 n3568 3.361e-02A M=8.345e-07
I3568 0 n3569 3.361e-02A M=6.322e-07
I3569 0 n3570 3.361e-02A M=1.114e-06
I3570 0 n3571 3.361e-02A M=1.205e-06
I3571 0 n3572 3.361e-02A M=1.251e-06
I3572 0 n3573 3.361e-02A M=2.637e-07
I3573 0 n3574 3.361e-02A M=4.824e-07
I3574 0 n3575 3.361e-02A M=6.628e-07
I3575 0 n3576 3.361e-02A M=9.062e-07
I3576 0 n3577 3.361e-02A M=9.680e-07
I3577 0 n3578 3.361e-02A M=6.220e-07
I3578 0 n3579 3.361e-02A M=1.318e-06
I3579 0 n3580 3.361e-02A M=1.269e-06
I3580 0 n3581 3.361e-02A M=8.664e-07
I3581 0 n3582 3.361e-02A M=9.764e-07
I3582 0 n3583 3.361e-02A M=2.039e-07
I3583 0 n3584 3.361e-02A M=1.362e-06
I3584 0 n3585 3.361e-02A M=1.858e-06
I3585 0 n3586 3.361e-02A M=6.656e-07
I3586 0 n3587 3.361e-02A M=8.165e-07
I3587 0 n3588 3.361e-02A M=7.933e-07
I3588 0 n3589 3.361e-02A M=1.183e-06
I3589 0 n3590 3.361e-02A M=1.706e-06
I3590 0 n3591 3.361e-02A M=1.444e-06
I3591 0 n3592 3.361e-02A M=1.495e-06
I3592 0 n3593 3.361e-02A M=1.759e-06
I3593 0 n3594 3.361e-02A M=1.413e-06
I3594 0 n3595 3.361e-02A M=4.286e-07
I3595 0 n3596 3.361e-02A M=1.285e-06
I3596 0 n3597 3.361e-02A M=2.806e-06
I3597 0 n3598 3.361e-02A M=8.495e-07
I3598 0 n3599 3.361e-02A M=1.073e-06
I3599 0 n3600 3.361e-02A M=8.035e-07
I3600 0 n3601 3.361e-02A M=6.542e-07
I3601 0 n3602 3.361e-02A M=6.276e-07
I3602 0 n3603 3.361e-02A M=1.561e-06
I3603 0 n3604 3.361e-02A M=9.641e-07
I3604 0 n3605 3.361e-02A M=8.403e-07
I3605 0 n3606 3.361e-02A M=1.072e-06
I3606 0 n3607 3.361e-02A M=1.011e-06
I3607 0 n3608 3.361e-02A M=8.701e-07
I3608 0 n3609 3.361e-02A M=1.191e-06
I3609 0 n3610 3.361e-02A M=8.743e-07
I3610 0 n3611 3.361e-02A M=2.543e-07
I3611 0 n3612 3.361e-02A M=1.302e-06
I3612 0 n3613 3.361e-02A M=4.432e-07
I3613 0 n3614 3.361e-02A M=1.542e-07
I3614 0 n3615 3.361e-02A M=2.613e-06
I3615 0 n3616 3.361e-02A M=3.373e-07
I3616 0 n3617 3.361e-02A M=6.871e-07
I3617 0 n3618 3.361e-02A M=7.901e-07
I3618 0 n3619 3.361e-02A M=1.175e-06
I3619 0 n3620 3.361e-02A M=5.834e-07
I3620 0 n3621 3.361e-02A M=5.379e-07
I3621 0 n3622 3.361e-02A M=6.775e-07
I3622 0 n3623 3.361e-02A M=6.263e-07
I3623 0 n3624 3.361e-02A M=1.496e-06
I3624 0 n3625 3.361e-02A M=1.579e-06
I3625 0 n3626 3.361e-02A M=2.819e-07
I3626 0 n3627 3.361e-02A M=1.627e-06
I3627 0 n3628 3.361e-02A M=3.135e-07
I3628 0 n3629 3.361e-02A M=3.588e-07
I3629 0 n3630 3.361e-02A M=6.379e-07
I3630 0 n3631 3.361e-02A M=5.745e-07
I3631 0 n3632 3.361e-02A M=3.903e-07
I3632 0 n3633 3.361e-02A M=1.052e-06
I3633 0 n3634 3.361e-02A M=2.176e-06
I3634 0 n3635 3.361e-02A M=1.286e-06
I3635 0 n3636 3.361e-02A M=9.360e-07
I3636 0 n3637 3.361e-02A M=5.289e-07
I3637 0 n3638 3.361e-02A M=9.777e-07
I3638 0 n3639 3.361e-02A M=1.263e-06
I3639 0 n3640 3.361e-02A M=6.518e-07
I3640 0 n3641 3.361e-02A M=1.013e-06
I3641 0 n3642 3.361e-02A M=9.030e-07
I3642 0 n3643 3.361e-02A M=1.000e-06
I3643 0 n3644 3.361e-02A M=1.066e-06
I3644 0 n3645 3.361e-02A M=9.494e-07
I3645 0 n3646 3.361e-02A M=8.755e-07
I3646 0 n3647 3.361e-02A M=1.094e-06
I3647 0 n3648 3.361e-02A M=1.267e-06
I3648 0 n3649 3.361e-02A M=7.411e-07
I3649 0 n3650 3.361e-02A M=8.164e-07
I3650 0 n3651 3.361e-02A M=1.320e-06
I3651 0 n3652 3.361e-02A M=9.501e-07
I3652 0 n3653 3.361e-02A M=8.165e-07
I3653 0 n3654 3.361e-02A M=5.036e-07
I3654 0 n3655 3.361e-02A M=8.015e-07
I3655 0 n3656 3.361e-02A M=1.366e-06
I3656 0 n3657 3.361e-02A M=8.999e-07
I3657 0 n3658 3.361e-02A M=5.180e-07
I3658 0 n3659 3.361e-02A M=3.751e-07
I3659 0 n3660 3.361e-02A M=4.227e-07
I3660 0 n3661 3.361e-02A M=4.283e-07
I3661 0 n3662 3.361e-02A M=1.656e-06
I3662 0 n3663 3.361e-02A M=5.555e-07
I3663 0 n3664 3.361e-02A M=1.055e-06
I3664 0 n3665 3.361e-02A M=9.698e-07
I3665 0 n3666 3.361e-02A M=7.029e-07
I3666 0 n3667 3.361e-02A M=2.396e-06
I3667 0 n3668 3.361e-02A M=8.458e-07
I3668 0 n3669 3.361e-02A M=1.745e-06
I3669 0 n3670 3.361e-02A M=9.766e-07
I3670 0 n3671 3.361e-02A M=1.787e-06
I3671 0 n3672 3.361e-02A M=5.659e-07
I3672 0 n3673 3.361e-02A M=1.170e-06
I3673 0 n3674 3.361e-02A M=7.940e-07
I3674 0 n3675 3.361e-02A M=8.162e-07
I3675 0 n3676 3.361e-02A M=8.300e-07
I3676 0 n3677 3.361e-02A M=7.528e-07
I3677 0 n3678 3.361e-02A M=1.633e-06
I3678 0 n3679 3.361e-02A M=8.258e-07
I3679 0 n3680 3.361e-02A M=1.171e-06
I3680 0 n3681 3.361e-02A M=6.355e-07
I3681 0 n3682 3.361e-02A M=3.364e-07
I3682 0 n3683 3.361e-02A M=2.264e-07
I3683 0 n3684 3.361e-02A M=7.555e-07
I3684 0 n3685 3.361e-02A M=1.155e-06
I3685 0 n3686 3.361e-02A M=2.897e-07
I3686 0 n3687 3.361e-02A M=6.324e-07
I3687 0 n3688 3.361e-02A M=2.077e-07
I3688 0 n3689 3.361e-02A M=1.111e-06
I3689 0 n3690 3.361e-02A M=8.593e-07
I3690 0 n3691 3.361e-02A M=1.691e-06
I3691 0 n3692 3.361e-02A M=3.398e-07
I3692 0 n3693 3.361e-02A M=1.509e-06
I3693 0 n3694 3.361e-02A M=8.456e-07
I3694 0 n3695 3.361e-02A M=1.476e-06
I3695 0 n3696 3.361e-02A M=2.403e-06
I3696 0 n3697 3.361e-02A M=1.030e-06
I3697 0 n3698 3.361e-02A M=2.367e-07
I3698 0 n3699 3.361e-02A M=9.434e-07
I3699 0 n3700 3.361e-02A M=7.311e-07
I3700 0 n3701 3.361e-02A M=8.188e-07
I3701 0 n3702 3.361e-02A M=4.997e-07
I3702 0 n3703 3.361e-02A M=1.271e-06
I3703 0 n3704 3.361e-02A M=6.334e-07
I3704 0 n3705 3.361e-02A M=1.029e-06
I3705 0 n3706 3.361e-02A M=3.424e-07
I3706 0 n3707 3.361e-02A M=8.759e-07
I3707 0 n3708 3.361e-02A M=6.741e-07
I3708 0 n3709 3.361e-02A M=2.050e-06
I3709 0 n3710 3.361e-02A M=8.945e-07
I3710 0 n3711 3.361e-02A M=9.582e-07
I3711 0 n3712 3.361e-02A M=8.029e-07
I3712 0 n3713 3.361e-02A M=1.159e-06
I3713 0 n3714 3.361e-02A M=5.949e-07
I3714 0 n3715 3.361e-02A M=2.587e-06
I3715 0 n3716 3.361e-02A M=1.456e-06
I3716 0 n3717 3.361e-02A M=2.625e-07
I3717 0 n3718 3.361e-02A M=2.430e-06
I3718 0 n3719 3.361e-02A M=7.714e-07
I3719 0 n3720 3.361e-02A M=8.536e-07
I3720 0 n3721 3.361e-02A M=2.497e-06
I3721 0 n3722 3.361e-02A M=5.500e-07
I3722 0 n3723 3.361e-02A M=1.118e-06
I3723 0 n3724 3.361e-02A M=1.922e-06
I3724 0 n3725 3.361e-02A M=4.843e-07
I3725 0 n3726 3.361e-02A M=1.442e-06
I3726 0 n3727 3.361e-02A M=1.487e-06
I3727 0 n3728 3.361e-02A M=4.958e-07
I3728 0 n3729 3.361e-02A M=8.478e-07
I3729 0 n3730 3.361e-02A M=7.523e-07
I3730 0 n3731 3.361e-02A M=1.085e-06
I3731 0 n3732 3.361e-02A M=6.988e-07
I3732 0 n3733 3.361e-02A M=6.509e-07
I3733 0 n3734 3.361e-02A M=2.483e-06
I3734 0 n3735 3.361e-02A M=1.758e-06
I3735 0 n3736 3.361e-02A M=9.130e-07
I3736 0 n3737 3.361e-02A M=4.440e-07
I3737 0 n3738 3.361e-02A M=9.703e-07
I3738 0 n3739 3.361e-02A M=6.794e-07
I3739 0 n3740 3.361e-02A M=5.190e-07
I3740 0 n3741 3.361e-02A M=1.230e-06
I3741 0 n3742 3.361e-02A M=1.347e-06
I3742 0 n3743 3.361e-02A M=2.322e-07
I3743 0 n3744 3.361e-02A M=3.729e-07
I3744 0 n3745 3.361e-02A M=7.807e-07
I3745 0 n3746 3.361e-02A M=5.555e-07
I3746 0 n3747 3.361e-02A M=1.194e-06
I3747 0 n3748 3.361e-02A M=1.160e-06
I3748 0 n3749 3.361e-02A M=2.453e-06
I3749 0 n3750 3.361e-02A M=6.547e-07
I3750 0 n3751 3.361e-02A M=1.437e-07
I3751 0 n3752 3.361e-02A M=1.727e-06
I3752 0 n3753 3.361e-02A M=1.105e-06
I3753 0 n3754 3.361e-02A M=1.151e-06
I3754 0 n3755 3.361e-02A M=7.075e-07
I3755 0 n3756 3.361e-02A M=4.709e-07
I3756 0 n3757 3.361e-02A M=6.466e-07
I3757 0 n3758 3.361e-02A M=9.032e-07
I3758 0 n3759 3.361e-02A M=1.097e-06
I3759 0 n3760 3.361e-02A M=4.878e-07
I3760 0 n3761 3.361e-02A M=1.006e-06
I3761 0 n3762 3.361e-02A M=6.838e-07
I3762 0 n3763 3.361e-02A M=1.582e-06
I3763 0 n3764 3.361e-02A M=7.305e-07
I3764 0 n3765 3.361e-02A M=3.445e-07
I3765 0 n3766 3.361e-02A M=3.228e-07
I3766 0 n3767 3.361e-02A M=1.579e-06
I3767 0 n3768 3.361e-02A M=1.870e-06
I3768 0 n3769 3.361e-02A M=1.546e-06
I3769 0 n3770 3.361e-02A M=1.247e-06
I3770 0 n3771 3.361e-02A M=5.771e-07
I3771 0 n3772 3.361e-02A M=8.279e-07
I3772 0 n3773 3.361e-02A M=6.017e-07
I3773 0 n3774 3.361e-02A M=1.147e-06
I3774 0 n3775 3.361e-02A M=2.479e-06
I3775 0 n3776 3.361e-02A M=1.225e-06
I3776 0 n3777 3.361e-02A M=3.666e-06
I3777 0 n3778 3.361e-02A M=1.502e-06
I3778 0 n3779 3.361e-02A M=4.181e-07
I3779 0 n3780 3.361e-02A M=1.308e-06
I3780 0 n3781 3.361e-02A M=2.553e-06
I3781 0 n3782 3.361e-02A M=1.705e-06
I3782 0 n3783 3.361e-02A M=6.911e-07
I3783 0 n3784 3.361e-02A M=1.318e-06
I3784 0 n3785 3.361e-02A M=1.251e-06
I3785 0 n3786 3.361e-02A M=1.960e-06
I3786 0 n3787 3.361e-02A M=2.378e-06
I3787 0 n3788 3.361e-02A M=8.510e-07
I3788 0 n3789 3.361e-02A M=7.216e-07
I3789 0 n3790 3.361e-02A M=1.877e-07
I3790 0 n3791 3.361e-02A M=4.995e-07
I3791 0 n3792 3.361e-02A M=2.938e-06
I3792 0 n3793 3.361e-02A M=1.545e-06
I3793 0 n3794 3.361e-02A M=1.158e-06
I3794 0 n3795 3.361e-02A M=9.355e-07
I3795 0 n3796 3.361e-02A M=7.078e-07
I3796 0 n3797 3.361e-02A M=1.438e-06
I3797 0 n3798 3.361e-02A M=9.696e-07
I3798 0 n3799 3.361e-02A M=2.716e-06
I3799 0 n3800 3.361e-02A M=1.022e-06
I3800 0 n3801 3.361e-02A M=1.447e-06
I3801 0 n3802 3.361e-02A M=7.202e-07
I3802 0 n3803 3.361e-02A M=1.342e-06
I3803 0 n3804 3.361e-02A M=1.302e-06
I3804 0 n3805 3.361e-02A M=5.343e-07
I3805 0 n3806 3.361e-02A M=1.045e-07
I3806 0 n3807 3.361e-02A M=1.800e-06
I3807 0 n3808 3.361e-02A M=1.811e-06
I3808 0 n3809 3.361e-02A M=3.795e-07
I3809 0 n3810 3.361e-02A M=1.179e-06
I3810 0 n3811 3.361e-02A M=1.098e-06
I3811 0 n3812 3.361e-02A M=7.647e-07
I3812 0 n3813 3.361e-02A M=5.347e-07
I3813 0 n3814 3.361e-02A M=1.030e-06
I3814 0 n3815 3.361e-02A M=1.066e-06
I3815 0 n3816 3.361e-02A M=2.039e-07
I3816 0 n3817 3.361e-02A M=4.828e-07
I3817 0 n3818 3.361e-02A M=2.026e-06
I3818 0 n3819 3.361e-02A M=1.570e-06
I3819 0 n3820 3.361e-02A M=8.063e-07
I3820 0 n3821 3.361e-02A M=1.157e-06
I3821 0 n3822 3.361e-02A M=4.548e-07
I3822 0 n3823 3.361e-02A M=4.584e-07
I3823 0 n3824 3.361e-02A M=2.085e-06
I3824 0 n3825 3.361e-02A M=1.605e-06
I3825 0 n3826 3.361e-02A M=4.210e-07
I3826 0 n3827 3.361e-02A M=9.730e-07
I3827 0 n3828 3.361e-02A M=8.246e-07
I3828 0 n3829 3.361e-02A M=9.755e-07
I3829 0 n3830 3.361e-02A M=9.656e-07
I3830 0 n3831 3.361e-02A M=8.125e-07
I3831 0 n3832 3.361e-02A M=1.443e-06
I3832 0 n3833 3.361e-02A M=6.724e-07
I3833 0 n3834 3.361e-02A M=3.696e-07
I3834 0 n3835 3.361e-02A M=8.609e-07
I3835 0 n3836 3.361e-02A M=1.286e-06
I3836 0 n3837 3.361e-02A M=1.003e-06
I3837 0 n3838 3.361e-02A M=1.209e-06
I3838 0 n3839 3.361e-02A M=5.160e-07
I3839 0 n3840 3.361e-02A M=9.438e-07
I3840 0 n3841 3.361e-02A M=5.285e-07
I3841 0 n3842 3.361e-02A M=9.412e-07
I3842 0 n3843 3.361e-02A M=5.619e-07
I3843 0 n3844 3.361e-02A M=6.681e-07
I3844 0 n3845 3.361e-02A M=7.623e-07
I3845 0 n3846 3.361e-02A M=3.175e-07
I3846 0 n3847 3.361e-02A M=1.671e-06
I3847 0 n3848 3.361e-02A M=8.044e-07
I3848 0 n3849 3.361e-02A M=1.320e-06
I3849 0 n3850 3.361e-02A M=1.322e-06
I3850 0 n3851 3.361e-02A M=1.278e-06
I3851 0 n3852 3.361e-02A M=3.744e-07
I3852 0 n3853 3.361e-02A M=8.123e-07
I3853 0 n3854 3.361e-02A M=1.884e-06
I3854 0 n3855 3.361e-02A M=1.474e-06
I3855 0 n3856 3.361e-02A M=5.409e-07
I3856 0 n3857 3.361e-02A M=9.930e-07
I3857 0 n3858 3.361e-02A M=6.365e-07
I3858 0 n3859 3.361e-02A M=3.776e-08
I3859 0 n3860 3.361e-02A M=3.613e-07
I3860 0 n3861 3.361e-02A M=8.328e-07
I3861 0 n3862 3.361e-02A M=1.127e-06
I3862 0 n3863 3.361e-02A M=2.099e-07
I3863 0 n3864 3.361e-02A M=5.383e-07
I3864 0 n3865 3.361e-02A M=1.315e-06
I3865 0 n3866 3.361e-02A M=1.629e-06
I3866 0 n3867 3.361e-02A M=3.564e-07
I3867 0 n3868 3.361e-02A M=1.356e-06
I3868 0 n3869 3.361e-02A M=1.950e-06
I3869 0 n3870 3.361e-02A M=9.083e-07
I3870 0 n3871 3.361e-02A M=9.430e-07
I3871 0 n3872 3.361e-02A M=2.075e-06
I3872 0 n3873 3.361e-02A M=1.049e-06
I3873 0 n3874 3.361e-02A M=1.628e-06
I3874 0 n3875 3.361e-02A M=8.192e-07
I3875 0 n3876 3.361e-02A M=1.089e-06
I3876 0 n3877 3.361e-02A M=9.792e-07
I3877 0 n3878 3.361e-02A M=8.124e-07
I3878 0 n3879 3.361e-02A M=6.025e-07
I3879 0 n3880 3.361e-02A M=8.938e-07
I3880 0 n3881 3.361e-02A M=7.428e-07
I3881 0 n3882 3.361e-02A M=7.821e-07
I3882 0 n3883 3.361e-02A M=1.380e-06
I3883 0 n3884 3.361e-02A M=1.034e-06
I3884 0 n3885 3.361e-02A M=2.630e-07
I3885 0 n3886 3.361e-02A M=1.012e-06
I3886 0 n3887 3.361e-02A M=6.967e-07
I3887 0 n3888 3.361e-02A M=4.540e-07
I3888 0 n3889 3.361e-02A M=6.820e-07
I3889 0 n3890 3.361e-02A M=4.847e-07
I3890 0 n3891 3.361e-02A M=1.088e-06
I3891 0 n3892 3.361e-02A M=7.831e-07
I3892 0 n3893 3.361e-02A M=7.094e-07
I3893 0 n3894 3.361e-02A M=6.013e-07
I3894 0 n3895 3.361e-02A M=5.032e-07
I3895 0 n3896 3.361e-02A M=1.083e-06
I3896 0 n3897 3.361e-02A M=6.876e-07
I3897 0 n3898 3.361e-02A M=9.702e-07
I3898 0 n3899 3.361e-02A M=1.018e-06
I3899 0 n3900 3.361e-02A M=1.779e-06
I3900 0 n3901 3.361e-02A M=1.252e-06
I3901 0 n3902 3.361e-02A M=1.160e-06
I3902 0 n3903 3.361e-02A M=1.187e-06
I3903 0 n3904 3.361e-02A M=1.442e-06
I3904 0 n3905 3.361e-02A M=2.253e-07
I3905 0 n3906 3.361e-02A M=7.124e-07
I3906 0 n3907 3.361e-02A M=3.710e-07
I3907 0 n3908 3.361e-02A M=9.550e-07
I3908 0 n3909 3.361e-02A M=5.417e-07
I3909 0 n3910 3.361e-02A M=6.207e-07
I3910 0 n3911 3.361e-02A M=5.088e-07
I3911 0 n3912 3.361e-02A M=7.641e-07
I3912 0 n3913 3.361e-02A M=2.786e-07
I3913 0 n3914 3.361e-02A M=6.048e-07
I3914 0 n3915 3.361e-02A M=5.120e-07
I3915 0 n3916 3.361e-02A M=2.000e-06
I3916 0 n3917 3.361e-02A M=9.889e-07
I3917 0 n3918 3.361e-02A M=9.928e-07
I3918 0 n3919 3.361e-02A M=7.103e-07
I3919 0 n3920 3.361e-02A M=1.135e-06
I3920 0 n3921 3.361e-02A M=6.284e-07
I3921 0 n3922 3.361e-02A M=1.019e-06
I3922 0 n3923 3.361e-02A M=8.489e-07
I3923 0 n3924 3.361e-02A M=1.004e-06
I3924 0 n3925 3.361e-02A M=1.484e-06
I3925 0 n3926 3.361e-02A M=8.006e-07
I3926 0 n3927 3.361e-02A M=6.419e-07
I3927 0 n3928 3.361e-02A M=3.753e-07
I3928 0 n3929 3.361e-02A M=5.239e-07
I3929 0 n3930 3.361e-02A M=2.094e-06
I3930 0 n3931 3.361e-02A M=9.051e-07
I3931 0 n3932 3.361e-02A M=3.897e-07
I3932 0 n3933 3.361e-02A M=2.878e-06
I3933 0 n3934 3.361e-02A M=1.507e-06
I3934 0 n3935 3.361e-02A M=9.366e-07
I3935 0 n3936 3.361e-02A M=6.612e-07
I3936 0 n3937 3.361e-02A M=1.956e-06
I3937 0 n3938 3.361e-02A M=1.135e-06
I3938 0 n3939 3.361e-02A M=1.520e-07
I3939 0 n3940 3.361e-02A M=1.601e-06
I3940 0 n3941 3.361e-02A M=8.622e-07
I3941 0 n3942 3.361e-02A M=1.365e-06
I3942 0 n3943 3.361e-02A M=4.352e-07
I3943 0 n3944 3.361e-02A M=1.051e-06
I3944 0 n3945 3.361e-02A M=9.823e-07
I3945 0 n3946 3.361e-02A M=2.581e-06
I3946 0 n3947 3.361e-02A M=7.096e-07
I3947 0 n3948 3.361e-02A M=1.792e-06
I3948 0 n3949 3.361e-02A M=3.447e-07
I3949 0 n3950 3.361e-02A M=2.303e-06
I3950 0 n3951 3.361e-02A M=1.836e-07
I3951 0 n1 3.361e-02A M=1.134e-06
I3952 0 n3953 3.361e-02A M=1.525e-06
I3953 0 n3954 3.361e-02A M=1.255e-06
I3954 0 n3955 3.361e-02A M=8.089e-07
I3955 0 n3956 3.361e-02A M=1.139e-06
I3956 0 n3957 3.361e-02A M=1.695e-06
I3957 0 n3958 3.361e-02A M=9.380e-07
I3958 0 n3959 3.361e-02A M=1.450e-06
I3959 0 n3960 3.361e-02A M=1.646e-06
I3960 0 n3961 3.361e-02A M=4.707e-07
I3961 0 n3962 3.361e-02A M=1.263e-06
I3962 0 n3963 3.361e-02A M=1.187e-06
I3963 0 n3964 3.361e-02A M=9.064e-07
I3964 0 n3965 3.361e-02A M=1.630e-06
I3965 0 n3966 3.361e-02A M=5.200e-07
I3966 0 n3967 3.361e-02A M=1.685e-06
I3967 0 n3968 3.361e-02A M=8.600e-07
I3968 0 n3969 3.361e-02A M=7.040e-07
I3969 0 n3970 3.361e-02A M=2.497e-06
I3970 0 n3971 3.361e-02A M=8.638e-07
I3971 0 n3972 3.361e-02A M=1.522e-06
I3972 0 n3973 3.361e-02A M=7.603e-07
I3973 0 n3974 3.361e-02A M=1.736e-06
I3974 0 n3975 3.361e-02A M=1.195e-06
I3975 0 n3976 3.361e-02A M=9.135e-07
I3976 0 n3977 3.361e-02A M=3.964e-07
I3977 0 n3978 3.361e-02A M=1.853e-07
I3978 0 n3979 3.361e-02A M=1.893e-06
I3979 0 n3980 3.361e-02A M=5.427e-07
I3980 0 n3981 3.361e-02A M=4.704e-07
I3981 0 n3982 3.361e-02A M=1.044e-06
I3982 0 n3983 3.361e-02A M=5.805e-07
I3983 0 n3984 3.361e-02A M=2.422e-06
I3984 0 n3985 3.361e-02A M=9.561e-07
I3985 0 n3986 3.361e-02A M=6.093e-07
I3986 0 n3987 3.361e-02A M=2.702e-06
I3987 0 n3988 3.361e-02A M=7.391e-07
I3988 0 n3989 3.361e-02A M=6.121e-07
I3989 0 n3990 3.361e-02A M=7.973e-07
I3990 0 n3991 3.361e-02A M=7.523e-07
I3991 0 n3992 3.361e-02A M=9.225e-07
I3992 0 n3993 3.361e-02A M=7.699e-07
I3993 0 n3994 3.361e-02A M=1.148e-07
I3994 0 n3995 3.361e-02A M=6.335e-07
I3995 0 n3996 3.361e-02A M=1.372e-06
I3996 0 n3997 3.361e-02A M=2.198e-06
I3997 0 n3998 3.361e-02A M=1.528e-06
I3998 0 n3999 3.361e-02A M=1.140e-06
I3999 0 n4000 3.361e-02A M=6.874e-07
I4000 0 n4001 3.361e-02A M=2.002e-07
I4001 0 n4002 3.361e-02A M=1.476e-06
I4002 0 n4003 3.361e-02A M=1.080e-06
I4003 0 n4004 3.361e-02A M=6.948e-07
I4004 0 n4005 3.361e-02A M=5.536e-07
I4005 0 n4006 3.361e-02A M=8.652e-07
I4006 0 n4007 3.361e-02A M=9.365e-07
I4007 0 n4008 3.361e-02A M=1.385e-06
I4008 0 n4009 3.361e-02A M=5.870e-07
I4009 0 n4010 3.361e-02A M=5.456e-07
I4010 0 n4011 3.361e-02A M=6.999e-07
I4011 0 n4012 3.361e-02A M=1.250e-06
I4012 0 n4013 3.361e-02A M=1.096e-06
I4013 0 n4014 3.361e-02A M=8.570e-07
I4014 0 n4015 3.361e-02A M=1.494e-06
I4015 0 n4016 3.361e-02A M=1.832e-06
I4016 0 n4017 3.361e-02A M=9.298e-07
I4017 0 n4018 3.361e-02A M=8.067e-07
I4018 0 n4019 3.361e-02A M=2.317e-07
I4019 0 n4020 3.361e-02A M=4.479e-07
I4020 0 n4021 3.361e-02A M=2.360e-06
I4021 0 n4022 3.361e-02A M=3.218e-06
I4022 0 n4023 3.361e-02A M=1.064e-06
I4023 0 n4024 3.361e-02A M=2.398e-06
I4024 0 n4025 3.361e-02A M=5.349e-07
I4025 0 n4026 3.361e-02A M=1.218e-06
I4026 0 n4027 3.361e-02A M=1.275e-06
I4027 0 n4028 3.361e-02A M=8.261e-07
I4028 0 n4029 3.361e-02A M=6.988e-07
I4029 0 n4030 3.361e-02A M=1.148e-06
I4030 0 n4031 3.361e-02A M=8.716e-07
I4031 0 n4032 3.361e-02A M=1.038e-06
I4032 0 n4033 3.361e-02A M=1.060e-06
I4033 0 n4034 3.361e-02A M=1.181e-06
I4034 0 n4035 3.361e-02A M=8.606e-07
I4035 0 n4036 3.361e-02A M=8.316e-07
I4036 0 n4037 3.361e-02A M=1.266e-06
I4037 0 n4038 3.361e-02A M=1.049e-06
I4038 0 n4039 3.361e-02A M=4.756e-07
I4039 0 n4040 3.361e-02A M=8.496e-07
I4040 0 n4041 3.361e-02A M=1.079e-06
I4041 0 n4042 3.361e-02A M=1.177e-06
I4042 0 n4043 3.361e-02A M=1.955e-06
I4043 0 n4044 3.361e-02A M=2.842e-07
I4044 0 n4045 3.361e-02A M=1.350e-06
I4045 0 n4046 3.361e-02A M=2.084e-06
I4046 0 n4047 3.361e-02A M=3.935e-07
I4047 0 n4048 3.361e-02A M=2.813e-06
I4048 0 n4049 3.361e-02A M=3.126e-07
I4049 0 n4050 3.361e-02A M=3.708e-07
I4050 0 n4051 3.361e-02A M=5.874e-07
I4051 0 n4052 3.361e-02A M=9.194e-07
I4052 0 n4053 3.361e-02A M=1.671e-06
I4053 0 n4054 3.361e-02A M=9.562e-07
I4054 0 n4055 3.361e-02A M=1.271e-06
I4055 0 n4056 3.361e-02A M=1.213e-06
I4056 0 n4057 3.361e-02A M=1.055e-06
I4057 0 n4058 3.361e-02A M=6.047e-07
I4058 0 n4059 3.361e-02A M=2.382e-06
I4059 0 n4060 3.361e-02A M=6.332e-07
I4060 0 n4061 3.361e-02A M=8.426e-07
I4061 0 n4062 3.361e-02A M=1.200e-06
I4062 0 n4063 3.361e-02A M=6.048e-07
I4063 0 n4064 3.361e-02A M=1.559e-06
I4064 0 n4065 3.361e-02A M=3.125e-07
I4065 0 n4066 3.361e-02A M=6.412e-07
I4066 0 n4067 3.361e-02A M=2.975e-07
I4067 0 n4068 3.361e-02A M=2.566e-06
I4068 0 n4069 3.361e-02A M=6.065e-07
I4069 0 n4070 3.361e-02A M=8.303e-07
I4070 0 n4071 3.361e-02A M=9.999e-07
I4071 0 n4072 3.361e-02A M=7.605e-07
I4072 0 n4073 3.361e-02A M=1.195e-06
I4073 0 n4074 3.361e-02A M=4.947e-07
I4074 0 n4075 3.361e-02A M=9.973e-07
I4075 0 n4076 3.361e-02A M=8.370e-07
I4076 0 n4077 3.361e-02A M=6.294e-07
I4077 0 n4078 3.361e-02A M=3.909e-07
I4078 0 n4079 3.361e-02A M=2.546e-06
I4079 0 n4080 3.361e-02A M=1.590e-06
I4080 0 n4081 3.361e-02A M=5.466e-07
I4081 0 n4082 3.361e-02A M=1.393e-06
I4082 0 n4083 3.361e-02A M=8.094e-07
I4083 0 n4084 3.361e-02A M=1.023e-06
I4084 0 n4085 3.361e-02A M=7.720e-07
I4085 0 n4086 3.361e-02A M=3.493e-07
I4086 0 n4087 3.361e-02A M=4.234e-07
I4087 0 n4088 3.361e-02A M=4.867e-07
I4088 0 n4089 3.361e-02A M=1.985e-06
I4089 0 n4090 3.361e-02A M=8.145e-07
I4090 0 n4091 3.361e-02A M=8.285e-07
I4091 0 n4092 3.361e-02A M=8.436e-07
I4092 0 n4093 3.361e-02A M=1.694e-06
I4093 0 n4094 3.361e-02A M=1.266e-06
I4094 0 n4095 3.361e-02A M=1.175e-06
I4095 0 n4096 3.361e-02A M=1.059e-06
I4096 0 n4097 3.361e-02A M=2.293e-06
I4097 0 n4098 3.361e-02A M=9.917e-07
I4098 0 n4099 3.361e-02A M=7.242e-07
I4099 0 n4100 3.361e-02A M=5.620e-07
I4100 0 n4101 3.361e-02A M=1.446e-06
I4101 0 n4102 3.361e-02A M=4.386e-07
I4102 0 n4103 3.361e-02A M=1.455e-06
I4103 0 n4104 3.361e-02A M=3.738e-07
I4104 0 n4105 3.361e-02A M=1.385e-06
I4105 0 n4106 3.361e-02A M=2.057e-06
I4106 0 n4107 3.361e-02A M=1.107e-06
I4107 0 n4108 3.361e-02A M=1.026e-06
I4108 0 n4109 3.361e-02A M=7.103e-07
I4109 0 n4110 3.361e-02A M=1.404e-06
I4110 0 n4111 3.361e-02A M=3.599e-07
I4111 0 n4112 3.361e-02A M=1.140e-06
I4112 0 n4113 3.361e-02A M=7.060e-07
I4113 0 n4114 3.361e-02A M=1.449e-06
I4114 0 n4115 3.361e-02A M=1.106e-06
I4115 0 n4116 3.361e-02A M=1.291e-06
I4116 0 n4117 3.361e-02A M=1.313e-06
I4117 0 n4118 3.361e-02A M=3.748e-07
I4118 0 n4119 3.361e-02A M=3.540e-07
I4119 0 n4120 3.361e-02A M=1.944e-06
I4120 0 n4121 3.361e-02A M=1.339e-06
I4121 0 n4122 3.361e-02A M=4.032e-07
I4122 0 n4123 3.361e-02A M=1.115e-06
I4123 0 n4124 3.361e-02A M=3.487e-07
I4124 0 n4125 3.361e-02A M=1.120e-06
I4125 0 n4126 3.361e-02A M=1.135e-06
I4126 0 n4127 3.361e-02A M=4.728e-07
I4127 0 n4128 3.361e-02A M=8.735e-07
I4128 0 n4129 3.361e-02A M=1.837e-06
I4129 0 n4130 3.361e-02A M=2.166e-06
I4130 0 n4131 3.361e-02A M=1.690e-06
I4131 0 n4132 3.361e-02A M=5.911e-07
I4132 0 n4133 3.361e-02A M=3.983e-07
I4133 0 n4134 3.361e-02A M=7.826e-07
I4134 0 n4135 3.361e-02A M=1.827e-06
I4135 0 n4136 3.361e-02A M=3.929e-07
I4136 0 n4137 3.361e-02A M=1.211e-06
I4137 0 n4138 3.361e-02A M=2.087e-06
I4138 0 n4139 3.361e-02A M=2.578e-06
I4139 0 n4140 3.361e-02A M=4.896e-07
I4140 0 n4141 3.361e-02A M=1.103e-06
I4141 0 n4142 3.361e-02A M=7.332e-07
I4142 0 n4143 3.361e-02A M=1.459e-06
I4143 0 n4144 3.361e-02A M=2.489e-06
I4144 0 n4145 3.361e-02A M=5.223e-07
I4145 0 n4146 3.361e-02A M=5.902e-07
I4146 0 n4147 3.361e-02A M=1.363e-06
I4147 0 n4148 3.361e-02A M=1.919e-06
I4148 0 n4149 3.361e-02A M=6.256e-07
I4149 0 n4150 3.361e-02A M=1.422e-06
I4150 0 n4151 3.361e-02A M=1.244e-06
I4151 0 n4152 3.361e-02A M=6.705e-07
I4152 0 n4153 3.361e-02A M=1.623e-06
I4153 0 n4154 3.361e-02A M=8.136e-07
I4154 0 n4155 3.361e-02A M=1.255e-06
I4155 0 n4156 3.361e-02A M=6.143e-07
I4156 0 n4157 3.361e-02A M=9.150e-07
I4157 0 n4158 3.361e-02A M=9.773e-07
I4158 0 n4159 3.361e-02A M=1.884e-06
I4159 0 n4160 3.361e-02A M=2.920e-07
I4160 0 n4161 3.361e-02A M=5.072e-07
I4161 0 n4162 3.361e-02A M=5.440e-07
I4162 0 n4163 3.361e-02A M=1.707e-06
I4163 0 n4164 3.361e-02A M=7.917e-07
I4164 0 n4165 3.361e-02A M=2.480e-06
I4165 0 n4166 3.361e-02A M=7.679e-07
I4166 0 n4167 3.361e-02A M=8.071e-07
I4167 0 n4168 3.361e-02A M=5.845e-07
I4168 0 n4169 3.361e-02A M=1.159e-06
I4169 0 n4170 3.361e-02A M=7.948e-07
I4170 0 n4171 3.361e-02A M=9.418e-07
I4171 0 n4172 3.361e-02A M=1.059e-06
I4172 0 n4173 3.361e-02A M=6.433e-07
I4173 0 n4174 3.361e-02A M=9.255e-07
I4174 0 n4175 3.361e-02A M=1.313e-06
I4175 0 n4176 3.361e-02A M=9.170e-07
I4176 0 n4177 3.361e-02A M=7.866e-07
I4177 0 n4178 3.361e-02A M=8.215e-07
I4178 0 n4179 3.361e-02A M=1.591e-06
I4179 0 n4180 3.361e-02A M=3.525e-07
I4180 0 n4181 3.361e-02A M=8.303e-07
I4181 0 n4182 3.361e-02A M=4.523e-07
I4182 0 n4183 3.361e-02A M=4.228e-07
I4183 0 n4184 3.361e-02A M=9.439e-07
I4184 0 n4185 3.361e-02A M=1.109e-06
I4185 0 n4186 3.361e-02A M=5.079e-07
I4186 0 n4187 3.361e-02A M=8.967e-07
I4187 0 n4188 3.361e-02A M=8.215e-07
I4188 0 n4189 3.361e-02A M=6.405e-07
I4189 0 n1 3.361e-02A M=1.048e-06
I4190 0 n4191 3.361e-02A M=9.232e-07
I4191 0 n4192 3.361e-02A M=1.488e-06
I4192 0 n4193 3.361e-02A M=1.138e-06
I4193 0 n4194 3.361e-02A M=1.069e-06
I4194 0 n4195 3.361e-02A M=1.183e-07
I4195 0 n4196 3.361e-02A M=2.495e-06
I4196 0 n4197 3.361e-02A M=4.611e-07
I4197 0 n4198 3.361e-02A M=5.078e-07
I4198 0 n4199 3.361e-02A M=1.599e-06
I4199 0 n4200 3.361e-02A M=8.638e-07
I4200 0 n4201 3.361e-02A M=6.423e-07
I4201 0 n4202 3.361e-02A M=6.893e-07
I4202 0 n4203 3.361e-02A M=7.532e-07
I4203 0 n4204 3.361e-02A M=5.643e-07
I4204 0 n4205 3.361e-02A M=1.390e-06
I4205 0 n4206 3.361e-02A M=4.057e-07
I4206 0 n4207 3.361e-02A M=5.832e-07
I4207 0 n4208 3.361e-02A M=4.457e-07
I4208 0 n4209 3.361e-02A M=2.666e-07
I4209 0 n4210 3.361e-02A M=9.526e-07
I4210 0 n4211 3.361e-02A M=2.191e-06
I4211 0 n4212 3.361e-02A M=1.060e-06
I4212 0 n4213 3.361e-02A M=7.373e-07
I4213 0 n4214 3.361e-02A M=4.472e-07
I4214 0 n4215 3.361e-02A M=3.838e-07
I4215 0 n4216 3.361e-02A M=2.414e-06
I4216 0 n4217 3.361e-02A M=8.533e-07
I4217 0 n4218 3.361e-02A M=7.939e-07
I4218 0 n4219 3.361e-02A M=1.650e-06
I4219 0 n4220 3.361e-02A M=6.948e-07
I4220 0 n4221 3.361e-02A M=5.896e-07
I4221 0 n4222 3.361e-02A M=9.310e-07
I4222 0 n4223 3.361e-02A M=3.161e-07
I4223 0 n4224 3.361e-02A M=5.248e-07
I4224 0 n4225 3.361e-02A M=1.365e-06
I4225 0 n4226 3.361e-02A M=6.717e-07
I4226 0 n4227 3.361e-02A M=1.635e-07
I4227 0 n4228 3.361e-02A M=9.423e-07
I4228 0 n4229 3.361e-02A M=7.847e-07
I4229 0 n4230 3.361e-02A M=1.110e-06
I4230 0 n4231 3.361e-02A M=8.525e-07
I4231 0 n4232 3.361e-02A M=1.025e-06
I4232 0 n4233 3.361e-02A M=4.814e-07
I4233 0 n4234 3.361e-02A M=4.058e-07
I4234 0 n4235 3.361e-02A M=1.738e-06
I4235 0 n4236 3.361e-02A M=8.729e-07
I4236 0 n4237 3.361e-02A M=6.838e-07
I4237 0 n4238 3.361e-02A M=2.495e-06
I4238 0 n4239 3.361e-02A M=8.585e-07
I4239 0 n4240 3.361e-02A M=1.069e-06
I4240 0 n4241 3.361e-02A M=1.140e-06
I4241 0 n4242 3.361e-02A M=8.617e-07
I4242 0 n4243 3.361e-02A M=2.667e-07
I4243 0 n4244 3.361e-02A M=3.775e-07
I4244 0 n4245 3.361e-02A M=8.489e-07
I4245 0 n4246 3.361e-02A M=8.519e-07
I4246 0 n4247 3.361e-02A M=8.189e-07
I4247 0 n4248 3.361e-02A M=6.930e-07
I4248 0 n4249 3.361e-02A M=1.373e-06
I4249 0 n4250 3.361e-02A M=8.628e-07
I4250 0 n4251 3.361e-02A M=9.185e-07
I4251 0 n4252 3.361e-02A M=1.102e-06
I4252 0 n4253 3.361e-02A M=4.924e-07
I4253 0 n4254 3.361e-02A M=5.864e-07
I4254 0 n4255 3.361e-02A M=1.413e-06
I4255 0 n4256 3.361e-02A M=1.292e-06
I4256 0 n4257 3.361e-02A M=4.708e-07
I4257 0 n4258 3.361e-02A M=7.233e-07
I4258 0 n4259 3.361e-02A M=1.170e-06
I4259 0 n4260 3.361e-02A M=9.257e-07
I4260 0 n4261 3.361e-02A M=1.796e-06
I4261 0 n4262 3.361e-02A M=1.851e-06
I4262 0 n4263 3.361e-02A M=1.084e-06
I4263 0 n4264 3.361e-02A M=6.369e-07
I4264 0 n4265 3.361e-02A M=7.541e-07
I4265 0 n4266 3.361e-02A M=1.747e-06
I4266 0 n4267 3.361e-02A M=1.829e-07
I4267 0 n4268 3.361e-02A M=6.147e-07
I4268 0 n4269 3.361e-02A M=1.382e-06
I4269 0 n4270 3.361e-02A M=1.043e-06
I4270 0 n4271 3.361e-02A M=6.632e-07
I4271 0 n4272 3.361e-02A M=2.035e-06
I4272 0 n4273 3.361e-02A M=8.499e-07
I4273 0 n4274 3.361e-02A M=1.730e-06
I4274 0 n4275 3.361e-02A M=1.061e-06
I4275 0 n4276 3.361e-02A M=3.174e-07
I4276 0 n4277 3.361e-02A M=9.379e-07
I4277 0 n4278 3.361e-02A M=1.003e-06
I4278 0 n4279 3.361e-02A M=1.464e-06
I4279 0 n4280 3.361e-02A M=7.483e-07
I4280 0 n4281 3.361e-02A M=1.687e-06
I4281 0 n4282 3.361e-02A M=1.092e-06
I4282 0 n4283 3.361e-02A M=8.773e-07
I4283 0 n4284 3.361e-02A M=9.578e-07
I4284 0 n4285 3.361e-02A M=1.307e-06
I4285 0 n4286 3.361e-02A M=3.727e-07
I4286 0 n4287 3.361e-02A M=2.431e-07
I4287 0 n4288 3.361e-02A M=1.487e-06
I4288 0 n4289 3.361e-02A M=3.472e-07
I4289 0 n4290 3.361e-02A M=8.070e-07
I4290 0 n4291 3.361e-02A M=1.004e-06
I4291 0 n4292 3.361e-02A M=1.109e-06
I4292 0 n4293 3.361e-02A M=1.617e-06
I4293 0 n4294 3.361e-02A M=3.929e-07
I4294 0 n4295 3.361e-02A M=1.030e-06
I4295 0 n4296 3.361e-02A M=9.951e-07
I4296 0 n4297 3.361e-02A M=3.791e-07
I4297 0 n4298 3.361e-02A M=5.411e-07
I4298 0 n4299 3.361e-02A M=3.892e-07
I4299 0 n4300 3.361e-02A M=1.971e-06
I4300 0 n4301 3.361e-02A M=1.276e-06
I4301 0 n4302 3.361e-02A M=1.726e-06
I4302 0 n4303 3.361e-02A M=1.181e-06
I4303 0 n4304 3.361e-02A M=1.665e-06
I4304 0 n4305 3.361e-02A M=1.452e-06
I4305 0 n4306 3.361e-02A M=2.394e-07
I4306 0 n4307 3.361e-02A M=5.411e-07
I4307 0 n4308 3.361e-02A M=8.108e-07
I4308 0 n4309 3.361e-02A M=5.124e-07
I4309 0 n4310 3.361e-02A M=1.016e-06
I4310 0 n4311 3.361e-02A M=1.096e-06
I4311 0 n4312 3.361e-02A M=7.745e-07
I4312 0 n4313 3.361e-02A M=1.343e-06
I4313 0 n4314 3.361e-02A M=1.650e-06
I4314 0 n4315 3.361e-02A M=2.876e-06
I4315 0 n4316 3.361e-02A M=1.062e-06
I4316 0 n4317 3.361e-02A M=6.877e-07
I4317 0 n4318 3.361e-02A M=5.937e-07
I4318 0 n4319 3.361e-02A M=7.740e-07
I4319 0 n4320 3.361e-02A M=6.598e-07
I4320 0 n4321 3.361e-02A M=3.790e-07
I4321 0 n4322 3.361e-02A M=5.738e-07
I4322 0 n4323 3.361e-02A M=2.108e-06
I4323 0 n4324 3.361e-02A M=5.369e-07
I4324 0 n4325 3.361e-02A M=1.344e-06
I4325 0 n4326 3.361e-02A M=8.138e-07
I4326 0 n4327 3.361e-02A M=1.313e-06
I4327 0 n4328 3.361e-02A M=8.785e-07
I4328 0 n4329 3.361e-02A M=7.887e-07
I4329 0 n4330 3.361e-02A M=1.709e-06
I4330 0 n1 3.361e-02A M=4.818e-07
I4331 0 n1 3.361e-02A M=8.180e-07
I4332 0 n4333 3.361e-02A M=6.799e-07
I4333 0 n4334 3.361e-02A M=1.051e-06
I4334 0 n4335 3.361e-02A M=5.873e-07
I4335 0 n4336 3.361e-02A M=1.073e-06
I4336 0 n4337 3.361e-02A M=7.384e-07
I4337 0 n4338 3.361e-02A M=1.312e-06
I4338 0 n1 3.361e-02A M=7.876e-07
I4339 0 n4340 3.361e-02A M=5.262e-07
I4340 0 n4341 3.361e-02A M=7.622e-07
I4341 0 n4342 3.361e-02A M=4.644e-07
I4342 0 n4343 3.361e-02A M=2.045e-06
I4343 0 n4344 3.361e-02A M=3.291e-06
I4344 0 n4345 3.361e-02A M=1.273e-06
I4345 0 n4346 3.361e-02A M=1.505e-06
I4346 0 n4347 3.361e-02A M=9.687e-07
I4347 0 n4348 3.361e-02A M=3.825e-07
I4348 0 n4349 3.361e-02A M=6.595e-07
I4349 0 n4350 3.361e-02A M=3.473e-07
I4350 0 n4351 3.361e-02A M=8.975e-07
I4351 0 n4352 3.361e-02A M=1.182e-06
I4352 0 n4353 3.361e-02A M=1.262e-06
I4353 0 n4354 3.361e-02A M=2.211e-06
I4354 0 n4355 3.361e-02A M=2.060e-06
I4355 0 n4356 3.361e-02A M=3.707e-07
I4356 0 n4357 3.361e-02A M=8.471e-07
I4357 0 n4358 3.361e-02A M=7.446e-07
I4358 0 n4359 3.361e-02A M=5.947e-07
I4359 0 n4360 3.361e-02A M=1.389e-06
I4360 0 n4361 3.361e-02A M=1.093e-06
I4361 0 n4362 3.361e-02A M=8.821e-07
I4362 0 n4363 3.361e-02A M=2.226e-06
I4363 0 n4364 3.361e-02A M=2.440e-06
I4364 0 n4365 3.361e-02A M=8.322e-07
I4365 0 n4366 3.361e-02A M=6.755e-07
I4366 0 n4367 3.361e-02A M=1.184e-06
I4367 0 n4368 3.361e-02A M=1.377e-06
I4368 0 n4369 3.361e-02A M=4.658e-07
I4369 0 n4370 3.361e-02A M=9.097e-07
I4370 0 n4371 3.361e-02A M=6.594e-07
I4371 0 n4372 3.361e-02A M=6.060e-07
I4372 0 n4373 3.361e-02A M=1.410e-06
I4373 0 n4374 3.361e-02A M=6.746e-07
I4374 0 n4375 3.361e-02A M=1.179e-06
I4375 0 n4376 3.361e-02A M=1.530e-06
I4376 0 n4377 3.361e-02A M=2.051e-07
I4377 0 n4378 3.361e-02A M=8.812e-07
I4378 0 n4379 3.361e-02A M=2.603e-06
I4379 0 n4380 3.361e-02A M=4.134e-07
I4380 0 n4381 3.361e-02A M=1.151e-06
I4381 0 n4382 3.361e-02A M=7.858e-07
I4382 0 n4383 3.361e-02A M=8.157e-07
I4383 0 n4384 3.361e-02A M=1.006e-06
I4384 0 n4385 3.361e-02A M=7.641e-07
I4385 0 n1 3.361e-02A M=7.157e-07
I4386 0 n4387 3.361e-02A M=1.172e-06
I4387 0 n4388 3.361e-02A M=7.395e-07
I4388 0 n4389 3.361e-02A M=7.918e-07
I4389 0 n4390 3.361e-02A M=1.484e-06
I4390 0 n4391 3.361e-02A M=1.088e-06
I4391 0 n4392 3.361e-02A M=2.196e-06
I4392 0 n4393 3.361e-02A M=2.890e-06
I4393 0 n4394 3.361e-02A M=1.694e-06
I4394 0 n4395 3.361e-02A M=4.613e-07
I4395 0 n4396 3.361e-02A M=6.283e-07
I4396 0 n4397 3.361e-02A M=6.655e-07
I4397 0 n4398 3.361e-02A M=2.150e-06
I4398 0 n4399 3.361e-02A M=2.153e-06
I4399 0 n4400 3.361e-02A M=1.474e-06
I4400 0 n4401 3.361e-02A M=8.503e-07
I4401 0 n4402 3.361e-02A M=1.852e-06
I4402 0 n4403 3.361e-02A M=1.347e-06
I4403 0 n4404 3.361e-02A M=3.539e-07
I4404 0 n4405 3.361e-02A M=3.538e-07
I4405 0 n4406 3.361e-02A M=6.409e-07
I4406 0 n4407 3.361e-02A M=9.869e-07
I4407 0 n4408 3.361e-02A M=6.869e-07
I4408 0 n4409 3.361e-02A M=1.075e-06
I4409 0 n4410 3.361e-02A M=1.377e-06
I4410 0 n4411 3.361e-02A M=3.502e-07
I4411 0 n4412 3.361e-02A M=3.620e-07
I4412 0 n4413 3.361e-02A M=1.201e-06
I4413 0 n4414 3.361e-02A M=7.283e-07
I4414 0 n4415 3.361e-02A M=1.257e-06
I4415 0 n4416 3.361e-02A M=5.114e-07
I4416 0 n4417 3.361e-02A M=9.447e-07
I4417 0 n4418 3.361e-02A M=1.026e-06
I4418 0 n4419 3.361e-02A M=1.807e-07
I4419 0 n4420 3.361e-02A M=1.168e-06
I4420 0 n4421 3.361e-02A M=9.629e-07
I4421 0 n4422 3.361e-02A M=3.128e-06
I4422 0 n4423 3.361e-02A M=6.792e-07
I4423 0 n4424 3.361e-02A M=5.093e-07
I4424 0 n4425 3.361e-02A M=5.670e-07
I4425 0 n4426 3.361e-02A M=1.612e-06
I4426 0 n4427 3.361e-02A M=1.621e-07
I4427 0 n4428 3.361e-02A M=3.540e-07
I4428 0 n4429 3.361e-02A M=4.925e-07
I4429 0 n4430 3.361e-02A M=8.668e-07
I4430 0 n4431 3.361e-02A M=1.126e-06
I4431 0 n4432 3.361e-02A M=2.066e-07
I4432 0 n4433 3.361e-02A M=9.135e-07
I4433 0 n4434 3.361e-02A M=1.220e-06
I4434 0 n4435 3.361e-02A M=1.255e-06
I4435 0 n4436 3.361e-02A M=7.393e-07
I4436 0 n4437 3.361e-02A M=1.668e-07
I4437 0 n4438 3.361e-02A M=1.809e-06
I4438 0 n4439 3.361e-02A M=7.077e-07
I4439 0 n4440 3.361e-02A M=1.328e-06
I4440 0 n4441 3.361e-02A M=4.566e-07
I4441 0 n4442 3.361e-02A M=3.957e-07
I4442 0 n4443 3.361e-02A M=7.970e-07
I4443 0 n4444 3.361e-02A M=1.316e-06
I4444 0 n4445 3.361e-02A M=1.205e-06
I4445 0 n4446 3.361e-02A M=1.257e-06
I4446 0 n4447 3.361e-02A M=6.599e-07
I4447 0 n4448 3.361e-02A M=5.796e-07
I4448 0 n4449 3.361e-02A M=8.215e-07
I4449 0 n4450 3.361e-02A M=3.691e-07
I4450 0 n4451 3.361e-02A M=2.042e-06
I4451 0 n4452 3.361e-02A M=1.088e-06
I4452 0 n4453 3.361e-02A M=7.657e-07
I4453 0 n4454 3.361e-02A M=4.744e-07
I4454 0 n4455 3.361e-02A M=1.649e-06
I4455 0 n4456 3.361e-02A M=1.778e-07
I4456 0 n4457 3.361e-02A M=2.251e-07
I4457 0 n4458 3.361e-02A M=9.499e-07
I4458 0 n4459 3.361e-02A M=8.332e-07
I4459 0 n4460 3.361e-02A M=1.340e-06
I4460 0 n4461 3.361e-02A M=1.050e-06
I4461 0 n4462 3.361e-02A M=3.449e-07
I4462 0 n4463 3.361e-02A M=1.620e-06
I4463 0 n4464 3.361e-02A M=1.048e-06
I4464 0 n4465 3.361e-02A M=1.069e-06
I4465 0 n4466 3.361e-02A M=9.725e-07
I4466 0 n4467 3.361e-02A M=2.680e-07
I4467 0 n4468 3.361e-02A M=6.168e-07
I4468 0 n4469 3.361e-02A M=5.317e-07
I4469 0 n4470 3.361e-02A M=1.215e-06
I4470 0 n4471 3.361e-02A M=9.827e-07
I4471 0 n4472 3.361e-02A M=7.004e-07
I4472 0 n4473 3.361e-02A M=2.665e-06
I4473 0 n4474 3.361e-02A M=8.190e-07
I4474 0 n4475 3.361e-02A M=9.317e-07
I4475 0 n4476 3.361e-02A M=5.397e-07
I4476 0 n4477 3.361e-02A M=4.978e-07
I4477 0 n4478 3.361e-02A M=8.607e-07
I4478 0 n4479 3.361e-02A M=1.070e-06
I4479 0 n4480 3.361e-02A M=1.575e-06
I4480 0 n4481 3.361e-02A M=4.924e-07
I4481 0 n4482 3.361e-02A M=5.499e-07
I4482 0 n4483 3.361e-02A M=1.463e-06
I4483 0 n4484 3.361e-02A M=8.438e-07
I4484 0 n4485 3.361e-02A M=7.316e-07
I4485 0 n4486 3.361e-02A M=2.182e-06
I4486 0 n4487 3.361e-02A M=1.050e-06
I4487 0 n4488 3.361e-02A M=7.267e-07
I4488 0 n4489 3.361e-02A M=9.928e-07
I4489 0 n4490 3.361e-02A M=4.149e-07
I4490 0 n4491 3.361e-02A M=9.077e-07
I4491 0 n4492 3.361e-02A M=9.199e-07
I4492 0 n4493 3.361e-02A M=6.912e-07
I4493 0 n4494 3.361e-02A M=4.884e-07
I4494 0 n4495 3.361e-02A M=1.855e-06
I4495 0 n4496 3.361e-02A M=8.807e-07
I4496 0 n4497 3.361e-02A M=5.235e-07
I4497 0 n4498 3.361e-02A M=1.913e-06
I4498 0 n4499 3.361e-02A M=7.979e-07
I4499 0 n4500 3.361e-02A M=1.572e-06
I4500 0 n4501 3.361e-02A M=1.324e-06
I4501 0 n4502 3.361e-02A M=1.156e-06
I4502 0 n4503 3.361e-02A M=2.222e-07
I4503 0 n4504 3.361e-02A M=1.514e-06
I4504 0 n4505 3.361e-02A M=5.984e-07
I4505 0 n4506 3.361e-02A M=7.083e-07
I4506 0 n4507 3.361e-02A M=1.454e-06
I4507 0 n4508 3.361e-02A M=7.352e-07
I4508 0 n4509 3.361e-02A M=6.859e-07
I4509 0 n4510 3.361e-02A M=1.279e-06
I4510 0 n4511 3.361e-02A M=1.580e-06
I4511 0 n4512 3.361e-02A M=6.058e-07
I4512 0 n4513 3.361e-02A M=5.350e-07
I4513 0 n4514 3.361e-02A M=5.929e-07
I4514 0 n4515 3.361e-02A M=1.549e-06
I4515 0 n4516 3.361e-02A M=7.770e-07
I4516 0 n4517 3.361e-02A M=6.097e-07
I4517 0 n4518 3.361e-02A M=5.069e-07
I4518 0 n4519 3.361e-02A M=1.736e-06
I4519 0 n4520 3.361e-02A M=8.891e-07
I4520 0 n4521 3.361e-02A M=1.903e-06
I4521 0 n4522 3.361e-02A M=4.467e-07
I4522 0 n4523 3.361e-02A M=9.193e-07
I4523 0 n4524 3.361e-02A M=6.443e-07
I4524 0 n4525 3.361e-02A M=1.203e-06
I4525 0 n4526 3.361e-02A M=7.676e-07
I4526 0 n4527 3.361e-02A M=2.064e-06
I4527 0 n4528 3.361e-02A M=8.549e-07
I4528 0 n4529 3.361e-02A M=1.221e-06
I4529 0 n4530 3.361e-02A M=1.613e-06
I4530 0 n1 3.361e-02A M=1.208e-06
I4531 0 n4532 3.361e-02A M=9.056e-07
I4532 0 n4533 3.361e-02A M=1.742e-06
I4533 0 n4534 3.361e-02A M=6.537e-07
I4534 0 n4535 3.361e-02A M=9.614e-07
I4535 0 n4536 3.361e-02A M=1.760e-07
I4536 0 n4537 3.361e-02A M=7.775e-07
I4537 0 n4538 3.361e-02A M=7.564e-07
I4538 0 n4539 3.361e-02A M=7.788e-07
I4539 0 n4540 3.361e-02A M=4.542e-07
I4540 0 n4541 3.361e-02A M=1.293e-06
I4541 0 n4542 3.361e-02A M=4.628e-07
I4542 0 n4543 3.361e-02A M=2.408e-06
I4543 0 n4544 3.361e-02A M=3.579e-07
I4544 0 n4545 3.361e-02A M=1.453e-06
I4545 0 n4546 3.361e-02A M=1.020e-06
I4546 0 n4547 3.361e-02A M=9.347e-07
I4547 0 n4548 3.361e-02A M=9.275e-07
I4548 0 n4549 3.361e-02A M=3.829e-07
I4549 0 n4550 3.361e-02A M=1.124e-06
I4550 0 n4551 3.361e-02A M=1.254e-06
I4551 0 n4552 3.361e-02A M=5.122e-07
I4552 0 n4553 3.361e-02A M=1.770e-06
I4553 0 n4554 3.361e-02A M=1.185e-06
I4554 0 n4555 3.361e-02A M=9.783e-07
I4555 0 n4556 3.361e-02A M=6.685e-07
I4556 0 n4557 3.361e-02A M=8.692e-07
I4557 0 n4558 3.361e-02A M=1.194e-06
I4558 0 n4559 3.361e-02A M=3.357e-07
I4559 0 n4560 3.361e-02A M=1.472e-06
I4560 0 n4561 3.361e-02A M=8.490e-07
I4561 0 n4562 3.361e-02A M=2.437e-07
I4562 0 n4563 3.361e-02A M=6.516e-07
I4563 0 n4564 3.361e-02A M=5.830e-07
I4564 0 n4565 3.361e-02A M=8.914e-07
I4565 0 n4566 3.361e-02A M=7.273e-07
I4566 0 n4567 3.361e-02A M=1.239e-06
I4567 0 n4568 3.361e-02A M=1.076e-06
I4568 0 n4569 3.361e-02A M=7.158e-07
I4569 0 n4570 3.361e-02A M=3.087e-07
I4570 0 n4571 3.361e-02A M=9.207e-07
I4571 0 n4572 3.361e-02A M=2.711e-06
I4572 0 n4573 3.361e-02A M=1.258e-06
I4573 0 n4574 3.361e-02A M=1.109e-06
I4574 0 n4575 3.361e-02A M=6.088e-07
I4575 0 n4576 3.361e-02A M=8.902e-07
I4576 0 n4577 3.361e-02A M=1.519e-06
I4577 0 n4578 3.361e-02A M=8.457e-07
I4578 0 n4579 3.361e-02A M=1.119e-06
I4579 0 n4580 3.361e-02A M=2.124e-06
I4580 0 n4581 3.361e-02A M=5.874e-07
I4581 0 n4582 3.361e-02A M=7.023e-07
I4582 0 n4583 3.361e-02A M=4.113e-07
I4583 0 n4584 3.361e-02A M=9.607e-07
I4584 0 n4585 3.361e-02A M=1.556e-06
I4585 0 n4586 3.361e-02A M=1.891e-06
I4586 0 n4587 3.361e-02A M=8.939e-07
I4587 0 n4588 3.361e-02A M=1.253e-06
I4588 0 n4589 3.361e-02A M=4.110e-07
I4589 0 n4590 3.361e-02A M=7.043e-07
I4590 0 n4591 3.361e-02A M=8.203e-07
I4591 0 n4592 3.361e-02A M=9.205e-07
I4592 0 n4593 3.361e-02A M=1.545e-06
I4593 0 n4594 3.361e-02A M=1.177e-06
I4594 0 n4595 3.361e-02A M=2.002e-06
I4595 0 n4596 3.361e-02A M=1.137e-06
I4596 0 n4597 3.361e-02A M=1.442e-06
I4597 0 n4598 3.361e-02A M=9.858e-07
I4598 0 n4599 3.361e-02A M=6.698e-07
I4599 0 n4600 3.361e-02A M=1.468e-06
I4600 0 n4601 3.361e-02A M=1.743e-07
I4601 0 n4602 3.361e-02A M=1.156e-06
I4602 0 n4603 3.361e-02A M=6.210e-07
I4603 0 n4604 3.361e-02A M=1.724e-06
I4604 0 n4605 3.361e-02A M=8.507e-07
I4605 0 n4606 3.361e-02A M=2.574e-06
I4606 0 n4607 3.361e-02A M=1.073e-06
I4607 0 n4608 3.361e-02A M=8.583e-07
I4608 0 n4609 3.361e-02A M=5.222e-07
I4609 0 n1 3.361e-02A M=1.412e-06
I4610 0 n4611 3.361e-02A M=1.053e-06
I4611 0 n4612 3.361e-02A M=1.019e-06
I4612 0 n4613 3.361e-02A M=1.371e-06
I4613 0 n4614 3.361e-02A M=1.233e-06
I4614 0 n4615 3.361e-02A M=9.963e-07
I4615 0 n4616 3.361e-02A M=2.111e-06
I4616 0 n4617 3.361e-02A M=7.486e-07
I4617 0 n4618 3.361e-02A M=2.933e-07
I4618 0 n4619 3.361e-02A M=1.033e-06
I4619 0 n4620 3.361e-02A M=5.758e-07
I4620 0 n4621 3.361e-02A M=4.930e-07
I4621 0 n4622 3.361e-02A M=1.230e-06
I4622 0 n4623 3.361e-02A M=8.840e-07
I4623 0 n4624 3.361e-02A M=5.672e-07
I4624 0 n4625 3.361e-02A M=1.028e-06
I4625 0 n4626 3.361e-02A M=7.985e-07
I4626 0 n4627 3.361e-02A M=2.937e-07
I4627 0 n4628 3.361e-02A M=7.059e-07
I4628 0 n4629 3.361e-02A M=9.912e-07
I4629 0 n4630 3.361e-02A M=8.790e-07
I4630 0 n4631 3.361e-02A M=1.360e-06
I4631 0 n4632 3.361e-02A M=7.005e-07
I4632 0 n4633 3.361e-02A M=1.428e-06
I4633 0 n4634 3.361e-02A M=4.700e-07
I4634 0 n4635 3.361e-02A M=1.087e-06
I4635 0 n4636 3.361e-02A M=7.478e-07
I4636 0 n4637 3.361e-02A M=9.424e-07
I4637 0 n4638 3.361e-02A M=3.143e-07
I4638 0 n4639 3.361e-02A M=5.717e-07
I4639 0 n4640 3.361e-02A M=1.499e-06
I4640 0 n4641 3.361e-02A M=4.347e-07
I4641 0 n4642 3.361e-02A M=3.311e-07
I4642 0 n4643 3.361e-02A M=7.428e-07
I4643 0 n4644 3.361e-02A M=2.913e-07
I4644 0 n4645 3.361e-02A M=4.348e-07
I4645 0 n4646 3.361e-02A M=9.540e-07
I4646 0 n4647 3.361e-02A M=1.716e-06
I4647 0 n4648 3.361e-02A M=9.178e-07
I4648 0 n4649 3.361e-02A M=9.487e-07
I4649 0 n4650 3.361e-02A M=1.302e-06
I4650 0 n4651 3.361e-02A M=4.838e-07
I4651 0 n4652 3.361e-02A M=1.122e-06
I4652 0 n4653 3.361e-02A M=1.279e-06
I4653 0 n4654 3.361e-02A M=1.907e-06
I4654 0 n4655 3.361e-02A M=7.492e-07
I4655 0 n4656 3.361e-02A M=6.288e-07
I4656 0 n4657 3.361e-02A M=5.471e-07
I4657 0 n4658 3.361e-02A M=3.988e-07
I4658 0 n4659 3.361e-02A M=7.652e-07
I4659 0 n4660 3.361e-02A M=4.826e-07
I4660 0 n4661 3.361e-02A M=8.577e-07
I4661 0 n4662 3.361e-02A M=2.752e-06
I4662 0 n4663 3.361e-02A M=9.810e-07
I4663 0 n4664 3.361e-02A M=8.048e-07
I4664 0 n4665 3.361e-02A M=1.123e-06
I4665 0 n4666 3.361e-02A M=6.877e-07
I4666 0 n1 3.361e-02A M=9.757e-07
I4667 0 n4668 3.361e-02A M=6.223e-07
I4668 0 n4669 3.361e-02A M=7.155e-07
I4669 0 n4670 3.361e-02A M=1.219e-06
I4670 0 n4671 3.361e-02A M=1.008e-06
I4671 0 n4672 3.361e-02A M=7.146e-07
I4672 0 n4673 3.361e-02A M=1.044e-06
I4673 0 n4674 3.361e-02A M=1.735e-06
I4674 0 n4675 3.361e-02A M=1.954e-06
I4675 0 n4676 3.361e-02A M=9.395e-07
I4676 0 n4677 3.361e-02A M=1.526e-06
I4677 0 n4678 3.361e-02A M=7.287e-07
I4678 0 n4679 3.361e-02A M=1.134e-07
I4679 0 n4680 3.361e-02A M=7.958e-07
I4680 0 n4681 3.361e-02A M=5.796e-07
I4681 0 n4682 3.361e-02A M=6.636e-07
I4682 0 n4683 3.361e-02A M=1.229e-06
I4683 0 n4684 3.361e-02A M=1.500e-06
I4684 0 n4685 3.361e-02A M=4.386e-07
I4685 0 n4686 3.361e-02A M=1.869e-06
I4686 0 n4687 3.361e-02A M=6.567e-07
I4687 0 n4688 3.361e-02A M=1.977e-06
I4688 0 n4689 3.361e-02A M=1.656e-06
I4689 0 n4690 3.361e-02A M=6.939e-07
I4690 0 n4691 3.361e-02A M=9.286e-07
I4691 0 n4692 3.361e-02A M=4.328e-07
I4692 0 n4693 3.361e-02A M=7.343e-07
I4693 0 n4694 3.361e-02A M=7.578e-07
I4694 0 n4695 3.361e-02A M=1.324e-06
I4695 0 n4696 3.361e-02A M=1.295e-06
I4696 0 n4697 3.361e-02A M=6.542e-07
I4697 0 n4698 3.361e-02A M=6.369e-07
I4698 0 n4699 3.361e-02A M=7.161e-07
I4699 0 n4700 3.361e-02A M=1.447e-06
I4700 0 n4701 3.361e-02A M=1.370e-06
I4701 0 n4702 3.361e-02A M=9.511e-07
I4702 0 n4703 3.361e-02A M=1.542e-06
I4703 0 n4704 3.361e-02A M=2.137e-06
I4704 0 n4705 3.361e-02A M=2.028e-06
I4705 0 n4706 3.361e-02A M=5.523e-07
I4706 0 n4707 3.361e-02A M=1.684e-06
I4707 0 n4708 3.361e-02A M=1.570e-06
I4708 0 n4709 3.361e-02A M=1.682e-06
I4709 0 n4710 3.361e-02A M=1.677e-06
I4710 0 n4711 3.361e-02A M=1.370e-06
I4711 0 n4712 3.361e-02A M=1.467e-06
I4712 0 n4713 3.361e-02A M=4.934e-07
I4713 0 n4714 3.361e-02A M=1.247e-06
I4714 0 n4715 3.361e-02A M=1.500e-06
I4715 0 n4716 3.361e-02A M=7.945e-07
I4716 0 n4717 3.361e-02A M=6.502e-07
I4717 0 n4718 3.361e-02A M=1.149e-06
I4718 0 n4719 3.361e-02A M=1.093e-06
I4719 0 n4720 3.361e-02A M=3.755e-07
I4720 0 n4721 3.361e-02A M=4.603e-07
I4721 0 n4722 3.361e-02A M=1.188e-06
I4722 0 n4723 3.361e-02A M=6.627e-07
I4723 0 n4724 3.361e-02A M=7.543e-07
I4724 0 n4725 3.361e-02A M=1.142e-06
I4725 0 n4726 3.361e-02A M=2.414e-07
I4726 0 n4727 3.361e-02A M=1.151e-06
I4727 0 n4728 3.361e-02A M=5.673e-07
I4728 0 n4729 3.361e-02A M=8.875e-07
I4729 0 n4730 3.361e-02A M=1.231e-06
I4730 0 n4731 3.361e-02A M=1.127e-06
I4731 0 n4732 3.361e-02A M=6.826e-07
I4732 0 n4733 3.361e-02A M=9.684e-07
I4733 0 n4734 3.361e-02A M=1.642e-06
I4734 0 n4735 3.361e-02A M=1.130e-06
I4735 0 n4736 3.361e-02A M=2.138e-07
I4736 0 n4737 3.361e-02A M=7.361e-07
I4737 0 n4738 3.361e-02A M=8.079e-07
I4738 0 n4739 3.361e-02A M=1.245e-06
I4739 0 n4740 3.361e-02A M=6.017e-07
I4740 0 n4741 3.361e-02A M=1.173e-06
I4741 0 n4742 3.361e-02A M=5.031e-07
I4742 0 n4743 3.361e-02A M=1.444e-06
I4743 0 n4744 3.361e-02A M=6.538e-07
I4744 0 n4745 3.361e-02A M=1.676e-06
I4745 0 n4746 3.361e-02A M=4.110e-07
I4746 0 n4747 3.361e-02A M=1.522e-06
I4747 0 n4748 3.361e-02A M=8.666e-07
I4748 0 n4749 3.361e-02A M=9.732e-07
I4749 0 n4750 3.361e-02A M=3.532e-07
I4750 0 n4751 3.361e-02A M=1.222e-06
I4751 0 n4752 3.361e-02A M=2.170e-06
I4752 0 n4753 3.361e-02A M=1.017e-06
I4753 0 n4754 3.361e-02A M=3.766e-07
I4754 0 n4755 3.361e-02A M=4.555e-07
I4755 0 n4756 3.361e-02A M=1.118e-06
I4756 0 n4757 3.361e-02A M=1.612e-06
I4757 0 n4758 3.361e-02A M=8.456e-07
I4758 0 n4759 3.361e-02A M=1.280e-06
I4759 0 n4760 3.361e-02A M=3.538e-07
I4760 0 n4761 3.361e-02A M=9.195e-07
I4761 0 n4762 3.361e-02A M=1.634e-06
I4762 0 n4763 3.361e-02A M=1.337e-06
I4763 0 n4764 3.361e-02A M=3.890e-07
I4764 0 n4765 3.361e-02A M=1.657e-06
I4765 0 n4766 3.361e-02A M=7.270e-07
I4766 0 n4767 3.361e-02A M=6.937e-07
I4767 0 n4768 3.361e-02A M=3.200e-07
I4768 0 n4769 3.361e-02A M=1.337e-06
I4769 0 n4770 3.361e-02A M=1.345e-06
I4770 0 n4771 3.361e-02A M=8.278e-07
I4771 0 n4772 3.361e-02A M=1.066e-06
I4772 0 n4773 3.361e-02A M=1.140e-06
I4773 0 n4774 3.361e-02A M=7.059e-07
I4774 0 n4775 3.361e-02A M=1.059e-06
I4775 0 n4776 3.361e-02A M=1.313e-06
I4776 0 n4777 3.361e-02A M=1.440e-06
I4777 0 n4778 3.361e-02A M=4.035e-07
I4778 0 n1 3.361e-02A M=3.751e-07
I4779 0 n4780 3.361e-02A M=1.271e-06
I4780 0 n4781 3.361e-02A M=7.076e-07
I4781 0 n4782 3.361e-02A M=7.602e-07
I4782 0 n4783 3.361e-02A M=9.778e-07
I4783 0 n4784 3.361e-02A M=9.722e-07
I4784 0 n4785 3.361e-02A M=7.447e-07
I4785 0 n4786 3.361e-02A M=5.884e-07
I4786 0 n4787 3.361e-02A M=4.085e-07
I4787 0 n4788 3.361e-02A M=8.302e-07
I4788 0 n4789 3.361e-02A M=2.072e-06
I4789 0 n4790 3.361e-02A M=8.547e-07
I4790 0 n4791 3.361e-02A M=1.188e-06
I4791 0 n4792 3.361e-02A M=2.215e-06
I4792 0 n4793 3.361e-02A M=2.420e-07
I4793 0 n4794 3.361e-02A M=1.245e-06
I4794 0 n4795 3.361e-02A M=4.390e-07
I4795 0 n4796 3.361e-02A M=4.431e-07
I4796 0 n4797 3.361e-02A M=1.104e-06
I4797 0 n4798 3.361e-02A M=1.274e-06
I4798 0 n4799 3.361e-02A M=2.887e-07
I4799 0 n4800 3.361e-02A M=2.443e-06
I4800 0 n4801 3.361e-02A M=6.392e-07
I4801 0 n4802 3.361e-02A M=1.761e-06
I4802 0 n4803 3.361e-02A M=2.469e-06
I4803 0 n4804 3.361e-02A M=7.483e-07
I4804 0 n4805 3.361e-02A M=1.412e-06
I4805 0 n4806 3.361e-02A M=1.193e-06
I4806 0 n4807 3.361e-02A M=1.771e-06
I4807 0 n1 3.361e-02A M=9.124e-07
I4808 0 n4809 3.361e-02A M=1.379e-06
I4809 0 n4810 3.361e-02A M=5.655e-07
I4810 0 n4811 3.361e-02A M=9.968e-07
I4811 0 n4812 3.361e-02A M=6.343e-07
I4812 0 n4813 3.361e-02A M=8.651e-07
I4813 0 n4814 3.361e-02A M=1.783e-06
I4814 0 n4815 3.361e-02A M=8.734e-07
I4815 0 n4816 3.361e-02A M=5.766e-07
I4816 0 n4817 3.361e-02A M=2.751e-07
I4817 0 n4818 3.361e-02A M=6.912e-07
I4818 0 n4819 3.361e-02A M=9.673e-07
I4819 0 n4820 3.361e-02A M=6.823e-07
I4820 0 n4821 3.361e-02A M=4.447e-07
I4821 0 n4822 3.361e-02A M=1.560e-06
I4822 0 n4823 3.361e-02A M=1.925e-06
I4823 0 n4824 3.361e-02A M=7.476e-07
I4824 0 n4825 3.361e-02A M=4.740e-07
I4825 0 n4826 3.361e-02A M=3.363e-07
I4826 0 n4827 3.361e-02A M=1.751e-06
I4827 0 n4828 3.361e-02A M=6.548e-07
I4828 0 n4829 3.361e-02A M=1.872e-07
I4829 0 n4830 3.361e-02A M=7.444e-07
I4830 0 n4831 3.361e-02A M=1.209e-06
I4831 0 n4832 3.361e-02A M=1.146e-06
I4832 0 n4833 3.361e-02A M=8.973e-07
I4833 0 n4834 3.361e-02A M=1.226e-06
I4834 0 n4835 3.361e-02A M=3.120e-07
I4835 0 n4836 3.361e-02A M=7.289e-07
I4836 0 n4837 3.361e-02A M=3.702e-07
I4837 0 n4838 3.361e-02A M=9.609e-07
I4838 0 n4839 3.361e-02A M=5.808e-07
I4839 0 n4840 3.361e-02A M=3.344e-07
I4840 0 n4841 3.361e-02A M=1.399e-06
I4841 0 n4842 3.361e-02A M=1.547e-06
I4842 0 n4843 3.361e-02A M=1.143e-06
I4843 0 n4844 3.361e-02A M=3.111e-07
I4844 0 n4845 3.361e-02A M=1.063e-06
I4845 0 n4846 3.361e-02A M=6.490e-07
I4846 0 n4847 3.361e-02A M=9.578e-07
I4847 0 n4848 2.976e-02A M=1.046e-06
I4848 0 n4849 2.976e-02A M=7.614e-07
I4849 0 n4850 2.976e-02A M=1.053e-06
I4850 0 n4851 2.976e-02A M=1.328e-06
I4851 0 n4852 2.976e-02A M=4.409e-07
I4852 0 n4853 2.976e-02A M=1.204e-06
I4853 0 n4854 2.976e-02A M=8.714e-07
I4854 0 n4855 2.976e-02A M=3.476e-07
I4855 0 n4856 2.976e-02A M=7.279e-07
I4856 0 n4857 2.976e-02A M=4.012e-06
I4857 0 n4858 2.976e-02A M=1.837e-06
I4858 0 n4859 2.976e-02A M=9.303e-07
I4859 0 n4860 2.976e-02A M=2.686e-07
I4860 0 n4861 2.976e-02A M=8.868e-07
I4861 0 n4862 2.976e-02A M=2.902e-07
I4862 0 n4863 2.976e-02A M=5.308e-07
I4863 0 n4864 2.976e-02A M=1.422e-06
I4864 0 n4865 2.976e-02A M=9.156e-07
I4865 0 n4866 2.976e-02A M=9.049e-07
I4866 0 n4867 2.976e-02A M=1.857e-06
I4867 0 n4868 2.976e-02A M=8.523e-07
I4868 0 n4869 2.976e-02A M=9.346e-07
I4869 0 n4870 2.976e-02A M=7.523e-07
I4870 0 n4871 2.976e-02A M=1.171e-06
I4871 0 n4872 2.976e-02A M=4.187e-07
I4872 0 n4873 2.976e-02A M=9.190e-07
I4873 0 n4874 2.976e-02A M=1.169e-06
I4874 0 n4875 2.976e-02A M=4.616e-07
I4875 0 n4876 2.976e-02A M=8.934e-07
I4876 0 n4877 2.976e-02A M=1.450e-06
I4877 0 n4878 2.976e-02A M=2.544e-07
I4878 0 n4879 2.976e-02A M=1.144e-06
I4879 0 n4880 2.976e-02A M=9.680e-07
I4880 0 n4881 2.976e-02A M=6.387e-07
I4881 0 n4882 2.976e-02A M=9.759e-07
I4882 0 n4883 2.976e-02A M=7.238e-07
I4883 0 n4884 2.976e-02A M=1.043e-06
I4884 0 n4885 2.976e-02A M=3.366e-07
I4885 0 n4886 2.976e-02A M=4.044e-07
I4886 0 n4887 2.976e-02A M=1.745e-06
I4887 0 n4888 2.976e-02A M=1.804e-06
I4888 0 n4889 2.976e-02A M=1.170e-06
I4889 0 n4890 2.976e-02A M=6.821e-07
I4890 0 n4891 2.976e-02A M=2.558e-07
I4891 0 n4892 2.976e-02A M=3.185e-07
I4892 0 n4893 2.976e-02A M=7.170e-07
I4893 0 n4894 2.976e-02A M=1.118e-06
I4894 0 n4895 2.976e-02A M=5.745e-07
I4895 0 n4896 2.976e-02A M=4.835e-07
I4896 0 n4897 2.976e-02A M=6.224e-07
I4897 0 n4898 2.976e-02A M=7.356e-07
I4898 0 n4899 2.976e-02A M=8.107e-07
I4899 0 n4900 2.976e-02A M=7.691e-07
I4900 0 n4901 2.976e-02A M=8.602e-07
I4901 0 n4902 2.976e-02A M=7.421e-07
I4902 0 n4903 2.976e-02A M=1.344e-06
I4903 0 n4904 2.976e-02A M=1.542e-06
I4904 0 n4905 2.976e-02A M=6.035e-07
I4905 0 n4906 2.976e-02A M=5.768e-07
I4906 0 n4907 2.976e-02A M=6.036e-07
I4907 0 n4908 2.976e-02A M=1.652e-06
I4908 0 n4909 2.976e-02A M=2.023e-06
I4909 0 n4910 2.976e-02A M=5.563e-07
I4910 0 n4911 2.976e-02A M=5.590e-07
I4911 0 n4912 2.976e-02A M=6.625e-07
I4912 0 n4913 2.976e-02A M=2.097e-06
I4913 0 n4914 2.976e-02A M=1.607e-06
I4914 0 n4915 2.976e-02A M=3.663e-07
I4915 0 n4916 2.976e-02A M=1.284e-06
I4916 0 n4917 2.976e-02A M=6.208e-07
I4917 0 n4918 2.976e-02A M=1.487e-06
I4918 0 n4919 2.976e-02A M=8.912e-07
I4919 0 n1 2.976e-02A M=3.125e-07
I4920 0 n4921 2.976e-02A M=2.055e-06
I4921 0 n4922 2.976e-02A M=8.014e-07
I4922 0 n4923 2.976e-02A M=1.056e-06
I4923 0 n4924 2.976e-02A M=1.310e-06
I4924 0 n4925 2.976e-02A M=7.943e-07
I4925 0 n4926 2.976e-02A M=5.858e-07
I4926 0 n4927 2.976e-02A M=7.364e-07
I4927 0 n4928 2.976e-02A M=8.525e-07
I4928 0 n4929 2.976e-02A M=7.454e-07
I4929 0 n4930 2.976e-02A M=1.269e-06
I4930 0 n4931 2.976e-02A M=2.875e-06
I4931 0 n4932 2.976e-02A M=1.105e-06
I4932 0 n4933 2.976e-02A M=1.558e-07
I4933 0 n4934 2.976e-02A M=1.888e-07
I4934 0 n4935 2.976e-02A M=6.545e-07
I4935 0 n4936 2.976e-02A M=6.274e-07
I4936 0 n4937 2.976e-02A M=2.607e-06
I4937 0 n4938 2.976e-02A M=1.343e-06
I4938 0 n4939 2.976e-02A M=1.062e-06
I4939 0 n4940 2.976e-02A M=6.856e-07
I4940 0 n4941 2.976e-02A M=1.025e-06
I4941 0 n4942 2.976e-02A M=1.246e-06
I4942 0 n4943 2.976e-02A M=1.295e-06
I4943 0 n4944 2.976e-02A M=1.016e-06
I4944 0 n4945 2.976e-02A M=9.476e-07
I4945 0 n4946 2.976e-02A M=2.738e-07
I4946 0 n4947 2.976e-02A M=4.281e-07
I4947 0 n4948 2.976e-02A M=4.377e-07
I4948 0 n4949 2.976e-02A M=2.578e-06
I4949 0 n4950 2.976e-02A M=5.885e-07
I4950 0 n4951 2.976e-02A M=7.572e-07
I4951 0 n4952 2.976e-02A M=9.881e-07
I4952 0 n4953 2.976e-02A M=1.886e-06
I4953 0 n4954 2.976e-02A M=3.354e-07
I4954 0 n4955 2.976e-02A M=1.720e-06
I4955 0 n4956 2.976e-02A M=7.478e-07
I4956 0 n4957 2.976e-02A M=2.388e-06
I4957 0 n4958 2.976e-02A M=7.157e-07
I4958 0 n4959 2.976e-02A M=8.521e-07
I4959 0 n4960 2.976e-02A M=3.183e-07
I4960 0 n4961 2.976e-02A M=4.207e-07
I4961 0 n4962 2.976e-02A M=1.446e-06
I4962 0 n4963 2.976e-02A M=3.635e-07
I4963 0 n4964 2.976e-02A M=8.401e-07
I4964 0 n4965 2.976e-02A M=2.220e-07
I4965 0 n4966 2.976e-02A M=1.910e-06
I4966 0 n4967 2.976e-02A M=1.832e-06
I4967 0 n4968 2.976e-02A M=1.112e-06
I4968 0 n4969 2.976e-02A M=1.503e-06
I4969 0 n4970 2.976e-02A M=8.235e-07
I4970 0 n4971 2.976e-02A M=3.260e-07
I4971 0 n4972 2.976e-02A M=8.690e-07
I4972 0 n4973 2.976e-02A M=8.397e-07
I4973 0 n4974 2.976e-02A M=9.962e-07
I4974 0 n4975 2.976e-02A M=1.055e-06
I4975 0 n4976 2.976e-02A M=9.329e-07
I4976 0 n4977 2.976e-02A M=5.377e-07
I4977 0 n4978 2.976e-02A M=1.724e-06
I4978 0 n4979 2.976e-02A M=1.343e-06
I4979 0 n4980 2.976e-02A M=1.334e-06
I4980 0 n4981 2.976e-02A M=1.202e-06
I4981 0 n4982 2.976e-02A M=2.907e-06
I4982 0 n4983 2.976e-02A M=8.334e-07
I4983 0 n4984 2.976e-02A M=1.427e-06
I4984 0 n4985 2.976e-02A M=3.703e-07
I4985 0 n4986 2.976e-02A M=9.487e-07
I4986 0 n4987 2.976e-02A M=1.121e-06
I4987 0 n4988 2.976e-02A M=2.594e-06
I4988 0 n4989 2.976e-02A M=7.244e-07
I4989 0 n4990 2.976e-02A M=9.051e-07
I4990 0 n4991 2.976e-02A M=1.321e-06
I4991 0 n4992 2.976e-02A M=1.421e-06
I4992 0 n4993 2.976e-02A M=2.648e-06
I4993 0 n4994 2.976e-02A M=1.101e-06
I4994 0 n4995 2.976e-02A M=9.097e-07
I4995 0 n4996 2.976e-02A M=1.831e-06
I4996 0 n1 2.976e-02A M=1.000e-06
I4997 0 n4998 2.976e-02A M=9.628e-07
I4998 0 n4999 2.976e-02A M=1.485e-06
I4999 0 n5000 2.976e-02A M=5.188e-07
I5000 0 n5001 2.976e-02A M=2.183e-06
I5001 0 n5002 2.976e-02A M=1.446e-06
I5002 0 n5003 2.976e-02A M=2.108e-06
I5003 0 n5004 2.976e-02A M=1.618e-06
I5004 0 n5005 2.976e-02A M=6.537e-07
I5005 0 n5006 2.976e-02A M=6.469e-07
I5006 0 n5007 2.976e-02A M=2.414e-06
I5007 0 n5008 2.976e-02A M=1.031e-06
I5008 0 n5009 2.976e-02A M=4.610e-07
I5009 0 n5010 2.976e-02A M=5.483e-07
I5010 0 n5011 2.976e-02A M=1.326e-06
I5011 0 n5012 2.976e-02A M=5.782e-07
I5012 0 n5013 2.976e-02A M=1.350e-06
I5013 0 n5014 2.976e-02A M=1.034e-06
I5014 0 n5015 2.976e-02A M=2.047e-06
I5015 0 n5016 2.976e-02A M=9.660e-07
I5016 0 n5017 2.976e-02A M=4.306e-07
I5017 0 n5018 2.976e-02A M=6.264e-07
I5018 0 n5019 2.976e-02A M=8.126e-07
I5019 0 n5020 2.976e-02A M=8.900e-07
I5020 0 n5021 2.976e-02A M=7.378e-07
I5021 0 n5022 2.976e-02A M=1.700e-07
I5022 0 n5023 2.976e-02A M=5.695e-07
I5023 0 n5024 2.976e-02A M=1.557e-06
I5024 0 n5025 2.976e-02A M=3.888e-07
I5025 0 n5026 2.976e-02A M=5.091e-07
I5026 0 n5027 2.976e-02A M=6.649e-07
I5027 0 n5028 2.976e-02A M=7.829e-07
I5028 0 n5029 2.976e-02A M=6.270e-07
I5029 0 n5030 2.976e-02A M=5.877e-07
I5030 0 n5031 2.976e-02A M=1.155e-06
I5031 0 n5032 2.976e-02A M=6.314e-07
I5032 0 n5033 2.976e-02A M=3.843e-07
I5033 0 n5034 2.976e-02A M=3.390e-07
I5034 0 n5035 2.976e-02A M=2.038e-06
I5035 0 n5036 2.976e-02A M=9.973e-07
I5036 0 n5037 2.976e-02A M=1.184e-06
I5037 0 n5038 2.976e-02A M=1.340e-06
I5038 0 n5039 2.976e-02A M=1.651e-07
I5039 0 n5040 2.976e-02A M=7.603e-07
I5040 0 n5041 2.976e-02A M=7.741e-07
I5041 0 n5042 2.976e-02A M=7.156e-07
I5042 0 n5043 2.976e-02A M=1.331e-06
I5043 0 n5044 2.976e-02A M=2.924e-07
I5044 0 n5045 2.976e-02A M=1.390e-06
I5045 0 n5046 2.976e-02A M=3.589e-07
I5046 0 n5047 2.976e-02A M=4.495e-07
I5047 0 n5048 2.976e-02A M=7.244e-07
I5048 0 n5049 2.976e-02A M=1.151e-06
I5049 0 n5050 2.976e-02A M=9.764e-07
I5050 0 n5051 2.976e-02A M=3.893e-07
I5051 0 n5052 2.976e-02A M=1.686e-06
I5052 0 n5053 2.976e-02A M=9.205e-07
I5053 0 n5054 2.976e-02A M=8.258e-07
I5054 0 n5055 2.976e-02A M=1.018e-06
I5055 0 n5056 2.976e-02A M=1.325e-06
I5056 0 n5057 2.976e-02A M=9.168e-07
I5057 0 n5058 2.976e-02A M=1.206e-06
I5058 0 n5059 2.976e-02A M=9.646e-07
I5059 0 n5060 2.976e-02A M=8.015e-07
I5060 0 n5061 2.976e-02A M=2.013e-06
I5061 0 n5062 2.976e-02A M=4.647e-07
I5062 0 n5063 2.976e-02A M=6.884e-07
I5063 0 n5064 2.976e-02A M=1.189e-06
I5064 0 n5065 2.976e-02A M=1.534e-06
I5065 0 n5066 2.976e-02A M=8.549e-07
I5066 0 n5067 2.976e-02A M=5.895e-07
I5067 0 n5068 2.976e-02A M=5.794e-07
I5068 0 n5069 2.976e-02A M=6.845e-07
I5069 0 n5070 2.976e-02A M=1.537e-06
I5070 0 n5071 2.976e-02A M=5.793e-07
I5071 0 n5072 2.976e-02A M=1.932e-06
I5072 0 n5073 2.976e-02A M=1.390e-06
I5073 0 n5074 2.976e-02A M=1.135e-06
I5074 0 n5075 2.976e-02A M=8.154e-07
I5075 0 n5076 2.976e-02A M=4.848e-07
I5076 0 n5077 2.976e-02A M=2.621e-07
I5077 0 n5078 2.976e-02A M=5.245e-07
I5078 0 n5079 2.976e-02A M=1.344e-06
I5079 0 n5080 2.976e-02A M=1.082e-06
I5080 0 n5081 2.976e-02A M=1.265e-06
I5081 0 n5082 2.976e-02A M=1.383e-06
I5082 0 n5083 2.976e-02A M=1.251e-06
I5083 0 n5084 2.976e-02A M=8.326e-07
I5084 0 n5085 2.976e-02A M=1.623e-06
I5085 0 n5086 2.976e-02A M=1.991e-06
I5086 0 n5087 2.976e-02A M=6.515e-07
I5087 0 n5088 2.976e-02A M=1.032e-06
I5088 0 n5089 2.976e-02A M=5.068e-07
I5089 0 n5090 2.976e-02A M=6.705e-07
I5090 0 n5091 2.976e-02A M=1.734e-06
I5091 0 n5092 2.976e-02A M=1.420e-06
I5092 0 n5093 2.976e-02A M=7.939e-07
I5093 0 n5094 2.976e-02A M=3.395e-07
I5094 0 n1 2.976e-02A M=4.032e-07
I5095 0 n5096 2.976e-02A M=8.039e-07
I5096 0 n5097 2.976e-02A M=3.698e-07
I5097 0 n5098 2.976e-02A M=4.993e-07
I5098 0 n5099 2.976e-02A M=1.188e-06
I5099 0 n5100 2.976e-02A M=1.595e-06
I5100 0 n5101 2.976e-02A M=1.940e-06
I5101 0 n5102 2.976e-02A M=9.582e-07
I5102 0 n5103 2.976e-02A M=1.187e-06
I5103 0 n5104 2.976e-02A M=6.970e-07
I5104 0 n5105 2.976e-02A M=1.021e-06
I5105 0 n5106 2.976e-02A M=6.657e-07
I5106 0 n5107 2.976e-02A M=7.126e-07
I5107 0 n5108 2.976e-02A M=1.190e-06
I5108 0 n5109 2.976e-02A M=5.948e-07
I5109 0 n5110 2.976e-02A M=5.510e-07
I5110 0 n5111 2.976e-02A M=1.929e-06
I5111 0 n5112 2.976e-02A M=3.678e-07
I5112 0 n5113 2.976e-02A M=9.511e-07
I5113 0 n5114 2.976e-02A M=1.214e-06
I5114 0 n5115 2.976e-02A M=8.266e-07
I5115 0 n5116 2.976e-02A M=7.226e-07
I5116 0 n5117 2.976e-02A M=4.822e-07
I5117 0 n5118 2.976e-02A M=8.821e-07
I5118 0 n5119 2.976e-02A M=1.099e-06
I5119 0 n5120 2.976e-02A M=3.654e-07
I5120 0 n5121 2.976e-02A M=1.129e-06
I5121 0 n5122 2.976e-02A M=8.076e-07
I5122 0 n5123 2.976e-02A M=1.746e-06
I5123 0 n5124 2.976e-02A M=1.308e-06
I5124 0 n5125 2.976e-02A M=8.004e-07
I5125 0 n5126 2.976e-02A M=2.776e-07
I5126 0 n5127 2.976e-02A M=1.133e-06
I5127 0 n5128 2.976e-02A M=1.324e-06
I5128 0 n5129 2.976e-02A M=1.443e-06
I5129 0 n5130 2.976e-02A M=7.094e-07
I5130 0 n5131 2.976e-02A M=8.073e-07
I5131 0 n5132 2.976e-02A M=1.303e-06
I5132 0 n5133 2.976e-02A M=1.423e-06
I5133 0 n5134 2.976e-02A M=9.717e-07
I5134 0 n5135 2.976e-02A M=2.361e-07
I5135 0 n5136 2.976e-02A M=2.498e-07
I5136 0 n5137 2.976e-02A M=7.545e-07
I5137 0 n5138 2.976e-02A M=1.070e-06
I5138 0 n5139 2.976e-02A M=7.045e-07
I5139 0 n5140 2.976e-02A M=6.116e-07
I5140 0 n5141 2.976e-02A M=4.974e-07
I5141 0 n5142 2.976e-02A M=1.427e-06
I5142 0 n5143 2.976e-02A M=8.906e-07
I5143 0 n5144 2.976e-02A M=1.208e-06
I5144 0 n5145 2.976e-02A M=9.229e-07
I5145 0 n5146 2.976e-02A M=1.438e-06
I5146 0 n5147 2.976e-02A M=1.562e-06
I5147 0 n5148 2.976e-02A M=1.409e-07
I5148 0 n5149 2.976e-02A M=1.176e-06
I5149 0 n5150 2.976e-02A M=9.290e-07
I5150 0 n5151 2.976e-02A M=2.235e-06
I5151 0 n5152 2.976e-02A M=1.107e-06
I5152 0 n5153 2.976e-02A M=4.809e-07
I5153 0 n5154 2.976e-02A M=1.253e-06
I5154 0 n5155 2.976e-02A M=2.488e-07
I5155 0 n5156 2.976e-02A M=1.777e-06
I5156 0 n5157 2.976e-02A M=7.559e-07
I5157 0 n5158 2.976e-02A M=1.003e-06
I5158 0 n5159 2.976e-02A M=6.154e-07
I5159 0 n5160 2.976e-02A M=5.843e-07
I5160 0 n5161 2.976e-02A M=4.649e-07
I5161 0 n5162 2.976e-02A M=4.749e-07
I5162 0 n5163 2.976e-02A M=8.593e-07
I5163 0 n5164 2.976e-02A M=1.167e-06
I5164 0 n5165 2.976e-02A M=1.137e-06
I5165 0 n5166 2.976e-02A M=3.195e-07
I5166 0 n5167 2.976e-02A M=8.925e-07
I5167 0 n5168 2.976e-02A M=5.451e-07
I5168 0 n5169 2.976e-02A M=1.183e-06
I5169 0 n5170 2.976e-02A M=1.144e-06
I5170 0 n5171 2.976e-02A M=3.620e-07
I5171 0 n5172 2.976e-02A M=4.163e-07
I5172 0 n5173 2.976e-02A M=9.836e-07
I5173 0 n5174 2.976e-02A M=7.003e-07
I5174 0 n5175 2.976e-02A M=6.543e-07
I5175 0 n5176 2.976e-02A M=1.220e-06
I5176 0 n5177 2.976e-02A M=3.973e-07
I5177 0 n5178 2.976e-02A M=5.614e-07
I5178 0 n5179 2.976e-02A M=4.510e-07
I5179 0 n5180 2.976e-02A M=1.485e-06
I5180 0 n5181 2.976e-02A M=1.469e-06
I5181 0 n5182 2.976e-02A M=9.666e-07
I5182 0 n5183 2.976e-02A M=6.918e-07
I5183 0 n5184 2.976e-02A M=1.922e-07
I5184 0 n5185 2.976e-02A M=7.631e-07
I5185 0 n5186 2.976e-02A M=1.296e-06
I5186 0 n5187 2.976e-02A M=1.404e-06
I5187 0 n5188 2.976e-02A M=8.764e-07
I5188 0 n5189 2.976e-02A M=3.220e-07
I5189 0 n5190 2.976e-02A M=1.118e-06
I5190 0 n5191 2.976e-02A M=3.030e-07
I5191 0 n5192 2.976e-02A M=7.597e-07
I5192 0 n5193 2.976e-02A M=3.521e-07
I5193 0 n5194 2.976e-02A M=1.369e-06
I5194 0 n5195 2.976e-02A M=4.260e-07
I5195 0 n5196 2.976e-02A M=1.192e-06
I5196 0 n5197 2.976e-02A M=1.150e-06
I5197 0 n5198 2.976e-02A M=2.148e-07
I5198 0 n5199 2.976e-02A M=2.094e-06
I5199 0 n5200 2.976e-02A M=3.264e-07
I5200 0 n5201 2.976e-02A M=4.653e-07
I5201 0 n5202 2.976e-02A M=6.667e-07
I5202 0 n5203 2.976e-02A M=2.075e-07
I5203 0 n5204 2.976e-02A M=1.607e-06
I5204 0 n5205 2.976e-02A M=1.069e-06
I5205 0 n5206 2.976e-02A M=8.965e-07
I5206 0 n5207 2.976e-02A M=7.218e-07
I5207 0 n5208 2.976e-02A M=1.173e-06
I5208 0 n5209 2.976e-02A M=1.344e-06
I5209 0 n1 2.976e-02A M=6.978e-07
I5210 0 n5211 2.976e-02A M=2.867e-06
I5211 0 n5212 2.976e-02A M=7.528e-07
I5212 0 n5213 2.976e-02A M=1.022e-06
I5213 0 n5214 2.976e-02A M=1.075e-06
I5214 0 n5215 2.976e-02A M=1.349e-06
I5215 0 n5216 2.976e-02A M=6.489e-07
I5216 0 n5217 2.976e-02A M=5.055e-07
I5217 0 n5218 2.976e-02A M=8.185e-07
I5218 0 n5219 2.976e-02A M=1.035e-06
I5219 0 n5220 2.976e-02A M=1.269e-06
I5220 0 n5221 2.976e-02A M=1.299e-06
I5221 0 n5222 2.976e-02A M=5.758e-07
I5222 0 n5223 2.976e-02A M=1.769e-06
I5223 0 n5224 2.976e-02A M=3.758e-07
I5224 0 n5225 2.976e-02A M=1.199e-06
I5225 0 n5226 2.976e-02A M=1.646e-07
I5226 0 n5227 2.976e-02A M=4.583e-07
I5227 0 n5228 2.976e-02A M=1.012e-06
I5228 0 n5229 2.976e-02A M=8.616e-07
I5229 0 n5230 2.976e-02A M=1.763e-07
I5230 0 n5231 2.976e-02A M=5.722e-07
I5231 0 n5232 2.976e-02A M=1.305e-07
I5232 0 n5233 2.976e-02A M=9.308e-07
I5233 0 n5234 2.976e-02A M=9.161e-07
I5234 0 n5235 2.976e-02A M=6.711e-07
I5235 0 n5236 2.976e-02A M=5.345e-07
I5236 0 n5237 2.976e-02A M=2.724e-07
I5237 0 n5238 2.976e-02A M=1.684e-06
I5238 0 n5239 2.976e-02A M=7.514e-07
I5239 0 n5240 2.976e-02A M=1.442e-06
I5240 0 n5241 2.976e-02A M=5.889e-07
I5241 0 n5242 2.976e-02A M=8.515e-07
I5242 0 n5243 2.976e-02A M=3.208e-07
I5243 0 n1 2.976e-02A M=1.390e-06
I5244 0 n5245 2.976e-02A M=4.197e-07
I5245 0 n5246 2.976e-02A M=2.239e-06
I5246 0 n5247 2.976e-02A M=1.161e-06
I5247 0 n5248 2.976e-02A M=7.479e-07
I5248 0 n5249 2.976e-02A M=5.327e-07
I5249 0 n5250 2.976e-02A M=6.708e-07
I5250 0 n5251 2.976e-02A M=1.242e-06
I5251 0 n5252 2.976e-02A M=2.784e-07
I5252 0 n5253 2.976e-02A M=2.420e-07
I5253 0 n5254 2.976e-02A M=1.748e-06
I5254 0 n5255 2.976e-02A M=1.052e-06
I5255 0 n5256 2.976e-02A M=2.003e-06
I5256 0 n5257 2.976e-02A M=1.570e-06
I5257 0 n5258 2.976e-02A M=7.546e-07
I5258 0 n5259 2.976e-02A M=4.515e-07
I5259 0 n5260 2.976e-02A M=1.214e-06
I5260 0 n5261 2.976e-02A M=8.871e-07
I5261 0 n5262 2.976e-02A M=6.020e-07
I5262 0 n5263 2.976e-02A M=1.205e-06
I5263 0 n5264 2.976e-02A M=4.606e-07
I5264 0 n5265 2.976e-02A M=1.702e-06
I5265 0 n5266 2.976e-02A M=6.798e-07
I5266 0 n5267 2.976e-02A M=6.368e-07
I5267 0 n5268 2.976e-02A M=2.154e-07
I5268 0 n5269 2.976e-02A M=2.515e-07
I5269 0 n5270 2.976e-02A M=1.283e-06
I5270 0 n5271 2.976e-02A M=8.802e-07
I5271 0 n5272 2.976e-02A M=3.179e-07
I5272 0 n5273 2.976e-02A M=2.547e-07
I5273 0 n5274 2.976e-02A M=1.325e-06
I5274 0 n5275 2.976e-02A M=1.716e-06
I5275 0 n5276 2.976e-02A M=3.952e-07
I5276 0 n5277 2.976e-02A M=1.055e-06
I5277 0 n5278 2.976e-02A M=1.097e-06
I5278 0 n5279 2.976e-02A M=1.306e-06
I5279 0 n5280 2.976e-02A M=1.798e-06
I5280 0 n5281 2.976e-02A M=5.670e-07
I5281 0 n5282 2.976e-02A M=8.507e-07
I5282 0 n5283 2.976e-02A M=9.775e-07
I5283 0 n5284 2.976e-02A M=2.364e-07
I5284 0 n5285 2.976e-02A M=9.483e-07
I5285 0 n5286 2.976e-02A M=1.045e-06
I5286 0 n5287 2.976e-02A M=8.461e-07
I5287 0 n5288 2.976e-02A M=5.995e-07
I5288 0 n5289 2.976e-02A M=7.001e-07
I5289 0 n5290 2.976e-02A M=2.833e-07
I5290 0 n5291 2.976e-02A M=1.314e-06
I5291 0 n5292 2.976e-02A M=1.332e-06
I5292 0 n5293 2.976e-02A M=1.404e-06
I5293 0 n5294 2.976e-02A M=1.043e-06
I5294 0 n5295 2.976e-02A M=9.204e-07
I5295 0 n5296 2.976e-02A M=1.416e-06
I5296 0 n5297 2.976e-02A M=2.117e-06
I5297 0 n5298 2.976e-02A M=2.144e-07
I5298 0 n5299 2.976e-02A M=7.369e-07
I5299 0 n5300 2.976e-02A M=9.461e-07
I5300 0 n5301 2.976e-02A M=5.026e-07
I5301 0 n5302 2.976e-02A M=5.388e-07
I5302 0 n5303 2.976e-02A M=2.453e-07
I5303 0 n5304 2.976e-02A M=5.823e-07
I5304 0 n5305 2.976e-02A M=6.598e-07
I5305 0 n5306 2.976e-02A M=3.787e-07
I5306 0 n5307 2.976e-02A M=9.436e-07
I5307 0 n5308 2.976e-02A M=6.058e-07
I5308 0 n5309 2.976e-02A M=2.696e-07
I5309 0 n5310 2.976e-02A M=8.503e-07
I5310 0 n5311 2.976e-02A M=1.564e-06
I5311 0 n5312 2.976e-02A M=1.801e-06
I5312 0 n5313 2.976e-02A M=7.214e-07
I5313 0 n5314 2.976e-02A M=1.308e-06
I5314 0 n5315 2.976e-02A M=5.606e-07
I5315 0 n5316 2.976e-02A M=6.878e-07
I5316 0 n5317 2.976e-02A M=6.703e-07
I5317 0 n5318 2.976e-02A M=1.387e-06
I5318 0 n5319 2.976e-02A M=1.089e-06
I5319 0 n5320 2.976e-02A M=4.618e-07
I5320 0 n5321 2.976e-02A M=2.499e-07
I5321 0 n5322 2.976e-02A M=7.210e-07
I5322 0 n5323 2.976e-02A M=7.848e-07
I5323 0 n5324 2.976e-02A M=1.477e-06
I5324 0 n5325 2.976e-02A M=8.349e-07
I5325 0 n5326 2.976e-02A M=3.935e-07
I5326 0 n5327 2.976e-02A M=1.227e-06
I5327 0 n5328 2.976e-02A M=2.139e-06
I5328 0 n5329 2.976e-02A M=3.723e-07
I5329 0 n5330 2.976e-02A M=1.248e-06
I5330 0 n5331 2.976e-02A M=9.141e-07
I5331 0 n5332 2.976e-02A M=5.783e-07
I5332 0 n5333 2.976e-02A M=2.254e-06
I5333 0 n5334 2.976e-02A M=3.276e-07
I5334 0 n5335 2.976e-02A M=1.578e-06
I5335 0 n5336 2.976e-02A M=3.298e-07
I5336 0 n5337 2.976e-02A M=1.061e-06
I5337 0 n5338 2.976e-02A M=9.671e-07
I5338 0 n5339 2.976e-02A M=1.295e-06
I5339 0 n5340 2.976e-02A M=1.299e-06
I5340 0 n5341 2.976e-02A M=1.155e-06
I5341 0 n5342 2.976e-02A M=7.233e-07
I5342 0 n5343 2.976e-02A M=5.343e-07
I5343 0 n5344 2.976e-02A M=4.430e-07
I5344 0 n5345 2.976e-02A M=7.275e-07
I5345 0 n5346 2.976e-02A M=9.684e-07
I5346 0 n5347 2.976e-02A M=8.046e-07
I5347 0 n5348 2.976e-02A M=1.688e-07
I5348 0 n5349 2.976e-02A M=9.796e-07
I5349 0 n5350 2.976e-02A M=1.060e-06
I5350 0 n5351 2.976e-02A M=8.965e-07
I5351 0 n5352 2.976e-02A M=2.814e-07
I5352 0 n5353 2.976e-02A M=4.814e-07
I5353 0 n5354 2.976e-02A M=8.295e-07
I5354 0 n5355 2.976e-02A M=1.094e-06
I5355 0 n5356 2.976e-02A M=9.000e-07
I5356 0 n5357 2.976e-02A M=4.412e-07
I5357 0 n5358 2.976e-02A M=1.352e-06
I5358 0 n5359 2.976e-02A M=1.342e-06
I5359 0 n5360 2.976e-02A M=4.872e-07
I5360 0 n5361 2.976e-02A M=1.045e-06
I5361 0 n5362 2.976e-02A M=9.111e-07
I5362 0 n5363 2.976e-02A M=1.313e-06
I5363 0 n5364 2.976e-02A M=1.540e-06
I5364 0 n5365 2.976e-02A M=1.236e-06
I5365 0 n5366 2.976e-02A M=2.400e-06
I5366 0 n5367 2.976e-02A M=1.760e-06
I5367 0 n5368 2.976e-02A M=6.904e-08
I5368 0 n5369 2.976e-02A M=1.772e-07
I5369 0 n5370 2.976e-02A M=8.096e-07
I5370 0 n5371 2.976e-02A M=2.098e-06
I5371 0 n5372 2.976e-02A M=8.861e-07
I5372 0 n5373 2.976e-02A M=1.494e-06
I5373 0 n5374 2.976e-02A M=6.265e-07
I5374 0 n5375 2.976e-02A M=2.348e-06
I5375 0 n5376 2.976e-02A M=5.884e-07
I5376 0 n5377 2.976e-02A M=1.762e-07
I5377 0 n5378 2.976e-02A M=5.182e-07
I5378 0 n5379 2.976e-02A M=8.774e-07
I5379 0 n5380 2.976e-02A M=1.027e-06
I5380 0 n5381 2.976e-02A M=4.558e-07
I5381 0 n5382 2.976e-02A M=7.521e-07
I5382 0 n5383 2.976e-02A M=6.567e-07
I5383 0 n5384 2.976e-02A M=9.371e-07
I5384 0 n5385 2.976e-02A M=2.434e-06
I5385 0 n5386 2.976e-02A M=7.716e-07
I5386 0 n5387 2.976e-02A M=6.949e-07
I5387 0 n5388 2.976e-02A M=1.036e-06
I5388 0 n5389 2.976e-02A M=9.503e-07
I5389 0 n5390 2.976e-02A M=7.684e-07
I5390 0 n5391 2.976e-02A M=2.349e-06
I5391 0 n5392 2.976e-02A M=9.470e-07
I5392 0 n5393 2.976e-02A M=4.759e-07
I5393 0 n5394 2.976e-02A M=6.734e-07
I5394 0 n5395 2.976e-02A M=5.288e-07
I5395 0 n5396 2.976e-02A M=7.910e-07
I5396 0 n5397 2.976e-02A M=5.639e-07
I5397 0 n5398 2.976e-02A M=8.941e-07
I5398 0 n5399 2.976e-02A M=3.689e-07
I5399 0 n5400 2.976e-02A M=9.194e-07
I5400 0 n5401 2.976e-02A M=1.105e-06
I5401 0 n5402 2.976e-02A M=2.506e-06
I5402 0 n5403 2.976e-02A M=2.284e-06
I5403 0 n5404 2.976e-02A M=1.371e-06
I5404 0 n5405 2.976e-02A M=5.407e-07
I5405 0 n5406 2.976e-02A M=1.207e-06
I5406 0 n5407 2.976e-02A M=1.161e-06
I5407 0 n5408 2.976e-02A M=7.868e-07
I5408 0 n5409 2.976e-02A M=8.129e-07
I5409 0 n5410 2.976e-02A M=1.307e-06
I5410 0 n5411 2.976e-02A M=1.326e-06
I5411 0 n5412 2.976e-02A M=1.189e-06
I5412 0 n5413 2.976e-02A M=3.866e-07
I5413 0 n5414 2.976e-02A M=1.176e-06
I5414 0 n5415 2.976e-02A M=1.427e-06
I5415 0 n5416 2.976e-02A M=1.846e-07
I5416 0 n5417 2.976e-02A M=7.639e-07
I5417 0 n5418 2.976e-02A M=7.399e-07
I5418 0 n5419 2.976e-02A M=2.045e-06
I5419 0 n5420 2.976e-02A M=1.555e-06
I5420 0 n5421 2.976e-02A M=8.036e-07
I5421 0 n5422 2.976e-02A M=4.920e-07
I5422 0 n5423 2.976e-02A M=5.411e-07
I5423 0 n5424 2.976e-02A M=7.185e-07
I5424 0 n5425 2.976e-02A M=4.957e-07
I5425 0 n5426 2.976e-02A M=5.996e-07
I5426 0 n5427 2.976e-02A M=1.281e-06
I5427 0 n5428 2.976e-02A M=1.467e-06
I5428 0 n5429 2.976e-02A M=9.382e-07
I5429 0 n5430 2.976e-02A M=6.983e-07
I5430 0 n5431 2.976e-02A M=1.168e-06
I5431 0 n5432 2.976e-02A M=1.242e-06
I5432 0 n5433 2.976e-02A M=1.219e-06
I5433 0 n5434 2.976e-02A M=1.208e-06
I5434 0 n5435 2.976e-02A M=5.811e-07
I5435 0 n5436 2.976e-02A M=8.932e-07
I5436 0 n5437 2.976e-02A M=1.111e-06
I5437 0 n5438 2.976e-02A M=1.640e-06
I5438 0 n5439 2.976e-02A M=5.352e-07
I5439 0 n5440 2.976e-02A M=2.452e-06
I5440 0 n5441 2.976e-02A M=3.886e-07
I5441 0 n5442 2.976e-02A M=9.856e-07
I5442 0 n5443 2.976e-02A M=1.556e-06
I5443 0 n5444 2.976e-02A M=1.191e-06
I5444 0 n5445 2.976e-02A M=4.370e-07
I5445 0 n5446 2.976e-02A M=8.786e-07
I5446 0 n5447 2.976e-02A M=8.432e-07
I5447 0 n5448 2.976e-02A M=6.067e-07
I5448 0 n5449 2.976e-02A M=1.462e-06
I5449 0 n5450 2.976e-02A M=7.166e-07
I5450 0 n5451 2.976e-02A M=3.072e-07
I5451 0 n5452 2.976e-02A M=1.574e-06
I5452 0 n5453 2.976e-02A M=9.093e-07
I5453 0 n5454 2.976e-02A M=2.891e-06
I5454 0 n5455 2.976e-02A M=7.072e-07
I5455 0 n5456 2.976e-02A M=1.291e-06
I5456 0 n5457 2.976e-02A M=1.569e-06
I5457 0 n5458 2.976e-02A M=1.815e-06
I5458 0 n5459 2.976e-02A M=1.368e-06
I5459 0 n5460 2.976e-02A M=6.825e-07
I5460 0 n5461 2.976e-02A M=5.995e-07
I5461 0 n5462 2.976e-02A M=1.598e-06
I5462 0 n1 2.976e-02A M=7.589e-07
I5463 0 n5464 2.976e-02A M=1.031e-06
I5464 0 n5465 2.976e-02A M=8.655e-07
I5465 0 n5466 2.976e-02A M=7.245e-07
I5466 0 n5467 2.976e-02A M=1.012e-06
I5467 0 n5468 2.976e-02A M=1.103e-06
I5468 0 n5469 2.976e-02A M=1.143e-06
I5469 0 n5470 2.976e-02A M=8.380e-07
I5470 0 n5471 2.976e-02A M=1.209e-06
I5471 0 n5472 2.976e-02A M=3.073e-07
I5472 0 n5473 2.976e-02A M=9.071e-07
I5473 0 n5474 2.976e-02A M=4.829e-07
I5474 0 n5475 2.976e-02A M=3.433e-07
I5475 0 n5476 2.976e-02A M=4.926e-07
I5476 0 n5477 2.976e-02A M=5.980e-07
I5477 0 n5478 2.976e-02A M=1.149e-06
I5478 0 n5479 2.976e-02A M=8.801e-07
I5479 0 n5480 2.976e-02A M=5.020e-07
I5480 0 n5481 2.976e-02A M=9.801e-07
I5481 0 n5482 2.976e-02A M=1.056e-06
I5482 0 n5483 2.976e-02A M=1.001e-06
I5483 0 n5484 2.976e-02A M=1.369e-06
I5484 0 n5485 2.976e-02A M=9.767e-07
I5485 0 n5486 2.976e-02A M=5.177e-07
I5486 0 n5487 2.976e-02A M=6.527e-07
I5487 0 n5488 2.976e-02A M=1.491e-06
I5488 0 n5489 2.976e-02A M=1.394e-06
I5489 0 n5490 2.976e-02A M=1.196e-06
I5490 0 n5491 2.976e-02A M=7.104e-07
I5491 0 n5492 2.976e-02A M=1.188e-06
I5492 0 n5493 2.976e-02A M=3.055e-07
I5493 0 n5494 2.976e-02A M=5.677e-07
I5494 0 n5495 2.976e-02A M=1.255e-06
I5495 0 n5496 2.976e-02A M=3.502e-07
I5496 0 n5497 2.976e-02A M=9.397e-07
I5497 0 n5498 2.976e-02A M=1.303e-06
I5498 0 n5499 2.976e-02A M=3.181e-06
I5499 0 n5500 2.976e-02A M=1.434e-06
I5500 0 n5501 2.976e-02A M=9.352e-07
I5501 0 n5502 2.976e-02A M=4.204e-07
I5502 0 n5503 2.976e-02A M=8.260e-07
I5503 0 n1 2.976e-02A M=5.417e-07
I5504 0 n5505 2.976e-02A M=2.153e-06
I5505 0 n5506 2.976e-02A M=2.956e-07
I5506 0 n5507 2.976e-02A M=1.670e-06
I5507 0 n5508 2.976e-02A M=7.773e-07
I5508 0 n5509 2.976e-02A M=7.023e-07
I5509 0 n5510 2.976e-02A M=4.563e-07
I5510 0 n5511 2.976e-02A M=8.592e-07
I5511 0 n5512 2.976e-02A M=5.534e-07
I5512 0 n5513 2.976e-02A M=6.994e-07
I5513 0 n5514 2.976e-02A M=1.165e-06
I5514 0 n5515 2.976e-02A M=1.376e-06
I5515 0 n5516 2.976e-02A M=2.477e-06
I5516 0 n5517 2.976e-02A M=6.183e-07
I5517 0 n5518 2.976e-02A M=6.515e-07
I5518 0 n5519 2.976e-02A M=7.284e-07
I5519 0 n5520 2.976e-02A M=1.541e-06
I5520 0 n5521 2.976e-02A M=1.510e-06
I5521 0 n5522 2.976e-02A M=1.160e-06
I5522 0 n5523 2.976e-02A M=8.133e-07
I5523 0 n1 2.976e-02A M=3.191e-07
I5524 0 n5525 2.976e-02A M=7.955e-07
I5525 0 n5526 2.976e-02A M=6.398e-07
I5526 0 n5527 2.976e-02A M=2.069e-06
I5527 0 n5528 2.976e-02A M=1.124e-06
I5528 0 n5529 2.976e-02A M=6.838e-07
I5529 0 n5530 2.976e-02A M=5.466e-07
I5530 0 n5531 2.976e-02A M=5.453e-07
I5531 0 n5532 2.976e-02A M=2.404e-06
I5532 0 n5533 2.976e-02A M=1.018e-06
I5533 0 n5534 2.976e-02A M=6.538e-07
I5534 0 n5535 2.976e-02A M=9.133e-07
I5535 0 n5536 2.976e-02A M=6.155e-07
I5536 0 n5537 2.976e-02A M=6.219e-07
I5537 0 n5538 2.976e-02A M=6.797e-07
I5538 0 n5539 2.976e-02A M=4.600e-07
I5539 0 n5540 2.976e-02A M=8.972e-07
I5540 0 n5541 2.976e-02A M=6.791e-07
I5541 0 n5542 2.976e-02A M=9.833e-07
I5542 0 n5543 2.976e-02A M=1.333e-06
I5543 0 n5544 2.976e-02A M=9.160e-07
I5544 0 n5545 2.976e-02A M=1.663e-06
I5545 0 n5546 2.976e-02A M=1.809e-06
I5546 0 n5547 2.976e-02A M=1.387e-06
I5547 0 n5548 2.976e-02A M=1.445e-06
I5548 0 n5549 2.976e-02A M=1.045e-06
I5549 0 n5550 2.976e-02A M=4.297e-07
I5550 0 n5551 2.976e-02A M=1.577e-06
I5551 0 n5552 2.976e-02A M=6.999e-07
I5552 0 n5553 2.976e-02A M=1.385e-06
I5553 0 n5554 2.976e-02A M=1.104e-06
I5554 0 n5555 2.976e-02A M=1.336e-06
I5555 0 n5556 2.976e-02A M=7.614e-07
I5556 0 n5557 2.976e-02A M=9.728e-07
I5557 0 n5558 2.976e-02A M=2.814e-06
I5558 0 n5559 2.976e-02A M=8.780e-07
I5559 0 n5560 2.976e-02A M=1.331e-06
I5560 0 n5561 2.976e-02A M=5.211e-07
I5561 0 n5562 2.976e-02A M=5.382e-07
I5562 0 n5563 2.976e-02A M=1.141e-06
I5563 0 n5564 2.976e-02A M=1.846e-06
I5564 0 n5565 2.976e-02A M=1.577e-06
I5565 0 n5566 2.976e-02A M=5.229e-07
I5566 0 n5567 2.976e-02A M=6.791e-07
I5567 0 n5568 2.976e-02A M=4.545e-07
I5568 0 n5569 2.976e-02A M=6.619e-07
I5569 0 n5570 2.976e-02A M=8.432e-07
I5570 0 n1 2.976e-02A M=2.994e-07
I5571 0 n5572 2.976e-02A M=1.733e-06
I5572 0 n5573 2.976e-02A M=1.706e-06
I5573 0 n5574 2.976e-02A M=8.488e-07
I5574 0 n5575 2.976e-02A M=1.342e-06
I5575 0 n5576 2.976e-02A M=1.296e-06
I5576 0 n5577 2.976e-02A M=1.460e-06
I5577 0 n5578 2.976e-02A M=7.540e-07
I5578 0 n5579 2.976e-02A M=5.345e-07
I5579 0 n5580 2.976e-02A M=5.001e-07
I5580 0 n5581 2.976e-02A M=1.115e-06
I5581 0 n5582 2.976e-02A M=7.876e-07
I5582 0 n5583 2.976e-02A M=1.537e-06
I5583 0 n5584 2.976e-02A M=4.665e-07
I5584 0 n5585 2.976e-02A M=1.319e-06
I5585 0 n5586 2.976e-02A M=8.413e-07
I5586 0 n5587 2.976e-02A M=1.448e-06
I5587 0 n5588 2.976e-02A M=7.847e-07
I5588 0 n5589 2.976e-02A M=2.008e-06
I5589 0 n5590 2.976e-02A M=6.705e-07
I5590 0 n5591 2.976e-02A M=1.168e-06
I5591 0 n5592 2.976e-02A M=1.038e-06
I5592 0 n5593 2.976e-02A M=1.961e-06
I5593 0 n5594 2.976e-02A M=1.069e-06
I5594 0 n5595 2.976e-02A M=1.100e-06
I5595 0 n5596 2.976e-02A M=4.956e-07
I5596 0 n5597 2.976e-02A M=3.639e-07
I5597 0 n5598 2.976e-02A M=1.180e-06
I5598 0 n5599 2.976e-02A M=9.677e-07
I5599 0 n5600 2.976e-02A M=1.276e-06
I5600 0 n5601 2.976e-02A M=1.326e-06
I5601 0 n5602 2.976e-02A M=4.969e-07
I5602 0 n1 2.976e-02A M=1.445e-06
I5603 0 n5604 2.976e-02A M=8.921e-07
I5604 0 n5605 2.976e-02A M=3.784e-07
I5605 0 n5606 2.976e-02A M=6.814e-07
I5606 0 n5607 2.976e-02A M=1.066e-06
I5607 0 n5608 2.976e-02A M=9.867e-07
I5608 0 n5609 2.976e-02A M=7.303e-07
I5609 0 n5610 2.976e-02A M=6.324e-07
I5610 0 n5611 2.976e-02A M=2.216e-06
I5611 0 n5612 2.976e-02A M=7.338e-07
I5612 0 n5613 2.976e-02A M=1.517e-07
I5613 0 n5614 2.976e-02A M=8.546e-07
I5614 0 n5615 2.976e-02A M=4.042e-07
I5615 0 n5616 2.976e-02A M=6.246e-07
I5616 0 n5617 2.976e-02A M=1.352e-06
I5617 0 n5618 2.976e-02A M=6.086e-07
I5618 0 n5619 2.976e-02A M=1.441e-06
I5619 0 n5620 2.976e-02A M=9.208e-07
I5620 0 n5621 2.976e-02A M=8.983e-07
I5621 0 n5622 2.976e-02A M=4.745e-07
I5622 0 n5623 2.976e-02A M=8.279e-07
I5623 0 n5624 2.976e-02A M=9.148e-07
I5624 0 n5625 2.976e-02A M=7.702e-07
I5625 0 n5626 2.976e-02A M=3.516e-07
I5626 0 n5627 2.976e-02A M=4.677e-07
I5627 0 n5628 2.976e-02A M=1.352e-06
I5628 0 n5629 2.976e-02A M=1.309e-06
I5629 0 n5630 2.976e-02A M=1.005e-06
I5630 0 n5631 2.976e-02A M=6.823e-07
I5631 0 n5632 2.976e-02A M=2.502e-07
I5632 0 n5633 2.976e-02A M=8.812e-07
I5633 0 n5634 2.976e-02A M=1.249e-06
I5634 0 n5635 2.976e-02A M=1.814e-06
I5635 0 n5636 2.976e-02A M=9.676e-07
I5636 0 n5637 2.976e-02A M=1.484e-06
I5637 0 n5638 2.976e-02A M=3.627e-07
I5638 0 n5639 2.976e-02A M=9.678e-07
I5639 0 n5640 2.976e-02A M=6.474e-07
I5640 0 n5641 2.976e-02A M=9.367e-07
I5641 0 n5642 2.976e-02A M=7.925e-07
I5642 0 n5643 2.976e-02A M=1.395e-06
I5643 0 n5644 2.976e-02A M=1.065e-06
I5644 0 n5645 2.976e-02A M=4.934e-07
I5645 0 n5646 2.976e-02A M=3.291e-07
I5646 0 n5647 2.976e-02A M=2.310e-07
I5647 0 n5648 2.976e-02A M=4.196e-07
I5648 0 n5649 2.976e-02A M=5.361e-07
I5649 0 n5650 2.976e-02A M=1.717e-06
I5650 0 n5651 2.976e-02A M=7.728e-07
I5651 0 n5652 2.976e-02A M=5.324e-07
I5652 0 n5653 2.976e-02A M=7.774e-07
I5653 0 n5654 2.976e-02A M=7.579e-07
I5654 0 n5655 2.976e-02A M=7.718e-07
I5655 0 n5656 2.976e-02A M=5.293e-07
I5656 0 n5657 2.976e-02A M=2.018e-06
I5657 0 n5658 2.976e-02A M=1.589e-06
I5658 0 n5659 2.976e-02A M=8.850e-07
I5659 0 n5660 2.976e-02A M=1.835e-06
I5660 0 n5661 2.976e-02A M=2.302e-06
I5661 0 n5662 2.976e-02A M=1.110e-06
I5662 0 n5663 2.976e-02A M=4.376e-07
I5663 0 n5664 2.976e-02A M=9.806e-07
I5664 0 n5665 2.976e-02A M=1.523e-06
I5665 0 n5666 2.976e-02A M=1.196e-06
I5666 0 n5667 2.976e-02A M=1.091e-06
I5667 0 n5668 2.976e-02A M=6.100e-07
I5668 0 n5669 2.976e-02A M=1.634e-06
I5669 0 n5670 2.976e-02A M=1.471e-06
I5670 0 n5671 2.976e-02A M=9.254e-07
I5671 0 n5672 2.976e-02A M=5.075e-07
I5672 0 n5673 2.976e-02A M=8.763e-07
I5673 0 n5674 2.976e-02A M=9.733e-07
I5674 0 n5675 2.976e-02A M=1.407e-06
I5675 0 n5676 2.976e-02A M=9.768e-07
I5676 0 n5677 2.976e-02A M=5.402e-07
I5677 0 n5678 2.976e-02A M=1.343e-06
I5678 0 n5679 2.976e-02A M=9.556e-07
I5679 0 n5680 2.976e-02A M=6.862e-07
I5680 0 n5681 2.976e-02A M=8.392e-07
I5681 0 n5682 2.976e-02A M=7.882e-07
I5682 0 n5683 2.976e-02A M=7.303e-07
I5683 0 n5684 2.976e-02A M=2.869e-07
I5684 0 n5685 2.976e-02A M=1.136e-06
I5685 0 n5686 2.976e-02A M=1.802e-07
I5686 0 n5687 2.976e-02A M=2.626e-06
I5687 0 n5688 2.976e-02A M=4.972e-07
I5688 0 n5689 2.976e-02A M=2.957e-07
I5689 0 n5690 2.976e-02A M=2.744e-06
I5690 0 n5691 2.976e-02A M=6.076e-07
I5691 0 n5692 2.976e-02A M=7.112e-07
I5692 0 n5693 2.976e-02A M=5.852e-07
I5693 0 n5694 2.976e-02A M=1.536e-06
I5694 0 n5695 2.976e-02A M=1.087e-06
I5695 0 n5696 2.976e-02A M=7.048e-07
I5696 0 n5697 2.976e-02A M=3.201e-07
I5697 0 n5698 2.976e-02A M=6.198e-07
I5698 0 n5699 2.976e-02A M=8.441e-07
I5699 0 n5700 2.976e-02A M=1.756e-06
I5700 0 n5701 2.976e-02A M=1.599e-06
I5701 0 n5702 2.976e-02A M=1.222e-06
I5702 0 n5703 2.976e-02A M=2.066e-06
I5703 0 n5704 2.976e-02A M=6.806e-07
I5704 0 n5705 2.976e-02A M=5.343e-07
I5705 0 n5706 2.976e-02A M=3.088e-07
I5706 0 n5707 2.976e-02A M=1.571e-06
I5707 0 n1 2.976e-02A M=3.653e-07
I5708 0 n5709 2.976e-02A M=4.882e-07
I5709 0 n5710 2.976e-02A M=1.516e-06
I5710 0 n5711 2.976e-02A M=2.485e-07
I5711 0 n5712 2.976e-02A M=4.497e-07
I5712 0 n5713 2.976e-02A M=1.633e-06
I5713 0 n5714 2.976e-02A M=1.865e-06
I5714 0 n5715 2.976e-02A M=1.613e-06
I5715 0 n5716 2.976e-02A M=6.100e-07
I5716 0 n5717 2.976e-02A M=9.517e-07
I5717 0 n5718 2.976e-02A M=6.287e-07
I5718 0 n5719 2.976e-02A M=1.092e-06
I5719 0 n5720 2.976e-02A M=3.753e-07
I5720 0 n5721 2.976e-02A M=9.269e-07
I5721 0 n5722 2.976e-02A M=8.185e-07
I5722 0 n5723 2.976e-02A M=1.600e-06
I5723 0 n5724 2.976e-02A M=7.491e-08
I5724 0 n5725 2.976e-02A M=8.243e-07
I5725 0 n5726 2.976e-02A M=9.301e-07
I5726 0 n5727 2.976e-02A M=2.606e-07
I5727 0 n5728 2.976e-02A M=5.763e-07
I5728 0 n5729 2.976e-02A M=1.192e-06
I5729 0 n5730 2.976e-02A M=1.084e-06
I5730 0 n5731 2.976e-02A M=8.984e-07
I5731 0 n5732 2.976e-02A M=2.472e-07
I5732 0 n5733 2.976e-02A M=8.375e-07
I5733 0 n5734 2.976e-02A M=5.209e-07
I5734 0 n5735 2.976e-02A M=7.979e-07
I5735 0 n5736 2.976e-02A M=1.354e-06
I5736 0 n5737 2.976e-02A M=1.391e-06
I5737 0 n5738 2.976e-02A M=1.469e-06
I5738 0 n5739 2.976e-02A M=5.304e-07
I5739 0 n5740 2.976e-02A M=4.282e-07
I5740 0 n5741 2.976e-02A M=1.202e-06
I5741 0 n5742 2.976e-02A M=5.365e-07
I5742 0 n5743 2.976e-02A M=8.106e-07
I5743 0 n5744 2.976e-02A M=1.441e-06
I5744 0 n5745 2.976e-02A M=4.367e-07
I5745 0 n5746 2.976e-02A M=1.802e-06
I5746 0 n5747 2.976e-02A M=2.020e-06
I5747 0 n5748 2.976e-02A M=9.502e-07
I5748 0 n5749 2.976e-02A M=1.548e-06
I5749 0 n5750 2.976e-02A M=5.643e-07
I5750 0 n5751 2.976e-02A M=4.087e-07
I5751 0 n5752 2.976e-02A M=1.127e-06
I5752 0 n5753 2.976e-02A M=5.888e-07
I5753 0 n5754 2.976e-02A M=1.886e-06
I5754 0 n5755 2.976e-02A M=2.997e-07
I5755 0 n5756 2.976e-02A M=7.040e-07
I5756 0 n5757 2.976e-02A M=1.480e-06
I5757 0 n5758 2.976e-02A M=9.274e-07
I5758 0 n5759 2.976e-02A M=1.091e-06
I5759 0 n5760 2.976e-02A M=9.908e-07
I5760 0 n5761 2.976e-02A M=7.545e-07
I5761 0 n5762 2.976e-02A M=2.226e-06
I5762 0 n5763 2.976e-02A M=6.223e-07
I5763 0 n5764 2.976e-02A M=5.412e-07
I5764 0 n5765 2.976e-02A M=1.073e-07
I5765 0 n5766 2.976e-02A M=7.808e-07
I5766 0 n5767 2.976e-02A M=9.668e-07
I5767 0 n5768 2.976e-02A M=2.168e-07
I5768 0 n5769 2.976e-02A M=3.047e-07
I5769 0 n5770 2.976e-02A M=1.494e-06
I5770 0 n5771 2.976e-02A M=1.696e-06
I5771 0 n5772 2.976e-02A M=1.032e-06
I5772 0 n5773 2.976e-02A M=6.535e-07
I5773 0 n5774 2.976e-02A M=7.477e-07
I5774 0 n5775 2.976e-02A M=2.059e-07
I5775 0 n5776 2.976e-02A M=5.453e-07
I5776 0 n5777 2.976e-02A M=3.987e-07
I5777 0 n5778 2.976e-02A M=1.159e-06
I5778 0 n5779 2.976e-02A M=1.162e-06
I5779 0 n5780 2.976e-02A M=3.714e-07
I5780 0 n5781 2.976e-02A M=4.329e-07
I5781 0 n5782 2.976e-02A M=5.782e-07
I5782 0 n5783 2.976e-02A M=3.619e-07
I5783 0 n5784 2.976e-02A M=1.104e-06
I5784 0 n5785 2.976e-02A M=9.505e-07
I5785 0 n5786 2.976e-02A M=1.170e-06
I5786 0 n5787 2.976e-02A M=1.532e-06
I5787 0 n5788 2.976e-02A M=8.691e-07
I5788 0 n5789 2.976e-02A M=1.754e-06
I5789 0 n5790 2.976e-02A M=9.321e-07
I5790 0 n5791 2.976e-02A M=1.749e-06
I5791 0 n5792 2.976e-02A M=1.051e-06
I5792 0 n5793 2.976e-02A M=6.825e-07
I5793 0 n5794 2.976e-02A M=1.389e-06
I5794 0 n5795 2.976e-02A M=1.418e-06
I5795 0 n5796 2.976e-02A M=9.042e-07
I5796 0 n5797 2.976e-02A M=1.181e-06
I5797 0 n5798 2.976e-02A M=2.137e-06
I5798 0 n5799 2.976e-02A M=8.245e-07
I5799 0 n5800 2.976e-02A M=1.181e-06
I5800 0 n5801 2.976e-02A M=5.116e-07
I5801 0 n5802 2.976e-02A M=5.745e-07
I5802 0 n5803 2.976e-02A M=4.088e-07
I5803 0 n5804 2.976e-02A M=7.103e-07
I5804 0 n5805 2.976e-02A M=1.962e-06
I5805 0 n5806 2.976e-02A M=1.530e-06
I5806 0 n5807 2.976e-02A M=1.520e-06
I5807 0 n5808 2.976e-02A M=1.107e-06
I5808 0 n5809 2.976e-02A M=1.366e-06
I5809 0 n5810 2.976e-02A M=4.332e-07
I5810 0 n5811 2.976e-02A M=4.474e-07
I5811 0 n5812 2.976e-02A M=8.070e-07
I5812 0 n5813 2.976e-02A M=3.197e-07
I5813 0 n5814 2.976e-02A M=6.854e-07
I5814 0 n5815 2.976e-02A M=6.664e-07
I5815 0 n5816 2.976e-02A M=4.168e-07
I5816 0 n5817 2.976e-02A M=1.405e-06
I5817 0 n5818 2.976e-02A M=1.825e-06
I5818 0 n5819 2.976e-02A M=1.978e-06
I5819 0 n5820 2.976e-02A M=1.613e-06
I5820 0 n5821 2.976e-02A M=1.039e-06
I5821 0 n5822 2.976e-02A M=1.048e-06
I5822 0 n5823 2.976e-02A M=7.762e-07
I5823 0 n5824 2.976e-02A M=5.464e-07
I5824 0 n5825 2.976e-02A M=2.096e-06
I5825 0 n5826 2.976e-02A M=2.287e-07
I5826 0 n5827 2.976e-02A M=1.415e-06
I5827 0 n5828 2.976e-02A M=9.594e-07
I5828 0 n5829 2.976e-02A M=8.186e-07
I5829 0 n5830 2.976e-02A M=1.723e-06
I5830 0 n5831 2.976e-02A M=2.427e-07
I5831 0 n5832 2.976e-02A M=1.653e-06
I5832 0 n5833 2.976e-02A M=1.894e-06
I5833 0 n5834 2.976e-02A M=2.374e-06
I5834 0 n5835 2.976e-02A M=3.895e-07
I5835 0 n5836 2.976e-02A M=5.180e-07
I5836 0 n5837 2.976e-02A M=9.015e-07
I5837 0 n5838 2.976e-02A M=6.468e-07
I5838 0 n5839 2.976e-02A M=1.327e-06
I5839 0 n5840 2.976e-02A M=9.656e-07
I5840 0 n5841 2.976e-02A M=5.730e-07
I5841 0 n5842 2.976e-02A M=1.673e-06
I5842 0 n5843 2.976e-02A M=1.038e-06
I5843 0 n5844 2.976e-02A M=1.590e-06
I5844 0 n5845 2.976e-02A M=1.027e-06
I5845 0 n5846 2.976e-02A M=1.815e-06
I5846 0 n5847 2.976e-02A M=1.006e-06
I5847 0 n5848 2.976e-02A M=1.988e-06
I5848 0 n5849 2.976e-02A M=9.804e-07
I5849 0 n5850 2.976e-02A M=1.605e-06
I5850 0 n5851 2.976e-02A M=8.210e-07
I5851 0 n5852 2.976e-02A M=1.379e-06
I5852 0 n5853 2.976e-02A M=1.937e-07
I5853 0 n5854 2.976e-02A M=1.036e-06
I5854 0 n5855 2.976e-02A M=1.080e-06
I5855 0 n5856 2.976e-02A M=4.808e-07
I5856 0 n5857 2.976e-02A M=9.662e-07
I5857 0 n5858 2.976e-02A M=1.009e-06
I5858 0 n5859 2.976e-02A M=1.559e-06
I5859 0 n5860 2.976e-02A M=8.079e-08
I5860 0 n5861 2.976e-02A M=8.616e-07
I5861 0 n5862 2.976e-02A M=1.090e-06
I5862 0 n5863 2.976e-02A M=1.590e-06
I5863 0 n5864 2.976e-02A M=2.496e-06
I5864 0 n5865 2.976e-02A M=1.683e-06
I5865 0 n5866 2.976e-02A M=1.304e-06
I5866 0 n5867 2.976e-02A M=2.170e-06
I5867 0 n5868 2.976e-02A M=9.652e-07
I5868 0 n5869 2.976e-02A M=7.275e-07
I5869 0 n5870 2.976e-02A M=1.672e-06
I5870 0 n5871 2.976e-02A M=8.758e-07
I5871 0 n5872 2.976e-02A M=4.816e-07
I5872 0 n5873 2.976e-02A M=4.797e-07
I5873 0 n5874 2.976e-02A M=7.951e-07
I5874 0 n5875 2.976e-02A M=9.659e-07
I5875 0 n5876 2.976e-02A M=9.033e-07
I5876 0 n5877 2.976e-02A M=7.426e-07
I5877 0 n5878 2.976e-02A M=4.183e-07
I5878 0 n5879 2.976e-02A M=4.619e-07
I5879 0 n5880 2.976e-02A M=1.668e-06
I5880 0 n5881 2.976e-02A M=9.980e-07
I5881 0 n5882 2.976e-02A M=1.551e-06
I5882 0 n5883 2.976e-02A M=1.524e-06
I5883 0 n5884 2.976e-02A M=4.383e-07
I5884 0 n5885 2.976e-02A M=7.039e-07
I5885 0 n5886 2.976e-02A M=8.816e-07
I5886 0 n5887 2.976e-02A M=9.779e-07
I5887 0 n5888 2.976e-02A M=8.115e-07
I5888 0 n5889 2.976e-02A M=6.475e-07
I5889 0 n5890 2.976e-02A M=1.237e-06
I5890 0 n5891 2.976e-02A M=3.868e-07
I5891 0 n5892 2.976e-02A M=9.896e-07
I5892 0 n5893 2.976e-02A M=1.110e-06
I5893 0 n5894 2.976e-02A M=5.005e-07
I5894 0 n5895 2.976e-02A M=1.536e-06
I5895 0 n5896 2.976e-02A M=1.293e-06
I5896 0 n5897 2.976e-02A M=1.555e-06
I5897 0 n5898 2.976e-02A M=7.891e-07
I5898 0 n5899 2.976e-02A M=3.538e-07
I5899 0 n5900 2.976e-02A M=8.610e-07
I5900 0 n5901 2.976e-02A M=9.009e-07
I5901 0 n5902 2.976e-02A M=3.957e-07
I5902 0 n5903 2.976e-02A M=6.258e-07
I5903 0 n5904 2.976e-02A M=1.578e-06
I5904 0 n5905 2.976e-02A M=7.278e-07
I5905 0 n5906 2.976e-02A M=2.015e-07
I5906 0 n5907 2.976e-02A M=2.207e-06
I5907 0 n5908 2.976e-02A M=9.813e-07
I5908 0 n5909 2.976e-02A M=7.120e-07
I5909 0 n1 2.976e-02A M=1.027e-06
I5910 0 n5911 2.976e-02A M=1.136e-06
I5911 0 n5912 2.976e-02A M=5.802e-08
I5912 0 n5913 2.976e-02A M=7.248e-07
I5913 0 n5914 2.976e-02A M=1.781e-06
I5914 0 n5915 2.976e-02A M=1.388e-06
I5915 0 n5916 2.976e-02A M=8.736e-07
I5916 0 n5917 2.976e-02A M=2.169e-06
I5917 0 n5918 2.976e-02A M=8.338e-07
I5918 0 n5919 2.976e-02A M=1.016e-06
I5919 0 n5920 2.976e-02A M=1.279e-06
I5920 0 n5921 2.976e-02A M=8.514e-07
I5921 0 n5922 2.976e-02A M=1.455e-06
I5922 0 n5923 2.976e-02A M=5.314e-07
I5923 0 n5924 2.976e-02A M=4.059e-07
I5924 0 n5925 2.976e-02A M=6.819e-07
I5925 0 n5926 2.976e-02A M=9.849e-07
I5926 0 n5927 2.976e-02A M=1.376e-06
I5927 0 n5928 2.976e-02A M=3.215e-07
I5928 0 n5929 2.976e-02A M=6.784e-07
I5929 0 n5930 2.976e-02A M=2.686e-07
I5930 0 n5931 2.976e-02A M=1.146e-06
I5931 0 n5932 2.976e-02A M=1.684e-06
I5932 0 n1 2.976e-02A M=1.412e-06
I5933 0 n5934 2.976e-02A M=8.425e-07
I5934 0 n5935 2.976e-02A M=1.325e-06
I5935 0 n5936 2.976e-02A M=4.340e-07
I5936 0 n5937 2.976e-02A M=1.190e-06
I5937 0 n5938 2.976e-02A M=1.778e-06
I5938 0 n5939 2.976e-02A M=4.648e-07
I5939 0 n5940 2.976e-02A M=1.469e-06
I5940 0 n5941 2.976e-02A M=6.708e-07
I5941 0 n5942 2.976e-02A M=4.447e-07
I5942 0 n5943 2.976e-02A M=7.645e-07
I5943 0 n5944 2.976e-02A M=1.066e-06
I5944 0 n5945 2.976e-02A M=1.030e-06
I5945 0 n5946 2.976e-02A M=1.649e-06
I5946 0 n5947 2.976e-02A M=7.442e-07
I5947 0 n5948 2.976e-02A M=6.225e-07
I5948 0 n5949 2.976e-02A M=8.243e-07
I5949 0 n5950 2.976e-02A M=1.135e-06
I5950 0 n5951 2.976e-02A M=1.636e-06
I5951 0 n5952 2.976e-02A M=7.468e-07
I5952 0 n5953 2.976e-02A M=1.659e-06
I5953 0 n5954 2.976e-02A M=6.575e-07
I5954 0 n5955 2.976e-02A M=8.868e-07
I5955 0 n5956 2.976e-02A M=5.622e-07
I5956 0 n5957 2.976e-02A M=1.438e-06
I5957 0 n5958 2.976e-02A M=1.240e-06
I5958 0 n5959 2.976e-02A M=1.266e-06
I5959 0 n5960 2.976e-02A M=7.156e-07
I5960 0 n5961 2.976e-02A M=4.957e-07
I5961 0 n5962 2.976e-02A M=3.352e-06
I5962 0 n5963 2.976e-02A M=1.554e-06
I5963 0 n5964 2.976e-02A M=1.513e-06
I5964 0 n5965 2.976e-02A M=7.027e-07
I5965 0 n5966 2.976e-02A M=3.919e-07
I5966 0 n5967 2.976e-02A M=1.350e-06
I5967 0 n5968 2.976e-02A M=7.114e-07
I5968 0 n5969 2.976e-02A M=3.768e-07
I5969 0 n5970 2.976e-02A M=1.258e-06
I5970 0 n5971 2.976e-02A M=9.144e-07
I5971 0 n5972 2.976e-02A M=2.857e-06
I5972 0 n5973 2.976e-02A M=6.271e-07
I5973 0 n5974 2.976e-02A M=6.788e-07
I5974 0 n5975 2.976e-02A M=8.066e-07
I5975 0 n5976 2.976e-02A M=9.573e-07
I5976 0 n5977 2.976e-02A M=9.825e-07
I5977 0 n5978 2.976e-02A M=4.999e-07
I5978 0 n5979 2.976e-02A M=5.826e-07
I5979 0 n5980 2.976e-02A M=2.104e-06
I5980 0 n5981 2.976e-02A M=6.339e-07
I5981 0 n5982 2.976e-02A M=9.897e-07
I5982 0 n5983 2.976e-02A M=1.049e-06
I5983 0 n5984 2.976e-02A M=7.634e-07
I5984 0 n5985 2.976e-02A M=1.385e-06
I5985 0 n5986 2.976e-02A M=5.255e-07
I5986 0 n5987 2.976e-02A M=1.235e-06
I5987 0 n5988 2.976e-02A M=4.323e-07
I5988 0 n5989 2.976e-02A M=6.926e-07
I5989 0 n5990 2.976e-02A M=6.565e-07
I5990 0 n5991 2.976e-02A M=9.406e-07
I5991 0 n5992 2.976e-02A M=2.549e-07
I5992 0 n5993 2.976e-02A M=2.837e-07
I5993 0 n5994 2.976e-02A M=9.192e-07
I5994 0 n5995 2.976e-02A M=1.246e-06
I5995 0 n5996 2.976e-02A M=5.610e-07
I5996 0 n5997 2.976e-02A M=1.129e-06
I5997 0 n5998 2.976e-02A M=5.633e-07
I5998 0 n5999 2.976e-02A M=5.025e-07
I5999 0 n6000 2.976e-02A M=1.026e-06
I6000 0 n6001 2.976e-02A M=1.889e-06
I6001 0 n6002 2.976e-02A M=1.249e-06
I6002 0 n6003 2.976e-02A M=6.767e-07
I6003 0 n6004 2.976e-02A M=1.042e-06
I6004 0 n6005 2.976e-02A M=5.617e-07
I6005 0 n6006 2.976e-02A M=8.100e-07
I6006 0 n6007 2.976e-02A M=1.126e-06
I6007 0 n6008 2.976e-02A M=6.967e-07
I6008 0 n6009 2.976e-02A M=1.172e-07
I6009 0 n6010 2.976e-02A M=1.187e-06
I6010 0 n6011 2.976e-02A M=5.798e-07
I6011 0 n6012 2.976e-02A M=8.565e-07
I6012 0 n6013 2.976e-02A M=1.379e-06
I6013 0 n6014 2.976e-02A M=1.316e-06
I6014 0 n6015 2.976e-02A M=1.868e-06
I6015 0 n6016 2.976e-02A M=6.620e-07
I6016 0 n6017 2.976e-02A M=2.196e-07
I6017 0 n6018 2.976e-02A M=1.411e-06
I6018 0 n6019 2.976e-02A M=1.418e-06
I6019 0 n6020 2.976e-02A M=9.521e-07
I6020 0 n6021 2.976e-02A M=6.190e-07
I6021 0 n6022 2.976e-02A M=3.840e-07
I6022 0 n6023 2.976e-02A M=2.041e-06
I6023 0 n6024 2.976e-02A M=9.165e-07
I6024 0 n6025 2.976e-02A M=8.202e-07
I6025 0 n6026 2.976e-02A M=1.388e-07
I6026 0 n6027 2.976e-02A M=8.540e-07
I6027 0 n6028 2.976e-02A M=1.570e-06
I6028 0 n6029 2.976e-02A M=9.443e-07
I6029 0 n6030 2.976e-02A M=1.631e-06
I6030 0 n6031 2.976e-02A M=3.222e-07
I6031 0 n6032 2.976e-02A M=2.519e-06
I6032 0 n6033 2.976e-02A M=4.803e-07
I6033 0 n6034 2.976e-02A M=1.230e-06
I6034 0 n6035 2.976e-02A M=4.788e-07
I6035 0 n6036 2.976e-02A M=4.684e-07
I6036 0 n6037 2.976e-02A M=7.227e-07
I6037 0 n6038 2.976e-02A M=4.136e-07
I6038 0 n6039 2.976e-02A M=1.142e-06
I6039 0 n6040 2.976e-02A M=1.114e-06
I6040 0 n6041 2.976e-02A M=2.065e-06
I6041 0 n1 2.976e-02A M=8.357e-07
I6042 0 n6043 2.976e-02A M=1.373e-06
I6043 0 n6044 2.976e-02A M=3.447e-07
I6044 0 n6045 2.976e-02A M=1.635e-06
I6045 0 n6046 2.976e-02A M=2.996e-06
I6046 0 n6047 2.976e-02A M=1.065e-06
I6047 0 n6048 2.976e-02A M=6.173e-07
I6048 0 n6049 2.976e-02A M=1.036e-06
I6049 0 n6050 2.976e-02A M=2.196e-06
I6050 0 n6051 2.976e-02A M=9.337e-07
I6051 0 n6052 2.976e-02A M=6.564e-07
I6052 0 n6053 2.976e-02A M=5.446e-07
I6053 0 n6054 2.976e-02A M=2.421e-06
I6054 0 n6055 2.976e-02A M=7.790e-07
I6055 0 n6056 2.976e-02A M=3.390e-06
I6056 0 n6057 2.976e-02A M=1.084e-06
I6057 0 n6058 2.976e-02A M=1.258e-06
I6058 0 n6059 2.976e-02A M=7.069e-07
I6059 0 n6060 2.976e-02A M=8.453e-07
I6060 0 n6061 2.976e-02A M=9.155e-07
I6061 0 n6062 2.976e-02A M=1.425e-06
I6062 0 n6063 2.976e-02A M=1.001e-06
I6063 0 n6064 2.976e-02A M=1.081e-06
I6064 0 n6065 2.976e-02A M=9.849e-07
I6065 0 n6066 2.976e-02A M=8.879e-07
I6066 0 n6067 2.976e-02A M=1.224e-06
I6067 0 n6068 2.976e-02A M=6.146e-07
I6068 0 n6069 2.976e-02A M=4.282e-07
I6069 0 n6070 2.976e-02A M=5.767e-07
I6070 0 n6071 2.976e-02A M=5.539e-07
I6071 0 n6072 2.976e-02A M=3.303e-07
I6072 0 n6073 2.976e-02A M=2.834e-07
I6073 0 n6074 2.976e-02A M=8.939e-07
I6074 0 n6075 2.976e-02A M=6.740e-07
I6075 0 n6076 2.976e-02A M=1.740e-06
I6076 0 n6077 2.976e-02A M=5.105e-07
I6077 0 n6078 2.976e-02A M=1.300e-06
I6078 0 n6079 2.976e-02A M=9.511e-07
I6079 0 n6080 2.976e-02A M=8.584e-07
I6080 0 n6081 2.976e-02A M=7.585e-07
I6081 0 n6082 2.976e-02A M=1.507e-06
I6082 0 n6083 2.976e-02A M=3.761e-07
I6083 0 n6084 2.976e-02A M=4.884e-07
I6084 0 n6085 2.976e-02A M=3.524e-07
I6085 0 n6086 2.976e-02A M=6.899e-07
I6086 0 n6087 2.976e-02A M=1.593e-07
I6087 0 n6088 2.976e-02A M=1.010e-06
I6088 0 n6089 2.976e-02A M=8.431e-07
I6089 0 n6090 2.976e-02A M=7.542e-07
I6090 0 n6091 2.976e-02A M=1.059e-06
I6091 0 n6092 2.976e-02A M=9.565e-07
I6092 0 n6093 2.976e-02A M=1.870e-06
I6093 0 n6094 2.976e-02A M=5.695e-07
I6094 0 n6095 2.976e-02A M=8.721e-07
I6095 0 n6096 2.976e-02A M=1.934e-06
I6096 0 n6097 2.976e-02A M=9.766e-07
I6097 0 n6098 2.976e-02A M=9.305e-07
I6098 0 n6099 2.976e-02A M=1.063e-06
I6099 0 n6100 2.976e-02A M=6.594e-07
I6100 0 n6101 2.976e-02A M=8.897e-07
I6101 0 n6102 2.976e-02A M=3.187e-07
I6102 0 n6103 2.976e-02A M=1.136e-06
I6103 0 n6104 2.976e-02A M=1.429e-06
I6104 0 n6105 2.976e-02A M=8.522e-07
I6105 0 n6106 2.976e-02A M=4.150e-07
I6106 0 n6107 2.976e-02A M=4.474e-07
I6107 0 n6108 2.976e-02A M=4.624e-07
I6108 0 n6109 2.976e-02A M=1.302e-06
I6109 0 n6110 2.976e-02A M=8.057e-07
I6110 0 n6111 2.976e-02A M=1.223e-07
I6111 0 n6112 2.976e-02A M=1.637e-06
I6112 0 n6113 2.976e-02A M=1.714e-06
I6113 0 n6114 2.976e-02A M=7.786e-07
I6114 0 n6115 2.976e-02A M=7.114e-07
I6115 0 n6116 2.976e-02A M=2.549e-07
I6116 0 n6117 2.976e-02A M=1.735e-06
I6117 0 n6118 2.976e-02A M=5.700e-07
I6118 0 n6119 2.976e-02A M=8.047e-07
I6119 0 n1 2.976e-02A M=1.593e-06
I6120 0 n6121 2.976e-02A M=7.764e-07
I6121 0 n6122 2.976e-02A M=8.460e-07
I6122 0 n6123 2.976e-02A M=8.480e-07
I6123 0 n6124 2.976e-02A M=1.723e-06
I6124 0 n6125 2.976e-02A M=2.619e-07
I6125 0 n6126 2.976e-02A M=5.305e-07
I6126 0 n6127 2.976e-02A M=1.785e-06
I6127 0 n6128 2.976e-02A M=1.733e-06
I6128 0 n6129 2.976e-02A M=1.160e-06
I6129 0 n6130 2.976e-02A M=9.293e-07
I6130 0 n6131 2.976e-02A M=1.993e-06
I6131 0 n6132 2.976e-02A M=1.290e-06
I6132 0 n6133 2.976e-02A M=3.094e-06
I6133 0 n6134 2.976e-02A M=1.524e-06
I6134 0 n6135 2.976e-02A M=1.491e-06
I6135 0 n6136 2.976e-02A M=9.753e-07
I6136 0 n6137 2.976e-02A M=1.288e-06
I6137 0 n6138 2.976e-02A M=1.510e-06
I6138 0 n6139 2.976e-02A M=1.088e-06
I6139 0 n6140 2.976e-02A M=5.954e-07
I6140 0 n6141 2.976e-02A M=6.073e-07
I6141 0 n6142 2.976e-02A M=9.430e-07
I6142 0 n6143 2.976e-02A M=1.319e-06
I6143 0 n6144 2.976e-02A M=2.496e-07
I6144 0 n6145 2.976e-02A M=2.484e-07
I6145 0 n6146 2.976e-02A M=8.105e-07
I6146 0 n6147 2.976e-02A M=1.172e-06
I6147 0 n6148 2.976e-02A M=1.108e-06
I6148 0 n6149 2.976e-02A M=6.767e-07
I6149 0 n6150 2.976e-02A M=4.744e-07
I6150 0 n6151 2.976e-02A M=8.493e-07
I6151 0 n6152 2.976e-02A M=7.010e-07
I6152 0 n6153 2.976e-02A M=3.023e-07
I6153 0 n6154 2.976e-02A M=1.622e-06
I6154 0 n6155 2.976e-02A M=2.300e-06
I6155 0 n6156 2.976e-02A M=7.398e-07
I6156 0 n6157 2.976e-02A M=9.660e-07
I6157 0 n6158 2.976e-02A M=1.347e-06
I6158 0 n6159 2.976e-02A M=1.372e-06
I6159 0 n6160 2.976e-02A M=8.318e-07
I6160 0 n6161 2.976e-02A M=1.561e-06
I6161 0 n6162 2.976e-02A M=1.505e-06
I6162 0 n6163 2.976e-02A M=4.520e-07
I6163 0 n6164 2.976e-02A M=7.555e-07
I6164 0 n6165 2.976e-02A M=6.706e-07
I6165 0 n6166 2.976e-02A M=1.544e-06
I6166 0 n6167 2.976e-02A M=7.001e-07
I6167 0 n6168 2.976e-02A M=9.994e-07
I6168 0 n6169 2.976e-02A M=1.313e-06
I6169 0 n6170 2.976e-02A M=7.440e-07
I6170 0 n6171 2.976e-02A M=8.998e-07
I6171 0 n6172 2.976e-02A M=1.667e-06
I6172 0 n6173 2.976e-02A M=1.813e-06
I6173 0 n6174 2.976e-02A M=6.986e-07
I6174 0 n1 2.976e-02A M=6.605e-07
I6175 0 n6176 2.976e-02A M=5.889e-07
I6176 0 n6177 2.976e-02A M=6.479e-07
I6177 0 n6178 2.976e-02A M=9.661e-07
I6178 0 n6179 2.976e-02A M=1.413e-06
I6179 0 n6180 2.976e-02A M=6.165e-07
I6180 0 n6181 2.976e-02A M=4.764e-07
I6181 0 n6182 2.976e-02A M=7.710e-07
I6182 0 n6183 2.976e-02A M=6.853e-07
I6183 0 n6184 2.976e-02A M=6.425e-07
I6184 0 n6185 2.976e-02A M=1.322e-06
I6185 0 n6186 2.976e-02A M=1.497e-06
I6186 0 n6187 2.976e-02A M=1.239e-06
I6187 0 n6188 2.976e-02A M=9.959e-07
I6188 0 n6189 2.976e-02A M=1.967e-06
I6189 0 n6190 2.976e-02A M=1.549e-07
I6190 0 n6191 2.976e-02A M=6.373e-07
I6191 0 n6192 2.976e-02A M=2.731e-07
I6192 0 n6193 2.976e-02A M=1.261e-06
I6193 0 n6194 2.976e-02A M=1.641e-06
I6194 0 n6195 2.976e-02A M=2.120e-07
I6195 0 n6196 2.976e-02A M=3.348e-07
I6196 0 n6197 2.976e-02A M=4.663e-07
I6197 0 n6198 2.976e-02A M=1.368e-06
I6198 0 n6199 2.976e-02A M=1.099e-06
I6199 0 n6200 2.976e-02A M=6.262e-07
I6200 0 n6201 2.976e-02A M=9.603e-07
I6201 0 n6202 2.976e-02A M=7.031e-07
I6202 0 n6203 2.976e-02A M=6.485e-07
I6203 0 n6204 2.976e-02A M=7.716e-07
I6204 0 n6205 2.976e-02A M=1.424e-06
I6205 0 n6206 2.976e-02A M=5.646e-07
I6206 0 n6207 2.976e-02A M=1.587e-06
I6207 0 n6208 2.976e-02A M=1.205e-06
I6208 0 n6209 2.976e-02A M=1.291e-06
I6209 0 n6210 2.976e-02A M=4.979e-07
I6210 0 n6211 2.976e-02A M=1.328e-06
I6211 0 n6212 2.976e-02A M=1.404e-07
I6212 0 n6213 2.976e-02A M=8.239e-07
I6213 0 n6214 2.976e-02A M=1.014e-06
I6214 0 n6215 2.976e-02A M=6.344e-08
I6215 0 n6216 2.976e-02A M=2.822e-07
I6216 0 n6217 2.976e-02A M=1.748e-06
I6217 0 n6218 2.976e-02A M=2.595e-07
I6218 0 n6219 2.976e-02A M=1.665e-06
I6219 0 n6220 2.976e-02A M=8.980e-07
I6220 0 n6221 2.976e-02A M=1.583e-06
I6221 0 n6222 2.976e-02A M=4.543e-07
I6222 0 n6223 2.976e-02A M=8.112e-07
I6223 0 n6224 2.976e-02A M=1.561e-06
I6224 0 n6225 2.976e-02A M=1.577e-06
I6225 0 n6226 2.976e-02A M=1.181e-06
I6226 0 n6227 2.976e-02A M=1.170e-06
I6227 0 n6228 2.976e-02A M=1.299e-06
I6228 0 n6229 2.976e-02A M=5.158e-07
I6229 0 n6230 2.976e-02A M=1.768e-06
I6230 0 n6231 2.976e-02A M=4.372e-07
I6231 0 n6232 2.976e-02A M=2.532e-07
I6232 0 n6233 2.976e-02A M=1.042e-06
I6233 0 n6234 2.976e-02A M=1.838e-06
I6234 0 n6235 2.976e-02A M=1.381e-06
I6235 0 n6236 2.976e-02A M=4.102e-07
I6236 0 n6237 2.976e-02A M=6.637e-07
I6237 0 n6238 2.976e-02A M=1.692e-06
I6238 0 n6239 2.976e-02A M=1.408e-06
I6239 0 n6240 2.976e-02A M=6.966e-07
I6240 0 n6241 2.976e-02A M=1.802e-06
I6241 0 n6242 2.976e-02A M=1.082e-06
I6242 0 n6243 2.976e-02A M=1.553e-06
I6243 0 n6244 2.976e-02A M=1.064e-06
I6244 0 n6245 2.976e-02A M=1.128e-06
I6245 0 n6246 2.976e-02A M=1.169e-06
I6246 0 n6247 2.976e-02A M=1.388e-06
I6247 0 n6248 2.976e-02A M=1.154e-06
I6248 0 n6249 2.976e-02A M=8.186e-07
I6249 0 n6250 2.976e-02A M=8.047e-07
I6250 0 n6251 2.976e-02A M=1.177e-06
I6251 0 n6252 2.976e-02A M=2.321e-06
I6252 0 n6253 2.976e-02A M=2.161e-06
I6253 0 n6254 2.976e-02A M=1.361e-06
I6254 0 n6255 2.976e-02A M=1.595e-06
I6255 0 n6256 2.976e-02A M=1.536e-06
I6256 0 n6257 2.976e-02A M=5.306e-07
I6257 0 n6258 2.976e-02A M=9.960e-07
I6258 0 n6259 2.976e-02A M=1.342e-06
I6259 0 n6260 2.976e-02A M=1.720e-06
I6260 0 n6261 2.976e-02A M=8.745e-07
I6261 0 n6262 2.976e-02A M=6.743e-07
I6262 0 n6263 2.976e-02A M=1.887e-06
I6263 0 n6264 2.976e-02A M=1.165e-06
I6264 0 n6265 2.976e-02A M=6.028e-07
I6265 0 n6266 2.976e-02A M=8.434e-07
I6266 0 n6267 2.976e-02A M=1.225e-06
I6267 0 n6268 2.976e-02A M=1.150e-06
I6268 0 n6269 2.976e-02A M=4.561e-07
I6269 0 n6270 2.976e-02A M=7.159e-07
I6270 0 n6271 2.976e-02A M=9.907e-07
I6271 0 n6272 2.976e-02A M=1.057e-06
I6272 0 n6273 2.976e-02A M=1.247e-06
I6273 0 n6274 2.976e-02A M=1.319e-06
I6274 0 n6275 2.976e-02A M=5.935e-07
I6275 0 n6276 2.976e-02A M=8.640e-07
I6276 0 n6277 2.976e-02A M=1.415e-06
I6277 0 n6278 2.976e-02A M=1.595e-07
I6278 0 n6279 2.976e-02A M=8.679e-07
I6279 0 n6280 2.976e-02A M=8.710e-07
I6280 0 n6281 2.976e-02A M=1.268e-06
I6281 0 n6282 2.976e-02A M=5.187e-07
I6282 0 n6283 2.976e-02A M=6.978e-07
I6283 0 n6284 2.976e-02A M=2.658e-07
I6284 0 n6285 2.976e-02A M=1.202e-06
I6285 0 n6286 2.976e-02A M=8.817e-07
I6286 0 n6287 2.976e-02A M=1.033e-06
I6287 0 n6288 2.976e-02A M=6.443e-07
I6288 0 n6289 2.976e-02A M=1.495e-06
I6289 0 n6290 2.976e-02A M=1.090e-06
I6290 0 n6291 2.976e-02A M=3.304e-07
I6291 0 n6292 2.976e-02A M=2.475e-06
I6292 0 n6293 2.976e-02A M=9.661e-07
I6293 0 n6294 2.976e-02A M=1.310e-06
I6294 0 n6295 2.976e-02A M=1.608e-06
I6295 0 n6296 2.976e-02A M=4.479e-07
I6296 0 n6297 2.976e-02A M=8.873e-07
I6297 0 n6298 2.976e-02A M=1.355e-06
I6298 0 n6299 2.976e-02A M=1.626e-06
I6299 0 n6300 2.976e-02A M=7.928e-07
I6300 0 n6301 2.976e-02A M=5.500e-07
I6301 0 n6302 2.976e-02A M=6.839e-07
I6302 0 n6303 2.976e-02A M=1.515e-06
I6303 0 n6304 2.976e-02A M=2.581e-06
I6304 0 n6305 2.976e-02A M=3.297e-07
I6305 0 n6306 2.976e-02A M=8.101e-07
I6306 0 n6307 2.976e-02A M=1.722e-06
I6307 0 n6308 2.976e-02A M=9.768e-07
I6308 0 n6309 2.976e-02A M=4.683e-07
I6309 0 n6310 2.976e-02A M=1.379e-06
I6310 0 n6311 2.976e-02A M=1.545e-07
I6311 0 n6312 2.976e-02A M=9.597e-07
I6312 0 n6313 2.976e-02A M=2.889e-07
I6313 0 n6314 2.976e-02A M=1.479e-06
I6314 0 n6315 2.976e-02A M=1.266e-06
I6315 0 n6316 2.976e-02A M=1.122e-06
I6316 0 n6317 2.976e-02A M=9.791e-07
I6317 0 n6318 2.976e-02A M=1.115e-06
I6318 0 n6319 2.976e-02A M=1.448e-06
I6319 0 n6320 2.976e-02A M=9.281e-07
I6320 0 n6321 2.976e-02A M=1.212e-06
I6321 0 n6322 2.976e-02A M=1.793e-06
I6322 0 n6323 2.976e-02A M=1.809e-06
I6323 0 n6324 2.976e-02A M=6.341e-07
I6324 0 n6325 2.976e-02A M=1.094e-06
I6325 0 n6326 2.976e-02A M=1.128e-06
I6326 0 n6327 2.976e-02A M=8.110e-07
I6327 0 n6328 2.976e-02A M=8.565e-07
I6328 0 n6329 2.976e-02A M=1.816e-06
I6329 0 n6330 2.976e-02A M=1.558e-06
I6330 0 n6331 2.976e-02A M=9.532e-07
I6331 0 n6332 2.976e-02A M=5.541e-07
I6332 0 n6333 2.976e-02A M=9.980e-07
I6333 0 n6334 2.976e-02A M=2.334e-07
I6334 0 n6335 2.976e-02A M=1.111e-06
I6335 0 n6336 2.976e-02A M=1.168e-06
I6336 0 n6337 2.976e-02A M=7.384e-07
I6337 0 n6338 2.976e-02A M=3.182e-07
I6338 0 n6339 2.976e-02A M=1.190e-06
I6339 0 n6340 2.976e-02A M=7.563e-07
I6340 0 n6341 2.976e-02A M=2.392e-06
I6341 0 n6342 2.976e-02A M=1.482e-06
I6342 0 n1 2.976e-02A M=1.145e-06
I6343 0 n6344 2.976e-02A M=9.208e-07
I6344 0 n6345 2.976e-02A M=6.689e-07
I6345 0 n6346 2.976e-02A M=5.136e-07
I6346 0 n6347 2.976e-02A M=2.520e-06
I6347 0 n6348 2.976e-02A M=7.361e-07
I6348 0 n6349 2.976e-02A M=1.121e-06
I6349 0 n6350 2.976e-02A M=1.058e-06
I6350 0 n6351 2.976e-02A M=9.083e-07
I6351 0 n6352 2.976e-02A M=9.816e-07
I6352 0 n6353 2.976e-02A M=1.221e-06
I6353 0 n6354 2.976e-02A M=4.309e-07
I6354 0 n6355 2.976e-02A M=4.629e-07
I6355 0 n6356 2.976e-02A M=1.481e-06
I6356 0 n6357 2.976e-02A M=2.264e-06
I6357 0 n6358 2.976e-02A M=1.075e-06
I6358 0 n6359 2.976e-02A M=6.103e-07
I6359 0 n6360 2.976e-02A M=1.155e-06
I6360 0 n6361 2.976e-02A M=1.139e-06
I6361 0 n6362 2.976e-02A M=1.133e-06
I6362 0 n6363 2.976e-02A M=1.509e-06
I6363 0 n6364 2.976e-02A M=1.010e-06
I6364 0 n6365 2.976e-02A M=8.119e-07
I6365 0 n6366 2.976e-02A M=4.466e-07
I6366 0 n6367 2.976e-02A M=7.454e-07
I6367 0 n6368 2.976e-02A M=1.536e-06
I6368 0 n6369 2.976e-02A M=1.667e-06
I6369 0 n6370 2.976e-02A M=2.094e-06
I6370 0 n6371 2.976e-02A M=1.110e-06
I6371 0 n6372 2.976e-02A M=1.012e-06
I6372 0 n6373 2.976e-02A M=1.167e-06
I6373 0 n6374 2.976e-02A M=9.281e-07
I6374 0 n6375 2.976e-02A M=1.079e-06
I6375 0 n6376 2.976e-02A M=8.413e-07
I6376 0 n6377 2.976e-02A M=1.485e-06
I6377 0 n6378 2.976e-02A M=2.556e-07
I6378 0 n6379 2.976e-02A M=3.278e-07
I6379 0 n6380 2.976e-02A M=2.121e-06
I6380 0 n6381 2.976e-02A M=1.135e-06
I6381 0 n6382 2.976e-02A M=9.497e-07
I6382 0 n6383 2.976e-02A M=6.847e-07
I6383 0 n6384 2.976e-02A M=5.834e-07
I6384 0 n6385 2.976e-02A M=8.812e-07
I6385 0 n6386 2.976e-02A M=6.801e-07
I6386 0 n6387 2.976e-02A M=8.076e-07
I6387 0 n6388 2.976e-02A M=1.256e-06
I6388 0 n6389 2.976e-02A M=1.872e-06
I6389 0 n6390 2.976e-02A M=8.114e-07
I6390 0 n6391 2.976e-02A M=7.371e-07
I6391 0 n6392 2.976e-02A M=8.133e-07
I6392 0 n6393 2.976e-02A M=3.980e-07
I6393 0 n6394 2.976e-02A M=7.114e-07
I6394 0 n6395 2.976e-02A M=8.750e-07
I6395 0 n6396 2.976e-02A M=1.263e-06
I6396 0 n6397 2.976e-02A M=1.317e-06
I6397 0 n6398 2.976e-02A M=1.237e-06
I6398 0 n6399 2.976e-02A M=5.676e-07
I6399 0 n6400 2.976e-02A M=5.533e-07
I6400 0 n6401 2.976e-02A M=4.578e-07
I6401 0 n6402 2.976e-02A M=6.405e-07
I6402 0 n6403 2.976e-02A M=1.461e-06
I6403 0 n6404 2.976e-02A M=2.800e-07
I6404 0 n6405 2.976e-02A M=1.059e-06
I6405 0 n6406 2.976e-02A M=1.987e-06
I6406 0 n6407 2.976e-02A M=1.999e-06
I6407 0 n6408 2.976e-02A M=2.123e-06
I6408 0 n6409 2.976e-02A M=1.184e-06
I6409 0 n6410 2.976e-02A M=9.703e-07
I6410 0 n6411 2.976e-02A M=9.881e-07
I6411 0 n6412 2.976e-02A M=7.483e-07
I6412 0 n6413 2.976e-02A M=5.563e-07
I6413 0 n6414 2.976e-02A M=1.327e-06
I6414 0 n6415 2.976e-02A M=2.124e-07
I6415 0 n6416 2.976e-02A M=4.599e-07
I6416 0 n6417 2.976e-02A M=3.359e-07
I6417 0 n6418 2.976e-02A M=1.189e-06
I6418 0 n6419 2.976e-02A M=8.087e-07
I6419 0 n6420 2.976e-02A M=6.376e-07
I6420 0 n6421 2.976e-02A M=3.815e-07
I6421 0 n6422 2.976e-02A M=1.080e-06
I6422 0 n6423 2.976e-02A M=5.153e-07
I6423 0 n6424 2.976e-02A M=9.426e-07
I6424 0 n6425 2.976e-02A M=4.241e-07
I6425 0 n6426 2.976e-02A M=2.259e-07
I6426 0 n6427 2.976e-02A M=1.924e-06
I6427 0 n6428 2.976e-02A M=1.140e-06
I6428 0 n6429 2.976e-02A M=1.666e-06
I6429 0 n6430 2.976e-02A M=9.277e-07
I6430 0 n6431 2.976e-02A M=1.106e-06
I6431 0 n6432 2.976e-02A M=6.130e-07
I6432 0 n6433 2.976e-02A M=8.986e-07
I6433 0 n6434 2.976e-02A M=1.146e-06
I6434 0 n6435 2.976e-02A M=1.061e-06
I6435 0 n6436 2.976e-02A M=1.356e-07
I6436 0 n6437 2.976e-02A M=1.674e-06
I6437 0 n6438 2.976e-02A M=7.925e-07
I6438 0 n6439 2.976e-02A M=6.762e-07
I6439 0 n6440 2.976e-02A M=5.100e-07
I6440 0 n6441 2.976e-02A M=6.300e-07
I6441 0 n6442 2.976e-02A M=1.332e-06
I6442 0 n6443 2.976e-02A M=2.293e-06
I6443 0 n6444 2.976e-02A M=7.740e-07
I6444 0 n6445 2.976e-02A M=9.385e-07
I6445 0 n6446 2.976e-02A M=7.981e-07
I6446 0 n6447 2.976e-02A M=6.534e-07
I6447 0 n6448 2.976e-02A M=1.156e-06
I6448 0 n6449 2.976e-02A M=8.883e-07
I6449 0 n6450 2.976e-02A M=2.438e-06
I6450 0 n6451 2.976e-02A M=1.242e-06
I6451 0 n6452 2.976e-02A M=7.908e-07
I6452 0 n6453 2.976e-02A M=1.806e-06
I6453 0 n6454 2.976e-02A M=4.154e-07
I6454 0 n6455 2.976e-02A M=1.064e-06
I6455 0 n6456 2.976e-02A M=1.200e-06
I6456 0 n6457 2.976e-02A M=8.263e-07
I6457 0 n6458 2.976e-02A M=4.122e-07
I6458 0 n6459 2.976e-02A M=1.861e-06
I6459 0 n6460 2.976e-02A M=3.327e-07
I6460 0 n6461 2.976e-02A M=1.120e-06
I6461 0 n6462 2.976e-02A M=2.261e-07
I6462 0 n6463 2.976e-02A M=1.999e-06
I6463 0 n6464 2.976e-02A M=4.307e-07
I6464 0 n6465 2.976e-02A M=2.762e-06
I6465 0 n6466 2.976e-02A M=7.413e-07
I6466 0 n6467 2.976e-02A M=9.771e-07
I6467 0 n6468 2.976e-02A M=1.227e-06
I6468 0 n6469 2.976e-02A M=8.842e-07
I6469 0 n1 2.976e-02A M=2.747e-07
I6470 0 n6471 2.976e-02A M=1.024e-06
I6471 0 n6472 2.976e-02A M=5.212e-07
I6472 0 n6473 2.976e-02A M=6.349e-07
I6473 0 n6474 2.976e-02A M=6.778e-07
I6474 0 n6475 2.976e-02A M=1.037e-06
I6475 0 n6476 2.976e-02A M=7.276e-07
I6476 0 n6477 2.976e-02A M=1.093e-06
I6477 0 n6478 2.976e-02A M=8.051e-07
I6478 0 n6479 2.976e-02A M=6.204e-07
I6479 0 n6480 2.976e-02A M=1.091e-06
I6480 0 n6481 2.976e-02A M=1.048e-06
I6481 0 n6482 2.976e-02A M=1.069e-06
I6482 0 n6483 2.976e-02A M=6.810e-07
I6483 0 n6484 2.976e-02A M=1.056e-06
I6484 0 n6485 2.976e-02A M=1.640e-06
I6485 0 n6486 2.976e-02A M=1.016e-06
I6486 0 n6487 2.976e-02A M=1.003e-06
I6487 0 n6488 2.976e-02A M=5.766e-07
I6488 0 n6489 2.976e-02A M=1.590e-06
I6489 0 n6490 2.976e-02A M=1.674e-06
I6490 0 n6491 2.976e-02A M=1.010e-06
I6491 0 n6492 2.976e-02A M=8.331e-07
I6492 0 n6493 2.976e-02A M=1.652e-06
I6493 0 n6494 2.976e-02A M=8.447e-07
I6494 0 n6495 2.976e-02A M=1.957e-06
I6495 0 n6496 2.976e-02A M=5.733e-07
I6496 0 n6497 2.976e-02A M=8.672e-07
I6497 0 n6498 2.976e-02A M=8.244e-07
I6498 0 n6499 2.976e-02A M=2.311e-07
I6499 0 n6500 2.976e-02A M=2.042e-06
I6500 0 n6501 2.976e-02A M=7.595e-07
I6501 0 n6502 2.976e-02A M=4.144e-07
I6502 0 n6503 2.976e-02A M=6.993e-07
I6503 0 n6504 2.976e-02A M=1.634e-06
I6504 0 n6505 2.976e-02A M=6.438e-07
I6505 0 n6506 2.976e-02A M=5.892e-07
I6506 0 n6507 2.976e-02A M=1.091e-06
I6507 0 n6508 2.976e-02A M=8.508e-07
I6508 0 n6509 2.976e-02A M=9.457e-07
I6509 0 n6510 2.976e-02A M=1.879e-06
I6510 0 n6511 2.976e-02A M=1.312e-06
I6511 0 n6512 2.976e-02A M=5.262e-07
I6512 0 n6513 2.976e-02A M=1.528e-06
I6513 0 n6514 2.976e-02A M=1.136e-06
I6514 0 n6515 2.976e-02A M=1.012e-06
I6515 0 n6516 2.976e-02A M=1.378e-06
I6516 0 n6517 2.976e-02A M=8.884e-07
I6517 0 n6518 2.976e-02A M=5.982e-07
I6518 0 n6519 2.976e-02A M=1.064e-06
I6519 0 n6520 2.976e-02A M=5.608e-07
I6520 0 n6521 2.976e-02A M=7.260e-07
I6521 0 n6522 2.976e-02A M=1.008e-06
I6522 0 n6523 2.976e-02A M=1.735e-06
I6523 0 n6524 2.976e-02A M=1.548e-06
I6524 0 n6525 2.976e-02A M=1.206e-06
I6525 0 n6526 2.976e-02A M=2.079e-06
I6526 0 n6527 2.976e-02A M=7.247e-07
I6527 0 n6528 2.976e-02A M=1.478e-06
I6528 0 n6529 2.976e-02A M=8.107e-07
I6529 0 n6530 2.976e-02A M=1.993e-06
I6530 0 n6531 2.976e-02A M=1.922e-06
I6531 0 n6532 2.976e-02A M=4.763e-07
I6532 0 n6533 2.976e-02A M=4.632e-07
I6533 0 n6534 2.976e-02A M=9.854e-07
I6534 0 n6535 2.976e-02A M=8.199e-07
I6535 0 n6536 2.976e-02A M=1.049e-06
I6536 0 n6537 2.976e-02A M=1.509e-06
I6537 0 n6538 2.976e-02A M=9.350e-07
I6538 0 n6539 2.976e-02A M=7.016e-07
I6539 0 n6540 2.976e-02A M=1.952e-06
I6540 0 n6541 2.976e-02A M=7.957e-07
I6541 0 n6542 2.976e-02A M=5.938e-07
I6542 0 n6543 2.976e-02A M=8.415e-07
I6543 0 n6544 2.976e-02A M=2.354e-06
I6544 0 n6545 2.976e-02A M=5.064e-07
I6545 0 n6546 2.976e-02A M=2.355e-07
I6546 0 n6547 2.976e-02A M=4.938e-07
I6547 0 n6548 2.976e-02A M=9.645e-07
I6548 0 n6549 2.976e-02A M=6.352e-07
I6549 0 n6550 2.976e-02A M=3.310e-07
I6550 0 n6551 2.976e-02A M=3.600e-07
I6551 0 n6552 2.976e-02A M=1.338e-06
I6552 0 n6553 2.976e-02A M=1.315e-06
I6553 0 n6554 2.976e-02A M=2.537e-07
I6554 0 n6555 2.976e-02A M=9.237e-07
I6555 0 n6556 2.976e-02A M=5.346e-07
I6556 0 n6557 2.976e-02A M=3.800e-07
I6557 0 n6558 2.976e-02A M=4.212e-07
I6558 0 n6559 2.976e-02A M=1.640e-06
I6559 0 n6560 2.976e-02A M=5.836e-07
I6560 0 n6561 2.976e-02A M=3.608e-07
I6561 0 n6562 2.976e-02A M=6.380e-07
I6562 0 n6563 2.976e-02A M=7.754e-07
I6563 0 n6564 2.976e-02A M=1.438e-06
I6564 0 n6565 2.976e-02A M=9.009e-07
I6565 0 n6566 2.976e-02A M=5.848e-07
I6566 0 n6567 2.976e-02A M=1.382e-06
I6567 0 n6568 2.976e-02A M=1.364e-06
I6568 0 n6569 2.976e-02A M=1.527e-06
I6569 0 n6570 2.976e-02A M=1.320e-06
I6570 0 n6571 2.976e-02A M=8.526e-07
I6571 0 n6572 2.976e-02A M=6.696e-07
I6572 0 n6573 2.976e-02A M=1.099e-06
I6573 0 n6574 2.976e-02A M=3.481e-07
I6574 0 n6575 2.976e-02A M=1.292e-06
I6575 0 n6576 2.976e-02A M=1.105e-06
I6576 0 n6577 2.976e-02A M=1.010e-06
I6577 0 n6578 2.976e-02A M=4.838e-07
I6578 0 n6579 2.976e-02A M=1.665e-06
I6579 0 n6580 2.976e-02A M=8.200e-07
I6580 0 n6581 2.976e-02A M=2.524e-07
I6581 0 n6582 2.976e-02A M=5.716e-07
I6582 0 n6583 2.976e-02A M=5.987e-07
I6583 0 n6584 2.976e-02A M=4.369e-07
I6584 0 n6585 2.976e-02A M=1.191e-06
I6585 0 n6586 2.976e-02A M=5.611e-07
I6586 0 n6587 2.976e-02A M=2.965e-07
I6587 0 n6588 2.976e-02A M=1.717e-06
I6588 0 n6589 2.976e-02A M=1.250e-06
I6589 0 n6590 2.976e-02A M=4.345e-07
I6590 0 n6591 2.976e-02A M=4.866e-07
I6591 0 n6592 2.976e-02A M=1.360e-06
I6592 0 n6593 2.976e-02A M=1.015e-06
I6593 0 n6594 2.976e-02A M=6.801e-07
I6594 0 n6595 2.976e-02A M=4.848e-07
I6595 0 n6596 2.976e-02A M=2.477e-06
I6596 0 n6597 2.976e-02A M=1.879e-06
I6597 0 n6598 2.976e-02A M=1.157e-06
I6598 0 n6599 2.976e-02A M=1.052e-06
I6599 0 n6600 2.976e-02A M=1.528e-06
I6600 0 n6601 2.976e-02A M=1.170e-06
I6601 0 n6602 2.976e-02A M=1.585e-06
I6602 0 n6603 2.976e-02A M=1.138e-06
I6603 0 n6604 2.976e-02A M=1.942e-06
I6604 0 n6605 2.976e-02A M=6.837e-07
I6605 0 n6606 2.976e-02A M=5.664e-07
I6606 0 n6607 2.976e-02A M=6.266e-07
I6607 0 n6608 2.976e-02A M=5.565e-07
I6608 0 n6609 2.976e-02A M=5.505e-07
I6609 0 n6610 2.976e-02A M=4.797e-07
I6610 0 n6611 2.976e-02A M=4.086e-07
I6611 0 n6612 2.976e-02A M=8.390e-07
I6612 0 n6613 2.976e-02A M=7.562e-07
I6613 0 n6614 2.976e-02A M=1.470e-06
I6614 0 n6615 2.976e-02A M=1.054e-06
I6615 0 n6616 2.976e-02A M=6.917e-07
I6616 0 n6617 2.976e-02A M=9.748e-07
I6617 0 n6618 2.976e-02A M=3.851e-07
I6618 0 n6619 2.976e-02A M=1.581e-06
I6619 0 n6620 2.976e-02A M=8.485e-07
I6620 0 n6621 2.976e-02A M=9.538e-07
I6621 0 n6622 2.976e-02A M=1.966e-07
I6622 0 n6623 2.976e-02A M=4.653e-07
I6623 0 n6624 2.976e-02A M=9.217e-07
I6624 0 n6625 2.976e-02A M=9.486e-07
I6625 0 n6626 2.976e-02A M=1.258e-06
I6626 0 n6627 2.976e-02A M=6.009e-07
I6627 0 n6628 2.976e-02A M=6.427e-07
I6628 0 n6629 2.976e-02A M=5.126e-07
I6629 0 n6630 2.976e-02A M=1.440e-06
I6630 0 n6631 2.976e-02A M=5.035e-07
I6631 0 n6632 2.976e-02A M=6.530e-07
I6632 0 n6633 2.976e-02A M=1.885e-06
I6633 0 n6634 2.976e-02A M=1.873e-06
I6634 0 n6635 2.976e-02A M=2.481e-07
I6635 0 n6636 2.976e-02A M=1.997e-06
I6636 0 n6637 2.976e-02A M=6.767e-07
I6637 0 n6638 2.976e-02A M=1.538e-06
I6638 0 n6639 2.976e-02A M=4.616e-07
I6639 0 n6640 2.976e-02A M=2.700e-07
I6640 0 n6641 2.976e-02A M=1.593e-06
I6641 0 n6642 2.976e-02A M=1.938e-06
I6642 0 n6643 2.976e-02A M=2.000e-06
I6643 0 n6644 2.976e-02A M=1.227e-06
I6644 0 n6645 2.976e-02A M=1.065e-06
I6645 0 n6646 2.976e-02A M=1.081e-06
I6646 0 n1 2.976e-02A M=5.536e-07
I6647 0 n6648 2.976e-02A M=1.252e-06
I6648 0 n6649 2.976e-02A M=8.564e-07
I6649 0 n6650 2.976e-02A M=1.150e-06
I6650 0 n6651 2.976e-02A M=1.717e-06
I6651 0 n6652 2.976e-02A M=2.947e-06
I6652 0 n6653 2.976e-02A M=5.658e-07
I6653 0 n6654 2.976e-02A M=1.269e-06
I6654 0 n6655 2.976e-02A M=7.774e-07
I6655 0 n6656 2.976e-02A M=1.496e-06
I6656 0 n6657 2.976e-02A M=7.571e-07
I6657 0 n6658 2.976e-02A M=1.200e-06
I6658 0 n6659 2.976e-02A M=3.567e-07
I6659 0 n6660 2.976e-02A M=2.503e-06
I6660 0 n6661 2.976e-02A M=1.417e-06
I6661 0 n6662 2.976e-02A M=1.034e-06
I6662 0 n6663 2.976e-02A M=1.457e-06
I6663 0 n6664 2.976e-02A M=1.057e-06
I6664 0 n6665 2.976e-02A M=4.464e-07
I6665 0 n6666 2.976e-02A M=1.548e-06
I6666 0 n6667 2.976e-02A M=1.083e-06
I6667 0 n6668 2.976e-02A M=1.007e-06
I6668 0 n6669 2.976e-02A M=2.258e-06
I6669 0 n6670 2.976e-02A M=4.813e-07
I6670 0 n6671 2.976e-02A M=9.900e-07
I6671 0 n6672 2.976e-02A M=6.013e-07
I6672 0 n6673 2.976e-02A M=4.423e-07
I6673 0 n6674 2.976e-02A M=2.703e-06
I6674 0 n6675 2.976e-02A M=1.750e-06
I6675 0 n6676 2.976e-02A M=7.992e-07
I6676 0 n6677 2.976e-02A M=5.602e-07
I6677 0 n6678 2.976e-02A M=1.699e-06
I6678 0 n6679 2.976e-02A M=1.861e-06
I6679 0 n6680 2.976e-02A M=9.573e-07
I6680 0 n6681 2.976e-02A M=5.364e-07
I6681 0 n6682 2.976e-02A M=9.004e-07
I6682 0 n6683 2.976e-02A M=8.500e-07
I6683 0 n6684 2.976e-02A M=4.327e-07
I6684 0 n6685 2.976e-02A M=2.130e-07
I6685 0 n6686 2.976e-02A M=7.854e-07
I6686 0 n6687 2.976e-02A M=7.085e-07
I6687 0 n6688 2.976e-02A M=2.551e-06
I6688 0 n6689 2.976e-02A M=1.386e-06
I6689 0 n6690 2.976e-02A M=9.354e-07
I6690 0 n6691 2.976e-02A M=1.202e-07
I6691 0 n6692 2.976e-02A M=8.412e-07
I6692 0 n6693 2.976e-02A M=7.471e-07
I6693 0 n6694 2.976e-02A M=1.902e-06
I6694 0 n6695 2.976e-02A M=1.375e-06
I6695 0 n6696 2.976e-02A M=4.524e-07
I6696 0 n6697 2.976e-02A M=8.529e-07
I6697 0 n6698 2.976e-02A M=1.991e-06
I6698 0 n6699 2.976e-02A M=8.797e-07
I6699 0 n6700 2.976e-02A M=3.279e-07
I6700 0 n6701 2.976e-02A M=6.935e-07
I6701 0 n6702 2.976e-02A M=4.993e-07
I6702 0 n6703 2.976e-02A M=5.364e-07
I6703 0 n6704 2.976e-02A M=5.881e-07
I6704 0 n6705 2.976e-02A M=8.583e-07
I6705 0 n6706 2.976e-02A M=2.827e-06
I6706 0 n6707 2.976e-02A M=8.344e-07
I6707 0 n6708 2.976e-02A M=6.138e-07
I6708 0 n6709 2.976e-02A M=1.999e-06
I6709 0 n6710 2.976e-02A M=1.247e-06
I6710 0 n6711 2.976e-02A M=1.482e-06
I6711 0 n6712 2.976e-02A M=6.313e-07
I6712 0 n6713 2.976e-02A M=1.742e-06
I6713 0 n6714 2.976e-02A M=1.448e-06
I6714 0 n6715 2.976e-02A M=8.041e-07
I6715 0 n6716 2.976e-02A M=1.071e-06
I6716 0 n6717 2.976e-02A M=2.937e-07
I6717 0 n6718 2.976e-02A M=1.688e-07
I6718 0 n6719 2.976e-02A M=4.896e-07
I6719 0 n6720 2.976e-02A M=5.290e-07
I6720 0 n6721 2.976e-02A M=7.135e-07
I6721 0 n6722 2.976e-02A M=6.118e-07
I6722 0 n6723 2.976e-02A M=7.680e-07
I6723 0 n6724 2.976e-02A M=2.670e-06
I6724 0 n6725 2.976e-02A M=6.224e-07
I6725 0 n6726 2.976e-02A M=6.563e-07
I6726 0 n6727 2.976e-02A M=5.911e-07
I6727 0 n6728 2.976e-02A M=7.429e-07
I6728 0 n6729 2.976e-02A M=8.701e-07
I6729 0 n6730 2.976e-02A M=1.141e-06
I6730 0 n6731 2.976e-02A M=1.554e-06
I6731 0 n6732 2.976e-02A M=8.146e-07
I6732 0 n6733 2.976e-02A M=7.921e-07
I6733 0 n6734 2.976e-02A M=1.223e-06
I6734 0 n6735 2.976e-02A M=7.561e-07
I6735 0 n6736 2.976e-02A M=4.134e-07
I6736 0 n6737 2.976e-02A M=3.686e-07
I6737 0 n6738 2.976e-02A M=6.335e-07
I6738 0 n6739 2.976e-02A M=3.718e-07
I6739 0 n6740 2.976e-02A M=1.189e-06
I6740 0 n6741 2.976e-02A M=8.153e-07
I6741 0 n6742 2.976e-02A M=7.430e-07
I6742 0 n6743 2.976e-02A M=1.129e-06
I6743 0 n6744 2.976e-02A M=9.255e-07
I6744 0 n6745 2.976e-02A M=5.497e-07
I6745 0 n6746 2.976e-02A M=6.985e-07
I6746 0 n6747 2.976e-02A M=1.098e-06
I6747 0 n6748 2.976e-02A M=4.024e-07
I6748 0 n6749 2.976e-02A M=9.304e-07
I6749 0 n6750 2.976e-02A M=8.235e-07
I6750 0 n6751 2.976e-02A M=1.855e-06
I6751 0 n6752 2.976e-02A M=2.591e-07
I6752 0 n6753 2.976e-02A M=8.525e-07
I6753 0 n6754 2.976e-02A M=3.428e-07
I6754 0 n6755 2.976e-02A M=5.755e-07
I6755 0 n6756 2.976e-02A M=4.975e-07
I6756 0 n6757 2.976e-02A M=8.460e-07
I6757 0 n6758 2.976e-02A M=7.740e-07
I6758 0 n6759 2.976e-02A M=9.007e-07
I6759 0 n6760 2.976e-02A M=1.117e-06
I6760 0 n6761 2.976e-02A M=5.144e-07
I6761 0 n6762 2.976e-02A M=7.848e-07
I6762 0 n6763 2.976e-02A M=8.832e-07
I6763 0 n6764 2.976e-02A M=1.253e-06
I6764 0 n6765 2.976e-02A M=1.653e-06
I6765 0 n6766 2.976e-02A M=5.606e-07
I6766 0 n6767 2.976e-02A M=9.906e-07
I6767 0 n6768 2.976e-02A M=8.795e-07
I6768 0 n6769 2.976e-02A M=1.351e-06
I6769 0 n6770 2.976e-02A M=1.423e-06
I6770 0 n6771 2.976e-02A M=8.477e-07
I6771 0 n6772 2.976e-02A M=6.827e-07
I6772 0 n6773 2.976e-02A M=9.882e-07
I6773 0 n6774 2.976e-02A M=7.507e-07
I6774 0 n6775 2.976e-02A M=7.080e-07
I6775 0 n6776 2.976e-02A M=8.368e-07
I6776 0 n6777 2.976e-02A M=9.572e-07
I6777 0 n6778 2.976e-02A M=8.325e-07
I6778 0 n6779 2.976e-02A M=1.366e-06
I6779 0 n6780 2.976e-02A M=1.513e-06
I6780 0 n6781 2.976e-02A M=9.063e-07
I6781 0 n6782 2.976e-02A M=2.042e-07
I6782 0 n6783 2.976e-02A M=7.354e-07
I6783 0 n6784 2.976e-02A M=2.516e-06
I6784 0 n6785 2.976e-02A M=5.206e-07
I6785 0 n6786 2.976e-02A M=1.300e-07
I6786 0 n6787 2.976e-02A M=4.601e-07
I6787 0 n6788 2.976e-02A M=4.960e-07
I6788 0 n6789 2.976e-02A M=1.991e-06
I6789 0 n6790 2.976e-02A M=9.159e-07
I6790 0 n6791 2.976e-02A M=1.384e-06
I6791 0 n6792 2.976e-02A M=2.237e-06
I6792 0 n6793 2.976e-02A M=7.658e-07
I6793 0 n6794 2.976e-02A M=8.507e-07
I6794 0 n6795 2.976e-02A M=1.354e-06
I6795 0 n6796 2.976e-02A M=8.910e-07
I6796 0 n6797 2.976e-02A M=1.462e-07
I6797 0 n6798 2.976e-02A M=5.764e-07
I6798 0 n6799 2.976e-02A M=3.318e-07
I6799 0 n6800 2.976e-02A M=8.248e-07
I6800 0 n6801 2.976e-02A M=7.684e-07
I6801 0 n6802 2.976e-02A M=1.244e-06
I6802 0 n6803 2.976e-02A M=1.062e-06
I6803 0 n6804 2.976e-02A M=1.513e-06
I6804 0 n6805 2.976e-02A M=1.310e-06
I6805 0 n6806 2.976e-02A M=2.320e-06
I6806 0 n6807 2.976e-02A M=8.625e-07
I6807 0 n6808 2.976e-02A M=6.042e-07
I6808 0 n6809 2.976e-02A M=5.931e-07
I6809 0 n6810 2.976e-02A M=1.007e-06
I6810 0 n6811 2.976e-02A M=1.314e-06
I6811 0 n6812 2.976e-02A M=2.274e-06
I6812 0 n6813 2.976e-02A M=6.624e-07
I6813 0 n6814 2.976e-02A M=1.207e-06
I6814 0 n6815 2.976e-02A M=1.091e-06
I6815 0 n6816 2.976e-02A M=2.120e-07
I6816 0 n6817 2.976e-02A M=8.122e-07
I6817 0 n6818 2.976e-02A M=5.828e-07
I6818 0 n6819 2.976e-02A M=5.995e-07
I6819 0 n6820 2.976e-02A M=6.214e-07
I6820 0 n6821 2.976e-02A M=1.437e-06
I6821 0 n6822 2.976e-02A M=1.465e-06
I6822 0 n6823 2.976e-02A M=3.887e-07
I6823 0 n6824 2.976e-02A M=1.526e-06
I6824 0 n6825 2.976e-02A M=9.028e-07
I6825 0 n6826 2.976e-02A M=1.032e-06
I6826 0 n6827 2.976e-02A M=6.258e-07
I6827 0 n6828 2.976e-02A M=6.318e-07
I6828 0 n6829 2.976e-02A M=8.051e-07
I6829 0 n6830 2.976e-02A M=1.034e-06
I6830 0 n6831 2.976e-02A M=8.445e-07
I6831 0 n6832 2.976e-02A M=2.865e-07
I6832 0 n6833 2.976e-02A M=1.209e-06
I6833 0 n6834 2.976e-02A M=1.522e-06
I6834 0 n6835 2.976e-02A M=8.150e-07
I6835 0 n6836 2.976e-02A M=4.158e-07
I6836 0 n6837 2.976e-02A M=1.098e-06
I6837 0 n6838 2.976e-02A M=1.197e-06
I6838 0 n6839 2.976e-02A M=1.194e-06
I6839 0 n6840 2.976e-02A M=1.814e-06
I6840 0 n6841 2.976e-02A M=1.090e-06
I6841 0 n6842 2.976e-02A M=1.495e-06
I6842 0 n6843 2.976e-02A M=1.121e-06
I6843 0 n6844 2.976e-02A M=4.681e-07
I6844 0 n6845 2.976e-02A M=4.058e-07
I6845 0 n6846 2.976e-02A M=1.167e-06
I6846 0 n6847 2.976e-02A M=1.236e-06
I6847 0 n6848 2.976e-02A M=1.140e-06
I6848 0 n6849 2.976e-02A M=1.801e-07
I6849 0 n6850 2.976e-02A M=7.520e-07
I6850 0 n6851 2.976e-02A M=5.091e-07
I6851 0 n6852 2.976e-02A M=3.926e-07
I6852 0 n6853 2.976e-02A M=9.244e-07
I6853 0 n6854 2.976e-02A M=3.374e-06
I6854 0 n6855 2.976e-02A M=7.713e-07
I6855 0 n6856 2.976e-02A M=1.424e-06
I6856 0 n6857 2.976e-02A M=1.650e-06
I6857 0 n6858 2.976e-02A M=1.404e-06
I6858 0 n6859 2.976e-02A M=1.038e-06
I6859 0 n6860 2.976e-02A M=9.372e-07
I6860 0 n6861 2.976e-02A M=1.914e-06
I6861 0 n6862 2.976e-02A M=5.576e-07
I6862 0 n6863 2.976e-02A M=9.290e-07
I6863 0 n6864 2.976e-02A M=5.137e-07
I6864 0 n6865 2.976e-02A M=7.042e-08
I6865 0 n6866 2.976e-02A M=4.628e-07
I6866 0 n6867 2.976e-02A M=6.348e-07
I6867 0 n6868 2.976e-02A M=1.329e-06
I6868 0 n6869 2.976e-02A M=2.812e-06
I6869 0 n6870 2.976e-02A M=5.195e-07
I6870 0 n6871 2.976e-02A M=3.099e-07
I6871 0 n6872 2.976e-02A M=7.729e-07
I6872 0 n6873 2.976e-02A M=1.243e-06
I6873 0 n6874 2.976e-02A M=8.202e-07
I6874 0 n6875 2.976e-02A M=5.241e-07
I6875 0 n6876 2.976e-02A M=1.061e-06
I6876 0 n6877 2.976e-02A M=7.334e-07
I6877 0 n6878 2.976e-02A M=7.541e-07
I6878 0 n6879 2.976e-02A M=1.136e-06
I6879 0 n6880 2.976e-02A M=1.182e-06
I6880 0 n6881 2.976e-02A M=4.630e-07
I6881 0 n6882 2.976e-02A M=8.095e-07
I6882 0 n6883 2.976e-02A M=4.492e-07
I6883 0 n6884 2.976e-02A M=7.642e-07
I6884 0 n6885 2.976e-02A M=2.118e-06
I6885 0 n6886 2.976e-02A M=1.326e-06
I6886 0 n6887 2.976e-02A M=7.498e-07
I6887 0 n6888 2.976e-02A M=1.483e-06
I6888 0 n6889 2.976e-02A M=1.071e-06
I6889 0 n6890 2.976e-02A M=6.602e-07
I6890 0 n6891 2.976e-02A M=1.185e-06
I6891 0 n6892 2.976e-02A M=2.535e-06
I6892 0 n6893 2.976e-02A M=3.702e-07
I6893 0 n6894 2.976e-02A M=8.358e-07
I6894 0 n6895 2.976e-02A M=8.962e-07
I6895 0 n6896 2.976e-02A M=8.031e-07
I6896 0 n6897 2.976e-02A M=2.255e-07
I6897 0 n6898 2.976e-02A M=2.504e-07
I6898 0 n6899 2.976e-02A M=5.770e-07
I6899 0 n6900 2.976e-02A M=6.353e-07
I6900 0 n6901 2.976e-02A M=7.280e-07
I6901 0 n6902 2.976e-02A M=2.172e-06
I6902 0 n6903 2.976e-02A M=8.278e-07
I6903 0 n6904 2.976e-02A M=8.967e-07
I6904 0 n6905 2.976e-02A M=1.500e-06
I6905 0 n6906 2.976e-02A M=7.494e-07
I6906 0 n6907 2.976e-02A M=1.143e-06
I6907 0 n6908 2.976e-02A M=1.431e-06
I6908 0 n6909 2.976e-02A M=1.183e-06
I6909 0 n6910 2.976e-02A M=1.159e-06
I6910 0 n6911 2.976e-02A M=7.997e-07
I6911 0 n6912 2.976e-02A M=1.849e-06
I6912 0 n6913 2.976e-02A M=2.945e-06
I6913 0 n6914 2.976e-02A M=1.238e-06
I6914 0 n6915 2.976e-02A M=1.489e-06
I6915 0 n6916 2.976e-02A M=9.382e-07
I6916 0 n6917 2.976e-02A M=7.988e-07
I6917 0 n6918 2.976e-02A M=3.017e-07
I6918 0 n6919 2.976e-02A M=1.063e-06
I6919 0 n6920 2.976e-02A M=7.082e-07
I6920 0 n6921 2.976e-02A M=1.545e-06
I6921 0 n6922 2.976e-02A M=4.670e-07
I6922 0 n6923 2.976e-02A M=1.002e-06
I6923 0 n6924 2.976e-02A M=8.202e-07
I6924 0 n6925 2.976e-02A M=1.161e-06
I6925 0 n6926 2.976e-02A M=1.543e-07
I6926 0 n6927 2.976e-02A M=4.467e-07
I6927 0 n6928 2.976e-02A M=5.007e-07
I6928 0 n6929 2.976e-02A M=1.435e-06
I6929 0 n6930 2.976e-02A M=3.219e-07
I6930 0 n6931 2.976e-02A M=1.438e-06
I6931 0 n6932 2.976e-02A M=6.053e-07
I6932 0 n6933 2.976e-02A M=2.308e-07
I6933 0 n6934 2.976e-02A M=2.245e-06
I6934 0 n6935 2.976e-02A M=1.206e-07
I6935 0 n6936 2.976e-02A M=5.972e-07
I6936 0 n6937 2.976e-02A M=1.300e-06
I6937 0 n6938 2.976e-02A M=1.481e-06
I6938 0 n6939 2.976e-02A M=1.486e-06
I6939 0 n6940 2.976e-02A M=1.263e-06
I6940 0 n6941 2.976e-02A M=7.115e-07
I6941 0 n6942 2.976e-02A M=3.629e-07
I6942 0 n6943 2.976e-02A M=1.258e-06
I6943 0 n6944 2.976e-02A M=5.553e-07
I6944 0 n6945 2.976e-02A M=7.323e-07
I6945 0 n6946 2.976e-02A M=1.418e-06
I6946 0 n6947 2.976e-02A M=6.412e-07
I6947 0 n6948 2.976e-02A M=5.113e-07
I6948 0 n6949 2.976e-02A M=1.235e-06
I6949 0 n6950 2.976e-02A M=7.348e-07
I6950 0 n6951 2.976e-02A M=7.974e-07
I6951 0 n6952 2.976e-02A M=4.211e-07
I6952 0 n6953 2.976e-02A M=2.143e-06
I6953 0 n6954 2.976e-02A M=5.467e-07
I6954 0 n6955 2.976e-02A M=1.097e-06
I6955 0 n6956 2.976e-02A M=1.490e-06
I6956 0 n6957 2.976e-02A M=1.288e-06
I6957 0 n6958 2.976e-02A M=6.000e-07
I6958 0 n6959 2.976e-02A M=6.940e-07
I6959 0 n6960 2.976e-02A M=1.335e-06
I6960 0 n6961 2.976e-02A M=1.461e-06
I6961 0 n6962 2.976e-02A M=9.446e-07
I6962 0 n6963 2.976e-02A M=3.583e-06
I6963 0 n6964 2.976e-02A M=8.129e-07
I6964 0 n6965 2.976e-02A M=4.043e-07
I6965 0 n6966 2.976e-02A M=5.735e-07
I6966 0 n1 2.976e-02A M=9.947e-07
I6967 0 n6968 2.976e-02A M=1.144e-06
I6968 0 n6969 2.976e-02A M=7.537e-07
I6969 0 n6970 2.976e-02A M=4.644e-07
I6970 0 n6971 2.976e-02A M=1.353e-06
I6971 0 n6972 2.976e-02A M=8.013e-07
I6972 0 n6973 2.976e-02A M=1.212e-06
I6973 0 n6974 2.976e-02A M=1.491e-06
I6974 0 n6975 2.976e-02A M=1.386e-06
I6975 0 n6976 2.976e-02A M=1.459e-06
I6976 0 n6977 2.976e-02A M=1.784e-06
I6977 0 n6978 2.976e-02A M=9.489e-07
I6978 0 n6979 2.976e-02A M=3.092e-06
I6979 0 n6980 2.976e-02A M=1.211e-06
I6980 0 n6981 2.976e-02A M=1.158e-06
I6981 0 n6982 2.976e-02A M=1.968e-07
I6982 0 n6983 2.976e-02A M=1.517e-06
I6983 0 n6984 2.976e-02A M=8.104e-07
I6984 0 n6985 2.976e-02A M=1.540e-06
I6985 0 n6986 2.976e-02A M=1.185e-06
I6986 0 n6987 2.976e-02A M=1.243e-06
I6987 0 n6988 2.976e-02A M=9.465e-07
I6988 0 n6989 2.976e-02A M=2.917e-07
I6989 0 n6990 2.976e-02A M=9.217e-07
I6990 0 n6991 2.976e-02A M=8.959e-07
I6991 0 n6992 2.976e-02A M=5.382e-07
I6992 0 n6993 2.976e-02A M=7.519e-07
I6993 0 n6994 2.976e-02A M=5.570e-07
I6994 0 n6995 2.976e-02A M=1.343e-06
I6995 0 n6996 2.976e-02A M=2.363e-06
I6996 0 n6997 2.976e-02A M=4.763e-07
I6997 0 n6998 2.976e-02A M=9.587e-07
I6998 0 n6999 2.976e-02A M=1.291e-06
I6999 0 n7000 2.976e-02A M=8.534e-07
I7000 0 n7001 2.976e-02A M=1.430e-06
I7001 0 n7002 2.976e-02A M=1.094e-06
I7002 0 n7003 2.976e-02A M=1.465e-06
I7003 0 n7004 2.976e-02A M=3.908e-07
I7004 0 n7005 2.976e-02A M=1.113e-06
I7005 0 n7006 2.976e-02A M=4.659e-07
I7006 0 n7007 2.976e-02A M=3.397e-07
I7007 0 n7008 2.976e-02A M=1.049e-06
I7008 0 n7009 2.976e-02A M=1.610e-06
I7009 0 n7010 2.976e-02A M=2.779e-07
I7010 0 n7011 2.976e-02A M=2.283e-06
I7011 0 n7012 2.976e-02A M=7.668e-07
I7012 0 n7013 2.976e-02A M=1.465e-06
I7013 0 n7014 2.976e-02A M=5.483e-07
I7014 0 n7015 2.976e-02A M=1.041e-06
I7015 0 n7016 2.976e-02A M=5.779e-07
I7016 0 n7017 2.976e-02A M=1.601e-06
I7017 0 n7018 2.976e-02A M=9.453e-07
I7018 0 n7019 2.976e-02A M=3.403e-07
I7019 0 n7020 2.976e-02A M=1.302e-06
I7020 0 n7021 2.976e-02A M=1.596e-06
I7021 0 n7022 2.976e-02A M=1.274e-06
I7022 0 n7023 2.976e-02A M=8.337e-07
I7023 0 n7024 2.976e-02A M=2.032e-06
I7024 0 n7025 2.976e-02A M=2.562e-06
I7025 0 n7026 2.976e-02A M=5.656e-07
I7026 0 n7027 2.976e-02A M=1.071e-06
I7027 0 n7028 2.976e-02A M=2.336e-07
I7028 0 n7029 2.976e-02A M=6.749e-07
I7029 0 n7030 2.976e-02A M=9.179e-07
I7030 0 n7031 2.976e-02A M=8.291e-07
I7031 0 n7032 2.976e-02A M=1.646e-06
I7032 0 n7033 2.976e-02A M=5.224e-07
I7033 0 n7034 2.976e-02A M=1.550e-06
I7034 0 n7035 2.976e-02A M=1.647e-06
I7035 0 n7036 2.976e-02A M=9.247e-07
I7036 0 n7037 2.976e-02A M=2.030e-06
I7037 0 n7038 2.976e-02A M=4.414e-07
I7038 0 n7039 2.976e-02A M=7.460e-07
I7039 0 n7040 2.976e-02A M=9.684e-07
I7040 0 n7041 2.976e-02A M=5.859e-07
I7041 0 n7042 2.976e-02A M=7.725e-07
I7042 0 n7043 2.976e-02A M=1.294e-06
I7043 0 n7044 2.976e-02A M=1.473e-06
I7044 0 n7045 2.976e-02A M=1.040e-06
I7045 0 n7046 2.976e-02A M=8.834e-07
I7046 0 n7047 2.976e-02A M=5.770e-07
I7047 0 n7048 2.976e-02A M=2.158e-06
I7048 0 n7049 2.976e-02A M=1.331e-06
I7049 0 n7050 2.976e-02A M=7.726e-07
I7050 0 n7051 2.976e-02A M=6.000e-07
I7051 0 n7052 2.976e-02A M=6.619e-07
I7052 0 n7053 2.976e-02A M=1.062e-06
I7053 0 n7054 2.976e-02A M=1.015e-06
I7054 0 n7055 2.976e-02A M=6.597e-07
I7055 0 n7056 2.976e-02A M=1.480e-06
I7056 0 n7057 2.976e-02A M=3.103e-07
I7057 0 n7058 2.976e-02A M=1.006e-06
I7058 0 n7059 2.976e-02A M=7.023e-07
I7059 0 n7060 2.976e-02A M=1.959e-06
I7060 0 n7061 2.976e-02A M=5.816e-07
I7061 0 n7062 2.976e-02A M=5.212e-07
I7062 0 n7063 2.976e-02A M=4.260e-07
I7063 0 n7064 2.976e-02A M=1.826e-07
I7064 0 n7065 2.976e-02A M=1.394e-06
I7065 0 n7066 2.976e-02A M=6.308e-07
I7066 0 n7067 2.976e-02A M=5.022e-07
I7067 0 n7068 2.976e-02A M=1.884e-06
I7068 0 n7069 2.976e-02A M=2.279e-07
I7069 0 n7070 2.976e-02A M=2.187e-06
I7070 0 n7071 2.976e-02A M=1.931e-06
I7071 0 n7072 2.976e-02A M=2.472e-06
I7072 0 n7073 2.976e-02A M=6.439e-07
I7073 0 n7074 2.976e-02A M=3.844e-07
I7074 0 n7075 2.976e-02A M=6.873e-07
I7075 0 n7076 2.976e-02A M=1.470e-07
I7076 0 n7077 2.976e-02A M=1.304e-06
I7077 0 n7078 2.976e-02A M=4.348e-07
I7078 0 n7079 2.976e-02A M=7.727e-07
I7079 0 n7080 2.976e-02A M=9.182e-07
I7080 0 n7081 2.976e-02A M=2.813e-07
I7081 0 n7082 2.976e-02A M=3.319e-07
I7082 0 n7083 2.976e-02A M=1.566e-06
I7083 0 n7084 2.976e-02A M=1.473e-06
I7084 0 n7085 2.976e-02A M=9.273e-07
I7085 0 n7086 2.976e-02A M=8.056e-07
I7086 0 n7087 2.976e-02A M=1.654e-06
I7087 0 n7088 2.976e-02A M=1.189e-06
I7088 0 n7089 2.976e-02A M=1.665e-06
I7089 0 n7090 2.976e-02A M=7.547e-07
I7090 0 n7091 2.976e-02A M=6.267e-07
I7091 0 n7092 2.976e-02A M=1.049e-06
I7092 0 n7093 2.976e-02A M=2.965e-07
I7093 0 n7094 2.976e-02A M=9.268e-07
I7094 0 n7095 2.976e-02A M=1.708e-06
I7095 0 n7096 2.976e-02A M=1.572e-06
I7096 0 n7097 2.976e-02A M=6.366e-07
I7097 0 n7098 2.976e-02A M=5.886e-07
I7098 0 n7099 2.976e-02A M=9.092e-07
I7099 0 n7100 2.976e-02A M=7.124e-07
I7100 0 n7101 2.976e-02A M=3.977e-07
I7101 0 n7102 2.976e-02A M=8.346e-07
I7102 0 n7103 2.976e-02A M=7.280e-07
I7103 0 n7104 2.976e-02A M=1.731e-06
I7104 0 n7105 2.976e-02A M=1.202e-06
I7105 0 n7106 2.976e-02A M=8.896e-07
I7106 0 n7107 2.976e-02A M=1.003e-06
I7107 0 n7108 2.976e-02A M=1.038e-06
I7108 0 n7109 2.976e-02A M=1.710e-06
I7109 0 n7110 2.976e-02A M=1.376e-06
I7110 0 n7111 2.976e-02A M=9.394e-07
I7111 0 n7112 2.976e-02A M=4.070e-07
I7112 0 n7113 2.976e-02A M=7.383e-07
I7113 0 n7114 2.976e-02A M=1.750e-06
I7114 0 n7115 2.976e-02A M=5.983e-07
I7115 0 n7116 2.976e-02A M=7.256e-07
I7116 0 n7117 2.976e-02A M=4.086e-07
I7117 0 n7118 2.976e-02A M=1.071e-06
I7118 0 n7119 2.976e-02A M=9.850e-07
I7119 0 n7120 2.976e-02A M=8.707e-07
I7120 0 n7121 2.976e-02A M=5.258e-07
I7121 0 n7122 2.976e-02A M=1.946e-06
I7122 0 n7123 2.976e-02A M=1.501e-06
I7123 0 n7124 2.976e-02A M=9.663e-07
I7124 0 n7125 2.976e-02A M=1.201e-06
I7125 0 n7126 2.976e-02A M=5.408e-07
I7126 0 n7127 2.976e-02A M=5.228e-07
I7127 0 n7128 2.976e-02A M=5.673e-07
I7128 0 n7129 2.976e-02A M=1.450e-06
I7129 0 n7130 2.976e-02A M=2.014e-06
I7130 0 n7131 2.976e-02A M=4.032e-07
I7131 0 n7132 2.976e-02A M=1.277e-06
I7132 0 n7133 2.976e-02A M=3.672e-07
I7133 0 n7134 2.976e-02A M=6.914e-07
I7134 0 n7135 2.976e-02A M=6.702e-07
I7135 0 n7136 2.976e-02A M=7.833e-07
I7136 0 n7137 2.976e-02A M=8.382e-07
I7137 0 n7138 2.976e-02A M=9.768e-07
I7138 0 n7139 2.976e-02A M=6.094e-07
I7139 0 n7140 2.976e-02A M=1.566e-06
I7140 0 n7141 2.976e-02A M=1.420e-06
I7141 0 n7142 2.976e-02A M=1.510e-06
I7142 0 n7143 2.976e-02A M=1.999e-06
I7143 0 n7144 2.976e-02A M=9.565e-07
I7144 0 n7145 2.976e-02A M=2.887e-06
I7145 0 n7146 2.976e-02A M=2.899e-06
I7146 0 n7147 2.976e-02A M=7.631e-07
I7147 0 n7148 2.976e-02A M=8.377e-07
I7148 0 n7149 2.976e-02A M=7.269e-07
I7149 0 n7150 2.976e-02A M=7.925e-08
I7150 0 n7151 2.976e-02A M=1.055e-06
I7151 0 n7152 2.976e-02A M=2.811e-07
I7152 0 n7153 2.976e-02A M=1.554e-06
I7153 0 n7154 2.976e-02A M=4.659e-07
I7154 0 n7155 2.976e-02A M=8.588e-07
I7155 0 n7156 2.976e-02A M=6.181e-07
I7156 0 n7157 2.976e-02A M=1.700e-06
I7157 0 n7158 2.976e-02A M=1.163e-06
I7158 0 n7159 2.976e-02A M=1.043e-06
I7159 0 n7160 2.976e-02A M=1.388e-06
I7160 0 n7161 2.976e-02A M=1.229e-06
I7161 0 n7162 2.976e-02A M=1.402e-06
I7162 0 n7163 2.976e-02A M=5.519e-07
I7163 0 n7164 2.976e-02A M=5.390e-07
I7164 0 n7165 2.976e-02A M=9.722e-07
I7165 0 n7166 2.976e-02A M=1.028e-06
I7166 0 n7167 2.976e-02A M=7.649e-07
I7167 0 n7168 2.976e-02A M=1.025e-06
I7168 0 n1 2.976e-02A M=2.157e-07
I7169 0 n7170 2.976e-02A M=6.130e-07
I7170 0 n7171 2.976e-02A M=4.804e-07
I7171 0 n7172 2.976e-02A M=4.851e-07
I7172 0 n7173 2.976e-02A M=9.342e-07
I7173 0 n7174 2.976e-02A M=6.431e-07
I7174 0 n7175 2.976e-02A M=1.863e-06
I7175 0 n7176 2.976e-02A M=1.040e-06
I7176 0 n7177 2.976e-02A M=2.819e-07
I7177 0 n7178 2.976e-02A M=2.412e-07
I7178 0 n7179 2.976e-02A M=1.141e-06
I7179 0 n7180 2.976e-02A M=2.357e-06
I7180 0 n7181 2.976e-02A M=7.857e-07
I7181 0 n7182 2.976e-02A M=6.407e-07
I7182 0 n7183 2.976e-02A M=1.955e-06
I7183 0 n7184 2.976e-02A M=6.504e-07
I7184 0 n7185 2.976e-02A M=3.403e-07
I7185 0 n7186 2.976e-02A M=7.053e-07
I7186 0 n7187 2.976e-02A M=7.651e-07
I7187 0 n7188 2.976e-02A M=1.448e-06
I7188 0 n7189 2.976e-02A M=1.513e-06
I7189 0 n7190 2.976e-02A M=1.313e-06
I7190 0 n7191 2.976e-02A M=1.129e-06
I7191 0 n7192 2.976e-02A M=1.855e-06
I7192 0 n7193 2.976e-02A M=4.948e-07
I7193 0 n7194 2.976e-02A M=9.615e-07
I7194 0 n7195 2.976e-02A M=1.969e-06
I7195 0 n7196 2.976e-02A M=1.127e-06
I7196 0 n7197 2.976e-02A M=1.328e-06
I7197 0 n7198 2.976e-02A M=1.405e-06
I7198 0 n7199 2.976e-02A M=3.735e-07
I7199 0 n7200 2.976e-02A M=1.830e-06
I7200 0 n7201 2.976e-02A M=4.236e-07
I7201 0 n7202 2.976e-02A M=6.751e-07
I7202 0 n7203 2.976e-02A M=4.161e-07
I7203 0 n7204 2.976e-02A M=1.953e-07
I7204 0 n7205 2.976e-02A M=1.256e-06
I7205 0 n7206 2.976e-02A M=7.722e-07
I7206 0 n7207 2.976e-02A M=9.701e-07
I7207 0 n7208 2.976e-02A M=1.554e-06
I7208 0 n7209 2.976e-02A M=8.120e-07
I7209 0 n7210 2.976e-02A M=1.195e-06
I7210 0 n7211 2.976e-02A M=4.135e-07
I7211 0 n7212 2.976e-02A M=1.245e-06
I7212 0 n7213 2.976e-02A M=5.599e-07
I7213 0 n7214 2.976e-02A M=2.744e-06
I7214 0 n7215 2.976e-02A M=2.750e-07
I7215 0 n7216 2.976e-02A M=1.457e-06
I7216 0 n7217 2.976e-02A M=1.643e-06
I7217 0 n7218 2.976e-02A M=7.085e-07
I7218 0 n7219 2.976e-02A M=1.601e-07
I7219 0 n7220 2.976e-02A M=4.437e-07
I7220 0 n7221 2.976e-02A M=1.671e-06
I7221 0 n7222 2.976e-02A M=6.532e-07
I7222 0 n7223 2.976e-02A M=1.304e-06
I7223 0 n7224 2.976e-02A M=8.250e-07
I7224 0 n7225 2.976e-02A M=9.751e-07
I7225 0 n7226 2.976e-02A M=2.748e-07
I7226 0 n7227 2.976e-02A M=1.723e-07
I7227 0 n7228 2.976e-02A M=5.698e-07
I7228 0 n7229 2.976e-02A M=3.792e-07
I7229 0 n7230 2.976e-02A M=1.195e-06
I7230 0 n7231 2.976e-02A M=1.618e-06
I7231 0 n7232 2.976e-02A M=4.217e-07
I7232 0 n7233 2.976e-02A M=1.027e-06
I7233 0 n7234 2.976e-02A M=1.191e-06
I7234 0 n7235 2.976e-02A M=7.241e-07
I7235 0 n7236 2.976e-02A M=8.282e-07
I7236 0 n7237 2.976e-02A M=1.365e-07
I7237 0 n7238 2.976e-02A M=1.038e-06
I7238 0 n7239 2.976e-02A M=7.584e-07
I7239 0 n7240 2.976e-02A M=5.862e-07
I7240 0 n7241 2.976e-02A M=3.322e-07
I7241 0 n7242 2.976e-02A M=7.144e-07
I7242 0 n7243 2.976e-02A M=1.668e-06
I7243 0 n7244 2.976e-02A M=1.887e-06
I7244 0 n7245 2.976e-02A M=5.332e-07
I7245 0 n7246 2.976e-02A M=1.044e-06
I7246 0 n7247 2.976e-02A M=8.767e-07
I7247 0 n7248 2.976e-02A M=7.168e-07
I7248 0 n7249 2.976e-02A M=9.362e-07
I7249 0 n7250 2.976e-02A M=1.955e-07
I7250 0 n7251 2.976e-02A M=7.274e-07
I7251 0 n7252 2.976e-02A M=1.132e-06
I7252 0 n7253 2.976e-02A M=4.233e-07
I7253 0 n7254 2.976e-02A M=7.261e-07
I7254 0 n7255 2.976e-02A M=3.955e-07
I7255 0 n7256 2.976e-02A M=1.073e-06
I7256 0 n7257 2.976e-02A M=1.116e-06
I7257 0 n7258 2.976e-02A M=2.573e-06
I7258 0 n7259 2.976e-02A M=5.721e-07
I7259 0 n7260 2.976e-02A M=4.995e-07
I7260 0 n7261 2.976e-02A M=1.318e-06
I7261 0 n7262 2.976e-02A M=4.409e-07
I7262 0 n7263 2.976e-02A M=2.338e-06
I7263 0 n7264 2.976e-02A M=2.512e-07
I7264 0 n7265 2.976e-02A M=9.688e-07
I7265 0 n7266 2.976e-02A M=2.193e-06
I7266 0 n7267 2.976e-02A M=1.596e-06
I7267 0 n7268 2.976e-02A M=1.262e-06
I7268 0 n7269 2.976e-02A M=5.034e-07
I7269 0 n7270 2.976e-02A M=7.614e-07
I7270 0 n7271 2.976e-02A M=1.059e-06
I7271 0 n7272 2.976e-02A M=7.370e-07
I7272 0 n7273 2.976e-02A M=6.558e-07
I7273 0 n7274 2.976e-02A M=6.700e-07
I7274 0 n7275 2.976e-02A M=1.008e-06
I7275 0 n7276 2.976e-02A M=7.501e-07
I7276 0 n7277 2.976e-02A M=7.231e-07
I7277 0 n7278 2.976e-02A M=1.271e-06
I7278 0 n7279 2.976e-02A M=7.572e-07
I7279 0 n7280 2.976e-02A M=3.924e-07
I7280 0 n7281 2.976e-02A M=1.288e-06
I7281 0 n7282 2.976e-02A M=2.309e-06
I7282 0 n7283 2.976e-02A M=1.534e-07
I7283 0 n7284 2.976e-02A M=7.591e-07
I7284 0 n7285 2.976e-02A M=2.274e-06
I7285 0 n7286 2.976e-02A M=4.608e-07
I7286 0 n7287 2.976e-02A M=2.044e-06
I7287 0 n7288 2.976e-02A M=8.991e-07
I7288 0 n7289 2.976e-02A M=1.070e-06
I7289 0 n7290 2.976e-02A M=7.958e-07
I7290 0 n7291 2.976e-02A M=8.421e-07
I7291 0 n7292 2.976e-02A M=8.275e-07
I7292 0 n7293 2.976e-02A M=1.405e-06
I7293 0 n7294 2.976e-02A M=1.352e-06
I7294 0 n7295 2.976e-02A M=8.157e-07
I7295 0 n7296 2.976e-02A M=1.919e-07
I7296 0 n7297 2.976e-02A M=2.770e-07
I7297 0 n7298 2.976e-02A M=8.808e-07
I7298 0 n7299 2.976e-02A M=4.074e-07
I7299 0 n7300 2.976e-02A M=8.466e-07
I7300 0 n7301 2.976e-02A M=9.741e-07
I7301 0 n7302 2.976e-02A M=7.697e-07
I7302 0 n1 2.976e-02A M=5.582e-07
I7303 0 n7304 2.976e-02A M=1.827e-06
I7304 0 n7305 2.976e-02A M=3.252e-07
I7305 0 n7306 2.976e-02A M=9.146e-07
I7306 0 n7307 2.976e-02A M=1.002e-06
I7307 0 n7308 2.976e-02A M=1.369e-06
I7308 0 n7309 2.976e-02A M=3.427e-07
I7309 0 n7310 2.976e-02A M=1.134e-06
I7310 0 n7311 2.976e-02A M=1.193e-06
I7311 0 n7312 2.976e-02A M=1.098e-06
I7312 0 n7313 2.976e-02A M=3.291e-07
I7313 0 n7314 2.976e-02A M=7.687e-07
I7314 0 n7315 2.976e-02A M=1.167e-06
I7315 0 n7316 2.976e-02A M=3.866e-07
I7316 0 n7317 2.976e-02A M=6.600e-07
I7317 0 n7318 2.976e-02A M=5.777e-07
I7318 0 n7319 2.976e-02A M=1.285e-06
I7319 0 n7320 2.976e-02A M=4.769e-07
I7320 0 n7321 2.976e-02A M=8.444e-07
I7321 0 n7322 2.976e-02A M=9.524e-07
I7322 0 n7323 2.976e-02A M=5.435e-07
I7323 0 n7324 2.976e-02A M=5.643e-07
I7324 0 n7325 2.976e-02A M=6.546e-07
I7325 0 n7326 2.976e-02A M=5.614e-07
I7326 0 n7327 2.976e-02A M=1.215e-06
I7327 0 n7328 2.976e-02A M=6.938e-07
I7328 0 n7329 2.976e-02A M=8.416e-07
I7329 0 n7330 2.976e-02A M=1.878e-06
I7330 0 n7331 2.976e-02A M=9.678e-07
I7331 0 n7332 2.976e-02A M=1.241e-06
I7332 0 n7333 2.976e-02A M=9.197e-07
I7333 0 n7334 2.976e-02A M=1.408e-06
I7334 0 n7335 2.976e-02A M=2.494e-07
I7335 0 n7336 2.976e-02A M=2.633e-07
I7336 0 n7337 2.976e-02A M=4.856e-07
I7337 0 n7338 2.976e-02A M=2.840e-06
I7338 0 n7339 2.976e-02A M=1.495e-06
I7339 0 n7340 2.976e-02A M=1.350e-06
I7340 0 n7341 2.976e-02A M=8.138e-07
I7341 0 n7342 2.976e-02A M=2.322e-07
I7342 0 n7343 2.976e-02A M=7.464e-07
I7343 0 n7344 2.976e-02A M=5.700e-07
I7344 0 n7345 2.976e-02A M=3.381e-07
I7345 0 n7346 2.976e-02A M=3.973e-07
I7346 0 n7347 2.976e-02A M=1.028e-06
I7347 0 n7348 2.976e-02A M=1.256e-06
I7348 0 n7349 2.976e-02A M=6.274e-07
I7349 0 n7350 2.976e-02A M=1.378e-06
I7350 0 n7351 2.976e-02A M=8.366e-07
I7351 0 n7352 2.976e-02A M=2.198e-06
I7352 0 n7353 2.976e-02A M=5.838e-07
I7353 0 n7354 2.976e-02A M=1.244e-06
I7354 0 n7355 2.976e-02A M=5.011e-07
I7355 0 n7356 2.976e-02A M=4.776e-07
I7356 0 n7357 2.976e-02A M=9.031e-07
I7357 0 n7358 2.976e-02A M=3.016e-07
I7358 0 n1 2.976e-02A M=1.692e-06
I7359 0 n7360 2.976e-02A M=3.038e-07
I7360 0 n7361 2.976e-02A M=1.520e-06
I7361 0 n7362 2.976e-02A M=5.084e-07
I7362 0 n7363 2.976e-02A M=1.454e-06
I7363 0 n7364 2.976e-02A M=1.436e-06
I7364 0 n7365 2.976e-02A M=1.165e-06
I7365 0 n7366 2.976e-02A M=4.343e-07
I7366 0 n7367 2.976e-02A M=8.132e-07
I7367 0 n7368 2.976e-02A M=6.955e-07
I7368 0 n7369 2.976e-02A M=9.732e-07
I7369 0 n7370 2.976e-02A M=1.566e-06
I7370 0 n7371 2.976e-02A M=1.732e-06
I7371 0 n7372 2.976e-02A M=7.832e-07
I7372 0 n7373 2.976e-02A M=2.188e-07
I7373 0 n7374 2.976e-02A M=1.016e-06
I7374 0 n7375 2.976e-02A M=8.235e-07
I7375 0 n7376 2.976e-02A M=5.771e-07
I7376 0 n7377 2.976e-02A M=6.190e-07
I7377 0 n7378 2.976e-02A M=1.513e-06
I7378 0 n7379 2.976e-02A M=8.198e-07
I7379 0 n7380 2.976e-02A M=1.421e-06
I7380 0 n7381 2.976e-02A M=1.052e-06
I7381 0 n7382 2.976e-02A M=1.065e-06
I7382 0 n7383 2.976e-02A M=1.871e-06
I7383 0 n7384 2.976e-02A M=8.737e-07
I7384 0 n7385 2.976e-02A M=8.845e-07
I7385 0 n7386 2.976e-02A M=5.056e-07
I7386 0 n7387 2.976e-02A M=1.211e-06
I7387 0 n7388 2.976e-02A M=4.795e-07
I7388 0 n7389 2.976e-02A M=5.676e-07
I7389 0 n7390 2.976e-02A M=2.304e-06
I7390 0 n7391 2.976e-02A M=1.222e-06
I7391 0 n7392 2.976e-02A M=1.118e-06
I7392 0 n7393 2.976e-02A M=2.474e-07
I7393 0 n7394 2.976e-02A M=3.583e-07
I7394 0 n7395 2.976e-02A M=1.240e-06
I7395 0 n7396 2.976e-02A M=7.290e-07
I7396 0 n7397 2.976e-02A M=1.382e-06
I7397 0 n7398 2.976e-02A M=1.176e-06
I7398 0 n7399 2.976e-02A M=6.219e-07
I7399 0 n7400 2.976e-02A M=1.348e-06
I7400 0 n7401 2.976e-02A M=1.185e-06
I7401 0 n7402 2.976e-02A M=9.452e-07
I7402 0 n7403 2.976e-02A M=1.178e-06
I7403 0 n7404 2.976e-02A M=2.067e-06
I7404 0 n7405 2.976e-02A M=8.935e-07
I7405 0 n7406 2.976e-02A M=1.506e-06
I7406 0 n7407 2.976e-02A M=9.980e-07
I7407 0 n7408 2.976e-02A M=4.620e-07
I7408 0 n7409 2.976e-02A M=1.189e-06
I7409 0 n7410 2.976e-02A M=5.474e-07
I7410 0 n7411 2.976e-02A M=5.839e-07
I7411 0 n7412 2.976e-02A M=4.622e-07
I7412 0 n7413 2.976e-02A M=7.976e-07
I7413 0 n7414 2.976e-02A M=9.684e-07
I7414 0 n7415 2.976e-02A M=8.500e-07
I7415 0 n7416 2.976e-02A M=1.001e-06
I7416 0 n7417 2.976e-02A M=1.287e-06
I7417 0 n7418 2.976e-02A M=7.768e-07
I7418 0 n7419 2.976e-02A M=1.273e-06
I7419 0 n7420 2.976e-02A M=9.609e-07
I7420 0 n7421 2.976e-02A M=3.158e-07
I7421 0 n7422 2.976e-02A M=3.483e-07
I7422 0 n7423 2.976e-02A M=4.498e-07
I7423 0 n7424 2.976e-02A M=1.500e-06
I7424 0 n7425 2.976e-02A M=1.452e-06
I7425 0 n7426 2.976e-02A M=1.680e-06
I7426 0 n7427 2.976e-02A M=2.822e-07
I7427 0 n7428 2.976e-02A M=6.494e-07
I7428 0 n7429 2.976e-02A M=3.633e-07
I7429 0 n7430 2.976e-02A M=2.643e-06
I7430 0 n7431 2.976e-02A M=9.018e-07
I7431 0 n7432 2.976e-02A M=7.036e-07
I7432 0 n7433 2.976e-02A M=1.018e-06
I7433 0 n7434 2.976e-02A M=6.292e-07
I7434 0 n7435 2.976e-02A M=7.245e-07
I7435 0 n7436 2.976e-02A M=1.430e-06
I7436 0 n7437 2.976e-02A M=7.339e-07
I7437 0 n7438 2.976e-02A M=6.708e-07
I7438 0 n7439 2.976e-02A M=4.812e-07
I7439 0 n7440 2.976e-02A M=1.634e-06
I7440 0 n7441 2.976e-02A M=1.640e-06
I7441 0 n7442 2.976e-02A M=6.083e-07
I7442 0 n7443 2.976e-02A M=4.836e-07
I7443 0 n7444 2.976e-02A M=5.349e-07
I7444 0 n7445 2.976e-02A M=9.998e-07
I7445 0 n7446 2.976e-02A M=2.013e-06
I7446 0 n7447 2.976e-02A M=8.874e-07
I7447 0 n7448 2.976e-02A M=2.197e-06
I7448 0 n7449 2.976e-02A M=2.239e-06
I7449 0 n7450 2.976e-02A M=9.020e-07
I7450 0 n7451 2.976e-02A M=8.751e-07
I7451 0 n7452 2.976e-02A M=1.687e-06
I7452 0 n7453 2.976e-02A M=4.882e-07
I7453 0 n7454 2.976e-02A M=1.472e-06
I7454 0 n7455 2.976e-02A M=7.809e-07
I7455 0 n7456 2.976e-02A M=1.658e-06
I7456 0 n7457 2.976e-02A M=5.311e-07
I7457 0 n7458 2.976e-02A M=8.339e-07
I7458 0 n7459 2.976e-02A M=7.621e-07
I7459 0 n7460 2.976e-02A M=7.168e-07
I7460 0 n7461 2.976e-02A M=4.730e-07
I7461 0 n7462 2.976e-02A M=1.337e-06
I7462 0 n7463 2.976e-02A M=1.249e-06
I7463 0 n7464 2.976e-02A M=1.161e-06
I7464 0 n7465 2.976e-02A M=2.178e-06
I7465 0 n7466 2.976e-02A M=7.020e-07
I7466 0 n7467 2.976e-02A M=7.818e-07
I7467 0 n7468 2.976e-02A M=1.127e-06
I7468 0 n7469 2.976e-02A M=1.060e-06
I7469 0 n7470 2.976e-02A M=5.639e-07
I7470 0 n7471 2.976e-02A M=7.437e-07
I7471 0 n7472 2.976e-02A M=8.445e-07
I7472 0 n7473 2.976e-02A M=1.233e-06
I7473 0 n7474 2.976e-02A M=1.093e-06
I7474 0 n7475 2.976e-02A M=6.380e-07
I7475 0 n7476 2.976e-02A M=5.688e-07
I7476 0 n7477 2.976e-02A M=7.709e-07
I7477 0 n7478 2.976e-02A M=1.573e-06
I7478 0 n7479 2.976e-02A M=1.461e-06
I7479 0 n7480 2.976e-02A M=8.074e-07
I7480 0 n7481 2.976e-02A M=9.682e-07
I7481 0 n7482 2.976e-02A M=8.159e-07
I7482 0 n7483 2.976e-02A M=9.980e-07
I7483 0 n7484 2.976e-02A M=1.150e-06
I7484 0 n7485 2.976e-02A M=5.322e-07
I7485 0 n7486 2.976e-02A M=8.742e-07
I7486 0 n7487 2.976e-02A M=8.402e-07
I7487 0 n7488 2.976e-02A M=1.196e-06
I7488 0 n7489 2.976e-02A M=8.114e-07
I7489 0 n7490 2.976e-02A M=1.231e-06
I7490 0 n7491 2.976e-02A M=5.834e-07
I7491 0 n7492 2.976e-02A M=3.995e-07
I7492 0 n7493 2.976e-02A M=1.013e-06
I7493 0 n7494 2.976e-02A M=1.430e-06
I7494 0 n7495 2.976e-02A M=8.803e-07
I7495 0 n7496 2.976e-02A M=1.011e-06
I7496 0 n7497 2.976e-02A M=9.533e-07
I7497 0 n7498 2.976e-02A M=1.042e-06
I7498 0 n7499 2.976e-02A M=1.331e-06
I7499 0 n7500 2.976e-02A M=5.227e-07
I7500 0 n7501 2.976e-02A M=1.380e-06
I7501 0 n7502 2.976e-02A M=4.645e-07
I7502 0 n7503 2.976e-02A M=1.558e-06
I7503 0 n7504 2.976e-02A M=4.918e-07
I7504 0 n7505 2.976e-02A M=1.587e-06
I7505 0 n7506 2.976e-02A M=1.501e-06
I7506 0 n7507 2.976e-02A M=4.070e-07
I7507 0 n7508 2.976e-02A M=1.098e-06
I7508 0 n7509 2.976e-02A M=7.549e-07
I7509 0 n7510 2.976e-02A M=1.974e-06
I7510 0 n7511 2.976e-02A M=1.581e-06
I7511 0 n7512 2.976e-02A M=7.516e-07
I7512 0 n7513 2.976e-02A M=1.538e-07
I7513 0 n7514 2.976e-02A M=1.302e-06
I7514 0 n1 2.976e-02A M=5.050e-07
I7515 0 n7516 2.976e-02A M=8.181e-07
I7516 0 n7517 2.976e-02A M=4.546e-07
I7517 0 n7518 2.976e-02A M=1.881e-06
I7518 0 n7519 2.976e-02A M=4.569e-07
I7519 0 n7520 2.976e-02A M=1.151e-06
I7520 0 n7521 2.976e-02A M=3.993e-07
I7521 0 n7522 2.976e-02A M=1.542e-06
I7522 0 n7523 2.976e-02A M=8.970e-07
I7523 0 n7524 2.976e-02A M=1.708e-06
I7524 0 n7525 2.976e-02A M=9.065e-07
I7525 0 n7526 2.976e-02A M=6.486e-07
I7526 0 n7527 2.976e-02A M=1.114e-06
I7527 0 n7528 2.976e-02A M=8.716e-07
I7528 0 n7529 2.976e-02A M=9.988e-07
I7529 0 n7530 2.976e-02A M=4.090e-07
I7530 0 n7531 2.976e-02A M=1.074e-06
I7531 0 n7532 2.976e-02A M=5.143e-07
I7532 0 n7533 2.976e-02A M=7.824e-07
I7533 0 n7534 2.976e-02A M=8.239e-07
I7534 0 n7535 2.976e-02A M=1.250e-06
I7535 0 n7536 2.976e-02A M=8.255e-07
I7536 0 n7537 2.976e-02A M=1.160e-06
I7537 0 n7538 2.976e-02A M=8.257e-07
I7538 0 n7539 2.976e-02A M=1.288e-06
I7539 0 n7540 2.976e-02A M=4.684e-07
I7540 0 n7541 2.976e-02A M=9.200e-07
I7541 0 n7542 2.976e-02A M=1.405e-06
I7542 0 n7543 2.976e-02A M=9.789e-07
I7543 0 n7544 2.976e-02A M=1.065e-06
I7544 0 n7545 2.976e-02A M=7.058e-07
I7545 0 n7546 2.976e-02A M=4.744e-07
I7546 0 n7547 2.976e-02A M=4.388e-07
I7547 0 n7548 2.976e-02A M=1.015e-06
I7548 0 n7549 2.976e-02A M=4.453e-07
I7549 0 n7550 2.976e-02A M=1.055e-06
I7550 0 n7551 2.976e-02A M=1.123e-06
I7551 0 n7552 2.976e-02A M=1.034e-06
I7552 0 n7553 2.976e-02A M=9.519e-07
I7553 0 n7554 2.976e-02A M=5.281e-07
I7554 0 n7555 2.976e-02A M=6.285e-07
I7555 0 n7556 2.976e-02A M=7.180e-07
I7556 0 n7557 2.976e-02A M=4.330e-07
I7557 0 n7558 2.976e-02A M=7.274e-07
I7558 0 n7559 2.976e-02A M=9.633e-07
I7559 0 n7560 2.976e-02A M=8.713e-07
I7560 0 n7561 2.976e-02A M=5.816e-07
I7561 0 n7562 2.976e-02A M=6.193e-07
I7562 0 n7563 2.976e-02A M=8.196e-07
I7563 0 n7564 2.976e-02A M=6.384e-07
I7564 0 n7565 2.976e-02A M=9.597e-07
I7565 0 n7566 2.976e-02A M=1.050e-06
I7566 0 n7567 2.976e-02A M=5.685e-07
I7567 0 n7568 2.976e-02A M=6.428e-07
I7568 0 n7569 2.976e-02A M=4.103e-07
I7569 0 n7570 2.976e-02A M=2.550e-07
I7570 0 n7571 2.976e-02A M=8.835e-07
I7571 0 n7572 2.976e-02A M=3.101e-07
I7572 0 n7573 2.976e-02A M=2.855e-06
I7573 0 n7574 2.976e-02A M=7.585e-07
I7574 0 n7575 2.976e-02A M=8.891e-07
I7575 0 n7576 2.976e-02A M=9.909e-07
I7576 0 n7577 2.976e-02A M=7.193e-07
I7577 0 n7578 2.976e-02A M=1.138e-06
I7578 0 n7579 2.976e-02A M=1.218e-06
I7579 0 n7580 2.976e-02A M=1.008e-06
I7580 0 n7581 2.976e-02A M=1.334e-06
I7581 0 n7582 2.976e-02A M=9.243e-07
I7582 0 n7583 2.976e-02A M=3.699e-07
I7583 0 n7584 2.976e-02A M=1.244e-06
I7584 0 n7585 2.976e-02A M=1.415e-06
I7585 0 n7586 2.976e-02A M=3.853e-07
I7586 0 n7587 2.976e-02A M=1.441e-07
I7587 0 n7588 2.976e-02A M=3.244e-07
I7588 0 n7589 2.976e-02A M=5.230e-07
I7589 0 n7590 2.976e-02A M=1.142e-06
I7590 0 n7591 2.976e-02A M=5.125e-07
I7591 0 n7592 2.976e-02A M=4.832e-07
I7592 0 n7593 2.976e-02A M=9.224e-07
I7593 0 n7594 2.976e-02A M=1.149e-06
I7594 0 n7595 2.976e-02A M=5.284e-07
I7595 0 n7596 2.976e-02A M=9.653e-07
I7596 0 n7597 2.976e-02A M=1.588e-06
I7597 0 n7598 2.976e-02A M=1.690e-06
I7598 0 n7599 2.976e-02A M=2.368e-06
I7599 0 n7600 2.976e-02A M=2.529e-06
I7600 0 n7601 2.976e-02A M=3.046e-07
I7601 0 n7602 2.976e-02A M=1.235e-06
I7602 0 n7603 2.976e-02A M=1.116e-06
I7603 0 n7604 2.976e-02A M=4.206e-07
I7604 0 n7605 2.976e-02A M=2.353e-06
I7605 0 n7606 2.976e-02A M=7.541e-07
I7606 0 n7607 2.976e-02A M=1.275e-06
I7607 0 n7608 2.976e-02A M=3.515e-07
I7608 0 n7609 2.976e-02A M=7.981e-07
I7609 0 n7610 2.976e-02A M=9.713e-07
I7610 0 n7611 2.976e-02A M=5.022e-07
I7611 0 n7612 2.976e-02A M=1.307e-06
I7612 0 n7613 2.976e-02A M=1.086e-06
I7613 0 n7614 2.976e-02A M=6.084e-07
I7614 0 n7615 2.976e-02A M=9.227e-07
I7615 0 n7616 2.976e-02A M=1.991e-06
I7616 0 n7617 2.976e-02A M=1.260e-06
I7617 0 n7618 2.976e-02A M=1.329e-06
I7618 0 n7619 2.976e-02A M=8.535e-07
I7619 0 n7620 2.976e-02A M=6.375e-07
I7620 0 n7621 2.976e-02A M=2.284e-06
I7621 0 n7622 2.976e-02A M=9.747e-07
I7622 0 n7623 2.976e-02A M=3.618e-07
I7623 0 n7624 2.976e-02A M=8.435e-07
I7624 0 n7625 2.976e-02A M=1.628e-06
I7625 0 n7626 2.976e-02A M=1.243e-06
I7626 0 n7627 2.976e-02A M=1.376e-06
I7627 0 n7628 2.976e-02A M=5.981e-07
I7628 0 n7629 2.976e-02A M=1.293e-06
I7629 0 n7630 2.976e-02A M=5.411e-07
I7630 0 n7631 2.976e-02A M=1.370e-06
I7631 0 n7632 2.976e-02A M=1.120e-06
I7632 0 n7633 2.976e-02A M=2.084e-06
I7633 0 n7634 2.976e-02A M=1.301e-06
I7634 0 n7635 2.976e-02A M=1.825e-06
I7635 0 n7636 2.976e-02A M=5.383e-07
I7636 0 n7637 2.976e-02A M=5.546e-07
I7637 0 n7638 2.976e-02A M=8.041e-07
I7638 0 n7639 2.976e-02A M=1.294e-06
I7639 0 n7640 2.976e-02A M=1.198e-06
I7640 0 n7641 2.976e-02A M=8.128e-07
I7641 0 n7642 2.976e-02A M=6.032e-07
I7642 0 n7643 2.976e-02A M=5.510e-07
I7643 0 n7644 2.976e-02A M=8.744e-07
I7644 0 n7645 2.976e-02A M=4.911e-07
I7645 0 n7646 2.976e-02A M=1.027e-06
I7646 0 n7647 2.976e-02A M=5.796e-07
I7647 0 n7648 2.976e-02A M=1.100e-06
I7648 0 n7649 2.976e-02A M=6.398e-07
I7649 0 n7650 2.976e-02A M=8.292e-07
I7650 0 n7651 2.976e-02A M=1.153e-06
I7651 0 n7652 2.976e-02A M=1.152e-06
I7652 0 n7653 2.976e-02A M=5.723e-07
I7653 0 n7654 2.976e-02A M=2.241e-06
I7654 0 n7655 2.976e-02A M=1.248e-06
I7655 0 n7656 2.976e-02A M=3.017e-07
I7656 0 n1 2.976e-02A M=6.673e-07
I7657 0 n7658 2.976e-02A M=1.191e-07
I7658 0 n7659 2.976e-02A M=1.161e-06
I7659 0 n7660 2.976e-02A M=1.148e-06
I7660 0 n7661 2.976e-02A M=2.136e-06
I7661 0 n7662 2.976e-02A M=1.077e-06
I7662 0 n1 2.976e-02A M=5.576e-07
I7663 0 n7664 2.976e-02A M=6.536e-07
I7664 0 n7665 2.976e-02A M=8.484e-07
I7665 0 n1 2.976e-02A M=9.278e-07
I7666 0 n7667 2.976e-02A M=1.564e-06
I7667 0 n7668 2.976e-02A M=1.658e-06
I7668 0 n7669 2.976e-02A M=4.194e-07
I7669 0 n7670 2.976e-02A M=3.392e-07
I7670 0 n7671 2.976e-02A M=1.062e-06
I7671 0 n1 2.976e-02A M=3.988e-07
I7672 0 n7673 2.976e-02A M=3.969e-07
I7673 0 n7674 2.976e-02A M=1.123e-06
I7674 0 n7675 2.976e-02A M=7.594e-07
I7675 0 n7676 2.976e-02A M=5.601e-07
I7676 0 n7677 2.976e-02A M=5.698e-07
I7677 0 n7678 2.976e-02A M=6.344e-07
I7678 0 n7679 2.976e-02A M=4.000e-07
I7679 0 n7680 2.976e-02A M=5.852e-07
I7680 0 n7681 2.976e-02A M=1.139e-06
I7681 0 n7682 2.976e-02A M=8.674e-07
I7682 0 n7683 2.976e-02A M=9.235e-07
I7683 0 n7684 2.976e-02A M=7.192e-07
I7684 0 n7685 2.976e-02A M=9.047e-07
I7685 0 n7686 2.976e-02A M=1.986e-06
I7686 0 n7687 2.976e-02A M=1.550e-06
I7687 0 n7688 2.976e-02A M=1.161e-06
I7688 0 n7689 2.976e-02A M=2.423e-07
I7689 0 n7690 2.976e-02A M=1.869e-07
I7690 0 n7691 2.976e-02A M=3.734e-07
I7691 0 n7692 2.976e-02A M=9.912e-07
I7692 0 n7693 2.976e-02A M=8.905e-07
I7693 0 n7694 2.976e-02A M=3.963e-07
I7694 0 n7695 2.976e-02A M=7.328e-07
I7695 0 n7696 2.976e-02A M=6.905e-07
I7696 0 n7697 2.976e-02A M=2.717e-07
I7697 0 n7698 2.976e-02A M=2.036e-06
I7698 0 n7699 2.976e-02A M=1.102e-06
I7699 0 n7700 2.976e-02A M=8.297e-07
I7700 0 n7701 2.976e-02A M=1.173e-06
I7701 0 n7702 2.976e-02A M=8.486e-07
I7702 0 n7703 2.976e-02A M=5.647e-07
I7703 0 n7704 2.976e-02A M=9.189e-07
I7704 0 n7705 2.976e-02A M=1.018e-06
I7705 0 n7706 2.976e-02A M=7.757e-07
I7706 0 n7707 2.976e-02A M=1.190e-06
I7707 0 n7708 2.976e-02A M=9.113e-07
I7708 0 n7709 2.976e-02A M=1.876e-06
I7709 0 n7710 2.976e-02A M=9.122e-07
I7710 0 n7711 2.976e-02A M=1.709e-06
I7711 0 n7712 2.976e-02A M=6.687e-07
I7712 0 n7713 2.976e-02A M=1.410e-06
I7713 0 n7714 2.976e-02A M=9.542e-07
I7714 0 n7715 2.976e-02A M=9.616e-07
I7715 0 n7716 2.976e-02A M=1.284e-06
I7716 0 n7717 2.976e-02A M=1.608e-06
I7717 0 n7718 2.976e-02A M=4.990e-07
I7718 0 n7719 2.976e-02A M=7.244e-07
I7719 0 n7720 2.976e-02A M=4.080e-07
I7720 0 n7721 2.976e-02A M=5.511e-07
I7721 0 n7722 2.976e-02A M=1.248e-06
I7722 0 n7723 2.976e-02A M=3.098e-06
I7723 0 n7724 2.976e-02A M=1.420e-06
I7724 0 n7725 2.976e-02A M=1.398e-06
I7725 0 n7726 2.976e-02A M=1.102e-06
I7726 0 n7727 2.976e-02A M=5.744e-07
I7727 0 n7728 2.976e-02A M=6.643e-07
I7728 0 n7729 2.976e-02A M=5.972e-07
I7729 0 n7730 2.976e-02A M=6.957e-08
I7730 0 n7731 2.976e-02A M=3.259e-07
I7731 0 n7732 2.976e-02A M=7.692e-07
I7732 0 n7733 2.976e-02A M=8.632e-07
I7733 0 n7734 2.976e-02A M=5.618e-07
I7734 0 n7735 2.976e-02A M=2.131e-06
I7735 0 n7736 2.976e-02A M=1.578e-06
I7736 0 n7737 2.976e-02A M=2.757e-06
I7737 0 n7738 2.976e-02A M=1.321e-06
I7738 0 n7739 2.976e-02A M=4.567e-07
I7739 0 n7740 2.976e-02A M=1.119e-06
I7740 0 n7741 2.976e-02A M=8.131e-07
I7741 0 n7742 2.976e-02A M=9.904e-07
I7742 0 n7743 2.976e-02A M=7.914e-07
I7743 0 n7744 2.976e-02A M=1.510e-06
I7744 0 n7745 2.976e-02A M=2.207e-06
I7745 0 n7746 2.976e-02A M=1.075e-06
I7746 0 n7747 2.976e-02A M=4.896e-07
I7747 0 n7748 2.976e-02A M=6.865e-07
I7748 0 n7749 2.976e-02A M=1.022e-06
I7749 0 n7750 2.976e-02A M=1.056e-06
I7750 0 n7751 2.976e-02A M=9.825e-07
I7751 0 n7752 2.976e-02A M=7.903e-07
I7752 0 n7753 2.976e-02A M=1.655e-06
I7753 0 n7754 2.976e-02A M=6.858e-07
I7754 0 n7755 2.976e-02A M=1.032e-06
I7755 0 n7756 2.976e-02A M=1.168e-06
I7756 0 n7757 2.976e-02A M=1.116e-06
I7757 0 n7758 2.976e-02A M=1.233e-06
I7758 0 n7759 2.976e-02A M=9.662e-07
I7759 0 n7760 2.976e-02A M=1.747e-06
I7760 0 n7761 2.976e-02A M=4.529e-07
I7761 0 n7762 2.976e-02A M=5.438e-07
I7762 0 n7763 2.976e-02A M=1.332e-06
I7763 0 n7764 2.976e-02A M=1.677e-06
I7764 0 n7765 2.976e-02A M=1.824e-06
I7765 0 n7766 2.976e-02A M=9.977e-07
I7766 0 n7767 2.976e-02A M=5.362e-07
I7767 0 n7768 2.976e-02A M=2.457e-07
I7768 0 n7769 2.976e-02A M=1.338e-06
I7769 0 n7770 2.976e-02A M=3.461e-07
I7770 0 n7771 2.976e-02A M=1.604e-06
I7771 0 n7772 2.976e-02A M=7.745e-07
I7772 0 n7773 2.976e-02A M=2.735e-07
I7773 0 n7774 2.976e-02A M=4.038e-07
I7774 0 n7775 2.976e-02A M=1.496e-06
I7775 0 n7776 2.976e-02A M=1.007e-06
I7776 0 n7777 2.976e-02A M=2.166e-06
I7777 0 n7778 2.976e-02A M=1.465e-06
I7778 0 n7779 2.976e-02A M=4.061e-07
I7779 0 n7780 2.976e-02A M=9.804e-07
I7780 0 n7781 2.976e-02A M=5.059e-07
I7781 0 n7782 2.976e-02A M=6.154e-07
I7782 0 n7783 2.976e-02A M=1.198e-06
I7783 0 n7784 2.976e-02A M=4.736e-07
I7784 0 n7785 2.976e-02A M=1.245e-06
I7785 0 n7786 2.976e-02A M=1.445e-06
I7786 0 n7787 2.976e-02A M=1.805e-06
I7787 0 n7788 2.976e-02A M=8.905e-07
I7788 0 n7789 2.976e-02A M=2.219e-06
I7789 0 n7790 2.976e-02A M=3.115e-07
I7790 0 n7791 2.976e-02A M=1.522e-07
I7791 0 n7792 2.976e-02A M=5.349e-07
I7792 0 n7793 2.976e-02A M=1.264e-06
I7793 0 n7794 2.976e-02A M=2.118e-07
I7794 0 n7795 2.976e-02A M=5.231e-07
I7795 0 n7796 2.976e-02A M=1.114e-06
I7796 0 n7797 2.976e-02A M=1.902e-06
I7797 0 n7798 2.976e-02A M=1.775e-06
I7798 0 n7799 2.976e-02A M=1.234e-06
I7799 0 n7800 2.976e-02A M=3.007e-07
I7800 0 n7801 2.976e-02A M=1.255e-06
I7801 0 n7802 2.976e-02A M=1.212e-06
I7802 0 n7803 2.976e-02A M=5.286e-07
I7803 0 n7804 2.976e-02A M=8.566e-07
I7804 0 n7805 2.976e-02A M=9.838e-07
I7805 0 n7806 2.976e-02A M=1.911e-06
I7806 0 n1 2.976e-02A M=3.627e-07
I7807 0 n7808 2.976e-02A M=2.222e-06
I7808 0 n7809 2.976e-02A M=4.761e-07
I7809 0 n7810 2.976e-02A M=1.605e-06
I7810 0 n7811 2.976e-02A M=1.464e-06
I7811 0 n7812 2.976e-02A M=7.727e-07
I7812 0 n7813 2.976e-02A M=9.829e-07
I7813 0 n7814 2.976e-02A M=9.861e-07
I7814 0 n7815 2.976e-02A M=3.563e-07
I7815 0 n7816 2.976e-02A M=4.682e-07
I7816 0 n7817 2.976e-02A M=8.995e-07
I7817 0 n7818 2.976e-02A M=2.375e-07
I7818 0 n7819 2.976e-02A M=6.766e-07
I7819 0 n7820 2.976e-02A M=1.255e-06
I7820 0 n7821 2.976e-02A M=4.247e-07
I7821 0 n7822 2.976e-02A M=8.593e-07
I7822 0 n7823 2.976e-02A M=6.122e-07
I7823 0 n7824 2.976e-02A M=4.446e-07
I7824 0 n7825 2.976e-02A M=1.516e-06
I7825 0 n1 2.976e-02A M=5.610e-07
I7826 0 n7827 2.976e-02A M=6.663e-07
I7827 0 n7828 2.976e-02A M=1.358e-06
I7828 0 n7829 2.976e-02A M=9.265e-07
I7829 0 n7830 2.976e-02A M=7.171e-07
I7830 0 n7831 2.976e-02A M=1.474e-06
I7831 0 n7832 2.976e-02A M=2.003e-06
I7832 0 n7833 2.976e-02A M=1.158e-06
I7833 0 n7834 2.976e-02A M=2.626e-07
I7834 0 n7835 2.976e-02A M=4.736e-07
I7835 0 n7836 2.976e-02A M=1.689e-06
I7836 0 n7837 2.976e-02A M=2.022e-06
I7837 0 n7838 2.976e-02A M=9.069e-07
I7838 0 n7839 2.976e-02A M=6.343e-07
I7839 0 n7840 2.976e-02A M=2.009e-06
I7840 0 n7841 2.976e-02A M=4.397e-07
I7841 0 n7842 2.976e-02A M=7.559e-07
I7842 0 n7843 2.976e-02A M=1.029e-06
I7843 0 n7844 2.976e-02A M=6.381e-07
I7844 0 n7845 2.976e-02A M=9.299e-07
I7845 0 n7846 2.976e-02A M=6.607e-07
I7846 0 n7847 2.976e-02A M=4.663e-07
I7847 0 n7848 2.976e-02A M=5.681e-07
I7848 0 n7849 2.976e-02A M=2.536e-06
I7849 0 n7850 2.976e-02A M=2.269e-06
I7850 0 n7851 2.976e-02A M=8.052e-07
I7851 0 n7852 2.976e-02A M=1.546e-06
I7852 0 n7853 2.976e-02A M=1.190e-06
I7853 0 n7854 2.976e-02A M=2.317e-06
I7854 0 n7855 2.976e-02A M=1.431e-06
I7855 0 n7856 2.976e-02A M=1.500e-06
I7856 0 n7857 2.976e-02A M=4.210e-07
I7857 0 n7858 2.976e-02A M=1.009e-06
I7858 0 n7859 2.976e-02A M=7.930e-07
I7859 0 n7860 2.976e-02A M=1.154e-06
I7860 0 n7861 2.976e-02A M=6.969e-07
I7861 0 n7862 2.976e-02A M=6.672e-07
I7862 0 n7863 2.976e-02A M=6.432e-07
I7863 0 n7864 2.976e-02A M=4.478e-07
I7864 0 n7865 2.976e-02A M=9.490e-07
I7865 0 n7866 2.976e-02A M=5.386e-07
I7866 0 n7867 2.976e-02A M=6.077e-07
I7867 0 n7868 2.976e-02A M=9.515e-07
I7868 0 n7869 2.976e-02A M=1.336e-06
I7869 0 n7870 2.976e-02A M=1.447e-06
I7870 0 n7871 2.976e-02A M=1.179e-06
I7871 0 n7872 2.976e-02A M=8.869e-07
I7872 0 n7873 2.976e-02A M=1.165e-06
I7873 0 n7874 2.976e-02A M=1.028e-06
I7874 0 n7875 2.976e-02A M=4.669e-07
I7875 0 n7876 2.976e-02A M=1.438e-06
I7876 0 n7877 2.976e-02A M=1.075e-06
I7877 0 n7878 2.976e-02A M=1.470e-06
I7878 0 n7879 2.976e-02A M=8.046e-07
I7879 0 n7880 2.976e-02A M=1.155e-06
I7880 0 n7881 2.976e-02A M=3.630e-07
I7881 0 n7882 2.976e-02A M=1.861e-06
I7882 0 n7883 2.976e-02A M=9.297e-07
I7883 0 n7884 2.976e-02A M=7.089e-07
I7884 0 n7885 2.976e-02A M=9.986e-07
I7885 0 n7886 2.976e-02A M=1.108e-06
I7886 0 n7887 2.976e-02A M=5.536e-07
I7887 0 n7888 2.976e-02A M=1.441e-06
I7888 0 n7889 2.976e-02A M=5.300e-07
I7889 0 n7890 2.976e-02A M=1.002e-06
I7890 0 n7891 2.976e-02A M=9.058e-07
I7891 0 n7892 2.976e-02A M=3.691e-07
I7892 0 n7893 2.976e-02A M=5.531e-07
I7893 0 n7894 2.976e-02A M=1.222e-06
I7894 0 n7895 2.976e-02A M=8.421e-07
I7895 0 n7896 2.976e-02A M=9.613e-07
I7896 0 n7897 2.976e-02A M=1.683e-06
I7897 0 n7898 2.976e-02A M=1.370e-06
I7898 0 n7899 2.976e-02A M=6.829e-07
I7899 0 n7900 2.976e-02A M=4.567e-07
I7900 0 n7901 2.976e-02A M=1.348e-06
I7901 0 n7902 2.976e-02A M=4.237e-07
I7902 0 n7903 2.976e-02A M=1.029e-06
I7903 0 n7904 2.976e-02A M=1.522e-06
I7904 0 n7905 2.976e-02A M=7.412e-07
I7905 0 n7906 2.976e-02A M=1.180e-06
I7906 0 n7907 2.976e-02A M=4.152e-07
I7907 0 n7908 2.976e-02A M=1.478e-06
I7908 0 n7909 2.976e-02A M=1.183e-06
I7909 0 n7910 2.976e-02A M=1.408e-06
I7910 0 n7911 2.976e-02A M=6.143e-07
I7911 0 n7912 2.976e-02A M=9.944e-07
I7912 0 n7913 2.976e-02A M=1.053e-06
I7913 0 n7914 2.976e-02A M=9.484e-07
I7914 0 n7915 2.976e-02A M=1.206e-06
I7915 0 n7916 2.976e-02A M=2.851e-08
I7916 0 n7917 2.976e-02A M=8.234e-07
I7917 0 n7918 2.976e-02A M=1.207e-06
I7918 0 n7919 2.976e-02A M=3.484e-07
I7919 0 n7920 2.976e-02A M=6.511e-07
I7920 0 n7921 2.976e-02A M=7.537e-07
I7921 0 n7922 2.976e-02A M=1.576e-06
I7922 0 n7923 2.976e-02A M=5.858e-07
I7923 0 n7924 2.976e-02A M=2.099e-06
I7924 0 n7925 2.976e-02A M=1.148e-06
I7925 0 n7926 2.976e-02A M=3.292e-07
I7926 0 n7927 2.976e-02A M=9.641e-07
I7927 0 n7928 2.976e-02A M=8.302e-07
I7928 0 n7929 2.976e-02A M=5.178e-07
I7929 0 n7930 2.976e-02A M=1.034e-06
I7930 0 n7931 2.976e-02A M=1.041e-06
I7931 0 n7932 2.976e-02A M=5.863e-07
I7932 0 n7933 2.976e-02A M=1.168e-06
I7933 0 n7934 2.976e-02A M=1.028e-06
I7934 0 n7935 2.976e-02A M=1.119e-06
I7935 0 n7936 2.976e-02A M=9.933e-07
I7936 0 n7937 2.976e-02A M=1.291e-06
I7937 0 n7938 2.976e-02A M=1.902e-06
I7938 0 n1 2.976e-02A M=8.455e-07
I7939 0 n7940 2.976e-02A M=4.854e-07
I7940 0 n7941 2.976e-02A M=7.771e-07
I7941 0 n7942 2.976e-02A M=1.853e-07
I7942 0 n7943 2.976e-02A M=4.712e-07
I7943 0 n7944 2.976e-02A M=4.998e-07
I7944 0 n7945 2.976e-02A M=1.876e-07
I7945 0 n7946 2.976e-02A M=6.624e-07
I7946 0 n7947 2.976e-02A M=1.038e-06
I7947 0 n7948 2.976e-02A M=1.052e-06
I7948 0 n7949 2.976e-02A M=1.082e-06
I7949 0 n7950 2.976e-02A M=8.409e-07
I7950 0 n7951 2.976e-02A M=1.255e-06
I7951 0 n7952 2.976e-02A M=6.414e-07
I7952 0 n7953 2.976e-02A M=5.953e-07
I7953 0 n7954 2.976e-02A M=1.434e-06
I7954 0 n7955 2.976e-02A M=4.020e-07
I7955 0 n7956 2.976e-02A M=8.956e-07
I7956 0 n7957 2.976e-02A M=8.795e-07
I7957 0 n7958 2.976e-02A M=6.071e-07
I7958 0 n7959 2.976e-02A M=1.215e-06
I7959 0 n7960 2.976e-02A M=9.190e-07
I7960 0 n7961 2.976e-02A M=8.318e-07
I7961 0 n7962 2.976e-02A M=6.217e-07
I7962 0 n7963 2.976e-02A M=8.332e-07
I7963 0 n7964 2.976e-02A M=6.619e-07
I7964 0 n7965 2.976e-02A M=3.967e-07
I7965 0 n7966 2.976e-02A M=1.776e-06
I7966 0 n7967 2.976e-02A M=5.473e-07
I7967 0 n7968 2.976e-02A M=1.459e-06
I7968 0 n7969 2.976e-02A M=1.249e-06
I7969 0 n7970 2.976e-02A M=7.431e-07
I7970 0 n7971 2.976e-02A M=4.115e-07
I7971 0 n7972 2.976e-02A M=3.317e-07
I7972 0 n7973 2.976e-02A M=1.122e-06
I7973 0 n7974 2.976e-02A M=1.035e-06
I7974 0 n7975 2.976e-02A M=6.196e-07
I7975 0 n7976 2.976e-02A M=1.062e-06
I7976 0 n7977 2.976e-02A M=1.007e-06
I7977 0 n7978 2.976e-02A M=6.824e-07
I7978 0 n7979 2.976e-02A M=4.080e-07
I7979 0 n7980 2.976e-02A M=4.399e-07
I7980 0 n7981 2.976e-02A M=1.112e-06
I7981 0 n7982 2.976e-02A M=6.414e-07
I7982 0 n7983 2.976e-02A M=1.472e-06
I7983 0 n7984 2.976e-02A M=4.651e-07
I7984 0 n7985 2.976e-02A M=5.185e-07
I7985 0 n7986 2.976e-02A M=2.676e-07
I7986 0 n7987 2.976e-02A M=3.398e-07
I7987 0 n7988 2.976e-02A M=8.779e-07
I7988 0 n7989 2.976e-02A M=7.090e-07
I7989 0 n7990 2.976e-02A M=1.219e-06
I7990 0 n7991 2.976e-02A M=1.244e-06
I7991 0 n7992 2.976e-02A M=6.295e-07
I7992 0 n7993 2.976e-02A M=8.855e-07
I7993 0 n7994 2.976e-02A M=1.120e-06
I7994 0 n7995 2.976e-02A M=5.021e-07
I7995 0 n7996 2.976e-02A M=6.254e-07
I7996 0 n7997 2.976e-02A M=1.191e-06
I7997 0 n7998 2.976e-02A M=5.113e-07
I7998 0 n7999 2.976e-02A M=1.622e-06
I7999 0 n8000 2.976e-02A M=7.915e-07
I8000 0 n8001 2.976e-02A M=4.627e-07
I8001 0 n8002 2.976e-02A M=1.489e-06
I8002 0 n8003 2.976e-02A M=1.173e-06
I8003 0 n8004 2.976e-02A M=1.410e-06
I8004 0 n8005 2.976e-02A M=6.948e-07
I8005 0 n8006 2.976e-02A M=1.344e-06
I8006 0 n8007 2.976e-02A M=3.262e-07
I8007 0 n8008 2.976e-02A M=1.383e-06
I8008 0 n8009 2.976e-02A M=1.623e-06
I8009 0 n8010 2.976e-02A M=1.485e-06
I8010 0 n8011 2.976e-02A M=5.388e-07
I8011 0 n8012 2.976e-02A M=1.351e-06
I8012 0 n8013 2.976e-02A M=1.350e-06
I8013 0 n8014 2.976e-02A M=7.921e-07
I8014 0 n8015 2.976e-02A M=4.867e-07
I8015 0 n8016 2.976e-02A M=3.358e-07
I8016 0 n8017 2.976e-02A M=1.300e-06
I8017 0 n8018 2.976e-02A M=1.254e-06
I8018 0 n8019 2.976e-02A M=7.777e-07
I8019 0 n8020 2.976e-02A M=9.437e-07
I8020 0 n8021 2.976e-02A M=6.240e-07
I8021 0 n8022 2.976e-02A M=7.386e-07
I8022 0 n8023 2.976e-02A M=1.213e-06
I8023 0 n8024 2.976e-02A M=3.256e-07
I8024 0 n8025 2.976e-02A M=1.201e-06
I8025 0 n8026 2.976e-02A M=7.565e-07
I8026 0 n8027 2.976e-02A M=2.179e-06
I8027 0 n8028 2.976e-02A M=1.486e-06
I8028 0 n8029 2.976e-02A M=2.182e-06
I8029 0 n8030 2.976e-02A M=3.756e-07
I8030 0 n8031 2.976e-02A M=1.009e-06
I8031 0 n8032 2.976e-02A M=1.223e-06
I8032 0 n8033 2.976e-02A M=4.855e-07
I8033 0 n8034 2.976e-02A M=1.871e-06
I8034 0 n8035 2.976e-02A M=1.497e-06
I8035 0 n8036 2.976e-02A M=9.460e-07
I8036 0 n8037 2.976e-02A M=1.566e-06
I8037 0 n8038 2.976e-02A M=1.242e-06
I8038 0 n8039 2.976e-02A M=3.360e-07
I8039 0 n8040 2.976e-02A M=1.614e-06
I8040 0 n8041 2.976e-02A M=8.769e-07
I8041 0 n8042 2.976e-02A M=6.633e-07
I8042 0 n8043 2.976e-02A M=7.020e-07
I8043 0 n8044 2.976e-02A M=5.206e-07
I8044 0 n8045 2.976e-02A M=1.167e-06
I8045 0 n8046 2.976e-02A M=1.883e-06
I8046 0 n8047 2.976e-02A M=4.481e-07
I8047 0 n8048 2.976e-02A M=1.423e-06
I8048 0 n8049 2.976e-02A M=9.216e-07
I8049 0 n8050 2.976e-02A M=3.392e-07
I8050 0 n8051 2.976e-02A M=1.533e-06
I8051 0 n8052 2.976e-02A M=9.892e-07
I8052 0 n8053 2.976e-02A M=1.238e-06
I8053 0 n8054 2.976e-02A M=2.761e-07
I8054 0 n8055 2.976e-02A M=9.362e-08
I8055 0 n8056 2.976e-02A M=7.718e-07
I8056 0 n8057 2.976e-02A M=1.331e-06
I8057 0 n8058 2.976e-02A M=1.058e-06
I8058 0 n8059 2.976e-02A M=1.064e-06
I8059 0 n8060 2.976e-02A M=7.125e-07
I8060 0 n8061 2.976e-02A M=8.303e-07
I8061 0 n8062 2.976e-02A M=1.606e-06
I8062 0 n8063 2.976e-02A M=5.895e-07
I8063 0 n8064 2.976e-02A M=2.873e-07
I8064 0 n8065 2.976e-02A M=4.793e-07
I8065 0 n8066 2.976e-02A M=1.860e-06
I8066 0 n8067 2.976e-02A M=9.930e-07
I8067 0 n8068 2.976e-02A M=1.104e-06
I8068 0 n8069 2.976e-02A M=7.210e-07
I8069 0 n8070 2.976e-02A M=3.556e-07
I8070 0 n8071 2.976e-02A M=2.005e-07
I8071 0 n8072 2.976e-02A M=1.023e-06
I8072 0 n8073 2.976e-02A M=4.102e-07
I8073 0 n8074 2.976e-02A M=8.362e-07
I8074 0 n8075 2.976e-02A M=8.057e-07
I8075 0 n8076 2.976e-02A M=1.030e-06
I8076 0 n8077 2.976e-02A M=8.188e-07
I8077 0 n8078 2.976e-02A M=1.053e-06
I8078 0 n8079 2.976e-02A M=1.648e-06
I8079 0 n8080 2.976e-02A M=1.209e-06
I8080 0 n8081 2.976e-02A M=1.597e-06
I8081 0 n8082 2.976e-02A M=6.713e-07
I8082 0 n8083 2.976e-02A M=1.366e-06
I8083 0 n8084 2.976e-02A M=9.593e-07
I8084 0 n8085 2.976e-02A M=7.823e-07
I8085 0 n8086 2.976e-02A M=6.863e-07
I8086 0 n8087 2.976e-02A M=1.430e-06
I8087 0 n8088 2.976e-02A M=5.645e-07
I8088 0 n8089 2.976e-02A M=2.105e-06
I8089 0 n8090 2.976e-02A M=1.359e-06
I8090 0 n8091 2.976e-02A M=1.475e-06
I8091 0 n8092 2.976e-02A M=7.592e-07
I8092 0 n8093 2.976e-02A M=8.607e-07
I8093 0 n8094 2.976e-02A M=6.221e-07
I8094 0 n8095 2.976e-02A M=1.683e-06
I8095 0 n8096 2.976e-02A M=9.482e-07
I8096 0 n8097 2.976e-02A M=1.499e-07
I8097 0 n8098 2.976e-02A M=5.174e-07
I8098 0 n8099 2.976e-02A M=3.083e-07
I8099 0 n8100 2.976e-02A M=8.234e-07
I8100 0 n8101 2.976e-02A M=1.549e-06
I8101 0 n8102 2.976e-02A M=1.190e-06
I8102 0 n8103 2.976e-02A M=7.780e-07
I8103 0 n8104 2.976e-02A M=7.054e-07
I8104 0 n8105 2.976e-02A M=7.703e-07
I8105 0 n8106 2.976e-02A M=9.988e-07
I8106 0 n8107 2.976e-02A M=5.761e-07
I8107 0 n8108 2.976e-02A M=1.921e-06
I8108 0 n8109 2.976e-02A M=9.327e-07
I8109 0 n8110 2.976e-02A M=1.493e-06
I8110 0 n8111 2.976e-02A M=9.993e-07
I8111 0 n8112 2.976e-02A M=6.825e-07
I8112 0 n8113 2.976e-02A M=6.481e-07
I8113 0 n8114 2.976e-02A M=3.010e-07
I8114 0 n8115 2.976e-02A M=1.539e-06
I8115 0 n8116 2.976e-02A M=4.940e-07
I8116 0 n8117 2.976e-02A M=1.732e-06
I8117 0 n8118 2.976e-02A M=1.652e-06
I8118 0 n8119 2.976e-02A M=1.002e-06
I8119 0 n8120 2.976e-02A M=1.376e-06
I8120 0 n8121 2.976e-02A M=1.812e-06
I8121 0 n8122 2.976e-02A M=1.012e-06
I8122 0 n8123 2.976e-02A M=4.968e-07
I8123 0 n8124 2.976e-02A M=9.051e-07
I8124 0 n8125 2.976e-02A M=6.042e-07
I8125 0 n8126 2.976e-02A M=1.319e-06
I8126 0 n8127 2.976e-02A M=1.109e-06
I8127 0 n8128 2.976e-02A M=1.366e-06
I8128 0 n8129 2.976e-02A M=1.278e-06
I8129 0 n8130 2.976e-02A M=1.646e-06
I8130 0 n8131 2.976e-02A M=3.926e-07
I8131 0 n8132 2.976e-02A M=1.849e-07
I8132 0 n8133 2.976e-02A M=5.811e-07
I8133 0 n8134 2.976e-02A M=7.916e-07
I8134 0 n8135 2.976e-02A M=7.805e-07
I8135 0 n8136 2.976e-02A M=1.022e-06
I8136 0 n8137 2.976e-02A M=3.020e-07
I8137 0 n8138 2.976e-02A M=1.423e-06
I8138 0 n8139 2.976e-02A M=7.098e-07
I8139 0 n8140 2.976e-02A M=1.232e-06
I8140 0 n8141 2.976e-02A M=9.960e-07
I8141 0 n8142 2.976e-02A M=2.998e-07
I8142 0 n8143 2.976e-02A M=1.152e-06
I8143 0 n8144 2.976e-02A M=9.159e-07
I8144 0 n8145 2.976e-02A M=5.629e-07
I8145 0 n8146 2.976e-02A M=2.398e-07
I8146 0 n8147 2.976e-02A M=1.397e-06
I8147 0 n8148 2.976e-02A M=6.326e-07
I8148 0 n8149 2.976e-02A M=8.175e-07
I8149 0 n8150 2.976e-02A M=8.541e-07
I8150 0 n8151 2.976e-02A M=9.879e-07
I8151 0 n8152 2.976e-02A M=1.232e-06
I8152 0 n8153 2.976e-02A M=2.055e-06
I8153 0 n8154 2.976e-02A M=1.192e-06
I8154 0 n8155 2.976e-02A M=1.217e-06
I8155 0 n8156 2.976e-02A M=5.826e-07
I8156 0 n8157 2.976e-02A M=1.226e-06
I8157 0 n8158 2.976e-02A M=9.656e-07
I8158 0 n8159 2.976e-02A M=1.122e-06
I8159 0 n8160 2.976e-02A M=5.119e-07
I8160 0 n8161 2.976e-02A M=8.551e-07
I8161 0 n8162 2.976e-02A M=1.261e-06
I8162 0 n8163 2.976e-02A M=3.068e-07
I8163 0 n8164 2.976e-02A M=6.763e-07
I8164 0 n8165 2.976e-02A M=6.280e-07
I8165 0 n8166 2.976e-02A M=6.969e-07
I8166 0 n8167 2.976e-02A M=1.924e-06
I8167 0 n8168 2.976e-02A M=1.109e-07
I8168 0 n8169 2.976e-02A M=1.057e-06
I8169 0 n8170 2.976e-02A M=1.138e-06
I8170 0 n8171 2.976e-02A M=1.380e-06
I8171 0 n8172 2.976e-02A M=2.041e-07
I8172 0 n8173 2.976e-02A M=8.880e-07
I8173 0 n8174 2.976e-02A M=1.316e-06
I8174 0 n8175 2.976e-02A M=9.538e-07
I8175 0 n8176 2.976e-02A M=1.061e-06
I8176 0 n8177 2.976e-02A M=1.092e-06
I8177 0 n8178 2.976e-02A M=1.308e-06
I8178 0 n8179 2.976e-02A M=5.974e-07
I8179 0 n8180 2.976e-02A M=8.163e-07
I8180 0 n8181 2.976e-02A M=5.807e-07
I8181 0 n8182 2.976e-02A M=9.041e-07
I8182 0 n8183 2.976e-02A M=1.577e-06
I8183 0 n8184 2.976e-02A M=1.774e-06
I8184 0 n8185 2.976e-02A M=4.401e-07
I8185 0 n8186 2.976e-02A M=5.740e-07
I8186 0 n8187 2.976e-02A M=1.697e-06
I8187 0 n8188 2.976e-02A M=1.428e-06
I8188 0 n8189 2.976e-02A M=9.402e-07
I8189 0 n8190 2.976e-02A M=8.040e-07
I8190 0 n8191 2.976e-02A M=3.503e-07
I8191 0 n8192 2.976e-02A M=8.223e-07
I8192 0 n8193 2.976e-02A M=5.379e-07
I8193 0 n8194 2.976e-02A M=2.291e-06
I8194 0 n8195 2.976e-02A M=3.980e-07
I8195 0 n8196 2.976e-02A M=2.072e-06
I8196 0 n8197 2.976e-02A M=4.762e-07
I8197 0 n8198 2.976e-02A M=6.692e-07
I8198 0 n8199 2.976e-02A M=1.039e-06
I8199 0 n8200 2.976e-02A M=9.675e-07
I8200 0 n8201 2.976e-02A M=4.992e-07
I8201 0 n8202 2.976e-02A M=1.396e-06
I8202 0 n8203 2.976e-02A M=2.398e-06
I8203 0 n8204 2.976e-02A M=1.077e-06
I8204 0 n8205 2.976e-02A M=6.006e-07
I8205 0 n8206 2.976e-02A M=1.047e-06
I8206 0 n8207 2.976e-02A M=1.601e-06
I8207 0 n8208 2.976e-02A M=6.009e-07
I8208 0 n8209 2.976e-02A M=2.195e-06
I8209 0 n8210 2.976e-02A M=7.265e-07
I8210 0 n8211 2.976e-02A M=2.782e-06
I8211 0 n8212 2.976e-02A M=1.275e-06
I8212 0 n8213 2.976e-02A M=4.230e-07
I8213 0 n8214 2.976e-02A M=1.691e-06
I8214 0 n8215 2.976e-02A M=7.046e-07
I8215 0 n8216 2.976e-02A M=1.608e-06
I8216 0 n8217 2.976e-02A M=1.866e-07
I8217 0 n8218 2.976e-02A M=4.917e-08
I8218 0 n8219 2.976e-02A M=5.441e-07
I8219 0 n8220 2.976e-02A M=1.230e-06
I8220 0 n8221 2.976e-02A M=2.032e-06
I8221 0 n8222 2.976e-02A M=1.357e-06
I8222 0 n8223 2.976e-02A M=7.357e-07
I8223 0 n8224 2.976e-02A M=8.597e-07
I8224 0 n8225 2.976e-02A M=8.222e-07
I8225 0 n8226 2.976e-02A M=6.762e-07
I8226 0 n8227 2.976e-02A M=6.390e-07
I8227 0 n8228 2.976e-02A M=4.982e-07
I8228 0 n8229 2.976e-02A M=4.149e-07
I8229 0 n8230 2.976e-02A M=4.051e-07
I8230 0 n8231 2.976e-02A M=1.072e-06
I8231 0 n8232 2.976e-02A M=1.004e-06
I8232 0 n8233 2.976e-02A M=2.312e-07
I8233 0 n8234 2.976e-02A M=1.426e-06
I8234 0 n8235 2.976e-02A M=8.799e-07
I8235 0 n8236 2.976e-02A M=1.027e-06
I8236 0 n8237 2.976e-02A M=1.091e-06
I8237 0 n8238 2.976e-02A M=2.104e-06
I8238 0 n8239 2.976e-02A M=9.711e-07
I8239 0 n8240 2.976e-02A M=1.332e-06
I8240 0 n8241 2.976e-02A M=5.763e-07
I8241 0 n8242 2.976e-02A M=1.637e-06
I8242 0 n8243 2.976e-02A M=9.211e-07
I8243 0 n8244 2.976e-02A M=5.966e-07
I8244 0 n8245 2.976e-02A M=1.446e-06
I8245 0 n8246 2.976e-02A M=7.274e-07
I8246 0 n8247 2.976e-02A M=5.752e-07
I8247 0 n8248 2.976e-02A M=5.628e-07
I8248 0 n8249 2.976e-02A M=1.776e-06
I8249 0 n8250 2.976e-02A M=6.455e-07
I8250 0 n8251 2.976e-02A M=2.080e-06
I8251 0 n8252 2.976e-02A M=6.941e-07
I8252 0 n8253 2.976e-02A M=6.554e-07
I8253 0 n8254 2.976e-02A M=8.357e-07
I8254 0 n8255 2.976e-02A M=7.659e-07
I8255 0 n8256 2.976e-02A M=7.018e-07
I8256 0 n8257 2.976e-02A M=1.717e-06
I8257 0 n8258 2.976e-02A M=5.295e-07
I8258 0 n8259 2.976e-02A M=2.127e-07
I8259 0 n8260 2.976e-02A M=1.462e-06
I8260 0 n8261 2.976e-02A M=1.221e-06
I8261 0 n8262 2.976e-02A M=1.404e-07
I8262 0 n8263 2.976e-02A M=1.779e-06
I8263 0 n8264 2.976e-02A M=9.885e-07
I8264 0 n8265 2.976e-02A M=5.906e-07
I8265 0 n8266 2.976e-02A M=1.097e-06
I8266 0 n8267 2.976e-02A M=2.135e-06
I8267 0 n8268 2.976e-02A M=7.794e-07
I8268 0 n8269 2.976e-02A M=2.273e-07
I8269 0 n8270 2.976e-02A M=7.562e-07
I8270 0 n8271 2.976e-02A M=1.009e-06
I8271 0 n8272 2.976e-02A M=1.077e-06
I8272 0 n8273 2.976e-02A M=1.897e-06
I8273 0 n8274 2.976e-02A M=4.341e-07
I8274 0 n8275 2.976e-02A M=1.435e-06
I8275 0 n8276 2.976e-02A M=1.296e-06
I8276 0 n8277 2.976e-02A M=8.529e-07
I8277 0 n8278 2.976e-02A M=1.005e-06
I8278 0 n8279 2.976e-02A M=1.847e-07
I8279 0 n8280 2.976e-02A M=3.579e-07
I8280 0 n8281 2.976e-02A M=8.749e-07
I8281 0 n8282 2.976e-02A M=9.731e-07
I8282 0 n8283 2.976e-02A M=1.260e-06
I8283 0 n8284 2.976e-02A M=1.347e-06
I8284 0 n8285 2.976e-02A M=6.752e-07
I8285 0 n8286 2.976e-02A M=5.426e-07
I8286 0 n8287 2.976e-02A M=9.413e-07
I8287 0 n8288 2.976e-02A M=8.981e-07
I8288 0 n8289 2.976e-02A M=5.531e-07
I8289 0 n8290 2.976e-02A M=6.316e-07
I8290 0 n8291 2.976e-02A M=9.583e-07
I8291 0 n8292 2.976e-02A M=1.059e-06
I8292 0 n8293 2.976e-02A M=1.306e-06
I8293 0 n8294 2.976e-02A M=4.084e-07
I8294 0 n8295 2.976e-02A M=7.025e-07
I8295 0 n8296 2.976e-02A M=2.998e-06
I8296 0 n8297 2.976e-02A M=9.305e-07
I8297 0 n8298 2.976e-02A M=2.316e-07
I8298 0 n8299 2.976e-02A M=1.640e-06
I8299 0 n8300 2.976e-02A M=5.490e-07
I8300 0 n8301 2.976e-02A M=1.508e-06
I8301 0 n8302 2.976e-02A M=5.213e-07
I8302 0 n8303 2.976e-02A M=5.682e-07
I8303 0 n8304 2.976e-02A M=5.614e-07
I8304 0 n8305 2.976e-02A M=1.520e-06
I8305 0 n8306 2.976e-02A M=3.270e-07
I8306 0 n8307 2.976e-02A M=1.247e-06
I8307 0 n8308 2.976e-02A M=7.401e-07
I8308 0 n8309 2.976e-02A M=8.496e-07
I8309 0 n8310 2.976e-02A M=6.512e-07
I8310 0 n8311 2.976e-02A M=4.617e-07
I8311 0 n8312 2.976e-02A M=2.019e-06
I8312 0 n8313 2.976e-02A M=7.104e-07
I8313 0 n8314 2.976e-02A M=1.328e-06
I8314 0 n8315 2.976e-02A M=4.541e-07
I8315 0 n8316 2.976e-02A M=1.714e-06
I8316 0 n8317 2.976e-02A M=8.444e-07
I8317 0 n8318 2.976e-02A M=7.923e-07
I8318 0 n8319 2.976e-02A M=7.954e-07
I8319 0 n8320 2.976e-02A M=8.273e-07
I8320 0 n8321 2.976e-02A M=1.487e-06
I8321 0 n8322 2.976e-02A M=6.010e-07
I8322 0 n8323 2.976e-02A M=1.705e-06
I8323 0 n8324 2.976e-02A M=1.100e-06
I8324 0 n8325 2.976e-02A M=6.657e-07
I8325 0 n8326 2.976e-02A M=2.807e-06
I8326 0 n8327 2.976e-02A M=8.329e-07
I8327 0 n8328 2.976e-02A M=1.310e-06
I8328 0 n8329 2.976e-02A M=8.375e-07
I8329 0 n8330 2.976e-02A M=8.945e-07
I8330 0 n8331 2.976e-02A M=9.520e-07
I8331 0 n8332 2.976e-02A M=4.570e-07
I8332 0 n8333 2.976e-02A M=1.328e-06
I8333 0 n8334 2.976e-02A M=2.020e-06
I8334 0 n8335 2.976e-02A M=1.295e-06
I8335 0 n1 2.976e-02A M=7.580e-07
I8336 0 n8337 2.976e-02A M=7.282e-07
I8337 0 n8338 2.976e-02A M=5.484e-07
I8338 0 n8339 2.976e-02A M=1.571e-06
I8339 0 n8340 2.976e-02A M=3.353e-07
I8340 0 n8341 2.976e-02A M=7.773e-07
I8341 0 n8342 2.976e-02A M=2.163e-06
I8342 0 n8343 2.976e-02A M=1.448e-06
I8343 0 n8344 2.976e-02A M=1.218e-06
I8344 0 n8345 2.976e-02A M=1.365e-06
I8345 0 n8346 2.976e-02A M=7.695e-07
I8346 0 n8347 2.976e-02A M=6.941e-07
I8347 0 n8348 2.976e-02A M=1.470e-06
I8348 0 n8349 2.976e-02A M=1.879e-06
I8349 0 n8350 2.976e-02A M=4.187e-07
I8350 0 n8351 2.976e-02A M=1.778e-06
I8351 0 n8352 2.976e-02A M=1.124e-06
I8352 0 n8353 2.976e-02A M=7.452e-07
I8353 0 n8354 2.976e-02A M=1.626e-06
I8354 0 n8355 2.976e-02A M=5.695e-07
I8355 0 n8356 2.976e-02A M=1.031e-06
I8356 0 n8357 2.976e-02A M=1.286e-06
I8357 0 n8358 2.976e-02A M=5.097e-07
I8358 0 n8359 2.976e-02A M=1.813e-06
I8359 0 n8360 2.976e-02A M=8.388e-07
I8360 0 n8361 2.976e-02A M=1.250e-06
I8361 0 n8362 2.976e-02A M=1.158e-06
I8362 0 n8363 2.976e-02A M=1.468e-06
I8363 0 n8364 2.976e-02A M=9.459e-07
I8364 0 n8365 2.976e-02A M=1.751e-06
I8365 0 n8366 2.976e-02A M=1.636e-06
I8366 0 n8367 2.976e-02A M=8.188e-07
I8367 0 n8368 2.976e-02A M=1.044e-06
I8368 0 n8369 2.976e-02A M=4.239e-07
I8369 0 n8370 2.976e-02A M=1.953e-06
I8370 0 n8371 2.976e-02A M=1.440e-06
I8371 0 n8372 2.976e-02A M=8.623e-07
I8372 0 n8373 2.976e-02A M=1.128e-06
I8373 0 n8374 2.976e-02A M=1.608e-06
I8374 0 n8375 2.976e-02A M=3.257e-07
I8375 0 n8376 2.976e-02A M=8.712e-07
I8376 0 n8377 2.976e-02A M=1.156e-07
I8377 0 n8378 2.976e-02A M=1.106e-06
I8378 0 n8379 2.976e-02A M=1.911e-06
I8379 0 n8380 2.976e-02A M=4.154e-07
I8380 0 n8381 2.976e-02A M=1.275e-06
I8381 0 n8382 2.976e-02A M=1.122e-06
I8382 0 n8383 2.976e-02A M=1.047e-06
I8383 0 n8384 2.976e-02A M=8.114e-07
I8384 0 n8385 2.976e-02A M=6.747e-07
I8385 0 n8386 2.976e-02A M=7.907e-07
I8386 0 n8387 2.976e-02A M=6.636e-07
I8387 0 n8388 2.976e-02A M=1.306e-06
I8388 0 n8389 2.976e-02A M=7.447e-07
I8389 0 n8390 2.976e-02A M=8.345e-07
I8390 0 n8391 2.976e-02A M=1.287e-06
I8391 0 n8392 2.976e-02A M=1.421e-06
I8392 0 n8393 2.976e-02A M=4.537e-07
I8393 0 n8394 2.976e-02A M=8.069e-07
I8394 0 n8395 2.976e-02A M=1.358e-06
I8395 0 n8396 2.976e-02A M=9.198e-07
I8396 0 n8397 2.976e-02A M=1.044e-06
I8397 0 n8398 2.976e-02A M=1.494e-06
I8398 0 n8399 2.976e-02A M=4.679e-07
I8399 0 n8400 2.976e-02A M=8.088e-07
I8400 0 n8401 2.976e-02A M=3.056e-07
I8401 0 n8402 2.976e-02A M=1.137e-06
I8402 0 n8403 2.976e-02A M=4.072e-07
I8403 0 n8404 2.976e-02A M=7.339e-07
I8404 0 n8405 2.976e-02A M=1.346e-06
I8405 0 n8406 2.976e-02A M=8.335e-07
I8406 0 n8407 2.976e-02A M=8.332e-07
I8407 0 n8408 2.976e-02A M=6.860e-07
I8408 0 n8409 2.976e-02A M=5.952e-07
I8409 0 n8410 2.976e-02A M=2.278e-06
I8410 0 n8411 2.976e-02A M=1.034e-06
I8411 0 n8412 2.976e-02A M=1.137e-06
I8412 0 n8413 2.976e-02A M=1.856e-06
I8413 0 n8414 2.976e-02A M=4.483e-07
I8414 0 n8415 2.976e-02A M=1.558e-06
I8415 0 n8416 2.976e-02A M=7.434e-07
I8416 0 n8417 2.976e-02A M=7.654e-07
I8417 0 n8418 2.976e-02A M=2.803e-07
I8418 0 n8419 2.976e-02A M=1.737e-06
I8419 0 n8420 2.976e-02A M=8.571e-07
I8420 0 n8421 2.976e-02A M=3.650e-07
I8421 0 n8422 2.976e-02A M=4.245e-07
I8422 0 n8423 2.976e-02A M=1.011e-06
I8423 0 n8424 2.976e-02A M=5.437e-07
I8424 0 n8425 2.976e-02A M=1.135e-06
I8425 0 n8426 2.976e-02A M=2.922e-07
I8426 0 n8427 2.976e-02A M=6.819e-07
I8427 0 n8428 2.976e-02A M=1.568e-06
I8428 0 n8429 2.976e-02A M=1.724e-06
I8429 0 n8430 2.976e-02A M=1.275e-06
I8430 0 n8431 2.976e-02A M=5.141e-07
I8431 0 n8432 2.976e-02A M=1.077e-06
I8432 0 n8433 2.976e-02A M=8.707e-07
I8433 0 n8434 2.976e-02A M=7.797e-07
I8434 0 n8435 2.976e-02A M=1.357e-06
I8435 0 n8436 2.976e-02A M=1.161e-06
I8436 0 n8437 2.976e-02A M=9.856e-07
I8437 0 n8438 2.976e-02A M=1.045e-06
I8438 0 n8439 2.976e-02A M=9.230e-07
I8439 0 n8440 2.976e-02A M=3.564e-07
I8440 0 n8441 2.976e-02A M=6.268e-07
I8441 0 n8442 2.976e-02A M=6.613e-07
I8442 0 n8443 2.976e-02A M=8.356e-07
I8443 0 n8444 2.976e-02A M=3.703e-06
I8444 0 n8445 2.976e-02A M=1.127e-06
I8445 0 n8446 2.976e-02A M=1.193e-06
I8446 0 n8447 2.976e-02A M=9.124e-07
I8447 0 n8448 2.976e-02A M=1.041e-06
I8448 0 n8449 2.976e-02A M=6.359e-07
I8449 0 n8450 2.976e-02A M=1.411e-06
I8450 0 n8451 2.976e-02A M=1.223e-06
I8451 0 n8452 2.976e-02A M=1.476e-06
I8452 0 n8453 2.976e-02A M=7.388e-07
I8453 0 n8454 2.976e-02A M=6.355e-07
I8454 0 n8455 2.976e-02A M=9.496e-07
I8455 0 n8456 2.976e-02A M=9.936e-07
I8456 0 n8457 2.976e-02A M=7.761e-07
I8457 0 n8458 2.976e-02A M=1.167e-06
I8458 0 n8459 2.976e-02A M=7.232e-07
I8459 0 n8460 2.976e-02A M=7.545e-07
I8460 0 n8461 2.976e-02A M=1.426e-06
I8461 0 n8462 2.976e-02A M=5.643e-07
I8462 0 n8463 2.976e-02A M=2.067e-06
I8463 0 n8464 2.976e-02A M=1.126e-06
I8464 0 n8465 2.976e-02A M=1.473e-06
I8465 0 n8466 2.976e-02A M=9.068e-07
I8466 0 n8467 2.976e-02A M=5.198e-07
I8467 0 n8468 2.976e-02A M=7.193e-07
I8468 0 n8469 2.976e-02A M=3.674e-07
I8469 0 n8470 2.976e-02A M=1.526e-06
I8470 0 n8471 2.976e-02A M=6.629e-07
I8471 0 n8472 2.976e-02A M=1.048e-06
I8472 0 n8473 2.976e-02A M=4.785e-07
I8473 0 n8474 2.976e-02A M=1.118e-06
I8474 0 n8475 2.976e-02A M=2.012e-06
I8475 0 n8476 2.976e-02A M=1.196e-06
I8476 0 n8477 2.976e-02A M=1.139e-06
I8477 0 n8478 2.976e-02A M=9.284e-07
I8478 0 n8479 2.976e-02A M=1.380e-06
I8479 0 n8480 2.976e-02A M=8.864e-07
I8480 0 n8481 2.976e-02A M=9.299e-07
I8481 0 n8482 2.976e-02A M=1.135e-06
I8482 0 n8483 2.976e-02A M=1.545e-06
I8483 0 n8484 2.976e-02A M=1.427e-06
I8484 0 n8485 2.976e-02A M=5.715e-07
I8485 0 n8486 2.976e-02A M=6.800e-07
I8486 0 n8487 2.976e-02A M=1.236e-06
I8487 0 n8488 2.976e-02A M=8.403e-07
I8488 0 n8489 2.976e-02A M=1.085e-06
I8489 0 n8490 2.976e-02A M=1.489e-06
I8490 0 n8491 2.976e-02A M=1.724e-06
I8491 0 n8492 2.976e-02A M=1.421e-06
I8492 0 n8493 2.976e-02A M=1.669e-06
I8493 0 n8494 2.976e-02A M=1.138e-06
I8494 0 n8495 2.976e-02A M=1.116e-06
I8495 0 n8496 2.976e-02A M=5.361e-07
I8496 0 n8497 2.976e-02A M=6.079e-07
I8497 0 n8498 2.976e-02A M=1.326e-06
I8498 0 n8499 2.976e-02A M=6.128e-07
I8499 0 n1 2.976e-02A M=3.641e-07
I8500 0 n8501 2.976e-02A M=6.395e-07
I8501 0 n8502 2.976e-02A M=1.210e-06
I8502 0 n8503 2.976e-02A M=1.207e-06
I8503 0 n8504 2.976e-02A M=5.439e-07
I8504 0 n8505 2.976e-02A M=1.924e-06
I8505 0 n8506 2.976e-02A M=1.474e-06
I8506 0 n8507 2.976e-02A M=1.262e-06
I8507 0 n8508 2.976e-02A M=4.675e-07
I8508 0 n8509 2.976e-02A M=1.409e-06
I8509 0 n8510 2.976e-02A M=7.203e-07
I8510 0 n8511 2.976e-02A M=4.354e-07
I8511 0 n8512 2.976e-02A M=1.179e-06
I8512 0 n8513 2.976e-02A M=3.753e-07
I8513 0 n8514 2.976e-02A M=8.431e-07
I8514 0 n8515 2.976e-02A M=7.982e-07
I8515 0 n8516 2.976e-02A M=2.148e-07
I8516 0 n8517 2.976e-02A M=7.741e-07
I8517 0 n8518 2.976e-02A M=5.689e-07
I8518 0 n8519 2.976e-02A M=4.964e-07
I8519 0 n8520 2.976e-02A M=7.436e-07
I8520 0 n8521 2.976e-02A M=1.890e-06
I8521 0 n8522 2.976e-02A M=1.400e-06
I8522 0 n8523 2.976e-02A M=5.859e-07
I8523 0 n8524 2.976e-02A M=1.062e-06
I8524 0 n8525 2.976e-02A M=1.300e-06
I8525 0 n8526 2.976e-02A M=1.558e-06
I8526 0 n8527 2.976e-02A M=1.355e-06
I8527 0 n8528 2.976e-02A M=1.621e-06
I8528 0 n8529 2.976e-02A M=1.741e-06
I8529 0 n8530 2.976e-02A M=7.159e-07
I8530 0 n8531 2.976e-02A M=6.573e-07
I8531 0 n8532 2.976e-02A M=9.314e-07
I8532 0 n8533 2.976e-02A M=6.240e-07
I8533 0 n8534 2.976e-02A M=1.377e-06
I8534 0 n8535 2.976e-02A M=1.628e-06
I8535 0 n8536 2.976e-02A M=9.093e-07
I8536 0 n8537 2.976e-02A M=2.763e-06
I8537 0 n8538 2.976e-02A M=9.538e-07
I8538 0 n8539 2.976e-02A M=1.412e-06
I8539 0 n8540 2.976e-02A M=3.315e-07
I8540 0 n8541 2.976e-02A M=5.841e-07
I8541 0 n8542 2.976e-02A M=1.327e-06
I8542 0 n8543 2.976e-02A M=1.243e-06
I8543 0 n8544 2.976e-02A M=1.109e-06
I8544 0 n8545 2.976e-02A M=1.447e-06
I8545 0 n8546 2.976e-02A M=3.683e-07
I8546 0 n8547 2.976e-02A M=2.888e-07
I8547 0 n8548 2.976e-02A M=8.267e-07
I8548 0 n8549 2.976e-02A M=4.284e-07
I8549 0 n8550 2.976e-02A M=2.490e-06
I8550 0 n8551 2.976e-02A M=6.979e-07
I8551 0 n8552 2.976e-02A M=4.526e-07
I8552 0 n8553 2.976e-02A M=1.427e-06
I8553 0 n8554 2.976e-02A M=6.424e-07
I8554 0 n1 2.976e-02A M=7.927e-07
I8555 0 n8556 2.976e-02A M=9.533e-07
I8556 0 n8557 2.976e-02A M=7.741e-07
I8557 0 n8558 2.976e-02A M=1.224e-06
I8558 0 n8559 2.976e-02A M=2.445e-06
I8559 0 n8560 2.976e-02A M=7.838e-07
I8560 0 n8561 2.976e-02A M=1.003e-06
I8561 0 n8562 2.976e-02A M=1.295e-06
I8562 0 n8563 2.976e-02A M=9.073e-07
I8563 0 n8564 2.976e-02A M=2.132e-06
I8564 0 n8565 2.976e-02A M=9.938e-07
I8565 0 n8566 2.976e-02A M=7.318e-07
I8566 0 n8567 2.976e-02A M=1.371e-06
I8567 0 n8568 2.976e-02A M=1.118e-06
I8568 0 n8569 2.976e-02A M=1.597e-06
I8569 0 n8570 2.976e-02A M=7.243e-07
I8570 0 n8571 2.976e-02A M=5.995e-07
I8571 0 n8572 2.976e-02A M=1.154e-06
I8572 0 n8573 2.976e-02A M=6.540e-07
I8573 0 n8574 2.976e-02A M=1.812e-06
I8574 0 n8575 2.976e-02A M=6.273e-07
I8575 0 n8576 2.976e-02A M=8.487e-07
I8576 0 n8577 2.976e-02A M=6.084e-07
I8577 0 n8578 2.976e-02A M=1.972e-06
I8578 0 n8579 2.976e-02A M=5.680e-07
I8579 0 n8580 2.976e-02A M=7.897e-07
I8580 0 n8581 2.976e-02A M=6.079e-07
I8581 0 n8582 2.976e-02A M=7.741e-07
I8582 0 n8583 2.976e-02A M=1.343e-06
I8583 0 n8584 2.976e-02A M=6.097e-07
I8584 0 n8585 2.976e-02A M=8.297e-07
I8585 0 n8586 2.976e-02A M=5.502e-07
I8586 0 n8587 2.976e-02A M=9.626e-07
I8587 0 n8588 2.976e-02A M=1.600e-06
I8588 0 n8589 2.976e-02A M=4.946e-07
I8589 0 n8590 2.976e-02A M=2.626e-07
I8590 0 n8591 2.976e-02A M=6.820e-07
I8591 0 n8592 2.976e-02A M=1.949e-06
I8592 0 n8593 2.976e-02A M=3.029e-07
I8593 0 n8594 2.976e-02A M=1.966e-06
I8594 0 n8595 2.976e-02A M=4.270e-07
I8595 0 n8596 2.976e-02A M=1.104e-06
I8596 0 n8597 2.976e-02A M=2.187e-07
I8597 0 n8598 2.976e-02A M=3.899e-07
I8598 0 n8599 2.976e-02A M=2.384e-06
I8599 0 n8600 2.976e-02A M=7.257e-07
I8600 0 n8601 2.976e-02A M=4.163e-07
I8601 0 n8602 2.976e-02A M=4.046e-07
I8602 0 n1 2.976e-02A M=1.378e-06
I8603 0 n8604 2.976e-02A M=7.068e-07
I8604 0 n8605 2.976e-02A M=8.184e-07
I8605 0 n8606 2.976e-02A M=1.381e-06
I8606 0 n8607 2.976e-02A M=1.388e-06
I8607 0 n8608 2.976e-02A M=6.637e-07
I8608 0 n8609 2.976e-02A M=2.686e-07
I8609 0 n8610 2.976e-02A M=1.634e-06
I8610 0 n8611 2.976e-02A M=1.245e-06
I8611 0 n8612 2.976e-02A M=6.811e-07
I8612 0 n8613 2.976e-02A M=9.537e-07
I8613 0 n8614 2.976e-02A M=3.403e-07
I8614 0 n8615 2.976e-02A M=9.037e-07
I8615 0 n8616 2.976e-02A M=8.665e-07
I8616 0 n8617 2.976e-02A M=7.988e-07
I8617 0 n8618 2.976e-02A M=5.663e-07
I8618 0 n8619 2.976e-02A M=1.240e-06
I8619 0 n8620 2.976e-02A M=2.017e-06
I8620 0 n8621 2.976e-02A M=1.224e-06
I8621 0 n8622 2.976e-02A M=1.047e-06
I8622 0 n8623 2.976e-02A M=8.764e-07
I8623 0 n8624 2.976e-02A M=1.901e-06
I8624 0 n8625 2.976e-02A M=1.940e-07
I8625 0 n8626 2.976e-02A M=4.094e-07
I8626 0 n8627 2.976e-02A M=9.609e-07
I8627 0 n8628 2.976e-02A M=1.360e-06
I8628 0 n8629 2.976e-02A M=1.043e-06
I8629 0 n8630 2.976e-02A M=1.561e-06
I8630 0 n8631 2.976e-02A M=8.270e-07
I8631 0 n8632 2.976e-02A M=1.492e-06
I8632 0 n8633 2.976e-02A M=9.758e-07
I8633 0 n8634 2.976e-02A M=5.700e-07
I8634 0 n8635 2.976e-02A M=7.943e-07
I8635 0 n8636 2.976e-02A M=7.884e-08
I8636 0 n8637 2.976e-02A M=8.708e-07
I8637 0 n8638 2.976e-02A M=1.231e-06
I8638 0 n8639 2.976e-02A M=5.934e-07
I8639 0 n8640 2.976e-02A M=8.490e-07
I8640 0 n8641 2.976e-02A M=5.933e-07
I8641 0 n8642 2.976e-02A M=1.299e-06
I8642 0 n8643 2.976e-02A M=4.241e-07
I8643 0 n8644 2.976e-02A M=7.564e-07
I8644 0 n8645 2.976e-02A M=1.169e-06
I8645 0 n8646 2.976e-02A M=1.258e-06
I8646 0 n8647 2.976e-02A M=1.027e-06
I8647 0 n8648 2.976e-02A M=6.677e-07
I8648 0 n8649 2.976e-02A M=2.551e-06
I8649 0 n8650 2.976e-02A M=1.090e-06
I8650 0 n8651 2.976e-02A M=7.045e-07
I8651 0 n8652 2.976e-02A M=1.018e-06
I8652 0 n8653 2.976e-02A M=1.529e-06
I8653 0 n8654 2.976e-02A M=9.381e-07
I8654 0 n8655 2.976e-02A M=2.773e-06
I8655 0 n8656 2.976e-02A M=1.484e-06
I8656 0 n8657 2.976e-02A M=1.414e-06
I8657 0 n8658 2.976e-02A M=8.773e-07
I8658 0 n8659 2.976e-02A M=4.288e-07
I8659 0 n8660 2.976e-02A M=2.052e-06
I8660 0 n8661 2.976e-02A M=1.040e-06
I8661 0 n8662 2.976e-02A M=2.408e-06
I8662 0 n8663 2.976e-02A M=1.295e-06
I8663 0 n8664 2.976e-02A M=7.860e-07
I8664 0 n8665 2.976e-02A M=1.703e-06
I8665 0 n8666 2.976e-02A M=9.438e-07
I8666 0 n8667 2.976e-02A M=2.915e-07
I8667 0 n8668 2.976e-02A M=2.466e-07
I8668 0 n8669 2.976e-02A M=8.897e-07
I8669 0 n8670 2.976e-02A M=1.644e-06
I8670 0 n8671 2.976e-02A M=1.426e-06
I8671 0 n8672 2.976e-02A M=9.967e-07
I8672 0 n8673 2.976e-02A M=1.155e-06
I8673 0 n8674 2.976e-02A M=1.001e-06
I8674 0 n8675 2.976e-02A M=1.053e-06
I8675 0 n8676 2.976e-02A M=8.792e-07
I8676 0 n8677 2.976e-02A M=6.576e-07
I8677 0 n8678 2.976e-02A M=9.566e-07
I8678 0 n8679 2.976e-02A M=1.663e-06
I8679 0 n1 2.976e-02A M=2.254e-06
I8680 0 n8681 2.976e-02A M=8.748e-07
I8681 0 n8682 2.976e-02A M=8.824e-07
I8682 0 n8683 2.976e-02A M=7.074e-07
I8683 0 n8684 2.976e-02A M=7.425e-07
I8684 0 n8685 2.976e-02A M=5.064e-07
I8685 0 n8686 2.976e-02A M=1.142e-06
I8686 0 n8687 2.976e-02A M=1.146e-06
I8687 0 n8688 2.976e-02A M=1.314e-06
I8688 0 n8689 2.976e-02A M=1.044e-06
I8689 0 n8690 2.976e-02A M=1.066e-06
I8690 0 n8691 2.976e-02A M=1.749e-06
I8691 0 n8692 2.976e-02A M=1.113e-06
I8692 0 n8693 2.976e-02A M=1.107e-06
I8693 0 n8694 2.976e-02A M=1.530e-06
I8694 0 n8695 2.976e-02A M=1.775e-07
I8695 0 n8696 2.976e-02A M=2.835e-06
I8696 0 n8697 2.976e-02A M=8.172e-07
I8697 0 n8698 2.976e-02A M=1.166e-06
I8698 0 n8699 2.976e-02A M=2.946e-06
I8699 0 n8700 2.976e-02A M=7.459e-07
I8700 0 n8701 2.976e-02A M=1.400e-06
I8701 0 n8702 2.976e-02A M=6.136e-07
I8702 0 n8703 2.976e-02A M=7.112e-07
I8703 0 n8704 2.976e-02A M=6.242e-07
I8704 0 n8705 2.976e-02A M=7.956e-07
I8705 0 n8706 2.976e-02A M=9.065e-07
I8706 0 n8707 2.976e-02A M=4.139e-07
I8707 0 n8708 2.976e-02A M=5.939e-07
I8708 0 n8709 2.976e-02A M=8.796e-07
I8709 0 n8710 2.976e-02A M=1.204e-06
I8710 0 n8711 2.976e-02A M=9.914e-07
I8711 0 n8712 2.976e-02A M=2.595e-06
I8712 0 n8713 2.976e-02A M=1.097e-06
I8713 0 n8714 2.976e-02A M=3.618e-07
I8714 0 n8715 2.976e-02A M=1.793e-06
I8715 0 n8716 2.976e-02A M=6.386e-07
I8716 0 n8717 2.976e-02A M=7.106e-07
I8717 0 n8718 2.976e-02A M=8.367e-07
I8718 0 n8719 2.976e-02A M=1.308e-06
I8719 0 n8720 2.976e-02A M=1.298e-06
I8720 0 n8721 2.976e-02A M=5.374e-07
I8721 0 n8722 2.976e-02A M=1.865e-06
I8722 0 n8723 2.976e-02A M=1.905e-06
I8723 0 n8724 2.976e-02A M=3.030e-06
I8724 0 n8725 2.976e-02A M=2.144e-06
I8725 0 n8726 2.976e-02A M=1.296e-06
I8726 0 n8727 2.976e-02A M=1.058e-06
I8727 0 n8728 2.976e-02A M=1.029e-06
I8728 0 n8729 2.976e-02A M=9.098e-07
I8729 0 n8730 2.976e-02A M=1.297e-06
I8730 0 n8731 2.976e-02A M=1.393e-06
I8731 0 n8732 2.976e-02A M=1.123e-06
I8732 0 n8733 2.976e-02A M=1.685e-07
I8733 0 n8734 2.976e-02A M=1.893e-06
I8734 0 n8735 2.976e-02A M=2.523e-07
I8735 0 n8736 2.976e-02A M=1.577e-06
I8736 0 n8737 2.976e-02A M=7.469e-07
I8737 0 n8738 2.976e-02A M=1.050e-06
I8738 0 n8739 2.976e-02A M=8.956e-07
I8739 0 n8740 2.976e-02A M=3.008e-07
I8740 0 n8741 2.976e-02A M=5.832e-07
I8741 0 n8742 2.976e-02A M=1.272e-06
I8742 0 n8743 2.976e-02A M=6.180e-07
I8743 0 n8744 2.976e-02A M=1.147e-06
I8744 0 n8745 2.976e-02A M=9.276e-07
I8745 0 n8746 2.976e-02A M=4.592e-07
I8746 0 n8747 2.976e-02A M=1.356e-06
I8747 0 n8748 2.976e-02A M=7.304e-07
I8748 0 n8749 2.976e-02A M=1.742e-06
I8749 0 n8750 2.976e-02A M=2.045e-06
I8750 0 n8751 2.976e-02A M=1.287e-06
I8751 0 n8752 2.976e-02A M=7.048e-07
I8752 0 n8753 2.976e-02A M=7.723e-07
I8753 0 n8754 2.976e-02A M=7.600e-07
I8754 0 n8755 2.976e-02A M=8.372e-07
I8755 0 n8756 2.976e-02A M=8.985e-07
I8756 0 n8757 2.976e-02A M=1.078e-06
I8757 0 n8758 2.976e-02A M=1.126e-06
I8758 0 n8759 2.976e-02A M=1.260e-06
I8759 0 n8760 2.976e-02A M=1.015e-06
I8760 0 n8761 2.976e-02A M=3.491e-07
I8761 0 n8762 2.976e-02A M=1.001e-06
I8762 0 n8763 2.976e-02A M=4.964e-07
I8763 0 n8764 2.976e-02A M=8.046e-07
I8764 0 n8765 2.976e-02A M=6.222e-07
I8765 0 n8766 2.976e-02A M=1.321e-06
I8766 0 n8767 2.976e-02A M=6.594e-07
I8767 0 n8768 2.976e-02A M=1.457e-06
I8768 0 n8769 2.976e-02A M=7.518e-07
I8769 0 n8770 2.976e-02A M=2.084e-07
I8770 0 n8771 2.976e-02A M=4.180e-07
I8771 0 n8772 2.976e-02A M=6.294e-07
I8772 0 n8773 2.976e-02A M=1.768e-06
I8773 0 n8774 2.976e-02A M=3.343e-07
I8774 0 n8775 2.976e-02A M=1.187e-06
I8775 0 n8776 2.976e-02A M=9.757e-07
I8776 0 n8777 2.976e-02A M=4.021e-07
I8777 0 n8778 2.976e-02A M=1.347e-06
I8778 0 n8779 2.976e-02A M=8.157e-07
I8779 0 n8780 2.976e-02A M=1.726e-06
I8780 0 n8781 2.976e-02A M=1.729e-06
I8781 0 n8782 2.976e-02A M=8.279e-07
I8782 0 n8783 2.976e-02A M=1.303e-06
I8783 0 n8784 2.976e-02A M=8.220e-07
I8784 0 n8785 2.976e-02A M=5.080e-07
I8785 0 n8786 2.976e-02A M=8.189e-07
I8786 0 n8787 2.976e-02A M=6.051e-07
I8787 0 n8788 2.976e-02A M=1.453e-06
I8788 0 n8789 2.976e-02A M=3.933e-07
I8789 0 n8790 2.976e-02A M=1.373e-06
I8790 0 n8791 2.976e-02A M=8.576e-07
I8791 0 n8792 2.976e-02A M=9.655e-07
I8792 0 n8793 2.976e-02A M=1.121e-06
I8793 0 n8794 2.976e-02A M=3.740e-07
I8794 0 n8795 2.976e-02A M=1.114e-06
I8795 0 n8796 2.976e-02A M=5.100e-07
I8796 0 n8797 2.976e-02A M=1.358e-06
I8797 0 n8798 2.976e-02A M=1.571e-06
I8798 0 n8799 2.976e-02A M=1.028e-06
I8799 0 n8800 2.976e-02A M=7.581e-07
I8800 0 n8801 2.976e-02A M=2.774e-06
I8801 0 n8802 2.976e-02A M=7.150e-07
I8802 0 n8803 2.976e-02A M=1.169e-06
I8803 0 n8804 2.976e-02A M=7.196e-07
I8804 0 n8805 2.976e-02A M=1.451e-06
I8805 0 n8806 2.976e-02A M=8.751e-07
I8806 0 n8807 2.976e-02A M=5.427e-07
I8807 0 n8808 2.976e-02A M=2.700e-07
I8808 0 n8809 2.976e-02A M=9.725e-07
I8809 0 n8810 2.976e-02A M=5.221e-07
I8810 0 n8811 2.976e-02A M=8.544e-07
I8811 0 n8812 2.976e-02A M=1.059e-06
I8812 0 n8813 2.976e-02A M=3.483e-07
I8813 0 n8814 2.976e-02A M=1.912e-06
I8814 0 n8815 2.976e-02A M=1.176e-06
I8815 0 n8816 2.976e-02A M=1.467e-06
I8816 0 n8817 2.976e-02A M=4.763e-07
I8817 0 n8818 2.976e-02A M=8.863e-07
I8818 0 n8819 2.976e-02A M=4.045e-07
I8819 0 n8820 2.976e-02A M=8.199e-07
I8820 0 n8821 2.976e-02A M=1.361e-06
I8821 0 n8822 2.976e-02A M=8.228e-07
I8822 0 n8823 2.976e-02A M=3.655e-07
I8823 0 n8824 2.976e-02A M=1.777e-06
I8824 0 n8825 2.976e-02A M=3.124e-07
I8825 0 n8826 2.976e-02A M=8.386e-07
I8826 0 n8827 2.976e-02A M=5.746e-07
I8827 0 n8828 2.976e-02A M=8.156e-07
I8828 0 n8829 2.976e-02A M=9.755e-07
I8829 0 n8830 2.976e-02A M=6.554e-07
I8830 0 n8831 2.976e-02A M=5.330e-07
I8831 0 n8832 2.976e-02A M=1.615e-06
I8832 0 n8833 2.976e-02A M=1.087e-06
I8833 0 n8834 2.976e-02A M=3.380e-07
I8834 0 n8835 2.976e-02A M=8.059e-07
I8835 0 n8836 2.976e-02A M=7.331e-07
I8836 0 n8837 2.976e-02A M=9.147e-07
I8837 0 n8838 2.976e-02A M=1.473e-06
I8838 0 n8839 2.976e-02A M=1.223e-06
I8839 0 n8840 2.976e-02A M=1.774e-06
I8840 0 n8841 2.976e-02A M=5.318e-07
I8841 0 n8842 2.976e-02A M=9.419e-07
I8842 0 n1 2.976e-02A M=1.409e-06
I8843 0 n8844 2.976e-02A M=1.585e-06
I8844 0 n8845 2.976e-02A M=9.685e-07
I8845 0 n8846 2.976e-02A M=9.943e-07
I8846 0 n8847 2.976e-02A M=9.164e-07
I8847 0 n8848 2.976e-02A M=5.550e-07
I8848 0 n8849 2.976e-02A M=1.298e-06
I8849 0 n8850 2.976e-02A M=1.351e-06
I8850 0 n8851 2.976e-02A M=7.609e-07
I8851 0 n8852 2.976e-02A M=1.249e-06
I8852 0 n8853 2.976e-02A M=1.083e-06
I8853 0 n8854 2.976e-02A M=1.021e-06
I8854 0 n8855 2.976e-02A M=1.521e-06
I8855 0 n8856 2.976e-02A M=7.684e-07
I8856 0 n8857 2.976e-02A M=8.424e-07
I8857 0 n8858 2.976e-02A M=1.623e-06
I8858 0 n8859 2.976e-02A M=1.616e-06
I8859 0 n8860 2.976e-02A M=9.313e-07
I8860 0 n8861 2.976e-02A M=5.559e-07
I8861 0 n8862 2.976e-02A M=9.609e-07
I8862 0 n8863 2.976e-02A M=1.257e-06
I8863 0 n8864 2.976e-02A M=2.931e-07
I8864 0 n8865 2.976e-02A M=1.501e-06
I8865 0 n8866 2.976e-02A M=8.047e-07
I8866 0 n8867 2.976e-02A M=1.412e-06
I8867 0 n8868 2.976e-02A M=1.268e-06
I8868 0 n8869 2.976e-02A M=1.230e-06
I8869 0 n8870 2.976e-02A M=1.241e-06
I8870 0 n8871 2.976e-02A M=6.378e-07
I8871 0 n8872 2.976e-02A M=1.112e-06
I8872 0 n8873 2.976e-02A M=1.221e-07
I8873 0 n8874 2.976e-02A M=1.165e-07
I8874 0 n8875 2.976e-02A M=7.613e-07
I8875 0 n8876 2.976e-02A M=8.237e-07
I8876 0 n8877 2.976e-02A M=8.698e-07
I8877 0 n8878 2.976e-02A M=9.569e-07
I8878 0 n8879 2.976e-02A M=4.140e-07
I8879 0 n8880 2.976e-02A M=8.338e-07
I8880 0 n8881 2.976e-02A M=1.003e-06
I8881 0 n8882 2.976e-02A M=1.025e-06
I8882 0 n8883 2.976e-02A M=8.868e-07
I8883 0 n8884 2.976e-02A M=2.821e-06
I8884 0 n8885 2.976e-02A M=3.296e-07
I8885 0 n8886 2.976e-02A M=1.504e-06
I8886 0 n8887 2.976e-02A M=5.538e-07
I8887 0 n8888 2.976e-02A M=6.406e-07
I8888 0 n8889 2.976e-02A M=5.921e-07
I8889 0 n8890 2.976e-02A M=2.608e-07
I8890 0 n8891 2.976e-02A M=1.761e-06
I8891 0 n8892 2.976e-02A M=6.937e-07
I8892 0 n8893 2.976e-02A M=8.129e-07
I8893 0 n8894 2.976e-02A M=7.372e-07
I8894 0 n8895 2.976e-02A M=5.805e-07
I8895 0 n8896 2.976e-02A M=1.670e-06
I8896 0 n8897 2.976e-02A M=6.345e-07
I8897 0 n8898 2.976e-02A M=2.142e-06
I8898 0 n8899 2.976e-02A M=9.214e-07
I8899 0 n8900 2.976e-02A M=1.203e-06
I8900 0 n8901 2.976e-02A M=1.260e-06
I8901 0 n8902 2.976e-02A M=9.908e-07
I8902 0 n8903 2.976e-02A M=2.469e-06
I8903 0 n8904 2.976e-02A M=9.955e-07
I8904 0 n8905 2.976e-02A M=6.653e-07
I8905 0 n8906 2.976e-02A M=6.382e-07
I8906 0 n8907 2.976e-02A M=8.489e-07
I8907 0 n8908 2.976e-02A M=1.120e-06
I8908 0 n8909 2.976e-02A M=1.202e-06
I8909 0 n8910 2.976e-02A M=1.033e-06
I8910 0 n8911 2.976e-02A M=9.804e-07
I8911 0 n8912 2.976e-02A M=1.646e-06
I8912 0 n8913 2.976e-02A M=2.431e-06
I8913 0 n8914 2.976e-02A M=1.145e-06
I8914 0 n8915 2.976e-02A M=1.019e-06
I8915 0 n8916 2.976e-02A M=4.440e-07
I8916 0 n8917 2.976e-02A M=9.123e-07
I8917 0 n8918 2.976e-02A M=4.410e-07
I8918 0 n8919 2.976e-02A M=1.759e-06
I8919 0 n8920 2.976e-02A M=6.015e-07
I8920 0 n8921 2.976e-02A M=1.571e-06
I8921 0 n8922 2.976e-02A M=8.554e-07
I8922 0 n8923 2.976e-02A M=7.187e-07
I8923 0 n8924 2.976e-02A M=8.595e-07
I8924 0 n8925 2.976e-02A M=6.887e-07
I8925 0 n1 2.976e-02A M=1.243e-06
I8926 0 n8927 2.976e-02A M=8.942e-07
I8927 0 n8928 2.976e-02A M=1.125e-06
I8928 0 n8929 2.976e-02A M=1.430e-06
I8929 0 n8930 2.976e-02A M=1.490e-06
I8930 0 n8931 2.976e-02A M=2.069e-06
I8931 0 n8932 2.976e-02A M=2.034e-06
I8932 0 n8933 2.976e-02A M=9.720e-07
I8933 0 n8934 2.976e-02A M=1.112e-06
I8934 0 n8935 2.976e-02A M=6.576e-07
I8935 0 n8936 2.976e-02A M=4.585e-07
I8936 0 n8937 2.976e-02A M=9.042e-07
I8937 0 n8938 2.976e-02A M=1.346e-06
I8938 0 n8939 2.976e-02A M=1.410e-06
I8939 0 n8940 2.976e-02A M=9.564e-07
I8940 0 n8941 2.976e-02A M=1.448e-06
I8941 0 n8942 2.976e-02A M=3.437e-07
I8942 0 n8943 2.976e-02A M=2.215e-06
I8943 0 n8944 2.976e-02A M=5.784e-07
I8944 0 n8945 2.976e-02A M=1.235e-06
I8945 0 n8946 2.976e-02A M=1.954e-06
I8946 0 n8947 2.976e-02A M=9.974e-07
I8947 0 n8948 2.976e-02A M=1.268e-06
I8948 0 n8949 2.976e-02A M=9.905e-07
I8949 0 n8950 2.976e-02A M=7.282e-07
I8950 0 n8951 2.976e-02A M=1.223e-06
I8951 0 n8952 2.976e-02A M=5.635e-07
I8952 0 n8953 2.976e-02A M=7.921e-07
I8953 0 n8954 2.976e-02A M=4.451e-07
I8954 0 n8955 2.976e-02A M=1.970e-06
I8955 0 n8956 2.976e-02A M=4.373e-07
I8956 0 n8957 2.976e-02A M=2.754e-07
I8957 0 n8958 2.976e-02A M=9.027e-07
I8958 0 n8959 2.976e-02A M=2.252e-07
I8959 0 n8960 2.976e-02A M=3.282e-06
I8960 0 n8961 2.976e-02A M=1.438e-06
I8961 0 n8962 2.976e-02A M=5.836e-07
I8962 0 n8963 2.976e-02A M=1.643e-06
I8963 0 n8964 2.976e-02A M=2.665e-06
I8964 0 n8965 2.976e-02A M=3.931e-07
I8965 0 n8966 2.976e-02A M=5.072e-07
I8966 0 n8967 2.976e-02A M=1.463e-06
I8967 0 n8968 2.976e-02A M=1.781e-06
I8968 0 n8969 2.976e-02A M=2.032e-06
I8969 0 n8970 2.976e-02A M=5.819e-07
I8970 0 n8971 2.976e-02A M=6.728e-07
I8971 0 n8972 2.976e-02A M=7.511e-07
I8972 0 n8973 2.976e-02A M=4.492e-07
I8973 0 n8974 2.976e-02A M=1.374e-06
I8974 0 n8975 2.976e-02A M=8.079e-07
I8975 0 n8976 2.976e-02A M=5.310e-07
I8976 0 n8977 2.976e-02A M=7.747e-07
I8977 0 n8978 2.976e-02A M=9.098e-07
I8978 0 n8979 2.976e-02A M=1.647e-06
I8979 0 n8980 2.976e-02A M=6.084e-07
I8980 0 n8981 2.976e-02A M=1.896e-06
I8981 0 n8982 2.976e-02A M=5.815e-07
I8982 0 n8983 2.976e-02A M=5.442e-07
I8983 0 n8984 2.976e-02A M=1.176e-06
I8984 0 n8985 2.976e-02A M=6.935e-07
I8985 0 n8986 2.976e-02A M=1.065e-06
I8986 0 n8987 2.976e-02A M=9.514e-07
I8987 0 n8988 2.976e-02A M=1.381e-06
I8988 0 n8989 2.976e-02A M=3.901e-07
I8989 0 n8990 2.976e-02A M=9.942e-07
I8990 0 n8991 2.976e-02A M=9.665e-07
I8991 0 n8992 2.976e-02A M=1.258e-06
I8992 0 n8993 2.976e-02A M=7.123e-07
I8993 0 n8994 2.976e-02A M=5.796e-07
I8994 0 n8995 2.976e-02A M=1.145e-06
I8995 0 n8996 2.976e-02A M=6.296e-07
I8996 0 n8997 2.976e-02A M=1.764e-06
I8997 0 n8998 2.976e-02A M=1.057e-06
I8998 0 n8999 2.976e-02A M=6.413e-07
I8999 0 n9000 2.976e-02A M=6.026e-07
I9000 0 n9001 2.976e-02A M=8.239e-07
I9001 0 n9002 2.976e-02A M=1.866e-06
I9002 0 n9003 2.976e-02A M=7.406e-07
I9003 0 n9004 2.976e-02A M=1.187e-06
I9004 0 n9005 2.976e-02A M=1.085e-06
I9005 0 n9006 2.976e-02A M=7.505e-07
I9006 0 n9007 2.976e-02A M=1.995e-06
I9007 0 n9008 2.976e-02A M=9.828e-07
I9008 0 n9009 2.976e-02A M=9.845e-07
I9009 0 n9010 2.976e-02A M=7.399e-07
I9010 0 n9011 2.976e-02A M=8.087e-07
I9011 0 n9012 2.976e-02A M=1.320e-06
I9012 0 n9013 2.976e-02A M=2.064e-06
I9013 0 n9014 2.976e-02A M=1.222e-06
I9014 0 n9015 2.976e-02A M=2.237e-07
I9015 0 n9016 2.976e-02A M=7.645e-07
I9016 0 n9017 2.976e-02A M=7.945e-07
I9017 0 n9018 2.976e-02A M=2.052e-06
I9018 0 n9019 2.976e-02A M=1.054e-06
I9019 0 n9020 2.976e-02A M=7.870e-07
I9020 0 n9021 2.976e-02A M=1.008e-06
I9021 0 n9022 2.976e-02A M=6.151e-07
I9022 0 n9023 2.976e-02A M=1.905e-06
I9023 0 n9024 2.976e-02A M=4.870e-07
I9024 0 n9025 2.976e-02A M=4.918e-07
I9025 0 n9026 2.976e-02A M=1.302e-06
I9026 0 n9027 2.976e-02A M=6.473e-07
I9027 0 n9028 2.976e-02A M=5.801e-07
I9028 0 n9029 2.976e-02A M=1.006e-06
I9029 0 n9030 2.976e-02A M=1.042e-06
I9030 0 n9031 2.976e-02A M=1.081e-06
I9031 0 n9032 2.976e-02A M=1.764e-06
I9032 0 n9033 2.976e-02A M=2.372e-06
I9033 0 n9034 2.976e-02A M=2.778e-06
I9034 0 n9035 2.976e-02A M=1.824e-06
I9035 0 n9036 2.976e-02A M=1.092e-06
I9036 0 n9037 2.976e-02A M=1.497e-06
I9037 0 n9038 2.976e-02A M=5.802e-07
I9038 0 n9039 2.976e-02A M=8.344e-07
I9039 0 n9040 2.976e-02A M=1.086e-06
I9040 0 n9041 2.976e-02A M=4.746e-07
I9041 0 n9042 2.976e-02A M=1.090e-06
I9042 0 n9043 2.976e-02A M=1.050e-06
I9043 0 n9044 2.976e-02A M=1.191e-06
I9044 0 n9045 2.976e-02A M=1.840e-06
I9045 0 n9046 2.976e-02A M=1.210e-06
I9046 0 n9047 2.976e-02A M=7.141e-07
I9047 0 n9048 2.976e-02A M=3.731e-07
I9048 0 n9049 2.976e-02A M=1.156e-06
I9049 0 n9050 2.976e-02A M=6.473e-07
I9050 0 n9051 2.976e-02A M=1.389e-06
I9051 0 n9052 2.976e-02A M=8.005e-07
I9052 0 n9053 2.976e-02A M=6.064e-07
I9053 0 n9054 2.976e-02A M=9.150e-07
I9054 0 n9055 2.976e-02A M=9.920e-07
I9055 0 n9056 2.976e-02A M=2.222e-06
I9056 0 n9057 2.976e-02A M=1.598e-06
I9057 0 n9058 2.976e-02A M=2.153e-06
I9058 0 n9059 2.976e-02A M=1.173e-06
I9059 0 n9060 2.976e-02A M=1.144e-06
I9060 0 n9061 2.976e-02A M=8.236e-07
I9061 0 n9062 2.976e-02A M=9.046e-07
I9062 0 n9063 2.976e-02A M=1.055e-06
I9063 0 n9064 2.976e-02A M=9.348e-07
I9064 0 n9065 2.976e-02A M=1.640e-06
I9065 0 n9066 2.976e-02A M=5.204e-07
I9066 0 n9067 2.976e-02A M=1.033e-06
I9067 0 n9068 2.976e-02A M=1.016e-06
I9068 0 n9069 2.976e-02A M=4.885e-07
I9069 0 n9070 2.976e-02A M=9.719e-07
I9070 0 n9071 2.976e-02A M=9.486e-07
I9071 0 n9072 2.976e-02A M=1.875e-07
I9072 0 n9073 2.976e-02A M=7.134e-07
I9073 0 n9074 2.976e-02A M=8.170e-07
I9074 0 n9075 2.976e-02A M=6.665e-07
I9075 0 n9076 2.976e-02A M=5.630e-07
I9076 0 n9077 2.976e-02A M=9.007e-07
I9077 0 n9078 2.976e-02A M=7.448e-07
I9078 0 n9079 2.976e-02A M=1.035e-06
I9079 0 n9080 2.976e-02A M=1.763e-06
I9080 0 n9081 2.976e-02A M=1.173e-06
I9081 0 n1 2.976e-02A M=9.370e-07
I9082 0 n9083 2.976e-02A M=6.217e-07
I9083 0 n9084 2.976e-02A M=4.770e-07
I9084 0 n9085 2.976e-02A M=1.312e-06
I9085 0 n9086 2.976e-02A M=7.326e-07
I9086 0 n9087 2.976e-02A M=7.066e-07
I9087 0 n9088 2.976e-02A M=1.615e-06
I9088 0 n9089 2.976e-02A M=1.514e-06
I9089 0 n9090 2.976e-02A M=9.708e-07
I9090 0 n9091 2.976e-02A M=5.126e-07
I9091 0 n9092 2.976e-02A M=4.423e-07
I9092 0 n9093 2.976e-02A M=7.587e-07
I9093 0 n9094 2.976e-02A M=1.859e-06
I9094 0 n9095 2.976e-02A M=1.779e-07
I9095 0 n9096 2.976e-02A M=7.933e-07
I9096 0 n9097 2.976e-02A M=8.364e-07
I9097 0 n9098 2.976e-02A M=9.857e-07
I9098 0 n9099 2.976e-02A M=1.232e-06
I9099 0 n9100 2.976e-02A M=1.204e-06
I9100 0 n9101 2.976e-02A M=2.840e-06
I9101 0 n9102 2.976e-02A M=5.841e-07
I9102 0 n9103 2.976e-02A M=2.478e-06
I9103 0 n9104 2.976e-02A M=4.680e-07
I9104 0 n9105 2.976e-02A M=2.315e-06
I9105 0 n9106 2.976e-02A M=1.483e-06
I9106 0 n9107 2.976e-02A M=1.380e-06
I9107 0 n9108 2.976e-02A M=1.184e-06
I9108 0 n9109 2.976e-02A M=1.093e-06
I9109 0 n9110 2.976e-02A M=1.111e-06
I9110 0 n9111 2.976e-02A M=6.597e-07
I9111 0 n9112 2.976e-02A M=2.559e-07
I9112 0 n9113 2.976e-02A M=5.110e-07
I9113 0 n9114 2.976e-02A M=1.655e-06
I9114 0 n9115 2.976e-02A M=1.036e-06
I9115 0 n9116 2.976e-02A M=6.803e-07
I9116 0 n9117 2.976e-02A M=4.589e-07
I9117 0 n9118 2.976e-02A M=3.260e-06
I9118 0 n9119 2.976e-02A M=6.220e-07
I9119 0 n9120 2.976e-02A M=1.499e-06
I9120 0 n9121 2.976e-02A M=6.944e-07
I9121 0 n9122 2.976e-02A M=1.475e-06
I9122 0 n9123 2.976e-02A M=5.548e-07
I9123 0 n9124 2.976e-02A M=1.175e-06
I9124 0 n9125 2.976e-02A M=3.769e-07
I9125 0 n9126 2.976e-02A M=2.746e-06
I9126 0 n9127 2.976e-02A M=1.436e-06
I9127 0 n9128 2.976e-02A M=9.416e-07
I9128 0 n9129 2.976e-02A M=6.171e-07
I9129 0 n9130 2.976e-02A M=7.856e-07
I9130 0 n9131 2.976e-02A M=1.264e-06
I9131 0 n9132 2.976e-02A M=9.014e-07
I9132 0 n9133 2.976e-02A M=1.325e-06
I9133 0 n9134 2.976e-02A M=5.441e-07
I9134 0 n9135 2.976e-02A M=4.225e-07
I9135 0 n9136 2.976e-02A M=1.005e-06
I9136 0 n9137 2.976e-02A M=6.365e-07
I9137 0 n1 2.976e-02A M=1.855e-06
I9138 0 n9139 2.976e-02A M=1.633e-06
I9139 0 n9140 2.976e-02A M=9.594e-07
I9140 0 n9141 2.976e-02A M=9.904e-07
I9141 0 n9142 2.976e-02A M=8.540e-07
I9142 0 n9143 2.976e-02A M=7.636e-07
I9143 0 n9144 2.976e-02A M=3.969e-07
I9144 0 n9145 2.976e-02A M=8.321e-07
I9145 0 n9146 2.976e-02A M=8.587e-07
I9146 0 n9147 2.976e-02A M=9.099e-07
I9147 0 n9148 2.976e-02A M=7.646e-07
I9148 0 n9149 2.976e-02A M=1.185e-06
I9149 0 n9150 2.976e-02A M=1.739e-06
I9150 0 n9151 2.976e-02A M=6.121e-07
I9151 0 n9152 2.976e-02A M=5.068e-07
I9152 0 n9153 2.976e-02A M=3.735e-07
I9153 0 n9154 2.976e-02A M=2.117e-06
I9154 0 n9155 2.976e-02A M=6.947e-07
I9155 0 n9156 2.976e-02A M=1.116e-06
I9156 0 n9157 2.976e-02A M=9.158e-07
I9157 0 n9158 2.976e-02A M=1.597e-06
I9158 0 n9159 2.976e-02A M=3.499e-07
I9159 0 n9160 2.976e-02A M=8.128e-07
I9160 0 n9161 2.976e-02A M=4.126e-07
I9161 0 n9162 2.976e-02A M=5.300e-07
I9162 0 n9163 2.976e-02A M=1.212e-06
I9163 0 n9164 2.976e-02A M=4.911e-07
I9164 0 n9165 2.976e-02A M=3.226e-07
I9165 0 n9166 2.976e-02A M=8.434e-07
I9166 0 n9167 2.976e-02A M=1.844e-06
I9167 0 n9168 2.976e-02A M=1.994e-06
I9168 0 n9169 2.976e-02A M=1.664e-06
I9169 0 n9170 2.976e-02A M=1.693e-07
I9170 0 n9171 2.976e-02A M=5.608e-07
I9171 0 n9172 2.976e-02A M=1.186e-06
I9172 0 n9173 2.976e-02A M=4.959e-07
I9173 0 n9174 2.976e-02A M=6.902e-07
I9174 0 n9175 2.976e-02A M=6.850e-07
I9175 0 n9176 2.976e-02A M=5.440e-07
I9176 0 n9177 2.976e-02A M=1.456e-06
I9177 0 n9178 2.976e-02A M=1.354e-06
I9178 0 n9179 2.976e-02A M=6.425e-07
I9179 0 n9180 2.976e-02A M=9.429e-07
I9180 0 n9181 2.976e-02A M=8.092e-07
I9181 0 n9182 2.976e-02A M=8.470e-07
I9182 0 n9183 2.976e-02A M=2.738e-07
I9183 0 n9184 2.976e-02A M=2.340e-07
I9184 0 n9185 2.976e-02A M=5.094e-07
I9185 0 n9186 2.976e-02A M=1.107e-06
I9186 0 n9187 2.976e-02A M=5.820e-07
I9187 0 n9188 2.976e-02A M=7.728e-07
I9188 0 n9189 2.976e-02A M=1.347e-06
I9189 0 n9190 2.976e-02A M=5.425e-07
I9190 0 n9191 2.976e-02A M=1.077e-06
I9191 0 n9192 2.976e-02A M=5.925e-07
I9192 0 n9193 2.976e-02A M=3.080e-07
I9193 0 n9194 2.976e-02A M=8.663e-07
I9194 0 n9195 2.976e-02A M=1.242e-07
I9195 0 n9196 2.976e-02A M=1.748e-07
I9196 0 n9197 2.976e-02A M=3.020e-07
I9197 0 n9198 2.976e-02A M=1.269e-06
I9198 0 n9199 2.976e-02A M=7.740e-07
I9199 0 n9200 2.976e-02A M=1.074e-06
I9200 0 n9201 2.976e-02A M=5.049e-07
I9201 0 n9202 2.976e-02A M=1.825e-06
I9202 0 n9203 2.976e-02A M=1.271e-06
I9203 0 n9204 2.976e-02A M=1.557e-06
I9204 0 n9205 2.976e-02A M=2.537e-06
I9205 0 n9206 2.976e-02A M=1.177e-06
I9206 0 n9207 2.976e-02A M=1.151e-06
I9207 0 n9208 2.976e-02A M=8.917e-07
I9208 0 n9209 2.976e-02A M=9.338e-07
I9209 0 n9210 2.976e-02A M=1.934e-06
I9210 0 n9211 2.976e-02A M=7.611e-07
I9211 0 n9212 2.976e-02A M=2.270e-06
I9212 0 n9213 2.976e-02A M=1.177e-06
I9213 0 n9214 2.976e-02A M=9.970e-07
I9214 0 n9215 2.976e-02A M=3.758e-07
I9215 0 n9216 2.976e-02A M=1.271e-06
I9216 0 n9217 2.976e-02A M=9.860e-07
I9217 0 n9218 2.976e-02A M=7.411e-07
I9218 0 n9219 2.976e-02A M=4.153e-07
I9219 0 n9220 2.976e-02A M=1.100e-06
I9220 0 n9221 2.976e-02A M=1.376e-06
I9221 0 n9222 2.976e-02A M=1.106e-06
I9222 0 n9223 2.976e-02A M=6.913e-07
I9223 0 n9224 2.976e-02A M=7.855e-07
I9224 0 n9225 2.976e-02A M=9.579e-07
I9225 0 n9226 2.976e-02A M=1.427e-07
I9226 0 n9227 2.976e-02A M=5.797e-07
I9227 0 n9228 2.976e-02A M=1.162e-06
I9228 0 n9229 2.976e-02A M=1.303e-06
I9229 0 n9230 2.976e-02A M=1.014e-06
I9230 0 n9231 2.976e-02A M=1.837e-06
I9231 0 n9232 2.976e-02A M=4.486e-07
I9232 0 n9233 2.976e-02A M=8.420e-07
I9233 0 n9234 2.976e-02A M=1.223e-06
I9234 0 n9235 2.976e-02A M=1.072e-06
I9235 0 n9236 2.976e-02A M=6.895e-07
I9236 0 n9237 2.976e-02A M=1.488e-06
I9237 0 n9238 2.976e-02A M=4.379e-07
I9238 0 n9239 2.976e-02A M=7.838e-07
I9239 0 n9240 2.976e-02A M=1.094e-06
I9240 0 n9241 2.976e-02A M=9.197e-07
I9241 0 n9242 2.976e-02A M=2.238e-07
I9242 0 n9243 2.976e-02A M=8.006e-07
I9243 0 n9244 2.976e-02A M=1.000e-06
I9244 0 n9245 2.976e-02A M=7.979e-07
I9245 0 n9246 2.976e-02A M=5.401e-07
I9246 0 n9247 2.976e-02A M=7.731e-07
I9247 0 n9248 2.976e-02A M=8.708e-07
I9248 0 n9249 2.976e-02A M=1.458e-06
I9249 0 n9250 2.976e-02A M=8.660e-07
I9250 0 n9251 2.976e-02A M=7.692e-07
I9251 0 n9252 2.976e-02A M=1.181e-06
I9252 0 n9253 2.976e-02A M=1.160e-06
I9253 0 n9254 2.976e-02A M=1.507e-06
I9254 0 n9255 2.976e-02A M=7.987e-07
I9255 0 n9256 2.976e-02A M=9.246e-07
I9256 0 n9257 2.976e-02A M=1.928e-06
I9257 0 n9258 2.976e-02A M=1.170e-06
I9258 0 n9259 2.976e-02A M=5.751e-07
I9259 0 n9260 2.976e-02A M=3.619e-07
I9260 0 n9261 2.976e-02A M=6.095e-07
I9261 0 n9262 2.976e-02A M=2.847e-07
I9262 0 n9263 2.976e-02A M=1.003e-06
I9263 0 n9264 2.976e-02A M=1.065e-06
I9264 0 n9265 2.976e-02A M=4.645e-07
I9265 0 n9266 2.976e-02A M=1.106e-06
I9266 0 n9267 2.976e-02A M=4.273e-07
I9267 0 n9268 2.976e-02A M=8.742e-07
I9268 0 n9269 2.976e-02A M=4.871e-07
I9269 0 n9270 2.976e-02A M=7.915e-07
I9270 0 n9271 2.976e-02A M=1.443e-06
I9271 0 n9272 2.976e-02A M=2.170e-06
I9272 0 n9273 2.976e-02A M=4.834e-07
I9273 0 n9274 2.976e-02A M=4.411e-07
I9274 0 n9275 2.976e-02A M=1.416e-06
I9275 0 n9276 2.976e-02A M=1.547e-06
I9276 0 n9277 2.976e-02A M=8.223e-07
I9277 0 n9278 2.976e-02A M=1.893e-07
I9278 0 n9279 2.976e-02A M=8.586e-07
I9279 0 n9280 2.976e-02A M=7.546e-07
I9280 0 n9281 2.976e-02A M=3.663e-07
I9281 0 n9282 2.976e-02A M=1.730e-06
I9282 0 n9283 2.976e-02A M=9.320e-07
I9283 0 n9284 2.976e-02A M=1.109e-06
I9284 0 n9285 2.976e-02A M=9.532e-07
I9285 0 n9286 2.976e-02A M=1.414e-06
I9286 0 n9287 2.976e-02A M=7.385e-07
I9287 0 n9288 2.976e-02A M=1.432e-06
I9288 0 n9289 2.976e-02A M=1.943e-06
I9289 0 n9290 2.976e-02A M=1.584e-06
I9290 0 n9291 2.976e-02A M=4.575e-07
I9291 0 n9292 2.976e-02A M=1.620e-06
I9292 0 n9293 2.976e-02A M=1.076e-06
I9293 0 n9294 2.976e-02A M=5.032e-07
I9294 0 n9295 2.976e-02A M=1.326e-06
I9295 0 n9296 2.976e-02A M=9.752e-07
I9296 0 n9297 2.976e-02A M=3.649e-07
I9297 0 n9298 2.976e-02A M=2.807e-06
I9298 0 n9299 2.976e-02A M=1.604e-06
I9299 0 n9300 2.976e-02A M=2.830e-07
I9300 0 n9301 2.976e-02A M=6.572e-07
I9301 0 n9302 2.976e-02A M=5.747e-07
I9302 0 n9303 2.976e-02A M=1.681e-06
I9303 0 n9304 2.976e-02A M=1.004e-06
I9304 0 n9305 2.976e-02A M=3.317e-07
I9305 0 n9306 2.976e-02A M=1.716e-06
I9306 0 n9307 2.976e-02A M=1.914e-06
I9307 0 n9308 2.976e-02A M=8.640e-07
I9308 0 n9309 2.976e-02A M=1.657e-06
I9309 0 n9310 2.976e-02A M=7.621e-07
I9310 0 n9311 2.976e-02A M=9.867e-07
I9311 0 n9312 2.976e-02A M=4.117e-07
I9312 0 n9313 2.976e-02A M=1.366e-06
I9313 0 n9314 2.976e-02A M=3.528e-07
I9314 0 n9315 2.976e-02A M=1.322e-06
I9315 0 n9316 2.976e-02A M=8.340e-07
I9316 0 n9317 2.976e-02A M=6.045e-07
I9317 0 n9318 2.976e-02A M=8.800e-07
I9318 0 n9319 2.976e-02A M=7.363e-07
I9319 0 n9320 2.976e-02A M=1.266e-06
I9320 0 n9321 2.976e-02A M=1.445e-06
I9321 0 n9322 2.976e-02A M=1.959e-06
I9322 0 n9323 2.976e-02A M=1.407e-06
I9323 0 n9324 2.976e-02A M=7.654e-07
I9324 0 n1 2.976e-02A M=9.194e-07
I9325 0 n9326 2.976e-02A M=5.794e-07
I9326 0 n9327 2.976e-02A M=1.413e-06
I9327 0 n9328 2.976e-02A M=5.108e-07
I9328 0 n9329 2.976e-02A M=4.352e-07
I9329 0 n9330 2.976e-02A M=2.216e-07
I9330 0 n9331 2.976e-02A M=5.426e-07
I9331 0 n9332 2.976e-02A M=1.917e-06
I9332 0 n9333 2.976e-02A M=1.038e-06
I9333 0 n9334 2.976e-02A M=6.376e-07
I9334 0 n9335 2.976e-02A M=3.560e-07
I9335 0 n9336 2.976e-02A M=1.352e-07
I9336 0 n9337 2.976e-02A M=4.764e-07
I9337 0 n9338 2.976e-02A M=1.040e-06
I9338 0 n9339 2.976e-02A M=1.784e-06
I9339 0 n9340 2.976e-02A M=3.271e-07
I9340 0 n9341 2.976e-02A M=3.134e-07
I9341 0 n9342 2.976e-02A M=2.185e-06
I9342 0 n9343 2.976e-02A M=2.946e-07
I9343 0 n9344 2.976e-02A M=1.260e-06
I9344 0 n9345 2.976e-02A M=1.001e-06
I9345 0 n9346 2.976e-02A M=1.429e-06
I9346 0 n9347 2.976e-02A M=1.361e-06
I9347 0 n9348 2.976e-02A M=4.281e-07
I9348 0 n9349 2.976e-02A M=1.296e-06
I9349 0 n9350 2.976e-02A M=6.922e-07
I9350 0 n9351 2.976e-02A M=6.154e-07
I9351 0 n9352 2.976e-02A M=6.006e-07
I9352 0 n9353 2.976e-02A M=8.781e-07
I9353 0 n9354 2.976e-02A M=1.306e-06
I9354 0 n9355 2.976e-02A M=1.285e-06
I9355 0 n9356 2.976e-02A M=6.447e-07
I9356 0 n9357 2.976e-02A M=2.246e-07
I9357 0 n9358 2.976e-02A M=7.244e-07
I9358 0 n9359 2.976e-02A M=7.382e-07
I9359 0 n9360 2.976e-02A M=5.200e-07
I9360 0 n9361 2.976e-02A M=8.816e-07
I9361 0 n9362 2.976e-02A M=4.203e-07
I9362 0 n9363 2.976e-02A M=6.849e-07
I9363 0 n9364 2.976e-02A M=9.534e-07
I9364 0 n9365 2.976e-02A M=1.670e-06
I9365 0 n9366 2.976e-02A M=1.254e-06
I9366 0 n9367 2.976e-02A M=5.298e-07
I9367 0 n9368 2.976e-02A M=9.960e-07
I9368 0 n9369 2.976e-02A M=1.227e-06
I9369 0 n9370 2.976e-02A M=1.460e-06
I9370 0 n9371 2.976e-02A M=4.797e-07
I9371 0 n9372 2.976e-02A M=4.509e-07
I9372 0 n9373 2.976e-02A M=1.497e-06
I9373 0 n9374 2.976e-02A M=5.381e-07
I9374 0 n9375 2.976e-02A M=1.034e-06
I9375 0 n9376 2.976e-02A M=4.288e-07
I9376 0 n9377 2.976e-02A M=8.231e-07
I9377 0 n9378 2.976e-02A M=1.783e-06
I9378 0 n9379 2.976e-02A M=1.662e-06
I9379 0 n9380 2.976e-02A M=1.190e-06
I9380 0 n9381 2.976e-02A M=7.706e-07
I9381 0 n9382 2.976e-02A M=2.200e-07
I9382 0 n9383 2.976e-02A M=8.227e-07
I9383 0 n9384 2.976e-02A M=6.616e-07
I9384 0 n9385 2.976e-02A M=5.589e-07
I9385 0 n9386 2.976e-02A M=1.075e-06
I9386 0 n9387 2.976e-02A M=1.821e-06
I9387 0 n9388 2.976e-02A M=2.202e-06
I9388 0 n9389 2.976e-02A M=6.938e-07
I9389 0 n9390 2.976e-02A M=5.198e-07
I9390 0 n9391 2.976e-02A M=7.991e-07
I9391 0 n9392 2.976e-02A M=5.208e-07
I9392 0 n9393 2.976e-02A M=1.003e-06
I9393 0 n9394 2.976e-02A M=7.983e-07
I9394 0 n9395 2.976e-02A M=5.863e-07
I9395 0 n9396 2.976e-02A M=2.169e-07
I9396 0 n9397 2.976e-02A M=2.355e-07
I9397 0 n9398 2.976e-02A M=2.596e-07
I9398 0 n9399 2.976e-02A M=3.143e-07
I9399 0 n9400 2.976e-02A M=1.151e-06
I9400 0 n9401 2.976e-02A M=7.042e-07
I9401 0 n9402 2.976e-02A M=7.218e-07
I9402 0 n9403 2.976e-02A M=7.292e-07
I9403 0 n9404 2.976e-02A M=5.938e-07
I9404 0 n9405 2.976e-02A M=1.936e-06
I9405 0 n9406 2.976e-02A M=7.133e-07
I9406 0 n9407 2.976e-02A M=9.208e-07
I9407 0 n9408 2.976e-02A M=1.420e-06
I9408 0 n9409 2.976e-02A M=1.093e-06
I9409 0 n9410 2.976e-02A M=4.933e-07
I9410 0 n9411 2.976e-02A M=7.933e-07
I9411 0 n9412 2.976e-02A M=1.038e-06
I9412 0 n9413 2.976e-02A M=1.623e-06
I9413 0 n9414 2.976e-02A M=3.005e-07
I9414 0 n9415 2.976e-02A M=6.112e-07
I9415 0 n9416 2.976e-02A M=1.242e-06
I9416 0 n9417 2.976e-02A M=1.571e-06
I9417 0 n9418 2.976e-02A M=2.266e-06
I9418 0 n9419 2.976e-02A M=1.034e-06
I9419 0 n9420 2.976e-02A M=7.575e-07
I9420 0 n9421 2.976e-02A M=6.052e-07
I9421 0 n9422 2.976e-02A M=8.355e-07
I9422 0 n9423 2.976e-02A M=9.919e-07
I9423 0 n9424 2.976e-02A M=7.359e-07
I9424 0 n9425 2.976e-02A M=1.493e-06
I9425 0 n9426 2.976e-02A M=2.462e-07
I9426 0 n9427 2.976e-02A M=5.893e-07
I9427 0 n9428 2.976e-02A M=4.235e-07
I9428 0 n9429 2.976e-02A M=7.408e-07
I9429 0 n9430 2.976e-02A M=5.185e-07
I9430 0 n9431 2.976e-02A M=6.979e-07
I9431 0 n9432 2.976e-02A M=8.173e-07
I9432 0 n9433 2.976e-02A M=1.193e-06
I9433 0 n9434 2.976e-02A M=8.609e-07
I9434 0 n9435 2.976e-02A M=1.429e-06
I9435 0 n9436 2.976e-02A M=3.458e-06
I9436 0 n9437 2.976e-02A M=1.120e-06
I9437 0 n9438 2.976e-02A M=1.146e-07
I9438 0 n9439 2.976e-02A M=8.051e-07
I9439 0 n9440 2.976e-02A M=1.068e-06
I9440 0 n9441 2.976e-02A M=7.821e-07
I9441 0 n9442 2.976e-02A M=3.458e-07
I9442 0 n9443 2.976e-02A M=1.338e-06
I9443 0 n9444 2.976e-02A M=1.536e-06
I9444 0 n9445 2.976e-02A M=2.610e-06
I9445 0 n9446 2.976e-02A M=1.369e-06
I9446 0 n9447 2.976e-02A M=6.551e-07
I9447 0 n9448 2.976e-02A M=9.482e-07
I9448 0 n9449 2.976e-02A M=1.038e-06
I9449 0 n9450 2.976e-02A M=1.521e-06
I9450 0 n9451 2.976e-02A M=2.089e-06
I9451 0 n9452 2.976e-02A M=1.398e-06
I9452 0 n9453 2.976e-02A M=1.007e-06
I9453 0 n9454 2.976e-02A M=6.556e-07
I9454 0 n9455 2.976e-02A M=1.641e-07
I9455 0 n9456 2.976e-02A M=1.272e-06
I9456 0 n9457 2.976e-02A M=4.481e-07
I9457 0 n9458 2.976e-02A M=9.561e-07
I9458 0 n9459 2.976e-02A M=3.976e-07
I9459 0 n9460 2.976e-02A M=5.475e-07
I9460 0 n9461 2.976e-02A M=1.143e-06
I9461 0 n9462 2.976e-02A M=1.515e-06
I9462 0 n9463 2.976e-02A M=7.430e-07
I9463 0 n9464 2.976e-02A M=1.416e-06
I9464 0 n9465 2.976e-02A M=1.050e-06
I9465 0 n9466 2.976e-02A M=4.960e-07
I9466 0 n9467 2.976e-02A M=4.925e-07
I9467 0 n9468 2.976e-02A M=7.081e-07
I9468 0 n9469 2.976e-02A M=1.526e-06
I9469 0 n9470 2.976e-02A M=8.594e-07
I9470 0 n9471 2.976e-02A M=1.062e-06
I9471 0 n9472 2.976e-02A M=1.281e-06
I9472 0 n9473 2.976e-02A M=7.555e-07
I9473 0 n9474 2.976e-02A M=7.517e-07
I9474 0 n9475 2.976e-02A M=9.537e-07
I9475 0 n9476 2.976e-02A M=5.160e-07
I9476 0 n9477 2.976e-02A M=6.872e-07
I9477 0 n9478 2.976e-02A M=3.708e-07
I9478 0 n9479 2.976e-02A M=1.022e-06
I9479 0 n9480 2.976e-02A M=1.646e-06
I9480 0 n9481 2.976e-02A M=1.643e-06
I9481 0 n9482 2.976e-02A M=6.375e-07
I9482 0 n9483 2.976e-02A M=9.534e-07
I9483 0 n9484 2.976e-02A M=2.337e-07
I9484 0 n9485 2.976e-02A M=9.238e-07
I9485 0 n9486 2.976e-02A M=6.732e-07
I9486 0 n9487 2.976e-02A M=1.816e-06
I9487 0 n9488 2.976e-02A M=7.160e-07
I9488 0 n9489 2.976e-02A M=6.668e-07
I9489 0 n9490 2.976e-02A M=1.067e-06
I9490 0 n9491 2.976e-02A M=1.108e-06
I9491 0 n9492 2.976e-02A M=4.998e-07
I9492 0 n9493 2.976e-02A M=1.928e-06
I9493 0 n9494 2.976e-02A M=1.155e-06
I9494 0 n9495 2.976e-02A M=1.040e-06
I9495 0 n9496 2.976e-02A M=6.379e-07
I9496 0 n9497 2.976e-02A M=6.973e-07
I9497 0 n9498 2.976e-02A M=3.038e-07
I9498 0 n9499 2.976e-02A M=7.334e-07
I9499 0 n9500 2.976e-02A M=1.474e-07
I9500 0 n9501 2.976e-02A M=3.476e-07
I9501 0 n9502 2.976e-02A M=6.793e-07
I9502 0 n9503 2.976e-02A M=1.510e-06
I9503 0 n9504 2.976e-02A M=3.998e-07
I9504 0 n9505 2.976e-02A M=8.567e-07
I9505 0 n9506 2.976e-02A M=1.991e-06
I9506 0 n9507 2.976e-02A M=1.582e-06
I9507 0 n9508 2.976e-02A M=6.213e-07
I9508 0 n9509 2.976e-02A M=5.476e-07
I9509 0 n9510 2.976e-02A M=4.532e-06
I9510 0 n1 2.976e-02A M=7.783e-07
I9511 0 n9512 2.976e-02A M=1.631e-06
I9512 0 n9513 2.976e-02A M=6.741e-07
I9513 0 n9514 2.976e-02A M=6.873e-07
I9514 0 n9515 2.976e-02A M=2.652e-06
I9515 0 n9516 2.976e-02A M=7.689e-07
I9516 0 n9517 2.976e-02A M=1.182e-06
I9517 0 n9518 2.976e-02A M=5.291e-07
I9518 0 n9519 2.976e-02A M=9.869e-07
I9519 0 n9520 2.976e-02A M=9.682e-07
I9520 0 n9521 2.976e-02A M=8.429e-07
I9521 0 n9522 2.976e-02A M=1.521e-06
I9522 0 n9523 2.976e-02A M=8.640e-07
I9523 0 n9524 2.976e-02A M=5.145e-07
I9524 0 n9525 2.976e-02A M=3.031e-06
I9525 0 n9526 2.976e-02A M=9.136e-07
I9526 0 n9527 2.976e-02A M=6.582e-07
I9527 0 n9528 2.976e-02A M=9.429e-07
I9528 0 n9529 2.976e-02A M=1.863e-06
I9529 0 n9530 2.976e-02A M=6.212e-07
I9530 0 n9531 2.976e-02A M=3.090e-07
I9531 0 n9532 2.976e-02A M=6.298e-07
I9532 0 n9533 2.976e-02A M=5.710e-07
I9533 0 n9534 2.976e-02A M=8.921e-07
I9534 0 n9535 2.976e-02A M=1.170e-06
I9535 0 n9536 2.976e-02A M=1.010e-06
I9536 0 n9537 2.976e-02A M=7.272e-07
I9537 0 n9538 2.976e-02A M=7.079e-07
I9538 0 n9539 2.976e-02A M=2.616e-07
I9539 0 n9540 2.976e-02A M=4.876e-07
I9540 0 n9541 2.976e-02A M=6.972e-07
I9541 0 n9542 2.976e-02A M=8.982e-07
I9542 0 n9543 2.976e-02A M=8.724e-07
I9543 0 n9544 2.976e-02A M=3.367e-07
I9544 0 n9545 2.976e-02A M=6.689e-07
I9545 0 n9546 2.976e-02A M=2.181e-06
I9546 0 n9547 2.976e-02A M=1.097e-06
I9547 0 n9548 2.976e-02A M=1.864e-06
I9548 0 n9549 2.976e-02A M=9.513e-07
I9549 0 n9550 2.976e-02A M=1.146e-06
I9550 0 n9551 2.976e-02A M=1.317e-06
I9551 0 n9552 2.976e-02A M=5.920e-07
I9552 0 n9553 2.976e-02A M=5.551e-07
I9553 0 n9554 2.976e-02A M=5.016e-07
I9554 0 n9555 2.976e-02A M=6.088e-07
I9555 0 n9556 2.976e-02A M=3.976e-07
I9556 0 n9557 2.976e-02A M=3.396e-07
I9557 0 n9558 2.976e-02A M=9.007e-07
I9558 0 n9559 2.976e-02A M=1.675e-06
I9559 0 n9560 2.976e-02A M=1.837e-06
I9560 0 n9561 2.976e-02A M=1.150e-06
I9561 0 n9562 2.976e-02A M=1.023e-06
I9562 0 n9563 2.976e-02A M=1.431e-06
I9563 0 n9564 2.976e-02A M=9.924e-07
I9564 0 n9565 2.976e-02A M=1.052e-06
I9565 0 n9566 2.976e-02A M=2.047e-06
I9566 0 n9567 2.976e-02A M=1.060e-06
I9567 0 n9568 2.976e-02A M=2.610e-06
I9568 0 n9569 2.976e-02A M=7.388e-07
I9569 0 n9570 2.976e-02A M=1.067e-06
I9570 0 n9571 2.976e-02A M=8.288e-07
I9571 0 n9572 2.976e-02A M=4.478e-07
I9572 0 n9573 2.976e-02A M=1.655e-06
I9573 0 n9574 2.976e-02A M=6.132e-07
I9574 0 n9575 2.976e-02A M=4.920e-07
I9575 0 n9576 2.976e-02A M=5.715e-07
I9576 0 n9577 2.976e-02A M=7.866e-07
I9577 0 n9578 2.976e-02A M=1.138e-06
I9578 0 n9579 2.976e-02A M=1.030e-06
I9579 0 n9580 2.976e-02A M=1.506e-06
I9580 0 n9581 2.976e-02A M=1.267e-06
I9581 0 n9582 2.976e-02A M=7.889e-07
I9582 0 n9583 2.976e-02A M=8.314e-07
I9583 0 n9584 2.976e-02A M=1.004e-06
I9584 0 n9585 2.976e-02A M=8.009e-07
I9585 0 n9586 2.976e-02A M=7.611e-07
I9586 0 n9587 2.976e-02A M=4.170e-07
I9587 0 n9588 2.976e-02A M=1.871e-06
I9588 0 n9589 2.976e-02A M=9.054e-07
I9589 0 n9590 2.976e-02A M=1.432e-06
I9590 0 n9591 2.976e-02A M=1.533e-06
I9591 0 n9592 2.976e-02A M=5.691e-07
I9592 0 n9593 2.976e-02A M=8.998e-07
I9593 0 n9594 2.976e-02A M=7.398e-07
I9594 0 n9595 2.976e-02A M=1.034e-06
I9595 0 n9596 2.976e-02A M=7.818e-07
I9596 0 n9597 2.976e-02A M=5.203e-07
I9597 0 n9598 2.976e-02A M=8.172e-07
I9598 0 n9599 2.976e-02A M=8.415e-07
I9599 0 n9600 2.976e-02A M=5.248e-07
I9600 0 n9601 2.976e-02A M=1.139e-06
I9601 0 n9602 2.976e-02A M=1.373e-06
I9602 0 n9603 2.976e-02A M=9.635e-07
I9603 0 n9604 2.976e-02A M=7.291e-07
I9604 0 n9605 2.976e-02A M=9.277e-07
I9605 0 n9606 2.976e-02A M=1.231e-06
I9606 0 n9607 2.976e-02A M=8.469e-07
I9607 0 n9608 2.976e-02A M=1.300e-06
I9608 0 n9609 2.976e-02A M=6.015e-07
I9609 0 n9610 2.976e-02A M=5.326e-07
I9610 0 n9611 2.976e-02A M=9.348e-07
I9611 0 n9612 2.976e-02A M=7.769e-07
I9612 0 n9613 2.976e-02A M=9.402e-07
I9613 0 n9614 2.976e-02A M=8.846e-07
I9614 0 n9615 2.976e-02A M=8.852e-07
I9615 0 n9616 2.976e-02A M=6.610e-07
I9616 0 n9617 2.976e-02A M=1.097e-06
I9617 0 n9618 2.976e-02A M=3.541e-07
I9618 0 n9619 2.976e-02A M=1.657e-06
I9619 0 n9620 2.976e-02A M=1.480e-06
I9620 0 n9621 2.976e-02A M=8.351e-07
I9621 0 n9622 2.976e-02A M=1.346e-06
I9622 0 n9623 2.976e-02A M=6.994e-07
I9623 0 n9624 2.976e-02A M=1.522e-06
I9624 0 n9625 2.976e-02A M=9.017e-07
I9625 0 n9626 2.976e-02A M=1.305e-06
I9626 0 n9627 2.976e-02A M=1.050e-06
I9627 0 n9628 2.976e-02A M=7.879e-07
I9628 0 n9629 2.976e-02A M=4.125e-07
I9629 0 n9630 2.976e-02A M=9.480e-07
I9630 0 n9631 2.976e-02A M=8.513e-07
I9631 0 n9632 2.976e-02A M=1.032e-06
I9632 0 n9633 2.976e-02A M=1.223e-06
I9633 0 n9634 2.976e-02A M=4.641e-07
I9634 0 n9635 2.976e-02A M=1.153e-06
I9635 0 n9636 2.976e-02A M=1.725e-06
I9636 0 n9637 2.976e-02A M=4.619e-07
I9637 0 n9638 2.976e-02A M=6.284e-07
I9638 0 n9639 2.976e-02A M=1.666e-07
I9639 0 n9640 2.976e-02A M=6.907e-07
I9640 0 n9641 2.976e-02A M=8.435e-07
I9641 0 n9642 2.976e-02A M=1.141e-06
I9642 0 n9643 2.976e-02A M=4.235e-07
I9643 0 n9644 2.976e-02A M=6.501e-07
I9644 0 n9645 2.976e-02A M=8.644e-07
I9645 0 n9646 2.976e-02A M=8.490e-07
I9646 0 n9647 2.976e-02A M=3.355e-07
I9647 0 n9648 2.976e-02A M=2.073e-07
I9648 0 n9649 2.976e-02A M=1.876e-06
I9649 0 n9650 2.976e-02A M=7.931e-07
I9650 0 n9651 2.976e-02A M=1.499e-06
I9651 0 n9652 2.976e-02A M=5.959e-07
I9652 0 n9653 2.976e-02A M=1.234e-06
I9653 0 n9654 2.976e-02A M=1.266e-07
I9654 0 n9655 2.976e-02A M=7.865e-07
I9655 0 n9656 2.976e-02A M=1.410e-06
I9656 0 n9657 2.976e-02A M=8.365e-07
I9657 0 n9658 2.976e-02A M=2.736e-07
I9658 0 n9659 2.976e-02A M=5.500e-07
I9659 0 n9660 2.976e-02A M=5.077e-07
I9660 0 n9661 2.976e-02A M=2.851e-06
I9661 0 n9662 2.976e-02A M=3.874e-07
I9662 0 n9663 2.976e-02A M=1.899e-07
I9663 0 n9664 2.976e-02A M=1.124e-06
I9664 0 n9665 2.976e-02A M=9.594e-07
I9665 0 n9666 2.976e-02A M=1.198e-06
I9666 0 n9667 2.976e-02A M=3.388e-07
I9667 0 n9668 2.976e-02A M=7.647e-07
I9668 0 n9669 2.976e-02A M=1.153e-06
I9669 0 n9670 2.976e-02A M=1.519e-06
I9670 0 n9671 2.976e-02A M=9.150e-07
I9671 0 n9672 2.976e-02A M=2.656e-07
I9672 0 n9673 2.976e-02A M=5.401e-07
I9673 0 n9674 2.976e-02A M=1.041e-06
I9674 0 n9675 2.976e-02A M=6.627e-07
I9675 0 n9676 2.976e-02A M=1.828e-06
I9676 0 n9677 2.976e-02A M=1.393e-06
I9677 0 n9678 2.976e-02A M=7.512e-07
I9678 0 n9679 2.976e-02A M=1.307e-06
I9679 0 n9680 2.976e-02A M=1.295e-06
I9680 0 n9681 2.976e-02A M=1.027e-06
I9681 0 n9682 2.976e-02A M=1.021e-06
I9682 0 n9683 2.976e-02A M=1.589e-06
I9683 0 n9684 2.976e-02A M=1.120e-06
I9684 0 n9685 2.976e-02A M=6.454e-07
I9685 0 n9686 2.976e-02A M=7.855e-07
I9686 0 n9687 2.976e-02A M=3.530e-07
I9687 0 n9688 2.976e-02A M=6.499e-07
I9688 0 n9689 2.976e-02A M=9.164e-07
I9689 0 n9690 2.976e-02A M=8.907e-07
I9690 0 n9691 2.976e-02A M=6.591e-07
I9691 0 n9692 2.976e-02A M=3.735e-07
I9692 0 n9693 2.976e-02A M=7.748e-07
I9693 0 n9694 4.100e-03A M=3.488e-07

*** resistors
R91t61 n92 n62 R=9.802e+00 
R114t47 n115 n48 R=2.214e+01 
R148t4 n149 n5 R=5.262e+00 
R148t54 n149 n55 R=1.025e+01 
R154t89 n155 n90 R=1.092e+01 
R161t54 n162 n55 R=4.059e+00 
R193t184 n194 n185 R=1.268e+01 
R208t124 n209 n125 R=1.145e+01 
R226t168 n227 n169 R=3.259e+00 
R236t158 n237 n159 R=1.068e+01 
R236t179 n237 n180 R=4.507e+00 
R254t243 n255 n244 R=1.020e+01 
R266t28 n267 n29 R=2.345e+00 
R271t119 n272 n120 R=5.524e+01 
R275t48 n276 n49 R=1.201e+02 
R289t46 n290 n47 R=4.972e+02 
R292t173 n293 n174 R=7.428e+00 
R297t255 n298 n256 R=9.683e+00 
R303t13 n304 n14 R=5.542e+00 
R306t20 n307 n21 R=3.258e+00 
R308t290 n309 n291 R=1.368e+01 
R320t144 n321 n145 R=4.093e+00 
R321t186 n322 n187 R=8.250e+00 
R321t319 n322 n320 R=2.126e+01 
R346t114 n347 n115 R=1.113e+01 
R360t185 n361 n186 R=7.830e+00 
R365t334 n366 n335 R=2.691e+00 
R367t51 n368 n52 R=7.159e+00 
R370t279 n371 n280 R=4.741e+00 
R373t199 n374 n200 R=8.201e+00 
R376t39 n377 n40 R=1.549e+01 
R377t270 n378 n271 R=3.204e+00 
R378t272 n379 n273 R=2.205e+01 
R380t240 n381 n241 R=3.615e+00 
R385t194 n386 n195 R=5.976e+00 
R389t347 n390 n348 R=9.605e+02 
R393t57 n394 n58 R=8.829e+00 
R409t274 n410 n275 R=1.240e+01 
R411t87 n412 n88 R=1.348e+01 
R418t390 n419 n391 R=5.832e+00 
R423t65 n424 n66 R=2.100e+01 
R428t188 n429 n189 R=4.805e+00 
R434t430 n435 n431 R=4.257e+01 
R435t147 n436 n148 R=3.040e+01 
R443t49 n444 n50 R=1.504e+01 
R445t133 n446 n134 R=5.721e+00 
R445t35 n446 n36 R=2.466e+01 
R454t133 n455 n134 R=1.241e+01 
R457t58 n458 n59 R=8.238e+00 
R460t64 n461 n65 R=6.569e+00 
R460t245 n461 n246 R=6.424e+00 
R465t129 n466 n130 R=6.121e+00 
R467t312 n468 n313 R=1.815e+02 
R473t406 n474 n407 R=9.158e+02 
R475t362 n476 n363 R=4.995e+00 
R477t281 n478 n282 R=4.245e+01 
R480t82 n481 n83 R=4.625e+00 
R485t332 n486 n333 R=4.958e+01 
R489t10 n490 n11 R=3.343e+01 
R492t314 n493 n315 R=3.382e+00 
R495t442 n496 n443 R=5.619e+00 
R503t396 n504 n397 R=1.617e+00 
R507t468 n508 n469 R=1.609e+01 
R521t466 n522 n467 R=4.863e+02 
R526t491 n527 n492 R=4.858e+00 
R528t70 n529 n71 R=4.125e+00 
R529t242 n530 n243 R=3.607e+00 
R531t101 n532 n102 R=9.725e+00 
R533t239 n534 n240 R=1.073e+01 
R534t185 n535 n186 R=4.121e+00 
R539t505 n540 n506 R=2.623e+00 
R543t418 n544 n419 R=1.030e+02 
R549t438 n550 n439 R=7.342e+00 
R550t373 n551 n374 R=1.199e+01 
R551t480 n552 n481 R=1.330e+01 
R558t383 n559 n384 R=5.747e+00 
R560t429 n561 n430 R=7.624e+00 
R564t6 n565 n7 R=1.342e+00 
R565t425 n566 n426 R=2.264e+00 
R566t520 n567 n521 R=8.489e+00 
R566t411 n567 n412 R=7.597e+00 
R580t271 n581 n272 R=9.493e+02 
R582t331 n583 n332 R=8.513e+01 
R582t75 n583 n76 R=8.369e+00 
R584t77 n585 n78 R=2.657e+01 
R584t272 n585 n273 R=1.696e+01 
R587t100 n588 n101 R=2.927e+01 
R589t31 n590 n32 R=6.163e+00 
R589t580 n590 n581 R=4.388e+00 
R592t318 n593 n319 R=4.378e+01 
R592t55 n593 n56 R=1.522e+01 
R595t393 n596 n394 R=4.406e+00 
R595t57 n596 n58 R=4.844e+00 
R596t587 n597 n588 R=1.187e+01 
R596t100 n597 n101 R=4.405e+00 
R599t458 n600 n459 R=6.369e+00 
R600t15 n601 n16 R=1.216e+01 
R601t496 n602 n497 R=6.962e+00 
R601t159 n602 n160 R=1.519e+01 
R606t382 n607 n383 R=2.229e+01 
R609t238 n610 n239 R=2.595e+00 
R610t141 n611 n142 R=2.077e+00 
R613t55 n614 n56 R=3.733e+00 
R619t581 n620 n582 R=5.664e+00 
R625t27 n626 n28 R=1.021e+01 
R627t292 n628 n293 R=1.557e+02 
R637t264 n638 n265 R=2.563e+00 
R641t412 n642 n413 R=1.950e+00 
R647t197 n648 n198 R=3.346e+00 
R649t17 n650 n18 R=1.366e+01 
R652t33 n653 n34 R=9.986e+00 
R656t188 n657 n189 R=1.061e+01 
R656t428 n657 n429 R=1.568e+01 
R658t454 n659 n455 R=2.549e+01 
R660t241 n661 n242 R=2.765e+01 
R662t284 n663 n285 R=1.073e+01 
R665t325 n666 n326 R=4.008e+01 
R666t311 n667 n312 R=1.464e+01 
R667t559 n668 n560 R=2.507e+01 
R671t358 n672 n359 R=7.140e+00 
R673t13 n674 n14 R=2.333e+00 
R677t213 n678 n214 R=2.481e+00 
R679t127 n680 n128 R=4.724e+00 
R680t528 n681 n529 R=3.794e+00 
R681t5 n682 n6 R=4.835e+00 
R683t551 n684 n552 R=4.976e+00 
R685t361 n686 n362 R=4.615e+00 
R685t488 n686 n489 R=1.376e+01 
R690t542 n691 n543 R=7.943e+01 
R693t659 n694 n660 R=5.229e+00 
R694t525 n695 n526 R=3.292e+00 
R697t545 n698 n546 R=4.030e+00 
R699t95 n700 n96 R=6.270e+00 
R707t623 n708 n624 R=3.299e+00 
R714t675 n715 n676 R=3.045e+00 
R714t41 n715 n42 R=6.561e+00 
R716t145 n717 n146 R=2.203e+01 
R718t172 n719 n173 R=4.559e+00 
R721t650 n722 n651 R=5.354e+00 
R721t203 n722 n204 R=1.407e+01 
R724t595 n725 n596 R=7.428e+00 
R724t393 n725 n394 R=1.031e+02 
R726t130 n727 n131 R=2.119e+01 
R729t359 n730 n360 R=1.368e+02 
R729t252 n730 n253 R=9.325e+00 
R730t271 n731 n272 R=8.692e+01 
R731t714 n732 n715 R=7.924e+01 
R731t412 n732 n413 R=1.887e+01 
R736t162 n737 n163 R=1.743e+01 
R738t183 n739 n184 R=6.360e+00 
R738t169 n739 n170 R=8.455e+00 
R740t633 n741 n634 R=1.329e+01 
R743t198 n744 n199 R=3.852e+00 
R745t686 n746 n687 R=2.999e+01 
R745t548 n746 n549 R=3.285e+01 
R747t576 n748 n577 R=3.385e+00 
R749t572 n750 n573 R=1.200e+01 
R751t175 n752 n176 R=5.584e+00 
R752t328 n753 n329 R=5.975e+00 
R754t641 n755 n642 R=3.384e+00 
R755t36 n756 n37 R=3.209e+00 
R758t52 n759 n53 R=1.047e+01 
R758t673 n759 n674 R=6.293e+00 
R758t13 n759 n14 R=1.735e+01 
R759t535 n760 n536 R=2.919e+00 
R762t436 n763 n437 R=3.229e+00 
R763t659 n764 n660 R=9.632e+00 
R764t671 n765 n672 R=3.823e+00 
R764t358 n765 n359 R=1.214e+01 
R767t45 n768 n46 R=3.891e+00 
R767t457 n768 n458 R=4.029e+00 
R772t194 n773 n195 R=5.778e+00 
R772t385 n773 n386 R=7.812e+00 
R773t53 n774 n54 R=5.310e+00 
R775t509 n776 n510 R=2.526e+01 
R779t444 n780 n445 R=2.096e+01 
R781t402 n782 n403 R=6.276e+00 
R782t512 n783 n513 R=1.592e+02 
R783t244 n784 n245 R=8.263e+00 
R785t541 n786 n542 R=7.775e+00 
R786t172 n787 n173 R=1.313e+01 
R790t598 n791 n599 R=2.650e+00 
R792t504 n793 n505 R=3.617e+00 
R792t713 n793 n714 R=6.380e+00 
R797t518 n798 n519 R=1.860e+00 
R798t500 n799 n501 R=2.139e+01 
R798t661 n799 n662 R=5.339e+00 
R799t6 n800 n7 R=1.727e+00 
R801t22 n802 n23 R=3.876e+00 
R803t26 n804 n27 R=1.237e+02 
R804t228 n805 n229 R=2.531e+01 
R805t495 n806 n496 R=4.604e+00 
R807t753 n808 n754 R=5.113e+00 
R813t688 n814 n689 R=7.346e+00 
R816t763 n817 n764 R=2.110e+01 
R816t659 n817 n660 R=3.334e+00 
R817t88 n818 n89 R=6.169e+00 
R817t14 n818 n15 R=3.787e+01 
R819t26 n820 n27 R=1.780e+01 
R821t609 n822 n610 R=4.229e+00 
R822t17 n823 n18 R=1.501e+01 
R823t460 n824 n461 R=1.050e+01 
R823t245 n824 n246 R=2.043e+01 
R829t332 n830 n333 R=1.130e+01 
R829t485 n830 n486 R=5.344e+00 
R833t724 n834 n725 R=1.361e+01 
R835t135 n836 n136 R=1.229e+02 
R838t372 n839 n373 R=5.127e+00 
R839t118 n840 n119 R=2.434e+00 
R839t266 n840 n267 R=1.601e+01 
R840t714 n841 n715 R=5.805e+00 
R840t731 n841 n732 R=3.516e+00 
R842t206 n843 n207 R=5.445e+00 
R843t209 n844 n210 R=3.365e+00 
R844t781 n845 n782 R=4.129e+00 
R844t402 n845 n403 R=5.225e+00 
R845t807 n846 n808 R=1.639e+01 
R845t753 n846 n754 R=3.164e+00 
R849t138 n850 n139 R=5.460e+00 
R850t666 n851 n667 R=4.995e+00 
R852t580 n853 n581 R=8.075e+00 
R852t589 n853 n590 R=8.120e+01 
R853t825 n854 n826 R=3.362e+00 
R857t583 n858 n584 R=1.568e+01 
R858t26 n859 n27 R=2.687e+00 
R858t803 n859 n804 R=2.245e+01 
R859t785 n860 n786 R=5.941e+00 
R860t386 n861 n387 R=5.509e+00 
R860t66 n861 n67 R=7.383e+00 
R861t435 n862 n436 R=3.077e+01 
R861t537 n862 n538 R=5.484e+00 
R862t411 n863 n412 R=1.075e+01 
R863t164 n864 n165 R=2.892e+01 
R863t487 n864 n488 R=8.434e+00 
R864t284 n865 n285 R=6.690e+00 
R868t441 n869 n442 R=5.341e+00 
R868t129 n869 n130 R=5.363e+00 
R868t465 n869 n466 R=4.895e+02 
R869t366 n870 n367 R=2.184e+01 
R869t247 n870 n248 R=5.563e+00 
R871t69 n872 n70 R=1.094e+01 
R872t295 n873 n296 R=3.459e+00 
R875t200 n876 n201 R=5.558e+00 
R878t117 n879 n118 R=8.058e+00 
R878t736 n879 n737 R=9.589e+01 
R879t390 n880 n391 R=6.852e+00 
R883t370 n884 n371 R=4.199e+00 
R883t392 n884 n393 R=2.289e+02 
R884t184 n885 n185 R=8.178e+00 
R884t193 n885 n194 R=4.446e+00 
R887t400 n888 n401 R=1.428e+01 
R890t155 n891 n156 R=1.062e+02 
R892t274 n893 n275 R=1.959e+01 
R892t409 n893 n410 R=1.770e+01 
R894t877 n895 n878 R=5.862e+00 
R897t42 n1 n43 R=3.704e+01 
R900t757 n901 n758 R=5.163e+00 
R901t750 n902 n751 R=2.853e+00 
R904t116 n905 n117 R=2.495e+02 
R904t292 n905 n293 R=2.028e+01 
R906t569 n907 n570 R=1.488e+01 
R909t441 n910 n442 R=3.565e+00 
R909t868 n910 n869 R=4.597e+01 
R910t485 n911 n486 R=6.384e+00 
R911t880 n912 n881 R=4.797e+00 
R912t695 n913 n696 R=7.903e+00 
R913t648 n914 n649 R=1.864e+01 
R915t599 n916 n600 R=2.037e+01 
R917t789 n918 n790 R=7.956e+00 
R922t392 n923 n393 R=7.765e+00 
R929t138 n930 n139 R=6.610e+00 
R931t135 n932 n136 R=1.728e+01 
R931t835 n932 n836 R=6.431e+00 
R934t49 n935 n50 R=5.320e+00 
R937t562 n938 n563 R=1.326e+01 
R938t596 n939 n597 R=1.590e+02 
R939t900 n940 n901 R=8.542e+01 
R941t531 n942 n532 R=2.482e+01 
R942t299 n943 n300 R=2.905e+00 
R942t221 n943 n222 R=4.219e+00 
R947t521 n948 n522 R=2.881e+01 
R947t466 n948 n467 R=3.590e+01 
R948t437 n949 n438 R=7.427e+00 
R950t559 n951 n560 R=2.380e+01 
R954t946 n955 n947 R=6.701e+01 
R955t809 n956 n810 R=1.306e+01 
R955t462 n956 n463 R=2.883e+00 
R957t351 n958 n352 R=4.871e+00 
R960t855 n961 n856 R=2.704e+00 
R961t440 n962 n441 R=1.238e+01 
R961t732 n962 n733 R=4.204e+00 
R967t707 n968 n708 R=2.579e+01 
R967t623 n968 n624 R=3.121e+00 
R968t608 n969 n609 R=4.385e+01 
R968t444 n969 n445 R=1.972e+01 
R969t737 n970 n738 R=7.403e+00 
R969t771 n970 n772 R=5.955e+00 
R970t4 n971 n5 R=8.064e+01 
R971t953 n972 n954 R=4.335e+01 
R972t139 n973 n140 R=7.785e+00 
R972t820 n973 n821 R=7.165e+00 
R973t324 n974 n325 R=4.259e+00 
R974t576 n975 n577 R=2.834e+00 
R975t889 n976 n890 R=3.081e+00 
R975t56 n976 n57 R=4.909e+01 
R976t76 n977 n77 R=4.228e+00 
R977t575 n978 n576 R=6.963e+00 
R977t393 n978 n394 R=1.062e+01 
R977t709 n978 n710 R=3.419e+01 
R979t860 n980 n861 R=5.681e+00 
R981t586 n982 n587 R=1.628e+01 
R984t248 n985 n249 R=5.548e+00 
R985t251 n986 n252 R=5.061e+01 
R987t399 n988 n400 R=6.540e+00 
R988t472 n989 n473 R=1.906e+01 
R990t943 n991 n944 R=7.198e+00 
R993t980 n994 n981 R=1.111e+01 
R995t461 n996 n462 R=2.307e+01 
R998t76 n999 n77 R=1.152e+01 
R998t456 n999 n457 R=9.249e+00 
R999t688 n1000 n689 R=2.265e+00 
R999t470 n1000 n471 R=1.255e+01 
R999t813 n1000 n814 R=5.391e+01 
R1005t388 n1006 n389 R=9.503e+01 
R1005t319 n1006 n320 R=3.721e+01 
R1006t972 n1007 n973 R=1.012e+01 
R1006t820 n1007 n821 R=1.092e+01 
R1007t630 n1008 n631 R=4.278e+01 
R1011t395 n1012 n396 R=2.367e+00 
R1015t11 n1016 n12 R=3.896e+00 
R1016t389 n1017 n390 R=9.383e+00 
R1016t582 n1017 n583 R=4.880e+00 
R1017t602 n1018 n603 R=7.792e+00 
R1018t992 n1019 n993 R=5.076e+00 
R1019t629 n1020 n630 R=1.764e+01 
R1019t72 n1020 n73 R=6.919e+00 
R1020t638 n1021 n639 R=6.038e+01 
R1022t206 n1023 n207 R=1.097e+01 
R1023t965 n1024 n966 R=1.192e+01 
R1026t226 n1027 n227 R=8.965e+00 
R1029t803 n1030 n804 R=4.633e+00 
R1036t1024 n1037 n1025 R=7.309e+00 
R1039t674 n1040 n675 R=4.667e+00 
R1040t490 n1041 n491 R=8.968e+00 
R1042t177 n1043 n178 R=4.626e+00 
R1044t403 n1045 n404 R=4.836e+00 
R1045t21 n1046 n22 R=5.660e+00 
R1046t408 n1047 n409 R=1.379e+01 
R1048t746 n1049 n747 R=3.406e+00 
R1048t168 n1049 n169 R=2.454e+00 
R1050t282 n1051 n283 R=9.268e+00 
R1051t501 n1052 n502 R=7.971e+00 
R1060t244 n1061 n245 R=1.182e+01 
R1060t783 n1061 n784 R=2.522e+00 
R1062t986 n1063 n987 R=5.933e+00 
R1066t333 n1067 n334 R=7.226e+00 
R1067t396 n1068 n397 R=4.407e+01 
R1067t503 n1068 n504 R=2.107e+01 
R1070t837 n1071 n838 R=5.102e+00 
R1070t537 n1071 n538 R=4.297e+00 
R1072t16 n1073 n17 R=3.283e+00 
R1074t980 n1075 n981 R=9.300e+00 
R1074t747 n1075 n748 R=2.194e+01 
R1075t333 n1076 n334 R=8.268e+00 
R1075t1066 n1076 n1067 R=5.192e+00 
R1077t547 n1078 n548 R=2.820e+00 
R1079t696 n1080 n697 R=8.429e+00 
R1081t542 n1082 n543 R=6.375e+02 
R1085t700 n1086 n701 R=3.403e+00 
R1086t1024 n1087 n1025 R=3.928e+00 
R1089t270 n1090 n271 R=3.660e+00 
R1090t488 n1091 n489 R=7.275e+00 
R1091t698 n1092 n699 R=1.260e+01 
R1091t497 n1092 n498 R=5.276e+00 
R1094t698 n1095 n699 R=2.795e+01 
R1095t605 n1096 n606 R=1.552e+01 
R1097t78 n1098 n79 R=9.225e+00 
R1097t1021 n1098 n1022 R=1.009e+01 
R1098t391 n1099 n392 R=1.456e+01 
R1099t29 n1100 n30 R=3.398e+01 
R1101t238 n1102 n239 R=2.447e+01 
R1102t895 n1103 n896 R=1.733e+00 
R1105t379 n1106 n380 R=4.943e+00 
R1107t1058 n1108 n1059 R=1.884e+01 
R1119t614 n1120 n615 R=4.542e+00 
R1123t925 n1124 n926 R=1.307e+02 
R1128t390 n1129 n391 R=5.975e+01 
R1128t879 n1129 n880 R=4.397e+01 
R1129t644 n1130 n645 R=8.780e+00 
R1130t164 n1131 n165 R=2.301e+02 
R1134t116 n1135 n117 R=2.606e+00 
R1136t399 n1137 n400 R=4.376e+00 
R1136t987 n1137 n988 R=1.017e+02 
R1137t587 n1138 n588 R=2.544e+01 
R1137t596 n1138 n597 R=6.088e+00 
R1140t678 n1141 n679 R=3.203e+01 
R1143t538 n1144 n539 R=1.105e+01 
R1144t136 n1145 n137 R=2.998e+00 
R1149t845 n1150 n846 R=8.966e+00 
R1149t807 n1150 n808 R=8.867e+00 
R1150t1115 n1151 n1116 R=4.443e+00 
R1153t234 n1154 n235 R=2.595e+03 
R1153t170 n1154 n171 R=1.131e+01 
R1154t1037 n1 n1038 R=6.330e+00 
R1155t1064 n1156 n1065 R=7.034e+00 
R1158t12 n1159 n13 R=1.013e+01 
R1160t332 n1161 n333 R=3.740e+00 
R1161t692 n1162 n1 R=1.458e+01 
R1161t706 n1162 n707 R=5.388e+00 
R1163t770 n1164 n771 R=4.100e+01 
R1164t290 n1165 n291 R=2.046e+01 
R1165t184 n1166 n185 R=3.832e+00 
R1165t193 n1166 n194 R=1.311e+01 
R1166t334 n1167 n335 R=2.427e+00 
R1168t1112 n1169 n1113 R=6.952e+00 
R1169t499 n1170 n500 R=3.564e+00 
R1170t269 n1171 n270 R=2.531e+00 
R1171t884 n1172 n885 R=1.021e+01 
R1172t335 n1173 n336 R=3.465e+01 
R1173t921 n1174 n922 R=2.368e+01 
R1174t1124 n1175 n1125 R=5.561e+00 
R1175t417 n1176 n418 R=4.586e+00 
R1176t881 n1177 n882 R=1.998e+01 
R1178t438 n1179 n439 R=2.606e+01 
R1178t549 n1179 n550 R=1.052e+01 
R1180t117 n1181 n118 R=5.025e+00 
R1181t1020 n1182 n1021 R=2.468e+01 
R1181t638 n1182 n639 R=3.434e+00 
R1185t493 n1186 n494 R=3.804e+00 
R1186t530 n1187 n531 R=3.795e+01 
R1188t1187 n1189 n1188 R=1.484e+01 
R1191t820 n1192 n821 R=2.657e+00 
R1192t1021 n1193 n1022 R=4.533e+00 
R1192t1097 n1193 n1098 R=4.614e+00 
R1194t309 n1195 n310 R=5.455e+00 
R1195t1084 n1196 n1085 R=1.736e+01 
R1197t1190 n1198 n1191 R=1.532e+01 
R1199t107 n1200 n108 R=7.722e+00 
R1200t281 n1201 n282 R=3.642e+00 
R1202t541 n1203 n542 R=5.490e+00 
R1204t1122 n1205 n1123 R=2.075e+01 
R1208t614 n1209 n615 R=5.491e+00 
R1208t1119 n1209 n1120 R=6.841e+00 
R1209t338 n1210 n339 R=5.413e+00 
R1210t791 n1211 n792 R=5.316e+00 
R1212t704 n1213 n705 R=5.208e+00 
R1212t363 n1213 n364 R=3.750e+00 
R1213t21 n1214 n22 R=1.727e+01 
R1213t1045 n1214 n1046 R=3.766e+00 
R1214t98 n1215 n99 R=5.272e+00 
R1215t1039 n1216 n1040 R=1.039e+01 
R1218t1056 n1219 n1057 R=1.824e+02 
R1218t746 n1219 n747 R=8.400e+00 
R1220t559 n1221 n560 R=4.308e+00 
R1220t667 n1221 n668 R=1.645e+02 
R1222t989 n1223 n990 R=5.080e+00 
R1223t478 n1224 n479 R=1.374e+01 
R1223t719 n1224 n720 R=1.148e+01 
R1224t433 n1225 n434 R=1.130e+01 
R1224t806 n1225 n807 R=8.428e+00 
R1225t953 n1226 n954 R=1.301e+00 
R1225t971 n1226 n972 R=1.148e+03 
R1226t705 n1227 n706 R=1.191e+01 
R1226t149 n1227 n150 R=9.347e+00 
R1227t1145 n1228 n1146 R=2.358e+01 
R1230t939 n1231 n940 R=9.189e+00 
R1231t857 n1232 n858 R=2.345e+00 
R1236t160 n1237 n161 R=2.891e+00 
R1238t290 n1239 n291 R=2.106e+01 
R1239t580 n1240 n581 R=5.923e+00 
R1240t1034 n1241 n1035 R=1.061e+02 
R1241t511 n1242 n512 R=4.511e+00 
R1241t557 n1242 n558 R=2.407e+00 
R1244t634 n1245 n635 R=7.713e+00 
R1248t718 n1249 n719 R=2.684e+00 
R1251t335 n1252 n336 R=1.803e+01 
R1253t804 n1254 n805 R=6.935e+00 
R1253t199 n1254 n200 R=4.222e+00 
R1253t373 n1254 n374 R=2.412e+01 
R1254t599 n1255 n600 R=2.853e+01 
R1254t915 n1255 n916 R=4.565e+00 
R1257t574 n1258 n575 R=1.344e+01 
R1258t124 n1259 n125 R=7.151e+00 
R1260t1249 n1261 n1250 R=1.473e+01 
R1261t225 n1262 n226 R=1.299e+01 
R1264t514 n1265 n515 R=4.929e+00 
R1265t522 n1266 n523 R=3.668e+00 
R1267t1242 n1268 n1243 R=2.553e+00 
R1267t76 n1268 n77 R=1.198e+01 
R1270t268 n1271 n269 R=2.450e+01 
R1272t1215 n1273 n1216 R=9.048e+00 
R1272t674 n1273 n675 R=5.354e+00 
R1272t1039 n1273 n1040 R=1.256e+01 
R1273t327 n1 n328 R=7.685e+01 
R1275t376 n1276 n377 R=2.622e+00 
R1275t39 n1276 n40 R=1.420e+01 
R1277t781 n1278 n782 R=3.604e+01 
R1277t844 n1278 n845 R=5.260e+00 
R1278t792 n1279 n793 R=2.585e+01 
R1278t1264 n1279 n1265 R=2.592e+01 
R1278t713 n1279 n714 R=5.253e+00 
R1279t614 n1280 n615 R=1.892e+01 
R1279t791 n1280 n792 R=4.344e+00 
R1281t738 n1282 n739 R=1.070e+01 
R1282t793 n1283 n794 R=2.438e+00 
R1283t916 n1284 n917 R=8.910e+00 
R1286t90 n1287 n91 R=3.434e+00 
R1287t892 n1288 n893 R=6.236e+00 
R1287t409 n1288 n410 R=5.483e+00 
R1288t345 n1289 n346 R=4.201e+02 
R1288t83 n1289 n84 R=1.382e+01 
R1291t104 n1292 n105 R=1.035e+01 
R1293t472 n1294 n473 R=5.658e+00 
R1294t855 n1295 n856 R=2.852e+00 
R1294t1221 n1295 n1222 R=9.580e+01 
R1295t786 n1296 n787 R=5.265e+00 
R1295t1031 n1296 n1032 R=3.172e+00 
R1296t330 n1297 n331 R=5.103e+00 
R1298t788 n1299 n789 R=5.735e+00 
R1299t378 n1300 n379 R=7.018e+01 
R1300t1210 n1301 n1211 R=9.793e+00 
R1301t352 n1302 n353 R=2.507e+02 
R1306t1004 n1307 n1005 R=8.410e+01 
R1308t731 n1309 n732 R=7.700e+00 
R1311t730 n1312 n731 R=1.507e+01 
R1312t220 n1313 n221 R=1.939e+00 
R1313t236 n1314 n237 R=2.902e+01 
R1313t158 n1314 n159 R=2.813e+00 
R1314t959 n1315 n960 R=4.304e+00 
R1316t162 n1317 n163 R=1.635e+02 
R1316t736 n1317 n737 R=5.415e+00 
R1316t878 n1317 n879 R=6.341e+00 
R1317t892 n1318 n893 R=1.028e+01 
R1320t178 n1321 n179 R=8.542e+00 
R1324t800 n1325 n801 R=9.401e+00 
R1326t665 n1327 n666 R=1.303e+02 
R1326t482 n1327 n483 R=1.153e+01 
R1326t993 n1327 n994 R=5.513e+00 
R1328t735 n1329 n736 R=4.547e+00 
R1329t1058 n1330 n1059 R=1.079e+02 
R1329t1107 n1330 n1108 R=4.194e+00 
R1330t1300 n1331 n1301 R=3.577e+00 
R1330t1279 n1331 n1280 R=1.131e+01 
R1330t791 n1331 n792 R=1.333e+01 
R1330t1210 n1331 n1211 R=8.909e+00 
R1331t1092 n1332 n1093 R=6.530e+00 
R1331t136 n1332 n137 R=2.493e+01 
R1331t1144 n1332 n1145 R=2.273e+02 
R1334t755 n1335 n756 R=3.573e+00 
R1335t988 n1336 n989 R=1.888e+01 
R1337t1277 n1338 n1278 R=1.420e+01 
R1338t23 n1339 n24 R=9.786e+00 
R1338t471 n1339 n472 R=4.256e+00 
R1340t675 n1341 n676 R=3.441e+01 
R1340t1164 n1341 n1165 R=1.009e+02 
R1344t740 n1345 n741 R=4.295e+00 
R1346t784 n1347 n785 R=5.394e+00 
R1347t1319 n1348 n1320 R=8.230e+00 
R1348t839 n1349 n840 R=1.095e+01 
R1348t266 n1349 n267 R=3.408e+01 
R1349t258 n1350 n259 R=3.392e+01 
R1350t872 n1351 n873 R=1.593e+01 
R1350t951 n1351 n952 R=7.668e+00 
R1352t454 n1353 n455 R=3.622e+00 
R1352t133 n1353 n134 R=2.950e+00 
R1353t60 n1354 n61 R=1.506e+01 
R1353t920 n1354 n921 R=1.306e+01 
R1354t1000 n1355 n1001 R=1.864e+01 
R1355t113 n1356 n114 R=3.269e+01 
R1355t585 n1356 n586 R=3.465e+01 
R1356t690 n1357 n691 R=1.402e+01 
R1356t259 n1357 n260 R=1.016e+01 
R1360t423 n1361 n424 R=4.065e+01 
R1365t392 n1366 n393 R=4.101e+01 
R1366t741 n1367 n742 R=2.277e+00 
R1367t1237 n1368 n1238 R=3.666e+00 
R1370t1035 n1371 n1036 R=3.418e+00 
R1372t695 n1373 n696 R=1.554e+01 
R1372t71 n1373 n72 R=4.982e+01 
R1374t68 n1375 n69 R=9.854e+00 
R1374t1311 n1375 n1312 R=6.302e+00 
R1374t271 n1375 n272 R=1.743e+01 
R1374t119 n1375 n120 R=7.270e+00 
R1378t1052 n1379 n1053 R=2.618e+00 
R1380t71 n1381 n72 R=1.418e+01 
R1382t619 n1383 n620 R=2.589e+00 
R1384t654 n1385 n655 R=4.300e+01 
R1386t730 n1387 n731 R=4.212e+00 
R1387t22 n1388 n23 R=7.022e+00 
R1388t1178 n1389 n1179 R=7.717e+01 
R1388t1145 n1389 n1146 R=4.754e+01 
R1389t1104 n1390 n1105 R=2.427e+01 
R1390t494 n1391 n495 R=4.569e+01 
R1392t976 n1393 n977 R=4.207e+00 
R1393t547 n1394 n548 R=7.374e+00 
R1393t1077 n1394 n1078 R=2.267e+01 
R1395t1298 n1396 n1299 R=2.529e+00 
R1396t796 n1397 n797 R=1.535e+01 
R1396t636 n1397 n637 R=5.538e+00 
R1402t224 n1403 n225 R=6.068e+00 
R1405t275 n1406 n276 R=1.014e+01 
R1405t59 n1406 n60 R=9.736e+00 
R1406t1206 n1407 n1207 R=9.575e+00 
R1409t1088 n1410 n1089 R=9.547e+00 
R1410t253 n1411 n254 R=4.596e+00 
R1412t960 n1413 n961 R=1.064e+01 
R1413t48 n1414 n49 R=1.016e+01 
R1413t600 n1414 n601 R=1.765e+01 
R1413t15 n1414 n16 R=3.641e+00 
R1414t696 n1415 n697 R=5.594e+00 
R1415t230 n1416 n231 R=7.126e+00 
R1418t545 n1419 n546 R=1.101e+02 
R1418t697 n1419 n698 R=8.838e+00 
R1418t633 n1419 n634 R=8.233e+00 
R1420t1244 n1421 n1245 R=2.213e+01 
R1420t634 n1421 n635 R=7.083e+01 
R1421t1415 n1422 n1416 R=5.754e+00 
R1424t584 n1425 n585 R=1.416e+01 
R1424t77 n1425 n78 R=2.342e+00 
R1426t866 n1427 n867 R=9.381e+00 
R1429t463 n1430 n464 R=4.073e+00 
R1430t938 n1431 n939 R=3.702e+00 
R1431t357 n1432 n358 R=9.558e+00 
R1432t1064 n1433 n1065 R=2.783e+00 
R1433t1265 n1434 n1266 R=5.516e+00 
R1433t1030 n1434 n1031 R=1.486e+01 
R1434t790 n1435 n791 R=4.169e+00 
R1434t1113 n1435 n1114 R=3.187e+00 
R1438t1142 n1439 n1143 R=8.997e+00 
R1439t402 n1440 n403 R=2.181e+00 
R1439t844 n1440 n845 R=1.044e+01 
R1439t1277 n1440 n1278 R=7.215e+01 
R1439t1337 n1440 n1338 R=2.464e+01 
R1441t1427 n1442 n1428 R=3.845e+00 
R1442t933 n1443 n934 R=7.298e+00 
R1443t1409 n1444 n1410 R=3.733e+01 
R1443t1210 n1444 n1211 R=7.986e+00 
R1443t791 n1444 n792 R=1.668e+01 
R1444t653 n1445 n654 R=3.136e+01 
R1445t725 n1446 n726 R=9.963e+00 
R1446t763 n1447 n764 R=9.883e+00 
R1446t693 n1447 n694 R=5.142e+01 
R1447t795 n1448 n796 R=3.719e+00 
R1448t430 n1449 n431 R=8.299e+00 
R1448t434 n1449 n435 R=3.625e+00 
R1449t264 n1450 n265 R=1.066e+01 
R1449t637 n1450 n638 R=9.612e+00 
R1451t83 n1452 n84 R=5.852e+01 
R1451t241 n1452 n242 R=2.361e+01 
R1451t5 n1452 n6 R=1.160e+01 
R1452t196 n1453 n197 R=4.411e+00 
R1453t935 n1454 n936 R=1.840e+00 
R1453t340 n1454 n341 R=3.534e+00 
R1454t293 n1455 n294 R=5.252e+01 
R1457t429 n1458 n430 R=1.431e+01 
R1457t800 n1458 n801 R=1.306e+01 
R1457t1324 n1458 n1325 R=5.910e+00 
R1458t1437 n1459 n1438 R=9.483e+00 
R1460t208 n1461 n209 R=7.895e+00 
R1461t1278 n1462 n1279 R=5.746e+00 
R1461t713 n1462 n714 R=2.263e+01 
R1464t376 n1465 n377 R=2.555e+02 
R1464t701 n1465 n702 R=2.987e+00 
R1464t39 n1465 n40 R=8.211e+00 
R1465t486 n1466 n487 R=6.397e+00 
R1466t102 n1467 n103 R=4.234e+00 
R1467t1002 n1468 n1003 R=7.907e+00 
R1467t547 n1468 n548 R=3.398e+01 
R1467t1415 n1468 n1416 R=1.076e+02 
R1467t1421 n1468 n1422 R=3.803e+00 
R1468t1116 n1469 n1117 R=1.958e+01 
R1469t1128 n1470 n1129 R=1.601e+01 
R1470t169 n1471 n170 R=2.040e+01 
R1471t1175 n1472 n1176 R=2.435e+01 
R1471t417 n1472 n418 R=2.860e+01 
R1475t73 n1476 n74 R=1.827e+01 
R1476t352 n1477 n353 R=6.890e+00 
R1478t420 n1479 n421 R=1.235e+01 
R1480t1360 n1481 n1361 R=7.817e+01 
R1481t1033 n1482 n1034 R=1.653e+01 
R1481t207 n1482 n208 R=1.889e+01 
R1482t56 n1483 n57 R=3.477e+00 
R1482t400 n1483 n401 R=3.941e+00 
R1483t461 n1484 n462 R=7.057e+01 
R1484t1383 n1 n1384 R=1.631e+01 
R1485t280 n1486 n281 R=8.498e+00 
R1486t1391 n1487 n1392 R=4.542e+00 
R1488t1159 n1489 n1160 R=6.572e+00 
R1489t1430 n1490 n1431 R=2.336e+01 
R1494t465 n1495 n466 R=1.015e+02 
R1494t297 n1495 n298 R=6.736e+01 
R1497t517 n1498 n518 R=7.530e+00 
R1497t261 n1498 n262 R=1.042e+02 
R1499t642 n1500 n643 R=3.718e+00 
R1501t803 n1502 n804 R=5.728e+00 
R1501t1029 n1502 n1030 R=6.997e+00 
R1504t197 n1505 n198 R=5.275e+00 
R1504t647 n1505 n648 R=9.676e+00 
R1506t124 n1507 n125 R=4.967e+00 
R1508t516 n1509 n517 R=2.751e+01 
R1509t777 n1510 n778 R=1.242e+01 
R1509t1417 n1510 n1418 R=1.032e+01 
R1509t211 n1510 n212 R=1.225e+01 
R1510t572 n1511 n573 R=2.885e+01 
R1515t1250 n1516 n1251 R=5.005e+00 
R1516t316 n1517 n317 R=7.746e+00 
R1518t855 n1519 n856 R=1.104e+03 
R1518t960 n1519 n961 R=6.118e+01 
R1518t1465 n1519 n1466 R=5.065e+03 
R1519t1416 n1520 n1417 R=2.889e+00 
R1519t877 n1520 n878 R=2.077e+02 
R1519t631 n1520 n632 R=5.631e+02 
R1525t716 n1526 n717 R=1.248e+01 
R1525t1194 n1526 n1195 R=9.305e+00 
R1525t145 n1526 n146 R=2.721e+00 
R1527t1107 n1528 n1108 R=2.251e+00 
R1528t145 n1529 n146 R=5.627e+00 
R1529t959 n1530 n960 R=1.941e+01 
R1529t1314 n1530 n1315 R=3.516e+00 
R1530t787 n1531 n788 R=5.240e+00 
R1530t1069 n1531 n1070 R=3.475e+00 
R1533t1023 n1534 n1024 R=2.896e+01 
R1533t965 n1534 n966 R=2.340e+00 
R1534t561 n1535 n562 R=2.863e+00 
R1535t261 n1536 n262 R=2.726e+00 
R1536t802 n1537 n803 R=2.476e+00 
R1541t470 n1542 n471 R=4.282e+00 
R1542t1495 n1543 n1496 R=5.120e+00 
R1543t1348 n1544 n1349 R=7.495e+00 
R1544t53 n1545 n54 R=1.193e+01 
R1545t466 n1546 n467 R=6.111e+00 
R1545t947 n1546 n948 R=8.296e+00 
R1546t430 n1547 n431 R=9.018e+00 
R1546t147 n1547 n148 R=3.266e+00 
R1549t1536 n1550 n1537 R=2.963e+02 
R1549t720 n1550 n721 R=5.861e+01 
R1549t802 n1550 n803 R=1.644e+01 
R1550t941 n1551 n942 R=9.369e+00 
R1550t101 n1551 n102 R=9.146e+00 
R1551t367 n1552 n368 R=2.534e+01 
R1552t1201 n1553 n1 R=6.010e+00 
R1552t398 n1553 n1 R=9.026e+00 
R1553t286 n1554 n287 R=8.666e+00 
R1556t214 n1557 n215 R=4.788e+00 
R1557t435 n1558 n436 R=1.798e+00 
R1557t919 n1558 n920 R=2.853e+01 
R1557t861 n1558 n862 R=1.034e+01 
R1558t265 n1559 n266 R=9.087e+00 
R1560t245 n1561 n246 R=1.482e+01 
R1562t810 n1563 n811 R=4.905e+00 
R1563t1493 n1564 n1494 R=1.011e+02 
R1563t728 n1564 n729 R=1.002e+01 
R1564t180 n1565 n181 R=3.781e+00 
R1565t753 n1566 n754 R=5.727e+00 
R1565t1361 n1566 n1362 R=4.256e+00 
R1566t1123 n1567 n1124 R=2.730e+01 
R1567t241 n1568 n242 R=5.358e+00 
R1567t660 n1568 n661 R=1.376e+01 
R1567t1451 n1568 n1452 R=5.225e+00 
R1567t1056 n1568 n1057 R=1.894e+01 
R1568t982 n1569 n983 R=2.542e+01 
R1569t837 n1570 n838 R=5.174e+00 
R1572t1388 n1573 n1389 R=1.107e+01 
R1573t369 n1574 n370 R=2.071e+01 
R1573t190 n1574 n191 R=2.217e+00 
R1574t835 n1575 n836 R=5.388e+00 
R1574t931 n1575 n932 R=1.064e+02 
R1576t695 n1577 n696 R=1.332e+01 
R1576t912 n1577 n913 R=1.196e+01 
R1578t312 n1579 n313 R=1.683e+01 
R1578t166 n1579 n167 R=8.431e+00 
R1579t766 n1580 n767 R=5.570e+00 
R1580t232 n1581 n233 R=2.408e+01 
R1583t1400 n1584 n1401 R=1.030e+01 
R1584t74 n1585 n75 R=2.762e+00 
R1586t1584 n1587 n1585 R=7.716e+01 
R1586t832 n1587 n833 R=1.210e+01 
R1587t742 n1588 n743 R=5.486e+00 
R1590t586 n1591 n587 R=2.159e+01 
R1591t1392 n1592 n1393 R=4.176e+00 
R1592t972 n1593 n973 R=1.482e+01 
R1592t820 n1593 n821 R=3.337e+01 
R1592t1191 n1593 n1192 R=9.665e+00 
R1592t681 n1593 n682 R=6.742e+01 
R1593t1490 n1594 n1491 R=2.066e+00 
R1594t469 n1595 n470 R=6.249e+00 
R1595t280 n1596 n281 R=2.680e+01 
R1595t1485 n1596 n1486 R=2.972e+00 
R1595t698 n1596 n699 R=6.989e+00 
R1597t69 n1598 n70 R=3.844e+01 
R1598t207 n1599 n208 R=9.994e+00 
R1601t873 n1602 n874 R=3.719e+01 
R1601t824 n1602 n825 R=2.126e+00 
R1603t234 n1604 n235 R=1.284e+01 
R1605t334 n1606 n335 R=6.532e+00 
R1606t1244 n1607 n1245 R=5.039e+00 
R1609t1531 n1610 n1532 R=6.537e+00 
R1610t1591 n1611 n1592 R=3.270e+00 
R1612t573 n1613 n574 R=1.208e+01 
R1615t1472 n1616 n1473 R=1.706e+01 
R1616t1360 n1617 n1361 R=2.058e+01 
R1622t1607 n1623 n1608 R=2.122e+01 
R1623t1187 n1624 n1188 R=7.955e+00 
R1623t1188 n1624 n1189 R=1.388e+01 
R1626t1419 n1627 n1420 R=9.715e+00 
R1627t1240 n1628 n1241 R=3.763e+01 
R1628t1094 n1629 n1095 R=4.290e+00 
R1629t167 n1630 n168 R=2.210e+00 
R1629t361 n1630 n362 R=3.423e+00 
R1630t629 n1631 n630 R=7.866e+00 
R1631t98 n1632 n99 R=1.261e+01 
R1631t1214 n1632 n1215 R=8.748e+00 
R1631t302 n1632 n303 R=1.272e+01 
R1634t865 n1635 n866 R=4.691e+00 
R1634t537 n1635 n538 R=3.087e+01 
R1634t861 n1635 n862 R=4.761e+00 
R1635t644 n1636 n645 R=5.029e+01 
R1635t1617 n1636 n1618 R=6.585e+00 
R1635t439 n1636 n440 R=3.038e+00 
R1636t340 n1637 n341 R=7.100e+00 
R1636t1453 n1637 n1454 R=6.256e+01 
R1636t935 n1637 n936 R=7.698e+01 
R1637t1200 n1638 n1201 R=3.625e+01 
R1639t483 n1640 n1 R=1.312e+01 
R1640t1191 n1641 n1192 R=9.783e+00 
R1640t681 n1641 n682 R=1.003e+01 
R1640t1592 n1641 n1593 R=3.381e+00 
R1642t328 n1643 n329 R=7.435e+01 
R1643t126 n1644 n127 R=2.878e+00 
R1643t1061 n1644 n1062 R=6.239e+00 
R1644t317 n1645 n318 R=3.664e+01 
R1645t678 n1646 n679 R=1.453e+01 
R1646t986 n1647 n987 R=2.166e+01 
R1646t1062 n1647 n1063 R=4.227e+00 
R1648t1110 n1649 n1111 R=3.070e+00 
R1648t1096 n1649 n1097 R=5.485e+00 
R1649t788 n1650 n789 R=6.844e+00 
R1650t1 n1651 n2 R=2.365e+01 
R1651t440 n1652 n441 R=3.871e+01 
R1655t273 n1656 n274 R=5.897e+00 
R1658t1239 n1659 n1240 R=5.913e+01 
R1658t927 n1659 n928 R=1.523e+00 
R1661t1597 n1662 n1598 R=9.582e+01 
R1662t353 n1663 n354 R=6.226e+00 
R1666t1019 n1667 n1020 R=7.745e+00 
R1667t717 n1668 n718 R=5.319e+00 
R1667t1106 n1668 n1107 R=2.022e+00 
R1669t1618 n1670 n1619 R=1.550e+00 
R1673t1627 n1674 n1628 R=5.623e+00 
R1673t114 n1674 n115 R=3.561e+01 
R1675t655 n1676 n656 R=1.144e+02 
R1676t1657 n1677 n1658 R=1.709e+01 
R1677t1211 n1678 n1212 R=3.709e+00 
R1677t317 n1678 n318 R=1.338e+01 
R1677t1548 n1678 n1549 R=3.362e+01 
R1680t1604 n1681 n1605 R=2.309e+00 
R1680t362 n1681 n363 R=2.207e+00 
R1681t1289 n1682 n1290 R=6.136e+01 
R1682t1147 n1683 n1148 R=3.611e+00 
R1682t484 n1683 n485 R=1.212e+01 
R1683t509 n1684 n510 R=9.532e+00 
R1683t769 n1684 n770 R=4.651e+00 
R1684t1558 n1685 n1559 R=2.310e+01 
R1685t1575 n1686 n1576 R=9.080e+00 
R1687t866 n1688 n867 R=1.056e+01 
R1688t40 n1689 n41 R=1.482e+01 
R1689t77 n1690 n78 R=1.513e+02 
R1691t373 n1692 n374 R=2.492e+01 
R1691t322 n1692 n323 R=1.123e+02 
R1694t522 n1695 n523 R=5.759e+00 
R1694t1265 n1695 n1266 R=4.693e+01 
R1694t1433 n1695 n1434 R=2.860e+01 
R1694t57 n1695 n58 R=2.449e+00 
R1695t283 n1696 n284 R=7.407e+00 
R1697t1220 n1698 n1221 R=1.939e+02 
R1698t1315 n1699 n1316 R=2.603e+00 
R1699t41 n1700 n42 R=1.240e+01 
R1702t499 n1703 n500 R=7.265e+00 
R1702t1169 n1703 n1170 R=4.148e+00 
R1703t1183 n1704 n1184 R=4.409e+00 
R1706t1290 n1707 n1291 R=9.622e+00 
R1707t587 n1708 n588 R=2.416e+02 
R1708t1626 n1 n1627 R=1.163e+02 
R1709t85 n1710 n86 R=1.191e+01 
R1709t1456 n1710 n1457 R=1.326e+01 
R1710t326 n1711 n327 R=6.625e+00 
R1710t486 n1711 n487 R=9.342e+00 
R1713t1401 n1714 n1402 R=6.984e+00 
R1714t1437 n1715 n1438 R=3.435e+01 
R1717t487 n1718 n488 R=7.878e+00 
R1718t1332 n1719 n1333 R=5.086e+00 
R1721t1679 n1722 n1680 R=7.815e+00 
R1722t1503 n1723 n1504 R=2.925e+00 
R1724t466 n1725 n467 R=3.227e+00 
R1724t521 n1725 n522 R=6.855e+00 
R1724t947 n1725 n948 R=2.649e+00 
R1725t737 n1726 n738 R=5.443e+01 
R1725t1700 n1726 n1701 R=7.415e+00 
R1725t404 n1726 n405 R=7.844e+00 
R1727t106 n1 n107 R=8.996e+01 
R1728t692 n1729 n1 R=5.121e+00 
R1728t1161 n1729 n1162 R=7.857e+00 
R1730t794 n1731 n795 R=3.801e+00 
R1731t966 n1732 n967 R=8.120e+00 
R1732t985 n1733 n986 R=4.187e+00 
R1733t276 n1734 n277 R=3.097e+00 
R1733t1054 n1734 n1055 R=1.436e+02 
R1734t310 n1735 n311 R=1.546e+01 
R1735t543 n1736 n544 R=7.487e+00 
R1736t994 n1737 n995 R=3.205e+00 
R1738t1108 n1739 n1109 R=6.935e+00 
R1739t1545 n1740 n1546 R=5.512e+01 
R1739t339 n1740 n340 R=1.587e+01 
R1740t105 n1741 n106 R=2.846e+00 
R1742t1224 n1743 n1225 R=1.592e+01 
R1744t79 n1745 n80 R=4.289e+00 
R1746t1502 n1747 n1503 R=1.742e+00 
R1748t39 n1749 n40 R=3.819e+01 
R1748t1454 n1749 n1455 R=2.181e+00 
R1751t249 n1752 n250 R=1.351e+01 
R1753t505 n1754 n506 R=2.690e+00 
R1754t1522 n1755 n1523 R=3.029e+01 
R1756t1027 n1757 n1028 R=6.234e+00 
R1758t1603 n1759 n1604 R=1.030e+01 
R1758t1153 n1759 n1154 R=1.969e+01 
R1758t1414 n1759 n1415 R=2.048e+00 
R1758t696 n1759 n697 R=4.003e+01 
R1759t1172 n1760 n1173 R=9.806e+00 
R1760t1146 n1761 n1147 R=1.975e+01 
R1760t1502 n1761 n1503 R=4.371e+01 
R1760t1746 n1761 n1747 R=3.895e+01 
R1762t518 n1763 n519 R=2.782e+01 
R1762t797 n1763 n798 R=1.962e+01 
R1762t227 n1763 n228 R=2.579e+01 
R1766t1638 n1767 n1639 R=8.099e+00 
R1766t1127 n1767 n1128 R=7.017e+01 
R1767t510 n1768 n511 R=1.963e+01 
R1767t123 n1768 n124 R=1.650e+02 
R1768t275 n1769 n276 R=1.120e+01 
R1768t48 n1769 n49 R=3.574e+00 
R1768t1413 n1769 n1414 R=1.155e+01 
R1768t600 n1769 n601 R=9.663e+00 
R1769t848 n1770 n849 R=4.035e+00 
R1770t1471 n1771 n1472 R=1.335e+02 
R1771t1194 n1772 n1195 R=1.224e+01 
R1771t1525 n1772 n1526 R=2.750e+01 
R1771t145 n1772 n146 R=1.531e+01 
R1771t309 n1772 n310 R=9.292e+00 
R1772t90 n1773 n91 R=8.244e+00 
R1772t1286 n1773 n1287 R=2.894e+01 
R1772t162 n1773 n163 R=9.915e+00 
R1773t1438 n1774 n1439 R=4.258e+00 
R1773t1237 n1774 n1238 R=4.833e+00 
R1773t1142 n1774 n1143 R=2.505e+01 
R1774t1637 n1775 n1638 R=3.650e+00 
R1775t201 n1776 n202 R=2.714e+00 
R1777t176 n1778 n177 R=8.323e+00 
R1780t215 n1781 n216 R=1.333e+01 
R1784t794 n1785 n795 R=8.881e+00 
R1785t1005 n1786 n1006 R=1.155e+01 
R1790t1690 n1791 n1691 R=5.789e+00 
R1791t779 n1792 n780 R=6.921e+00 
R1791t1083 n1792 n1084 R=1.959e+01 
R1791t1343 n1792 n1344 R=4.453e+00 
R1792t779 n1793 n780 R=1.788e+01 
R1792t1343 n1793 n1344 R=6.815e+00 
R1792t1791 n1793 n1792 R=2.086e+01 
R1793t126 n1794 n127 R=2.849e+01 
R1793t1643 n1794 n1644 R=1.136e+01 
R1795t1173 n1796 n1174 R=3.381e+00 
R1796t30 n1797 n31 R=7.926e+00 
R1797t1416 n1798 n1417 R=7.971e+00 
R1797t1519 n1798 n1520 R=1.548e+02 
R1799t1615 n1800 n1616 R=4.740e+00 
R1800t1335 n1801 n1336 R=7.425e+00 
R1802t203 n1803 n204 R=2.677e+00 
R1803t1065 n1804 n1066 R=4.085e+00 
R1805t653 n1806 n654 R=1.985e+01 
R1806t1551 n1807 n1552 R=1.401e+01 
R1807t432 n1808 n433 R=5.974e+00 
R1808t765 n1809 n766 R=7.216e+00 
R1812t1645 n1813 n1646 R=7.755e+02 
R1814t1713 n1815 n1714 R=1.874e+00 
R1817t918 n1818 n919 R=6.975e+00 
R1817t1535 n1818 n1536 R=6.548e+00 
R1820t1141 n1821 n1142 R=1.190e+03 
R1821t1795 n1822 n1796 R=1.705e+01 
R1823t120 n1824 n121 R=1.013e+01 
R1825t362 n1826 n363 R=3.184e+01 
R1828t1234 n1829 n1235 R=1.982e+01 
R1828t1617 n1829 n1618 R=3.538e+00 
R1829t500 n1830 n501 R=7.355e+00 
R1829t798 n1830 n799 R=9.526e+00 
R1829t1583 n1830 n1584 R=5.316e+00 
R1832t313 n1833 n314 R=6.559e+01 
R1833t512 n1834 n513 R=3.310e+00 
R1833t782 n1834 n783 R=5.580e+00 
R1834t455 n1835 n456 R=3.974e+01 
R1836t964 n1837 n965 R=5.463e+01 
R1836t998 n1837 n999 R=4.033e+00 
R1837t955 n1838 n956 R=4.072e+00 
R1837t809 n1838 n810 R=6.203e+00 
R1839t1084 n1 n1085 R=8.940e+00 
R1840t1700 n1841 n1701 R=1.281e+01 
R1844t222 n1845 n223 R=3.552e+01 
R1845t1496 n1846 n1497 R=2.205e+00 
R1845t1066 n1846 n1067 R=4.874e+00 
R1847t1628 n1848 n1629 R=7.069e+00 
R1848t768 n1849 n769 R=3.035e+00 
R1850t1478 n1851 n1479 R=3.447e+00 
R1850t246 n1851 n247 R=5.310e+01 
R1850t420 n1851 n421 R=6.416e+00 
R1851t910 n1852 n911 R=2.057e+01 
R1852t18 n1853 n19 R=1.959e+00 
R1852t1641 n1853 n1642 R=2.368e+00 
R1853t876 n1854 n877 R=6.806e+00 
R1856t1647 n1857 n1648 R=3.408e+01 
R1858t125 n1859 n126 R=5.338e+00 
R1859t1522 n1860 n1523 R=1.582e+02 
R1860t1585 n1861 n1586 R=2.546e+00 
R1861t361 n1862 n362 R=4.522e+00 
R1861t1629 n1862 n1630 R=1.631e+01 
R1862t1263 n1863 n1264 R=6.887e+00 
R1862t338 n1863 n339 R=7.292e+00 
R1863t1624 n1864 n1625 R=1.628e+01 
R1863t223 n1864 n224 R=1.766e+01 
R1863t347 n1864 n348 R=2.593e+01 
R1864t1714 n1865 n1715 R=3.185e+01 
R1864t1437 n1865 n1438 R=3.124e+00 
R1864t1458 n1865 n1459 R=1.105e+01 
R1865t234 n1866 n235 R=7.459e+00 
R1865t1153 n1866 n1154 R=1.405e+01 
R1866t1385 n1867 n1386 R=2.494e+00 
R1867t752 n1868 n753 R=7.348e+00 
R1867t504 n1868 n505 R=3.480e+00 
R1868t1341 n1869 n1342 R=3.689e+01 
R1868t366 n1869 n367 R=7.548e+00 
R1869t1472 n1870 n1473 R=6.405e+00 
R1874t834 n1875 n835 R=3.368e+00 
R1876t1038 n1877 n1039 R=3.423e+01 
R1877t238 n1878 n239 R=1.455e+01 
R1877t609 n1878 n610 R=7.435e+00 
R1877t821 n1878 n822 R=4.926e+01 
R1879t578 n1880 n579 R=2.308e+00 
R1879t870 n1880 n871 R=4.348e+00 
R1880t506 n1881 n507 R=1.671e+01 
R1880t1284 n1881 n1285 R=6.558e+00 
R1881t1572 n1882 n1573 R=7.643e+00 
R1882t936 n1883 n937 R=4.560e+00 
R1883t91 n1884 n92 R=1.157e+01 
R1883t901 n1884 n902 R=1.946e+01 
R1883t750 n1884 n751 R=5.793e+00 
R1884t422 n1885 n423 R=1.346e+01 
R1885t1005 n1886 n1006 R=5.425e+00 
R1885t388 n1886 n389 R=3.748e+00 
R1887t1489 n1888 n1490 R=3.134e+00 
R1887t1430 n1888 n1431 R=7.166e+00 
R1887t938 n1888 n939 R=1.692e+01 
R1888t455 n1889 n456 R=5.651e+00 
R1889t42 n1 n43 R=1.053e+01 
R1893t338 n1894 n339 R=8.086e+00 
R1893t1209 n1894 n1210 R=3.594e+00 
R1894t1605 n1895 n1606 R=1.372e+01 
R1895t437 n1896 n438 R=4.693e+01 
R1895t1008 n1896 n1009 R=2.063e+00 
R1897t416 n1898 n417 R=2.196e+00 
R1900t1608 n1901 n1609 R=6.875e+00 
R1901t263 n1902 n264 R=1.327e+01 
R1902t813 n1903 n814 R=4.617e+00 
R1902t617 n1903 n618 R=1.499e+01 
R1903t1876 n1904 n1877 R=5.593e+00 
R1905t294 n1906 n295 R=2.281e+00 
R1905t1820 n1906 n1821 R=1.292e+01 
R1906t648 n1907 n649 R=3.288e+00 
R1906t913 n1907 n914 R=4.120e+00 
R1907t399 n1908 n400 R=2.893e+01 
R1908t453 n1909 n454 R=1.031e+01 
R1908t415 n1909 n416 R=1.189e+02 
R1909t275 n1910 n276 R=4.362e+00 
R1909t48 n1910 n49 R=1.210e+01 
R1910t535 n1911 n536 R=2.725e+00 
R1911t37 n1912 n38 R=1.646e+01 
R1912t1104 n1913 n1105 R=1.744e+01 
R1914t1497 n1915 n1498 R=7.233e+00 
R1914t1738 n1915 n1739 R=1.246e+01 
R1917t216 n1918 n217 R=5.033e+00 
R1917t356 n1918 n357 R=9.650e+00 
R1918t503 n1919 n504 R=6.184e+00 
R1919t1744 n1920 n1745 R=3.218e+00 
R1920t701 n1921 n702 R=3.169e+01 
R1921t252 n1922 n253 R=3.928e+00 
R1921t729 n1922 n730 R=1.972e+01 
R1922t601 n1923 n602 R=1.930e+01 
R1922t496 n1923 n497 R=4.679e+00 
R1924t989 n1925 n990 R=5.663e+00 
R1924t1222 n1925 n1223 R=1.480e+01 
R1925t1776 n1926 n1777 R=4.364e+00 
R1926t328 n1927 n329 R=3.178e+01 
R1926t752 n1927 n753 R=1.411e+01 
R1926t1867 n1927 n1868 R=2.429e+02 
R1926t651 n1927 n652 R=1.046e+01 
R1927t458 n1928 n459 R=1.698e+01 
R1928t288 n1929 n289 R=4.853e+00 
R1929t856 n1930 n857 R=1.313e+01 
R1930t1631 n1931 n1632 R=6.267e+00 
R1930t302 n1931 n303 R=7.168e+00 
R1931t47 n1932 n48 R=2.226e+00 
R1931t114 n1932 n115 R=4.443e+00 
R1932t203 n1933 n204 R=8.422e+00 
R1932t1802 n1933 n1803 R=8.107e+00 
R1933t1834 n1934 n1835 R=3.832e+01 
R1933t1739 n1934 n1740 R=2.251e+01 
R1934t167 n1935 n168 R=1.808e+01 
R1934t1629 n1935 n1630 R=1.371e+01 
R1934t361 n1935 n362 R=1.846e+01 
R1934t685 n1935 n686 R=1.526e+01 
R1935t1381 n1936 n1382 R=4.109e+00 
R1937t193 n1938 n194 R=7.600e+00 
R1937t1165 n1938 n1166 R=3.077e+01 
R1938t1100 n1939 n1101 R=5.782e+00 
R1938t914 n1939 n915 R=1.411e+01 
R1940t1025 n1941 n1026 R=1.042e+01 
R1941t1390 n1942 n1391 R=4.750e+00 
R1942t387 n1943 n388 R=4.502e+00 
R1942t1456 n1943 n1457 R=4.739e+00 
R1944t1744 n1945 n1745 R=4.120e+00 
R1944t1919 n1945 n1920 R=4.856e+00 
R1948t638 n1949 n639 R=3.620e+00 
R1950t1303 n1951 n1304 R=6.576e+00 
R1952t1710 n1953 n1711 R=7.818e+00 
R1952t326 n1953 n327 R=2.706e+01 
R1954t1093 n1955 n1094 R=2.023e+00 
R1955t1049 n1956 n1050 R=8.115e+00 
R1956t221 n1957 n222 R=6.845e+00 
R1957t1539 n1958 n1540 R=3.172e+01 
R1957t962 n1958 n963 R=2.233e+01 
R1960t983 n1961 n984 R=2.469e+00 
R1961t728 n1962 n729 R=4.756e+00 
R1962t1746 n1963 n1747 R=7.150e+00 
R1962t1760 n1963 n1761 R=9.938e+00 
R1963t948 n1964 n949 R=2.196e+00 
R1964t474 n1965 n475 R=4.095e+00 
R1967t1090 n1968 n1091 R=5.023e+00 
R1968t1401 n1969 n1402 R=4.023e+01 
R1969t1681 n1970 n1682 R=4.533e+00 
R1970t456 n1971 n457 R=6.623e+00 
R1973t50 n1974 n51 R=3.160e+00 
R1974t1131 n1975 n1132 R=3.009e+00 
R1975t459 n1976 n460 R=1.511e+01 
R1976t1400 n1977 n1401 R=9.260e+00 
R1976t661 n1977 n662 R=6.796e+00 
R1977t1033 n1978 n1034 R=3.982e+00 
R1977t1481 n1978 n1482 R=1.750e+01 
R1977t481 n1978 n482 R=7.924e+00 
R1979t856 n1980 n857 R=1.436e+01 
R1979t1929 n1980 n1930 R=2.761e+00 
R1980t1607 n1981 n1608 R=9.969e+00 
R1980t1622 n1981 n1623 R=9.402e+00 
R1980t1716 n1981 n1717 R=1.180e+01 
R1981t742 n1982 n743 R=3.740e+00 
R1981t1587 n1982 n1588 R=1.124e+02 
R1982t1335 n1983 n1336 R=3.034e+00 
R1982t1800 n1983 n1801 R=2.714e+02 
R1982t988 n1983 n989 R=1.423e+01 
R1983t1229 n1984 n1230 R=2.122e+01 
R1985t972 n1986 n973 R=1.495e+01 
R1985t1006 n1986 n1007 R=2.465e+00 
R1985t139 n1986 n140 R=4.947e+00 
R1986t929 n1987 n930 R=2.433e+01 
R1986t697 n1987 n698 R=6.339e+02 
R1987t936 n1988 n937 R=8.116e+00 
R1988t1685 n1989 n1686 R=6.175e+00 
R1988t1032 n1989 n1033 R=1.027e+02 
R1989t577 n1990 n578 R=6.397e+00 
R1989t873 n1990 n874 R=2.002e+01 
R1991t1598 n1992 n1599 R=6.468e+00 
R1992t40 n1993 n41 R=5.114e+00 
R1993t1369 n1994 n1370 R=3.691e+00 
R1995t990 n1996 n991 R=4.113e+00 
R1995t943 n1996 n944 R=9.500e+00 
R1995t131 n1996 n132 R=3.911e+00 
R1999t1214 n2000 n1215 R=5.788e+01 
R2000t350 n2001 n351 R=2.602e+01 
R2001t1463 n2002 n1464 R=9.019e+00 
R2002t345 n2003 n346 R=9.246e+00 
R2004t463 n2005 n464 R=9.336e+00 
R2004t1429 n2005 n1430 R=3.095e+01 
R2005t104 n2006 n105 R=8.694e+00 
R2006t1984 n2007 n1985 R=3.235e+00 
R2007t733 n2008 n734 R=2.104e+00 
R2009t810 n2010 n811 R=2.594e+00 
R2009t1562 n2010 n1563 R=1.204e+01 
R2009t439 n2010 n440 R=3.878e+01 
R2010t347 n2011 n348 R=4.532e+02 
R2010t1863 n2011 n1864 R=7.599e+00 
R2011t1503 n2012 n1504 R=2.945e+01 
R2011t1722 n2012 n1723 R=1.922e+01 
R2012t885 n2013 n886 R=1.601e+01 
R2015t1577 n2016 n1578 R=2.122e+01 
R2016t733 n2017 n734 R=4.786e+00 
R2016t1589 n2017 n1590 R=4.162e+00 
R2017t1428 n2018 n1429 R=5.709e+00 
R2018t477 n2019 n478 R=9.291e+00 
R2019t1664 n2020 n1665 R=4.622e+00 
R2022t735 n2023 n736 R=2.117e+01 
R2022t1328 n2023 n1329 R=6.476e+00 
R2024t946 n2025 n947 R=2.050e+00 
R2024t954 n2025 n955 R=3.275e+00 
R2025t723 n2026 n724 R=1.893e+01 
R2026t306 n2027 n307 R=7.653e+00 
R2027t536 n2028 n537 R=3.001e+01 
R2028t855 n2029 n856 R=6.221e+00 
R2028t1518 n2029 n1519 R=3.068e+00 
R2028t1294 n2029 n1295 R=1.803e+01 
R2030t594 n2031 n595 R=1.152e+01 
R2031t1754 n2032 n1755 R=8.458e+00 
R2033t196 n2034 n197 R=9.953e+00 
R2035t1937 n2036 n1938 R=2.810e+00 
R2036t459 n2037 n460 R=6.789e+00 
R2036t793 n2037 n794 R=1.004e+01 
R2042t620 n2043 n621 R=3.080e+00 
R2043t1757 n2044 n1758 R=1.176e+01 
R2044t309 n2045 n310 R=1.223e+01 
R2045t350 n2046 n351 R=3.757e+00 
R2047t1812 n2048 n1813 R=3.916e+00 
R2047t1645 n2048 n1646 R=7.666e+00 
R2049t1190 n2050 n1191 R=3.264e+00 
R2050t1285 n2051 n1286 R=2.644e+01 
R2050t1226 n2051 n1227 R=1.285e+01 
R2050t149 n2051 n150 R=2.691e+00 
R2051t529 n2052 n530 R=8.531e+00 
R2052t1593 n2053 n1594 R=4.278e+00 
R2053t898 n2054 n899 R=1.890e+01 
R2053t656 n2054 n657 R=3.054e+00 
R2054t1293 n2055 n1294 R=6.384e+00 
R2054t1740 n2055 n1741 R=2.201e+01 
R2054t105 n2055 n106 R=1.861e+01 
R2054t70 n2055 n71 R=2.909e+02 
R2055t250 n2056 n251 R=3.823e+00 
R2056t581 n2057 n582 R=3.961e+00 
R2059t945 n2060 n946 R=6.188e+00 
R2060t122 n2061 n123 R=5.142e+00 
R2061t1034 n2062 n1035 R=3.584e+00 
R2062t1676 n2063 n1677 R=2.883e+01 
R2064t1014 n2065 n1015 R=2.069e+01 
R2065t766 n2066 n767 R=1.128e+01 
R2066t1459 n2067 n1460 R=9.524e+00 
R2068t1950 n2069 n1951 R=4.794e+00 
R2068t1303 n2069 n1304 R=1.444e+01 
R2071t643 n2072 n644 R=6.625e+00 
R2073t1886 n2074 n1887 R=1.118e+01 
R2074t1178 n2075 n1179 R=3.163e+01 
R2074t1388 n2075 n1389 R=2.625e+00 
R2074t1227 n2075 n1228 R=5.621e+00 
R2074t1145 n2075 n1146 R=5.669e+00 
R2075t210 n2076 n211 R=8.377e+00 
R2076t657 n2077 n658 R=3.874e+00 
R2077t136 n2078 n137 R=2.539e+00 
R2078t224 n2079 n225 R=8.931e+00 
R2078t1325 n2079 n1326 R=9.196e+00 
R2078t1915 n2079 n1916 R=2.968e+00 
R2078t1055 n2079 n1056 R=1.895e+01 
R2079t1085 n2080 n1086 R=8.181e+00 
R2080t1248 n2081 n1249 R=3.951e+01 
R2080t327 n2081 n328 R=4.464e+01 
R2081t1967 n2082 n1968 R=1.778e+01 
R2082t642 n2083 n643 R=1.883e+01 
R2082t1088 n2083 n1089 R=2.685e+01 
R2083t814 n2084 n815 R=7.429e+00 
R2084t99 n2085 n100 R=1.496e+01 
R2085t1384 n2086 n1385 R=3.375e+00 
R2086t1893 n2087 n1894 R=3.763e+00 
R2087t1828 n2088 n1829 R=1.999e+01 
R2087t1617 n2088 n1618 R=1.021e+01 
R2087t1635 n2088 n1636 R=1.660e+01 
R2087t644 n2088 n645 R=3.219e+00 
R2087t1129 n2088 n1130 R=1.990e+01 
R2088t1740 n2089 n1741 R=4.031e+00 
R2088t105 n2089 n106 R=2.560e+01 
R2089t401 n2090 n402 R=9.548e+01 
R2092t1858 n2093 n1859 R=3.048e+00 
R2094t1373 n2095 n1374 R=2.358e+01 
R2097t223 n2098 n224 R=3.324e+00 
R2097t1863 n2098 n1864 R=1.274e+02 
R2098t730 n2099 n731 R=8.216e+01 
R2098t271 n2099 n272 R=3.516e+00 
R2099t952 n2100 n953 R=5.244e+01 
R2099t768 n2100 n769 R=1.599e+01 
R2099t1848 n2100 n1849 R=8.486e+00 
R2100t154 n2101 n155 R=8.233e+01 
R2100t1777 n2101 n1778 R=9.937e+00 
R2101t817 n2102 n818 R=2.002e+00 
R2101t14 n2102 n15 R=3.049e+01 
R2103t474 n2104 n475 R=1.005e+01 
R2103t400 n2104 n401 R=4.378e+00 
R2103t1482 n2104 n1483 R=8.821e+01 
R2104t235 n2105 n236 R=1.179e+01 
R2104t1720 n2105 n1721 R=8.294e+00 
R2105t1141 n2106 n1142 R=1.365e+01 
R2105t669 n2106 n670 R=3.061e+01 
R2105t1903 n2106 n1904 R=1.263e+01 
R2106t2105 n2107 n2106 R=1.414e+02 
R2106t669 n2107 n670 R=2.976e+00 
R2107t1327 n2108 n1328 R=4.007e+00 
R2107t639 n2108 n640 R=3.904e+00 
R2108t1742 n2109 n1743 R=3.133e+00 
R2108t1224 n2109 n1225 R=1.275e+02 
R2110t1246 n2111 n1247 R=2.152e+01 
R2111t1148 n2112 n1149 R=4.831e+00 
R2111t720 n2112 n721 R=1.914e+00 
R2111t1549 n2112 n1550 R=6.942e+01 
R2112t712 n2113 n713 R=7.563e+00 
R2112t403 n2113 n404 R=8.021e+01 
R2114t362 n2115 n363 R=3.576e+01 
R2114t475 n2115 n476 R=5.352e+00 
R2114t1680 n2115 n1681 R=2.491e+01 
R2116t1287 n2117 n1288 R=1.200e+01 
R2116t113 n2117 n114 R=2.929e+00 
R2116t1355 n2117 n1356 R=1.451e+01 
R2117t1246 n2118 n1247 R=5.772e+00 
R2117t2110 n2118 n2111 R=3.172e+01 
R2118t1462 n2119 n1463 R=4.097e+00 
R2118t732 n2119 n733 R=1.259e+01 
R2118t961 n2119 n962 R=9.352e+00 
R2118t440 n2119 n441 R=1.034e+01 
R2120t1741 n2121 n1742 R=2.488e+00 
R2122t1259 n2123 n1260 R=5.359e+01 
R2123t399 n2124 n400 R=2.520e+01 
R2123t987 n2124 n988 R=5.772e+00 
R2124t1487 n2125 n1488 R=4.937e+00 
R2125t670 n2126 n671 R=3.410e+01 
R2126t637 n2127 n638 R=1.535e+00 
R2126t1449 n2127 n1450 R=5.920e+01 
R2127t336 n2128 n337 R=6.503e+00 
R2127t1817 n2128 n1818 R=2.605e+00 
R2127t918 n2128 n919 R=1.820e+02 
R2128t1286 n2129 n1287 R=8.786e+00 
R2128t2119 n2129 n2120 R=2.522e+00 
R2129t654 n2130 n655 R=4.853e+00 
R2130t1570 n2131 n1571 R=7.407e+00 
R2132t1611 n2133 n1612 R=2.477e+01 
R2133t234 n2134 n235 R=4.229e+00 
R2133t1865 n2134 n1866 R=4.596e+01 
R2134t1020 n2135 n1021 R=6.166e+00 
R2134t638 n2135 n639 R=4.315e+00 
R2135t1510 n2136 n1511 R=3.338e+00 
R2136t1972 n2137 n1973 R=6.390e+00 
R2138t983 n2139 n984 R=1.199e+02 
R2138t1960 n2139 n1961 R=6.948e+00 
R2138t994 n2139 n995 R=4.663e+00 
R2139t1943 n2140 n1944 R=3.555e+00 
R2142t1760 n2143 n1761 R=7.299e+00 
R2143t423 n2144 n424 R=7.976e+00 
R2143t65 n2144 n66 R=5.886e+00 
R2144t471 n2145 n472 R=4.228e+00 
R2145t709 n2146 n710 R=4.027e+00 
R2147t25 n2148 n26 R=2.276e+01 
R2147t93 n2148 n94 R=1.179e+01 
R2148t1443 n2149 n1444 R=9.184e+00 
R2149t1764 n2150 n1765 R=3.141e+01 
R2150t594 n2151 n595 R=3.040e+00 
R2151t207 n2152 n208 R=1.327e+01 
R2151t1481 n2152 n1482 R=1.118e+02 
R2152t1493 n2153 n1494 R=1.078e+01 
R2153t830 n2154 n831 R=3.117e+00 
R2153t516 n2154 n517 R=4.217e+00 
R2153t1508 n2154 n1509 R=5.107e+00 
R2154t1620 n2155 n1621 R=1.957e+03 
R2155t233 n2156 n234 R=1.123e+01 
R2156t1168 n2157 n1169 R=3.652e+01 
R2156t282 n2157 n283 R=1.038e+01 
R2157t938 n2158 n939 R=9.751e+00 
R2157t596 n2158 n597 R=5.274e+00 
R2157t1137 n2158 n1138 R=1.126e+01 
R2158t1447 n2159 n1448 R=3.574e+00 
R2159t451 n2160 n452 R=4.181e+00 
R2160t95 n2161 n96 R=2.694e+01 
R2162t2109 n2163 n2110 R=1.117e+01 
R2163t32 n2164 n33 R=1.673e+01 
R2164t1181 n2165 n1182 R=4.072e+00 
R2166t1820 n2167 n1821 R=5.758e+00 
R2166t1905 n2167 n1906 R=3.211e+00 
R2167t1765 n2168 n1766 R=7.692e+00 
R2167t1806 n2168 n1807 R=1.699e+01 
R2168t1775 n2169 n1776 R=1.026e+02 
R2168t201 n2169 n202 R=1.138e+01 
R2168t967 n2169 n968 R=3.494e+00 
R2169t523 n2170 n524 R=4.150e+00 
R2170t377 n2171 n378 R=5.223e+01 
R2170t155 n2171 n156 R=6.150e+00 
R2171t1751 n2172 n1752 R=2.018e+01 
R2173t652 n2174 n653 R=6.028e+00 
R2174t1494 n2175 n1495 R=3.502e+01 
R2174t255 n2175 n256 R=6.610e+00 
R2174t297 n2175 n298 R=2.650e+00 
R2175t215 n2176 n216 R=4.265e+00 
R2175t1780 n2176 n1781 R=2.583e+00 
R2176t1176 n2177 n1177 R=6.283e+01 
R2176t1691 n2177 n1692 R=5.597e+00 
R2176t1111 n2177 n1112 R=2.213e+00 
R2177t1176 n2178 n1177 R=3.416e+00 
R2177t63 n2178 n64 R=4.709e+00 
R2178t287 n2179 n288 R=2.504e+01 
R2179t1674 n2180 n1675 R=3.132e+00 
R2180t311 n2181 n312 R=4.381e+01 
R2181t411 n2182 n412 R=6.677e+01 
R2181t566 n2182 n567 R=4.653e+00 
R2183t1801 n2184 n1802 R=3.850e+01 
R2183t1370 n2184 n1371 R=3.514e+01 
R2184t1520 n2185 n1521 R=2.634e+00 
R2186t1817 n2187 n1818 R=2.512e+01 
R2186t1535 n2187 n1536 R=1.768e+01 
R2187t2185 n2188 n2186 R=3.539e+00 
R2188t1305 n2189 n1306 R=8.590e+00 
R2191t1929 n2192 n1930 R=2.899e+01 
R2191t1687 n2192 n1688 R=6.923e+00 
R2192t191 n2193 n192 R=1.148e+01 
R2192t1753 n2193 n1754 R=2.488e+01 
R2192t505 n2193 n506 R=2.005e+01 
R2194t744 n2195 n745 R=4.190e+02 
R2195t126 n2196 n127 R=1.584e+02 
R2195t1643 n2196 n1644 R=7.971e+00 
R2195t1061 n2196 n1062 R=4.702e+00 
R2199t19 n2200 n20 R=3.064e+00 
R2199t1036 n2200 n1037 R=2.924e+00 
R2201t1899 n2202 n1900 R=1.591e+01 
R2201t1663 n2202 n1664 R=4.311e+00 
R2202t504 n2203 n505 R=3.795e+00 
R2202t792 n2203 n793 R=6.678e+01 
R2202t713 n2203 n714 R=6.575e+00 
R2203t1636 n2204 n1637 R=3.290e+00 
R2203t340 n2204 n341 R=4.253e+00 
R2204t1417 n2205 n1418 R=7.641e+00 
R2206t1776 n2207 n1777 R=6.524e+00 
R2207t487 n2208 n488 R=9.814e+01 
R2207t1347 n2208 n1348 R=9.860e+00 
R2207t1717 n2208 n1718 R=9.668e+00 
R2208t2136 n2209 n2137 R=2.793e+00 
R2209t1243 n2210 n1244 R=3.636e+01 
R2210t1158 n2211 n1159 R=6.923e+00 
R2211t2140 n2212 n2141 R=5.108e+00 
R2212t1696 n2213 n1697 R=1.187e+01 
R2213t2017 n2214 n2018 R=6.739e+00 
R2213t1053 n2214 n1054 R=6.052e+00 
R2215t330 n2216 n331 R=2.570e+01 
R2216t705 n2217 n706 R=7.737e+00 
R2218t2146 n2219 n2147 R=3.892e+00 
R2219t316 n2220 n317 R=2.826e+00 
R2219t1516 n2220 n1517 R=3.691e+01 
R2219t1299 n2220 n1300 R=1.884e+02 
R2220t570 n2221 n571 R=2.198e+00 
R2221t1274 n2222 n1275 R=1.427e+01 
R2221t1049 n2222 n1050 R=5.919e+00 
R2222t869 n2223 n870 R=3.409e+00 
R2223t380 n2224 n381 R=1.846e+01 
R2224t2065 n2225 n2066 R=5.811e+01 
R2226t1808 n2227 n1809 R=1.496e+01 
R2227t33 n2228 n34 R=4.113e+00 
R2227t170 n2228 n171 R=4.553e+00 
R2229t1864 n2230 n1865 R=6.549e+00 
R2229t1714 n2230 n1715 R=2.639e+00 
R2229t705 n2230 n706 R=1.067e+01 
R2230t1289 n2231 n1290 R=7.346e+00 
R2231t1395 n2232 n1396 R=2.097e+01 
R2231t1298 n2232 n1299 R=1.054e+02 
R2231t788 n2232 n789 R=8.790e+01 
R2231t1975 n2232 n1976 R=4.475e+00 
R2231t343 n2232 n344 R=2.390e+00 
R2234t366 n2235 n367 R=2.985e+00 
R2234t2130 n2235 n2131 R=3.059e+01 
R2235t2182 n2236 n2183 R=5.755e+02 
R2236t2150 n2237 n2151 R=1.899e+01 
R2236t2030 n2237 n2031 R=3.268e+00 
R2236t594 n2237 n595 R=4.109e+00 
R2237t970 n2238 n971 R=1.276e+01 
R2237t484 n2238 n485 R=5.840e+00 
R2238t1729 n2239 n1730 R=4.637e+00 
R2239t878 n2240 n879 R=6.792e+00 
R2240t2105 n2241 n2106 R=1.029e+01 
R2241t22 n2242 n23 R=5.347e+00 
R2241t1387 n2242 n1388 R=1.378e+01 
R2243t280 n2244 n281 R=5.248e+02 
R2243t1485 n2244 n1486 R=6.812e+00 
R2244t1983 n2245 n1984 R=6.867e+00 
R2244t1943 n2245 n1944 R=1.567e+01 
R2245t645 n2246 n646 R=1.723e+00 
R2246t1203 n2247 n1204 R=3.738e+00 
R2247t1670 n2248 n1671 R=8.151e+00 
R2248t1163 n2249 n1164 R=9.700e+00 
R2249t1672 n2250 n1673 R=1.733e+00 
R2250t1121 n2251 n1122 R=8.705e+00 
R2251t284 n2252 n285 R=2.483e+00 
R2253t22 n2254 n23 R=1.212e+01 
R2253t2241 n2254 n2242 R=7.700e+00 
R2253t801 n2254 n802 R=1.254e+01 
R2254t1129 n2255 n1130 R=6.511e+00 
R2256t2023 n2257 n2024 R=1.631e+01 
R2256t1884 n2257 n1885 R=5.057e+00 
R2256t342 n2257 n343 R=7.105e+00 
R2257t2217 n2258 n2218 R=4.460e+01 
R2258t60 n2259 n61 R=6.672e+00 
R2258t1318 n2259 n1319 R=1.357e+02 
R2259t1175 n2260 n1176 R=4.091e+01 
R2260t1397 n2261 n1398 R=4.292e+00 
R2261t1146 n2262 n1147 R=3.828e+01 
R2261t1502 n2262 n1503 R=2.226e+01 
R2261t1760 n2262 n1761 R=3.337e+00 
R2262t216 n2263 n217 R=8.164e+00 
R2262t1917 n2263 n1918 R=8.053e+00 
R2262t356 n2263 n357 R=4.186e+00 
R2263t217 n2264 n218 R=3.749e+01 
R2263t1634 n2264 n1635 R=4.580e+00 
R2264t600 n2265 n601 R=1.428e+01 
R2264t15 n2265 n16 R=3.588e+01 
R2264t1309 n2265 n1310 R=6.421e+00 
R2265t1900 n2266 n1901 R=7.993e+00 
R2267t316 n2268 n317 R=5.207e+00 
R2267t1516 n2268 n1517 R=2.496e+00 
R2268t2048 n2269 n2049 R=9.253e+00 
R2269t224 n2270 n225 R=2.627e+00 
R2269t2078 n2270 n2079 R=1.494e+03 
R2269t1055 n2270 n1056 R=3.124e+00 
R2270t1946 n2271 n1947 R=3.327e+00 
R2270t519 n2271 n520 R=9.134e+00 
R2274t2230 n2275 n2231 R=1.959e+01 
R2274t499 n2275 n500 R=7.096e+00 
R2275t76 n2276 n77 R=9.560e+00 
R2275t976 n2276 n977 R=6.947e+00 
R2275t1392 n2276 n1393 R=6.955e+00 
R2275t456 n2276 n457 R=4.201e+00 
R2275t998 n2276 n999 R=7.856e+00 
R2276t1694 n2277 n1695 R=8.057e+00 
R2276t522 n2277 n523 R=5.209e+00 
R2278t1170 n2279 n1171 R=1.782e+01 
R2278t269 n2279 n270 R=7.867e+00 
R2279t429 n2280 n430 R=7.740e+00 
R2279t560 n2280 n561 R=2.422e+01 
R2280t472 n2281 n473 R=2.485e+01 
R2280t1293 n2281 n1294 R=2.041e+01 
R2280t2109 n2281 n2110 R=4.032e+00 
R2281t257 n2282 n258 R=5.718e+00 
R2282t2208 n2283 n2209 R=6.048e+01 
R2282t1139 n2283 n1140 R=2.428e+00 
R2283t470 n2284 n471 R=2.837e+00 
R2283t999 n2284 n1000 R=2.148e+00 
R2284t329 n2285 n330 R=6.524e+00 
R2284t442 n2285 n443 R=7.729e+00 
R2285t449 n2286 n450 R=3.093e+00 
R2287t848 n2288 n849 R=9.049e+00 
R2288t171 n2289 n172 R=1.256e+01 
R2289t2052 n2290 n2053 R=5.517e+00 
R2290t906 n2291 n907 R=7.121e+00 
R2291t383 n2292 n384 R=4.240e+01 
R2291t558 n2292 n559 R=1.175e+01 
R2291t476 n2292 n477 R=1.630e+01 
R2292t106 n2293 n107 R=8.720e+00 
R2293t1983 n2294 n1984 R=5.662e+00 
R2293t2244 n2294 n2245 R=1.194e+01 
R2294t2286 n2295 n2287 R=7.759e+00 
R2295t21 n2296 n22 R=5.806e+00 
R2295t1045 n2296 n1046 R=4.949e+01 
R2295t1479 n2296 n1480 R=2.511e+00 
R2296t823 n2297 n824 R=1.657e+01 
R2296t245 n2297 n246 R=1.792e+00 
R2297t506 n2298 n507 R=1.044e+01 
R2297t605 n2298 n606 R=2.592e+01 
R2297t1880 n2298 n1881 R=4.298e+00 
R2298t2093 n2299 n2094 R=7.131e+00 
R2299t2030 n2300 n2031 R=7.902e+00 
R2299t2236 n2300 n2237 R=5.629e+02 
R2300t318 n2301 n319 R=1.574e+02 
R2301t1930 n2302 n1931 R=1.114e+01 
R2302t1182 n2303 n1183 R=2.243e+01 
R2303t2021 n2304 n2022 R=1.123e+01 
R2304t727 n2305 n728 R=3.126e+00 
R2305t397 n2306 n398 R=2.550e+01 
R2305t722 n2306 n723 R=1.088e+01 
R2306t770 n2307 n771 R=4.170e+00 
R2306t1163 n2307 n1164 R=2.235e+02 
R2307t2013 n2308 n2014 R=5.996e+01 
R2307t1385 n2308 n1386 R=4.261e+00 
R2308t960 n2309 n961 R=3.604e+00 
R2308t1518 n2309 n1519 R=1.891e+01 
R2308t1412 n2309 n1413 R=1.245e+01 
R2308t1465 n2309 n1466 R=2.083e+01 
R2311t664 n2312 n665 R=1.948e+00 
R2313t19 n2314 n20 R=8.065e+00 
R2314t1898 n2315 n1899 R=4.652e+00 
R2315t1824 n2316 n1825 R=2.034e+00 
R2315t2094 n2316 n2095 R=6.624e+00 
R2316t1125 n2317 n1126 R=1.618e+01 
R2318t1245 n2319 n1246 R=1.027e+01 
R2319t1327 n2320 n1328 R=8.442e+00 
R2319t2107 n2320 n2108 R=1.133e+01 
R2320t523 n2321 n524 R=6.237e+00 
R2320t916 n2321 n917 R=6.340e+00 
R2322t822 n2323 n823 R=3.976e+01 
R2324t1160 n2325 n1161 R=1.123e+01 
R2325t368 n2326 n369 R=5.182e+00 
R2326t337 n2327 n338 R=2.324e+01 
R2327t1611 n2328 n1612 R=1.612e+01 
R2327t771 n2328 n772 R=3.315e+01 
R2328t1149 n2329 n1150 R=1.455e+01 
R2331t108 n2332 n109 R=3.682e+00 
R2332t812 n2333 n813 R=8.417e+00 
R2332t349 n2333 n350 R=5.478e+00 
R2332t1693 n2333 n1694 R=2.937e+01 
R2334t1968 n2335 n1969 R=3.114e+00 
R2335t1163 n2336 n1164 R=6.690e+00 
R2336t2332 n2337 n2333 R=7.332e+00 
R2336t349 n2337 n350 R=9.169e+00 
R2338t164 n2339 n165 R=2.292e+00 
R2338t1130 n2339 n1131 R=4.250e+00 
R2338t863 n2339 n864 R=4.187e+00 
R2339t1208 n2340 n1209 R=7.065e+00 
R2339t1119 n2340 n1120 R=1.078e+01 
R2340t1323 n2341 n1324 R=4.082e+00 
R2342t1342 n2343 n1343 R=2.753e+02 
R2343t1173 n2344 n1174 R=2.943e+00 
R2343t1795 n2344 n1796 R=2.380e+01 
R2344t2126 n2345 n2127 R=4.362e+00 
R2344t1449 n2345 n1450 R=2.335e+01 
R2344t1850 n2345 n1851 R=1.121e+01 
R2344t246 n2345 n247 R=2.669e+00 
R2345t78 n2346 n79 R=6.638e+00 
R2345t1097 n2346 n1098 R=1.403e+01 
R2345t1021 n2346 n1022 R=9.219e+01 
R2346t117 n2347 n118 R=7.024e+01 
R2347t2200 n2348 n2201 R=2.576e+01 
R2347t2242 n2348 n2243 R=9.418e+00 
R2348t513 n2349 n514 R=1.208e+01 
R2348t387 n2349 n388 R=1.016e+01 
R2349t622 n2350 n623 R=5.662e+00 
R2349t2147 n2350 n2148 R=5.092e+00 
R2350t1632 n2351 n1633 R=2.690e+00 
R2350t7 n2351 n8 R=7.608e+00 
R2351t1887 n2352 n1888 R=2.237e+01 
R2351t938 n2352 n939 R=6.049e+00 
R2352t563 n2353 n564 R=5.278e+00 
R2352t1984 n2353 n1985 R=6.863e+01 
R2354t370 n2355 n371 R=4.885e+00 
R2354t279 n2355 n280 R=3.158e+01 
R2355t670 n2356 n671 R=1.519e+01 
R2355t391 n2356 n392 R=1.082e+01 
R2356t231 n2357 n1 R=4.373e+00 
R2359t294 n2360 n295 R=6.672e+00 
R2359t1130 n2360 n1131 R=9.588e+01 
R2359t164 n2360 n165 R=3.229e+01 
R2360t1990 n2361 n1991 R=6.740e+00 
R2360t2301 n2361 n2302 R=6.501e+00 
R2363t263 n2364 n264 R=4.864e+00 
R2363t702 n2364 n703 R=5.980e+00 
R2364t1741 n2365 n1742 R=7.705e+00 
R2364t2120 n2365 n2121 R=5.625e+00 
R2365t409 n2366 n410 R=1.442e+01 
R2366t2239 n2367 n2240 R=5.042e+00 
R2366t878 n2367 n879 R=1.695e+01 
R2366t1461 n2367 n1462 R=6.839e+01 
R2368t841 n2369 n842 R=4.415e+00 
R2370t635 n2371 n636 R=1.363e+01 
R2370t540 n2371 n541 R=6.817e+00 
R2371t267 n2372 n268 R=1.056e+01 
R2371t1202 n2372 n1203 R=2.227e+01 
R2371t2011 n2372 n2012 R=7.554e+00 
R2372t1359 n2373 n1360 R=7.424e+01 
R2373t2081 n2374 n2082 R=5.896e+01 
R2375t1759 n2376 n1760 R=1.170e+01 
R2375t1172 n2376 n1173 R=8.641e+00 
R2379t1189 n2380 n1190 R=4.880e+00 
R2379t395 n2380 n396 R=1.565e+01 
R2380t1945 n2381 n1946 R=4.769e+00 
R2380t240 n2381 n241 R=9.528e+00 
R2381t607 n2382 n608 R=7.563e+00 
R2381t1529 n2382 n1530 R=5.276e+00 
R2382t2267 n2383 n2268 R=1.135e+01 
R2382t316 n2383 n317 R=1.139e+01 
R2382t2219 n2383 n2220 R=5.533e+00 
R2383t470 n2384 n471 R=2.518e+02 
R2383t2283 n2384 n2284 R=4.897e+00 
R2383t999 n2384 n1000 R=6.949e+01 
R2384t509 n2385 n510 R=2.659e+00 
R2384t1683 n2385 n1684 R=3.074e+01 
R2385t880 n2386 n881 R=6.516e+00 
R2385t767 n2386 n768 R=9.654e+00 
R2385t457 n2386 n458 R=1.760e+01 
R2386t434 n2387 n435 R=4.158e+00 
R2386t430 n2387 n431 R=1.282e+01 
R2387t2018 n2388 n2019 R=3.425e+01 
R2387t2356 n2388 n2357 R=1.094e+01 
R2387t706 n2388 n707 R=8.477e+00 
R2388t1968 n2389 n1969 R=2.057e+01 
R2388t2334 n2389 n2335 R=1.139e+02 
R2389t318 n2390 n319 R=1.584e+01 
R2389t2300 n2390 n2301 R=1.520e+00 
R2389t613 n2390 n614 R=1.989e+01 
R2391t1723 n2392 n1724 R=3.754e+00 
R2391t841 n2392 n842 R=2.345e+01 
R2391t1978 n2392 n1979 R=3.633e+00 
R2392t1936 n2393 n1937 R=3.060e+03 
R2392t1927 n2393 n1928 R=2.537e+01 
R2392t2005 n2393 n2006 R=1.557e+01 
R2392t104 n2393 n105 R=8.704e+01 
R2393t680 n2394 n681 R=2.448e+00 
R2394t1641 n2395 n1642 R=2.712e+00 
R2396t1512 n2397 n1513 R=2.222e+00 
R2397t5 n2398 n6 R=1.340e+01 
R2397t1451 n2398 n1452 R=1.814e+01 
R2397t241 n2398 n242 R=2.723e+00 
R2397t681 n2398 n682 R=1.598e+01 
R2398t502 n2399 n503 R=4.407e+01 
R2398t1158 n2399 n1159 R=5.954e+00 
R2398t12 n2399 n13 R=3.296e+00 
R2400t1316 n2401 n1317 R=1.172e+01 
R2401t1348 n2402 n1349 R=6.165e+00 
R2401t1543 n2402 n1544 R=2.700e+00 
R2401t266 n2402 n267 R=1.736e+01 
R2402t181 n2403 n182 R=2.372e+00 
R2404t1073 n2405 n1074 R=5.615e+02 
R2405t1302 n2406 n1303 R=9.762e+00 
R2406t773 n2407 n774 R=4.395e+00 
R2406t53 n2407 n54 R=4.904e+00 
R2407t1835 n2408 n1836 R=1.980e+00 
R2407t2140 n2408 n2141 R=3.022e+00 
R2408t2148 n2409 n2149 R=3.335e+00 
R2408t1443 n2409 n1444 R=9.438e+00 
R2408t791 n2409 n792 R=2.007e+01 
R2409t858 n2410 n859 R=4.521e+01 
R2409t26 n2410 n27 R=9.160e+00 
R2410t253 n2411 n254 R=1.416e+01 
R2411t1731 n2412 n1732 R=5.305e+00 
R2411t966 n2412 n967 R=1.174e+01 
R2412t256 n2413 n257 R=1.106e+01 
R2413t616 n2414 n617 R=7.401e+00 
R2414t1936 n2415 n1937 R=1.040e+01 
R2415t1961 n2416 n1962 R=6.297e+00 
R2415t728 n2416 n729 R=1.951e+01 
R2416t1514 n2417 n1515 R=6.095e+00 
R2418t102 n2419 n103 R=1.452e+01 
R2418t1390 n2419 n1391 R=6.485e+00 
R2419t1940 n2420 n1941 R=1.924e+01 
R2419t1025 n2420 n1026 R=7.710e+00 
R2420t1532 n2421 n1533 R=3.699e+00 
R2422t2141 n2423 n2142 R=5.663e+00 
R2422t365 n2423 n366 R=7.360e+01 
R2423t971 n2424 n972 R=6.349e+01 
R2423t1225 n2424 n1226 R=8.022e+00 
R2423t546 n2424 n547 R=1.294e+02 
R2423t109 n2424 n110 R=3.958e+01 
R2426t554 n2427 n555 R=8.912e+00 
R2427t207 n2428 n208 R=2.154e+01 
R2428t1880 n2429 n1881 R=6.849e+00 
R2428t1284 n2429 n1285 R=5.489e+00 
R2429t2324 n2430 n2325 R=4.671e+00 
R2429t296 n2430 n297 R=6.828e+00 
R2430t2268 n2431 n2269 R=5.929e+01 
R2432t2194 n2433 n2195 R=7.182e+00 
R2432t744 n2433 n745 R=1.042e+01 
R2433t243 n2434 n244 R=8.829e+00 
R2433t254 n2434 n255 R=6.832e+00 
R2433t860 n2434 n861 R=4.386e+00 
R2434t1168 n2435 n1169 R=2.279e+01 
R2434t2156 n2435 n2157 R=4.488e+00 
R2434t282 n2435 n283 R=1.811e+01 
R2434t1050 n2435 n1051 R=3.533e+00 
R2435t1040 n2436 n1041 R=2.564e+01 
R2436t2362 n2437 n2363 R=6.541e+00 
R2436t449 n2437 n450 R=1.299e+01 
R2437t606 n2438 n607 R=2.245e+01 
R2437t1826 n2438 n1827 R=1.826e+01 
R2438t2301 n2439 n2302 R=9.843e+00 
R2438t1930 n2439 n1931 R=6.643e+00 
R2438t1631 n2439 n1632 R=1.789e+01 
R2441t365 n2442 n366 R=1.117e+01 
R2441t334 n2442 n335 R=8.057e+01 
R2442t1500 n2443 n1501 R=1.710e+01 
R2443t1403 n2444 n1404 R=1.677e+00 
R2444t2321 n2445 n2322 R=5.505e+00 
R2445t940 n2446 n941 R=1.041e+01 
R2445t1987 n2446 n1988 R=1.676e+01 
R2445t936 n2446 n937 R=5.983e+00 
R2446t1625 n1 n1626 R=6.790e+00 
R2447t969 n2448 n970 R=9.212e+00 
R2448t1189 n2449 n1190 R=4.575e+01 
R2449t1934 n2450 n1935 R=1.253e+01 
R2449t305 n2450 n306 R=5.449e+00 
R2449t685 n2450 n686 R=3.860e+00 
R2450t1551 n2451 n1552 R=9.472e+00 
R2450t1806 n2451 n1807 R=1.195e+01 
R2450t824 n2451 n825 R=8.591e+00 
R2450t2167 n2451 n2168 R=8.512e+00 
R2454t508 n2455 n509 R=7.004e+00 
R2454t1444 n2455 n1445 R=8.938e+00 
R2455t212 n2456 n213 R=9.568e+01 
R2456t1393 n2457 n1394 R=7.751e+00 
R2457t2150 n2458 n2151 R=2.663e+01 
R2457t2236 n2458 n2237 R=4.604e+00 
R2457t2299 n2458 n2300 R=4.507e+00 
R2458t1112 n2459 n1113 R=8.408e+00 
R2458t1437 n2459 n1438 R=4.478e+00 
R2459t172 n2460 n173 R=8.525e+00 
R2459t786 n2460 n787 R=7.103e+00 
R2459t718 n2460 n719 R=3.995e+01 
R2459t1031 n2460 n1032 R=4.600e+00 
R2459t1295 n2460 n1296 R=1.529e+02 
R2460t611 n2461 n612 R=8.061e+00 
R2460t1474 n2461 n1475 R=6.306e+01 
R2461t628 n2462 n629 R=1.867e+01 
R2461t1446 n2462 n1447 R=1.023e+01 
R2461t195 n2462 n196 R=3.425e+01 
R2462t1297 n2463 n1298 R=2.725e+01 
R2462t679 n2463 n680 R=8.991e+00 
R2462t127 n2463 n128 R=1.707e+01 
R2463t301 n2464 n302 R=5.316e+00 
R2465t442 n2466 n443 R=4.207e+02 
R2465t805 n2466 n806 R=4.355e+00 
R2465t495 n2466 n496 R=3.394e+01 
R2466t2249 n2467 n2250 R=2.128e+01 
R2467t1854 n2468 n1855 R=6.371e+00 
R2467t1167 n2468 n1168 R=5.172e+00 
R2468t2173 n2469 n2174 R=4.439e+00 
R2468t652 n2469 n653 R=6.797e+00 
R2468t33 n2469 n34 R=7.600e+00 
R2468t2227 n2469 n2228 R=4.297e+00 
R2469t1206 n2470 n1207 R=3.288e+01 
R2469t353 n2470 n354 R=7.143e+00 
R2469t1662 n2470 n1663 R=3.269e+00 
R2470t1754 n2471 n1755 R=5.828e+00 
R2470t2031 n2471 n2032 R=2.831e+01 
R2470t1124 n2471 n1125 R=1.148e+02 
R2471t787 n2472 n788 R=1.386e+01 
R2472t305 n2473 n306 R=6.753e+00 
R2472t2449 n2473 n2450 R=6.328e+00 
R2472t685 n2473 n686 R=1.398e+02 
R2472t488 n2473 n489 R=3.708e+00 
R2473t891 n2474 n892 R=5.273e+00 
R2473t548 n2474 n549 R=3.525e+01 
R2474t1969 n2475 n1970 R=3.733e+00 
R2474t2187 n2475 n2188 R=7.233e+00 
R2476t987 n2477 n988 R=4.004e+00 
R2476t1136 n2477 n1137 R=1.285e+01 
R2477t1071 n2478 n1072 R=4.197e+00 
R2478t2441 n2479 n2442 R=1.884e+01 
R2479t531 n2480 n532 R=4.774e+00 
R2479t941 n2480 n942 R=3.944e+00 
R2479t101 n2480 n102 R=6.625e+00 
R2479t1550 n2480 n1551 R=1.263e+01 
R2480t1288 n2481 n1289 R=5.689e+01 
R2483t1147 n2484 n1148 R=3.836e+01 
R2483t1682 n2484 n1683 R=9.033e+00 
R2483t484 n2484 n485 R=7.166e+00 
R2484t1578 n2485 n1579 R=5.366e+00 
R2485t1506 n2486 n1507 R=6.810e+00 
R2487t1315 n2488 n1316 R=1.451e+01 
R2487t1698 n2488 n1699 R=3.514e+01 
R2487t671 n2488 n672 R=4.262e+00 
R2488t126 n2489 n127 R=3.069e+01 
R2488t2195 n2489 n2196 R=5.745e+00 
R2489t102 n2490 n103 R=4.587e+00 
R2489t2488 n2490 n2489 R=1.163e+02 
R2490t588 n2491 n589 R=2.666e+01 
R2490t374 n2491 n375 R=8.274e+00 
R2491t181 n2492 n182 R=3.006e+00 
R2491t2402 n2492 n2403 R=2.621e+01 
R2491t2076 n2492 n2077 R=3.427e+00 
R2493t140 n2494 n141 R=1.674e+02 
R2493t1778 n2494 n1779 R=4.262e+00 
R2494t1669 n2495 n1670 R=9.198e+01 
R2494t1618 n2495 n1619 R=1.988e+01 
R2495t2327 n2496 n2328 R=1.653e+01 
R2496t2122 n2497 n2123 R=2.921e+00 
R2496t924 n2497 n925 R=1.507e+01 
R2497t627 n2498 n628 R=6.668e+00 
R2499t1049 n2500 n1050 R=2.285e+01 
R2499t348 n2500 n349 R=1.648e+01 
R2500t614 n2501 n615 R=1.666e+02 
R2500t1279 n2501 n1280 R=5.887e+00 
R2500t1119 n2501 n1120 R=7.860e+00 
R2501t1324 n2502 n1325 R=6.604e+00 
R2502t1552 n2503 n1553 R=4.252e+01 
R2502t1201 n2503 n1 R=6.370e+00 
R2503t1884 n2504 n1885 R=6.205e+01 
R2503t2256 n2504 n2257 R=5.839e+00 
R2503t2023 n2504 n2024 R=8.452e+00 
R2504t854 n2505 n855 R=9.912e+00 
R2505t1080 n2506 n1081 R=7.894e+00 
R2506t1084 n2507 n1085 R=1.063e+01 
R2506t1839 n2507 n1 R=4.571e+00 
R2506t1670 n2507 n1671 R=2.979e+00 
R2507t983 n2508 n984 R=9.507e+00 
R2508t826 n2509 n827 R=1.026e+01 
R2509t832 n2510 n833 R=3.443e+00 
R2510t975 n2511 n976 R=5.539e+00 
R2510t1060 n2511 n1061 R=8.025e+00 
R2510t783 n2511 n784 R=1.848e+01 
R2511t224 n2512 n225 R=3.389e+01 
R2511t2078 n2512 n2079 R=6.045e+00 
R2511t1325 n2512 n1326 R=4.292e+00 
R2512t1752 n2513 n1753 R=6.763e+01 
R2513t1661 n2514 n1662 R=1.085e+01 
R2514t1277 n2515 n1278 R=4.883e+00 
R2514t1337 n2515 n1338 R=6.226e+00 
R2514t2019 n2515 n2020 R=5.882e+00 
R2515t1699 n2516 n1700 R=7.696e+00 
R2516t169 n2517 n170 R=2.207e+01 
R2516t738 n2517 n739 R=4.718e+00 
R2516t183 n2517 n184 R=3.746e+01 
R2517t2162 n2518 n2163 R=1.085e+03 
R2517t1740 n2518 n1741 R=1.377e+02 
R2519t1228 n2520 n1229 R=4.050e+00 
R2520t2339 n2521 n2340 R=1.366e+01 
R2520t624 n2521 n625 R=4.366e+00 
R2521t390 n2522 n391 R=3.762e+00 
R2521t1357 n2522 n1358 R=2.892e+01 
R2522t2121 n2523 n2122 R=1.041e+01 
R2523t199 n2524 n200 R=1.154e+01 
R2524t489 n2525 n490 R=2.998e+00 
R2525t83 n2526 n84 R=1.241e+01 
R2525t1892 n2526 n1893 R=1.966e+01 
R2528t1938 n2529 n1939 R=2.457e+00 
R2529t62 n2530 n63 R=2.256e+00 
R2531t1399 n2532 n1400 R=2.195e+01 
R2531t1730 n2532 n1731 R=5.431e+00 
R2531t130 n2532 n131 R=4.171e+00 
R2532t383 n2533 n384 R=4.852e+01 
R2532t2291 n2533 n2292 R=3.230e+00 
R2533t1354 n2534 n1355 R=1.036e+01 
R2533t1000 n2534 n1001 R=4.194e+00 
R2533t81 n2534 n82 R=1.266e+01 
R2535t364 n2536 n365 R=6.473e+00 
R2537t177 n2538 n178 R=7.016e+01 
R2537t1042 n2538 n1043 R=3.110e+00 
R2538t371 n2539 n372 R=3.220e+00 
R2539t1912 n2540 n1913 R=5.544e+00 
R2540t2509 n2541 n2510 R=4.932e+00 
R2541t2513 n2542 n2514 R=2.125e+00 
R2541t1597 n2542 n1598 R=4.722e+00 
R2541t1661 n2542 n1662 R=1.139e+01 
R2542t195 n2543 n196 R=3.703e+00 
R2544t1334 n2545 n1335 R=4.736e+01 
R2547t1646 n2548 n1647 R=1.893e+01 
R2548t53 n2549 n54 R=2.598e+01 
R2549t2527 n2550 n2528 R=4.534e+00 
R2550t2510 n2551 n2511 R=1.025e+02 
R2550t783 n2551 n784 R=3.049e+00 
R2551t2328 n2552 n2329 R=4.616e+00 
R2551t163 n2552 n164 R=1.342e+01 
R2552t971 n2553 n972 R=2.214e+01 
R2552t916 n2553 n917 R=2.162e+01 
R2553t1249 n2554 n1250 R=7.967e+00 
R2554t68 n2555 n69 R=3.826e+00 
R2554t119 n2555 n120 R=2.961e+00 
R2554t1374 n2555 n1375 R=3.499e+01 
R2556t1068 n2557 n1069 R=7.436e+00 
R2557t1891 n2558 n1892 R=6.777e+00 
R2557t2535 n2558 n2536 R=2.706e+00 
R2559t1838 n2560 n1839 R=2.716e+01 
R2560t1577 n2561 n1578 R=3.881e+00 
R2561t2122 n2562 n2123 R=5.126e+00 
R2561t2496 n2562 n2497 R=3.266e+02 
R2561t1259 n2562 n1260 R=3.480e+00 
R2563t1656 n2564 n1657 R=7.893e+00 
R2563t1185 n2564 n1186 R=8.866e+00 
R2564t601 n2565 n602 R=7.171e+01 
R2565t1116 n2566 n1117 R=5.620e+00 
R2565t1468 n2566 n1469 R=2.895e+01 
R2566t2212 n2567 n2213 R=1.118e+01 
R2567t444 n2568 n445 R=2.974e+01 
R2567t968 n2568 n969 R=1.582e+01 
R2568t1912 n2569 n1913 R=1.431e+01 
R2568t2539 n2569 n2540 R=4.780e+00 
R2568t1104 n2569 n1105 R=5.710e+00 
R2570t1652 n2571 n1653 R=1.435e+01 
R2571t1084 n1 n1085 R=3.724e+00 
R2572t586 n2573 n587 R=1.572e+01 
R2572t1590 n2573 n1591 R=5.989e+00 
R2572t2542 n2573 n2543 R=6.382e+00 
R2573t785 n2574 n786 R=4.480e+00 
R2573t859 n2574 n860 R=1.305e+01 
R2573t541 n2574 n542 R=3.843e+00 
R2574t2230 n2575 n2231 R=4.815e+00 
R2575t1076 n2576 n1077 R=5.031e+00 
R2576t2333 n2577 n2334 R=6.414e+01 
R2576t719 n2577 n720 R=4.107e+00 
R2577t1662 n2578 n1663 R=2.852e+02 
R2577t1473 n2578 n1474 R=2.323e+01 
R2577t1751 n2578 n1752 R=5.188e+00 
R2577t2171 n2578 n2172 R=4.303e+00 
R2578t1243 n2579 n1244 R=3.347e+00 
R2578t2209 n2579 n2210 R=4.630e+00 
R2578t94 n2579 n95 R=5.158e+00 
R2579t2048 n2580 n2049 R=1.409e+01 
R2579t526 n2580 n527 R=1.662e+01 
R2580t345 n2581 n346 R=2.444e+00 
R2581t1514 n2582 n1515 R=2.343e+01 
R2581t243 n2582 n244 R=4.761e+00 
R2582t341 n2583 n342 R=9.409e+00 
R2583t2115 n2584 n2116 R=2.664e+01 
R2583t1508 n2584 n1509 R=2.808e+00 
R2583t516 n2584 n517 R=1.452e+01 
R2584t2182 n2585 n2183 R=2.257e+00 
R2584t399 n2585 n400 R=1.423e+01 
R2584t2123 n2585 n2124 R=1.957e+00 
R2586t14 n2587 n15 R=2.719e+00 
R2587t2263 n2588 n2264 R=7.397e+00 
R2587t1634 n2588 n1635 R=9.555e+00 
R2588t1859 n2589 n1860 R=2.758e+01 
R2588t1754 n2589 n1755 R=5.029e+00 
R2588t2470 n2589 n2471 R=8.714e+00 
R2588t1124 n2589 n1125 R=1.005e+01 
R2589t1112 n2590 n1113 R=4.467e+00 
R2589t1168 n2590 n1169 R=7.819e+00 
R2589t2458 n2590 n2459 R=1.470e+01 
R2589t1050 n2590 n1051 R=6.832e+01 
R2589t2434 n2590 n2435 R=3.433e+00 
R2590t187 n2591 n188 R=2.131e+02 
R2591t394 n2592 n395 R=4.598e+00 
R2592t1283 n2593 n1284 R=4.797e+00 
R2592t953 n2593 n954 R=1.772e+01 
R2592t971 n2593 n972 R=3.694e+01 
R2593t1280 n2594 n1281 R=4.145e+00 
R2596t551 n2597 n552 R=1.373e+01 
R2596t2102 n2597 n2103 R=5.275e+00 
R2598t1787 n2599 n1788 R=4.841e+00 
R2599t1385 n2600 n1386 R=1.626e+02 
R2601t1276 n2602 n1277 R=2.994e+00 
R2602t2262 n2603 n2263 R=1.290e+01 
R2602t216 n2603 n217 R=6.278e+00 
R2603t403 n2604 n404 R=1.208e+01 
R2603t1044 n2604 n1045 R=2.494e+00 
R2603t712 n2604 n713 R=6.131e+00 
R2603t2112 n2604 n2113 R=1.089e+01 
R2605t1575 n2606 n1576 R=9.190e+00 
R2605t1856 n2606 n1857 R=3.061e+00 
R2608t255 n2609 n256 R=8.112e+00 
R2610t2502 n1 n2503 R=2.176e+01 
R2611t1878 n2612 n1879 R=1.200e+01 
R2612t1365 n2613 n1366 R=6.079e+00 
R2612t1993 n2613 n1994 R=6.138e+00 
R2613t31 n2614 n32 R=3.647e+00 
R2614t2214 n2615 n2215 R=2.138e+01 
R2614t1 n2615 n2 R=4.972e+01 
R2614t1625 n2615 n1626 R=4.318e+00 
R2615t743 n2616 n744 R=4.068e+02 
R2615t385 n2616 n386 R=1.800e+01 
R2616t2045 n2617 n2046 R=5.405e+00 
R2616t2000 n2617 n2001 R=4.173e+00 
R2616t350 n2617 n351 R=3.071e+01 
R2617t393 n2618 n394 R=3.023e+00 
R2617t724 n2618 n725 R=8.153e+00 
R2617t977 n2618 n978 R=2.282e+01 
R2619t1681 n2620 n1682 R=1.786e+01 
R2619t1969 n2620 n1970 R=5.178e+01 
R2620t1719 n2621 n1720 R=4.144e+00 
R2622t2208 n2623 n2209 R=5.768e+00 
R2622t2282 n2623 n2283 R=1.312e+01 
R2622t1139 n2623 n1140 R=1.538e+01 
R2625t2507 n2626 n2508 R=8.544e+00 
R2625t983 n2626 n984 R=3.409e+00 
R2625t1570 n2626 n1571 R=4.214e+00 
R2627t2090 n2628 n2091 R=3.671e+00 
R2627t107 n2628 n108 R=5.325e+00 
R2628t433 n2629 n434 R=1.179e+01 
R2629t2442 n2630 n2443 R=6.657e+00 
R2630t1904 n2631 n1905 R=3.566e+00 
R2631t2432 n2632 n2433 R=5.319e+00 
R2631t744 n2632 n745 R=3.327e+00 
R2632t1614 n2633 n1615 R=2.079e+01 
R2633t631 n2634 n632 R=3.731e+01 
R2633t1513 n2634 n1514 R=1.914e+01 
R2634t1874 n2635 n1875 R=4.080e+01 
R2635t359 n2636 n360 R=6.548e+00 
R2635t1782 n2636 n1783 R=6.521e+01 
R2638t1592 n2639 n1593 R=2.945e+00 
R2638t2480 n2639 n2481 R=1.849e+00 
R2639t1794 n2640 n1795 R=5.889e+00 
R2640t540 n2641 n541 R=1.749e+01 
R2641t2365 n2642 n2366 R=1.377e+01 
R2642t2350 n2643 n2351 R=1.227e+01 
R2642t7 n2643 n8 R=5.422e+00 
R2643t1186 n2644 n1187 R=1.658e+01 
R2644t2612 n2645 n2613 R=2.692e+01 
R2645t2037 n2646 n2038 R=2.598e+00 
R2647t2192 n2648 n2193 R=5.614e+00 
R2647t191 n2648 n192 R=1.135e+01 
R2647t202 n2648 n203 R=4.147e+00 
R2648t1491 n2649 n1492 R=1.759e+01 
R2649t1841 n2650 n1842 R=1.307e+01 
R2650t138 n2651 n139 R=7.148e+00 
R2650t929 n2651 n930 R=1.284e+01 
R2651t565 n2652 n566 R=5.720e+00 
R2651t425 n2652 n426 R=1.581e+01 
R2651t843 n2652 n844 R=2.428e+01 
R2652t1368 n2653 n1369 R=2.127e+01 
R2652t1799 n2653 n1800 R=2.539e+01 
R2654t1636 n2655 n1637 R=4.251e+01 
R2654t2203 n2655 n2204 R=3.999e+00 
R2655t812 n2656 n813 R=7.933e+00 
R2655t498 n2656 n499 R=1.337e+01 
R2655t349 n2656 n350 R=8.921e+00 
R2655t2332 n2656 n2333 R=1.814e+01 
R2656t2040 n2657 n2041 R=2.255e+00 
R2657t2626 n2658 n2627 R=8.811e+00 
R2657t219 n2658 n220 R=6.743e+00 
R2658t2458 n2659 n2459 R=4.137e+00 
R2658t2589 n2659 n2590 R=2.264e+01 
R2658t1437 n2659 n1438 R=1.116e+01 
R2658t1714 n2659 n1715 R=1.424e+01 
R2658t1050 n2659 n1051 R=2.916e+01 
R2659t1674 n2660 n1675 R=2.083e+01 
R2660t2464 n2661 n2465 R=5.124e+01 
R2660t15 n2661 n16 R=6.770e+00 
R2660t1413 n2661 n1414 R=2.481e+01 
R2662t304 n2663 n305 R=4.780e+00 
R2663t1306 n2664 n1307 R=3.294e+00 
R2663t1004 n2664 n1005 R=2.975e+00 
R2665t1003 n2666 n1004 R=3.174e+01 
R2665t2189 n2666 n2190 R=1.531e+01 
R2666t511 n2667 n512 R=2.060e+00 
R2666t1902 n2667 n1903 R=2.507e+00 
R2667t1762 n2668 n1763 R=2.056e+01 
R2667t181 n2668 n182 R=5.838e+00 
R2667t2402 n2668 n2403 R=7.418e+01 
R2667t645 n2668 n646 R=6.664e+00 
R2668t1206 n2669 n1207 R=1.724e+01 
R2668t405 n2669 n406 R=7.445e+01 
R2670t2211 n2671 n2212 R=5.632e+00 
R2671t811 n2672 n812 R=2.482e+01 
R2672t1851 n2673 n1852 R=4.023e+01 
R2672t910 n2673 n911 R=4.277e+00 
R2672t485 n2673 n486 R=1.256e+01 
R2674t189 n2675 n190 R=8.977e+00 
R2675t509 n2676 n510 R=7.147e+00 
R2675t775 n2676 n776 R=4.273e+00 
R2676t2193 n2677 n2194 R=6.699e+01 
R2676t2223 n2677 n2224 R=1.956e+01 
R2676t380 n2677 n381 R=8.011e+00 
R2676t240 n2677 n241 R=1.279e+01 
R2677t1575 n2678 n1576 R=2.111e+01 
R2677t2605 n2678 n2606 R=9.011e+00 
R2677t1856 n2678 n1857 R=1.033e+01 
R2678t2093 n2679 n2094 R=1.139e+01 
R2678t2163 n2679 n2164 R=1.051e+01 
R2679t1286 n2680 n1287 R=1.806e+01 
R2679t1772 n2680 n1773 R=6.332e+00 
R2679t2128 n2680 n2129 R=2.666e+00 
R2680t672 n2681 n673 R=3.681e+00 
R2681t62 n2682 n63 R=2.852e+02 
R2681t2529 n2682 n2530 R=2.835e+01 
R2682t2657 n2683 n2658 R=3.402e+01 
R2682t2626 n2683 n2627 R=1.446e+01 
R2683t166 n2684 n167 R=3.151e+00 
R2685t2240 n2686 n2241 R=1.944e+00 
R2685t2545 n2686 n2546 R=5.385e+00 
R2685t1903 n2686 n1904 R=7.146e+00 
R2685t2105 n2686 n2106 R=4.448e+01 
R2686t2192 n2687 n2193 R=1.236e+01 
R2686t2647 n2687 n2648 R=1.405e+02 
R2686t873 n2687 n874 R=2.523e+00 
R2687t511 n2688 n512 R=5.659e+00 
R2687t1241 n2688 n1242 R=4.439e+00 
R2687t813 n2688 n814 R=2.600e+01 
R2687t1902 n2688 n1903 R=6.167e+01 
R2687t2666 n2688 n2667 R=2.095e+01 
R2688t2092 n2689 n2093 R=2.144e+01 
R2689t1843 n2690 n1844 R=4.867e+01 
R2689t691 n2690 n692 R=1.161e+01 
R2690t2177 n2691 n2178 R=6.192e+00 
R2690t63 n2691 n64 R=5.810e+00 
R2691t854 n2692 n855 R=3.454e+00 
R2692t841 n2693 n842 R=2.528e+00 
R2692t2391 n2693 n2392 R=4.142e+01 
R2693t948 n2694 n949 R=2.699e+02 
R2694t138 n2695 n139 R=1.588e+02 
R2694t849 n2695 n850 R=3.254e+00 
R2695t2317 n2696 n2318 R=6.422e+00 
R2695t1427 n2696 n1428 R=1.365e+01 
R2696t450 n2697 n451 R=3.983e+00 
R2697t1438 n2698 n1439 R=1.921e+01 
R2697t1773 n2698 n1774 R=5.771e+00 
R2697t2420 n2698 n2421 R=5.728e+00 
R2698t2669 n2699 n2670 R=1.790e+00 
R2699t2295 n2700 n2296 R=2.456e+02 
R2701t459 n2702 n460 R=2.004e+01 
R2701t1649 n2702 n1650 R=4.115e+00 
R2701t2036 n2702 n2037 R=2.749e+00 
R2702t727 n2703 n728 R=5.502e+01 
R2702t2032 n2703 n2033 R=2.495e+00 
R2702t1458 n2703 n1459 R=5.264e+01 
R2703t2486 n2704 n2487 R=8.819e+00 
R2704t458 n2705 n459 R=3.690e+01 
R2704t599 n2705 n600 R=3.712e+00 
R2704t915 n2705 n916 R=4.476e+01 
R2705t2567 n2706 n2568 R=7.518e+00 
R2705t182 n2706 n183 R=4.716e+00 
R2706t1569 n2707 n1570 R=2.475e+00 
R2707t944 n2708 n945 R=1.594e+01 
R2707t506 n2708 n507 R=9.931e+00 
R2707t131 n2708 n132 R=3.102e+02 
R2708t1200 n2709 n1201 R=1.175e+01 
R2708t281 n2709 n282 R=1.295e+01 
R2709t71 n2710 n72 R=1.822e+02 
R2709t687 n2710 n688 R=1.573e+01 
R2709t1380 n2710 n1381 R=4.475e+00 
R2710t1822 n2711 n1823 R=2.632e+00 
R2710t1384 n2711 n1385 R=9.728e+00 
R2711t242 n2712 n243 R=9.612e+00 
R2712t1213 n2713 n1214 R=1.359e+01 
R2714t952 n2715 n953 R=3.474e+00 
R2715t2362 n2716 n2363 R=5.334e+01 
R2715t2436 n2716 n2437 R=8.224e+00 
R2715t151 n2716 n152 R=8.442e+00 
R2716t1012 n2717 n1013 R=8.937e+00 
R2716t1250 n2717 n1251 R=4.776e+00 
R2717t2536 n2718 n2537 R=3.573e+00 
R2717t564 n2718 n565 R=9.094e+00 
R2718t556 n2719 n557 R=9.442e+00 
R2719t2233 n2720 n2234 R=1.134e+02 
R2720t593 n2721 n594 R=2.246e+00 
R2722t1182 n2723 n1183 R=7.435e+00 
R2722t2302 n2723 n2303 R=2.076e+00 
R2723t749 n2724 n750 R=6.970e+00 
R2724t536 n2725 n537 R=3.998e+00 
R2724t2027 n2725 n2028 R=1.046e+01 
R2725t1016 n2726 n1017 R=6.590e+00 
R2725t389 n2726 n390 R=3.941e+00 
R2726t1621 n2727 n1622 R=6.334e+00 
R2727t1779 n2728 n1 R=2.345e+01 
R2729t826 n2730 n827 R=1.868e+01 
R2729t875 n2730 n876 R=2.140e+01 
R2730t115 n2731 n116 R=7.335e+00 
R2730t1359 n2731 n1360 R=5.643e+00 
R2731t832 n2732 n833 R=5.377e+00 
R2731t1586 n2732 n1587 R=1.400e+01 
R2732t1553 n2733 n1554 R=1.266e+01 
R2733t38 n2734 n39 R=4.938e+01 
R2734t323 n2735 n324 R=4.183e+01 
R2734t79 n2735 n80 R=5.428e+01 
R2734t1744 n2735 n1745 R=3.076e+02 
R2734t1919 n2735 n1920 R=8.505e+00 
R2735t2636 n2736 n2637 R=2.795e+01 
R2735t2233 n2736 n2234 R=3.574e+00 
R2735t2719 n2736 n2720 R=7.523e+01 
R2737t1807 n2738 n1808 R=8.901e+00 
R2738t262 n2739 n263 R=3.306e+01 
R2739t701 n2740 n702 R=4.021e+02 
R2739t293 n2740 n294 R=1.225e+01 
R2742t1490 n2743 n1491 R=8.719e+00 
R2742t2630 n2743 n2631 R=7.389e+00 
R2742t1904 n2743 n1905 R=2.962e+00 
R2743t2437 n2744 n2438 R=3.721e+00 
R2744t141 n2745 n142 R=4.213e+01 
R2744t610 n2745 n611 R=7.810e+00 
R2744t2604 n2745 n2605 R=2.750e+01 
R2745t1302 n2746 n1303 R=2.317e+01 
R2746t966 n2747 n967 R=4.977e+00 
R2746t729 n2747 n730 R=6.762e+01 
R2746t359 n2747 n360 R=1.159e+01 
R2746t2411 n2747 n2412 R=4.713e+00 
R2747t1118 n1 n1119 R=4.170e+00 
R2749t2378 n2750 n2379 R=2.730e+01 
R2750t896 n2751 n897 R=2.979e+01 
R2751t2679 n2752 n2680 R=8.908e+00 
R2751t162 n2752 n163 R=8.984e+00 
R2752t794 n2753 n795 R=3.013e+01 
R2752t585 n2753 n586 R=6.976e+00 
R2753t167 n2754 n168 R=2.723e+00 
R2753t1934 n2754 n1935 R=6.624e+01 
R2755t115 n2756 n116 R=7.731e+00 
R2755t1819 n2756 n1820 R=4.884e+00 
R2755t1359 n2756 n1360 R=8.792e+00 
R2755t2730 n2756 n2731 R=5.027e+00 
R2756t2149 n2757 n2150 R=3.507e+00 
R2756t1764 n2757 n1765 R=5.252e+00 
R2757t2233 n2758 n2234 R=9.884e+00 
R2757t2636 n2758 n2637 R=1.834e+01 
R2758t931 n2759 n932 R=5.964e+02 
R2758t1574 n2759 n1575 R=5.073e+01 
R2759t1333 n2760 n1334 R=1.281e+01 
R2759t1856 n2760 n1857 R=1.813e+02 
R2759t2605 n2760 n2606 R=3.177e+00 
R2761t220 n2762 n221 R=2.593e+00 
R2762t820 n2763 n821 R=4.033e+01 
R2762t2599 n2763 n2600 R=3.949e+01 
R2763t1614 n2764 n1615 R=6.142e+01 
R2763t2632 n2764 n2633 R=3.521e+00 
R2763t552 n2764 n553 R=3.283e+01 
R2764t2358 n2765 n2359 R=7.405e+00 
R2765t1775 n2766 n1776 R=4.721e+00 
R2765t2168 n2766 n2169 R=8.595e+01 
R2767t2095 n2768 n2096 R=4.291e+01 
R2768t1631 n2769 n1632 R=2.103e+01 
R2768t302 n2769 n303 R=5.182e+00 
R2768t1801 n2769 n1802 R=2.693e+00 
R2769t2640 n2770 n2641 R=3.252e+01 
R2770t801 n2771 n802 R=6.395e+01 
R2770t22 n2771 n23 R=1.034e+01 
R2770t1387 n2771 n1388 R=6.637e+00 
R2771t2458 n2772 n2459 R=7.395e+01 
R2771t1196 n2772 n1197 R=3.942e+00 
R2771t1458 n2772 n1459 R=4.212e+00 
R2771t1437 n2772 n1438 R=1.296e+01 
R2773t1460 n2774 n1461 R=2.109e+01 
R2773t1520 n2774 n1521 R=9.057e+00 
R2774t2337 n2775 n2338 R=3.624e+00 
R2774t1498 n2775 n1499 R=4.338e+00 
R2775t1488 n2776 n1489 R=7.078e+00 
R2776t1312 n2777 n1313 R=1.842e+01 
R2777t687 n2778 n688 R=3.049e+00 
R2777t2709 n2778 n2710 R=1.620e+01 
R2778t1742 n2779 n1743 R=7.280e+00 
R2778t1235 n2779 n1236 R=5.081e+00 
R2778t1224 n2779 n1225 R=3.633e+01 
R2779t2086 n2780 n2087 R=4.951e+00 
R2779t1893 n2780 n1894 R=1.958e+01 
R2780t776 n2781 n777 R=2.678e+00 
R2781t2544 n2782 n2545 R=5.393e+00 
R2781t1626 n2782 n1627 R=4.950e+00 
R2784t121 n2785 n122 R=5.685e+00 
R2785t1957 n2786 n1958 R=7.193e+00 
R2785t2251 n2786 n2252 R=4.355e+00 
R2785t284 n2786 n285 R=8.503e+01 
R2785t662 n2786 n663 R=3.242e+02 
R2785t1539 n2786 n1540 R=6.768e+00 
R2786t786 n2787 n787 R=6.209e+00 
R2786t859 n2787 n860 R=2.016e+03 
R2786t172 n2787 n173 R=5.411e+01 
R2788t815 n2789 n816 R=1.115e+01 
R2788t1807 n2789 n1808 R=9.844e+00 
R2788t432 n2789 n433 R=4.579e+00 
R2789t34 n2790 n35 R=6.250e+00 
R2791t820 n2792 n821 R=6.266e+00 
R2791t2762 n2792 n2763 R=7.329e+00 
R2792t1763 n2793 n1764 R=1.710e+00 
R2792t1599 n2793 n1600 R=1.139e+01 
R2793t442 n2794 n443 R=2.040e+01 
R2794t1362 n2795 n1363 R=2.235e+01 
R2794t2382 n2795 n2383 R=1.611e+01 
R2794t1269 n2795 n1270 R=1.142e+01 
R2795t2212 n2796 n2213 R=3.453e+01 
R2795t1696 n2796 n1697 R=1.309e+01 
R2795t348 n2796 n349 R=1.903e+01 
R2795t2499 n2796 n2500 R=6.157e+00 
R2796t96 n2797 n97 R=2.782e+00 
R2796t155 n2797 n156 R=2.730e+01 
R2797t2218 n2798 n2219 R=4.309e+00 
R2798t774 n2799 n775 R=5.411e+00 
R2798t2029 n2799 n2030 R=4.580e+00 
R2798t1282 n2799 n1283 R=2.674e+02 
R2799t1651 n2800 n1652 R=3.760e+00 
R2800t2427 n2801 n2428 R=1.620e+01 
R2800t207 n2801 n208 R=2.964e+00 
R2800t2151 n2801 n2152 R=6.010e+00 
R2801t2265 n2802 n2266 R=2.894e+00 
R2801t1688 n2802 n1689 R=2.543e+01 
R2801t40 n2802 n41 R=1.495e+01 
R2801t1992 n2802 n1993 R=4.279e+00 
R2802t907 n2803 n908 R=1.903e+01 
R2802t251 n2803 n252 R=7.506e+01 
R2803t2362 n2804 n2363 R=1.477e+00 
R2803t2715 n2804 n2716 R=2.665e+01 
R2803t173 n2804 n174 R=2.316e+00 
R2804t1877 n2805 n1878 R=2.725e+00 
R2806t2193 n2807 n2194 R=7.116e+00 
R2807t1510 n2808 n1511 R=8.695e+00 
R2808t1242 n2809 n1243 R=7.393e+01 
R2808t1267 n2809 n1268 R=2.140e+00 
R2809t1588 n2810 n1589 R=5.925e+00 
R2810t1175 n2811 n1176 R=7.974e+01 
R2810t2259 n2811 n2260 R=2.511e+00 
R2810t417 n2811 n418 R=8.614e+00 
R2811t631 n2812 n632 R=8.220e+00 
R2811t2633 n2812 n2634 R=2.424e+00 
R2811t1513 n2812 n1514 R=7.139e+01 
R2812t2312 n2813 n2313 R=1.661e+01 
R2812t1199 n2813 n1200 R=1.038e+01 
R2813t476 n2814 n477 R=6.017e+00 
R2813t2260 n2814 n2261 R=4.049e+00 
R2813t1397 n2814 n1398 R=2.892e+01 
R2814t2316 n2815 n2317 R=1.132e+01 
R2815t2580 n2816 n2581 R=9.514e+01 
R2815t139 n2816 n140 R=5.470e+02 
R2816t542 n2817 n543 R=1.547e+01 
R2818t2234 n2819 n2235 R=3.931e+01 
R2818t366 n2819 n367 R=6.797e+00 
R2818t211 n2819 n212 R=1.853e+01 
R2818t1947 n2819 n1948 R=4.597e+00 
R2820t886 n2821 n887 R=1.856e+01 
R2820t2688 n2821 n2689 R=7.094e+01 
R2821t1034 n2822 n1035 R=9.337e+01 
R2821t1240 n2822 n1241 R=1.894e+01 
R2821t2061 n2822 n2062 R=2.950e+00 
R2822t554 n2823 n555 R=1.215e+01 
R2822t142 n2823 n143 R=4.850e+00 
R2823t1545 n2824 n1546 R=9.176e+00 
R2823t466 n2824 n467 R=2.327e+01 
R2824t2313 n2825 n2314 R=1.227e+01 
R2825t726 n2826 n727 R=3.339e+00 
R2826t814 n2827 n815 R=4.068e+00 
R2826t2083 n2827 n2084 R=5.780e+00 
R2827t2497 n2828 n2498 R=2.805e+00 
R2827t1087 n2828 n1088 R=8.539e+00 
R2828t2164 n2829 n2165 R=6.810e+00 
R2830t2636 n2831 n2637 R=2.237e+00 
R2830t2757 n2831 n2758 R=3.344e+00 
R2830t2735 n2831 n2736 R=1.913e+01 
R2830t2233 n2831 n2234 R=7.352e+00 
R2831t2382 n2832 n2383 R=1.422e+02 
R2831t2790 n2832 n2791 R=5.983e+00 
R2831t2326 n2832 n2327 R=3.856e+01 
R2832t2775 n2833 n2776 R=5.643e+00 
R2833t1380 n2834 n1381 R=4.018e+00 
R2833t930 n2834 n931 R=6.945e+00 
R2834t1344 n2835 n1345 R=9.008e+00 
R2834t1843 n2835 n1844 R=1.154e+01 
R2836t1131 n2837 n1132 R=8.348e+01 
R2836t1302 n2837 n1303 R=1.905e+01 
R2837t1280 n2838 n1281 R=2.543e+01 
R2837t1358 n2838 n1359 R=4.178e+00 
R2838t1484 n2839 n1 R=4.816e+00 
R2839t1990 n2840 n1991 R=4.069e+01 
R2839t1339 n2840 n1340 R=3.008e+01 
R2840t761 n2841 n762 R=5.421e+01 
R2840t1421 n2841 n1422 R=1.723e+02 
R2841t23 n2842 n24 R=7.866e+00 
R2841t1338 n2842 n1339 R=1.506e+01 
R2841t471 n2842 n472 R=1.828e+01 
R2841t2144 n2842 n2145 R=8.257e+00 
R2842t2585 n2843 n2586 R=1.205e+01 
R2843t2034 n2844 n2035 R=9.145e+00 
R2844t2780 n2845 n2781 R=1.194e+02 
R2845t1615 n2846 n1616 R=2.234e+01 
R2845t1799 n2846 n1800 R=4.338e+00 
R2845t2652 n2846 n2653 R=1.501e+01 
R2846t2528 n2847 n2529 R=1.143e+01 
R2846t1938 n2847 n1939 R=8.775e+01 
R2846t1100 n2847 n1101 R=4.202e+00 
R2846t872 n2847 n873 R=2.806e+01 
R2846t295 n2847 n296 R=2.990e+00 
R2847t1439 n2848 n1440 R=4.129e+00 
R2847t1652 n2848 n1653 R=7.032e+00 
R2849t1385 n2850 n1386 R=3.085e+01 
R2850t1087 n1 n1088 R=3.651e+00 
R2851t1638 n2852 n1639 R=4.679e+00 
R2851t2100 n2852 n2101 R=1.007e+01 
R2851t1777 n2852 n1778 R=6.009e+00 
R2852t420 n2853 n421 R=1.337e+01 
R2853t452 n2854 n453 R=2.248e+02 
R2853t796 n2854 n797 R=6.872e+00 
R2855t1602 n2856 n1603 R=2.763e+02 
R2856t1971 n2857 n1972 R=1.998e+01 
R2856t708 n2857 n709 R=2.905e+01 
R2857t101 n2858 n102 R=5.822e+00 
R2858t2284 n2859 n2285 R=4.097e+00 
R2858t442 n2859 n443 R=4.227e+01 
R2858t2793 n2859 n2794 R=3.032e+00 
R2859t1376 n2860 n1377 R=1.760e+00 
R2860t2525 n2861 n2526 R=8.512e+00 
R2860t1288 n2861 n1289 R=1.976e+01 
R2860t345 n2861 n346 R=1.482e+01 
R2860t2002 n2861 n2003 R=5.754e+00 
R2861t2632 n2862 n2633 R=8.439e+00 
R2861t1614 n2862 n1615 R=2.605e+00 
R2863t2192 n2864 n2193 R=6.087e+00 
R2863t2686 n2864 n2687 R=7.550e+00 
R2863t505 n2864 n506 R=6.210e+00 
R2863t539 n2864 n540 R=2.048e+01 
R2864t2222 n2865 n2223 R=1.547e+02 
R2864t1341 n2865 n1342 R=3.989e+00 
R2864t1231 n2865 n1232 R=2.858e+00 
R2865t968 n2866 n969 R=8.914e+00 
R2865t608 n2866 n609 R=4.101e+00 
R2866t1385 n2867 n1386 R=7.261e+00 
R2866t2307 n2867 n2308 R=6.937e+00 
R2866t2599 n2867 n2600 R=5.695e+00 
R2866t2762 n2867 n2763 R=7.164e+00 
R2868t2641 n2869 n2642 R=1.240e+02 
R2868t1041 n2869 n1042 R=3.337e+01 
R2869t2417 n1 n2418 R=2.884e+00 
R2870t1212 n2871 n1213 R=6.069e+00 
R2870t363 n2871 n364 R=8.474e+00 
R2870t2033 n2871 n2034 R=7.114e+01 
R2870t2142 n2871 n2143 R=3.623e+00 
R2871t2538 n2872 n2539 R=3.439e+00 
R2871t2247 n2872 n2248 R=1.417e+01 
R2872t1883 n2873 n1884 R=3.402e+01 
R2873t1939 n2874 n1940 R=9.674e+00 
R2873t127 n2874 n128 R=4.398e+00 
R2873t2656 n2874 n2657 R=2.422e+01 
R2873t2040 n2874 n2041 R=5.452e+00 
R2873t2358 n2874 n2359 R=4.190e+01 
R2874t1806 n2875 n1807 R=6.171e+01 
R2875t629 n2876 n630 R=2.997e+01 
R2876t2442 n2877 n2443 R=7.006e+00 
R2876t2629 n2877 n2630 R=1.042e+01 
R2877t177 n2878 n178 R=1.480e+01 
R2877t2537 n2878 n2538 R=6.166e+00 
R2878t1636 n2879 n1637 R=1.456e+01 
R2879t1258 n2880 n1259 R=8.751e+00 
R2879t1716 n2880 n1717 R=5.688e+00 
R2879t1980 n2880 n1981 R=5.119e+00 
R2879t1622 n2880 n1623 R=2.885e+02 
R2880t359 n2881 n360 R=5.902e+00 
R2880t2635 n2881 n2636 R=7.695e+01 
R2882t2606 n2883 n2607 R=4.756e+01 
R2882t1623 n2883 n1624 R=1.146e+01 
R2882t1188 n2883 n1189 R=1.625e+01 
R2883t2566 n2884 n2567 R=6.573e+00 
R2884t2588 n2885 n2589 R=1.034e+01 
R2884t1559 n2885 n1560 R=1.936e+02 
R2884t1174 n2885 n1175 R=5.920e+00 
R2884t1124 n2885 n1125 R=5.893e+00 
R2886t1654 n2887 n1655 R=1.106e+01 
R2887t2527 n2888 n2528 R=5.373e+00 
R2887t2549 n2888 n2550 R=1.258e+01 
R2888t45 n2889 n46 R=2.882e+01 
R2888t544 n2889 n545 R=1.553e+01 
R2889t1101 n2890 n1102 R=1.259e+02 
R2889t2264 n2890 n2265 R=1.392e+01 
R2889t1309 n2890 n1310 R=8.744e+00 
R2890t1206 n2891 n1207 R=1.016e+01 
R2890t2469 n2891 n2470 R=8.299e+00 
R2890t2426 n2891 n2427 R=3.942e+00 
R2890t353 n2891 n354 R=1.186e+02 
R2891t715 n2892 n716 R=6.546e+00 
R2892t1909 n2893 n1910 R=4.588e+00 
R2892t48 n2893 n49 R=4.563e+00 
R2894t2544 n2895 n2545 R=1.692e+01 
R2895t229 n2896 n230 R=6.483e+00 
R2896t1215 n2897 n1216 R=1.912e+01 
R2896t524 n2897 n525 R=3.210e+01 
R2897t1744 n2898 n1745 R=2.119e+01 
R2897t1944 n2898 n1945 R=1.049e+03 
R2897t2894 n2898 n2895 R=4.688e+00 
R2898t342 n2899 n343 R=1.764e+00 
R2899t833 n2900 n834 R=1.730e+01 
R2901t1195 n2902 n1196 R=1.602e+01 
R2902t979 n2903 n980 R=1.485e+01 
R2902t860 n2903 n861 R=5.232e+01 
R2902t2433 n2903 n2434 R=5.439e+00 
R2902t243 n2903 n244 R=1.547e+01 
R2903t2200 n2904 n2201 R=4.825e+00 
R2903t1260 n2904 n1261 R=5.268e+00 
R2904t341 n2905 n342 R=3.660e+01 
R2904t2582 n2905 n2583 R=6.342e+00 
R2905t1788 n2906 n1789 R=2.389e+00 
R2906t2126 n2907 n2127 R=8.213e+01 
R2906t637 n2907 n638 R=1.415e+01 
R2906t264 n2907 n265 R=2.461e+01 
R2906t1416 n2907 n1417 R=4.983e+00 
R2906t1519 n2907 n1520 R=1.613e+01 
R2906t877 n2907 n878 R=7.157e+00 
R2907t1505 n2908 n1506 R=1.827e+00 
R2907t2767 n2908 n2768 R=5.503e+00 
R2909t1735 n2910 n1736 R=4.578e+00 
R2909t543 n2910 n544 R=6.062e+01 
R2910t1257 n2911 n1258 R=4.250e+01 
R2912t759 n2913 n760 R=9.177e+00 
R2912t1594 n2913 n1595 R=1.009e+01 
R2913t1674 n2914 n1675 R=8.063e+00 
R2914t606 n2915 n607 R=2.342e+01 
R2915t2333 n2916 n2334 R=9.032e+00 
R2915t1364 n2916 n1365 R=7.104e+00 
R2916t735 n2917 n736 R=6.274e+00 
R2916t2721 n2917 n2722 R=2.141e+01 
R2916t163 n2917 n164 R=1.191e+01 
R2917t2478 n2918 n2479 R=1.062e+01 
R2918t461 n2919 n462 R=1.553e+01 
R2918t2114 n2919 n2115 R=1.100e+01 
R2918t995 n2919 n996 R=4.480e+00 
R2919t561 n2920 n562 R=5.425e+00 
R2920t736 n2921 n737 R=2.491e+00 
R2920t878 n2921 n879 R=2.213e+01 
R2920t2239 n2921 n2240 R=4.232e+00 
R2922t1346 n2923 n1347 R=5.356e+00 
R2922t784 n2923 n785 R=5.401e+01 
R2923t1890 n2924 n1891 R=4.080e+00 
R2923t1608 n2924 n1609 R=5.553e+00 
R2924t407 n2925 n408 R=2.652e+01 
R2924t1795 n2925 n1796 R=1.158e+02 
R2925t727 n2926 n728 R=2.786e+01 
R2925t2304 n2926 n2305 R=1.374e+01 
R2926t2298 n2927 n2299 R=3.879e+01 
R2926t2093 n2927 n2094 R=4.869e+00 
R2927t510 n2928 n511 R=4.099e+00 
R2928t2194 n2929 n2195 R=7.264e+00 
R2929t1480 n2930 n1481 R=1.044e+02 
R2929t65 n2930 n66 R=2.479e+00 
R2930t908 n2931 n909 R=3.894e+00 
R2931t2881 n2932 n2882 R=6.903e+00 
R2932t769 n2933 n770 R=5.321e+00 
R2932t2783 n2933 n2784 R=7.370e+00 
R2933t1990 n2934 n1991 R=6.046e+01 
R2933t2360 n2934 n2361 R=1.046e+02 
R2933t2301 n2934 n2302 R=2.922e+02 
R2934t2325 n2935 n2326 R=7.140e+02 
R2934t134 n2935 n135 R=2.205e+00 
R2935t2442 n2936 n2443 R=3.173e+01 
R2935t2293 n2936 n2294 R=1.349e+01 
R2935t2629 n2936 n2630 R=1.231e+01 
R2936t1873 n2937 n1874 R=9.345e+00 
R2937t1343 n2938 n1344 R=7.092e+00 
R2937t1792 n2938 n1793 R=4.707e+00 
R2938t428 n2939 n429 R=1.060e+01 
R2938t1477 n2939 n1478 R=3.834e+00 
R2940t663 n2941 n664 R=6.763e+00 
R2942t2777 n2943 n2778 R=3.422e+00 
R2942t687 n2943 n688 R=3.918e+01 
R2944t2848 n2945 n2849 R=5.558e+01 
R2945t2939 n2946 n2940 R=6.015e+00 
R2946t2829 n2947 n2830 R=5.678e+00 
R2947t2840 n2948 n2841 R=3.675e+00 
R2947t761 n2948 n762 R=2.065e+01 
R2948t339 n2949 n340 R=2.606e+00 
R2948t1739 n2949 n1740 R=2.446e+00 
R2948t1545 n2949 n1546 R=7.429e+00 
R2949t1466 n2950 n1467 R=3.141e+00 
R2950t186 n2951 n187 R=1.708e+01 
R2950t321 n2951 n322 R=3.096e+00 
R2950t1785 n2951 n1786 R=4.563e+00 
R2950t2071 n2951 n2072 R=5.249e+00 
R2951t58 n2952 n59 R=5.354e+00 
R2951t457 n2952 n458 R=1.073e+01 
R2951t767 n2952 n768 R=4.424e+01 
R2951t45 n2952 n46 R=7.335e+00 
R2952t1867 n2953 n1868 R=2.139e+01 
R2953t2667 n2954 n2668 R=4.832e+01 
R2953t645 n2954 n646 R=3.982e+00 
R2953t2245 n2954 n2246 R=1.310e+01 
R2954t2709 n2955 n2710 R=7.564e+00 
R2955t1373 n2956 n1374 R=2.271e+01 
R2956t2341 n2957 n2342 R=3.230e+00 
R2957t1549 n2958 n1550 R=3.642e+00 
R2957t567 n2958 n568 R=4.856e+00 
R2958t2673 n2959 n2674 R=2.564e+01 
R2959t854 n2960 n855 R=4.867e+00 
R2959t2504 n2960 n2505 R=2.951e+01 
R2960t161 n2961 n162 R=1.202e+03 
R2960t1682 n2961 n1683 R=5.160e+01 
R2960t2736 n2961 n2737 R=8.345e+00 
R2961t2002 n2962 n2003 R=3.663e+00 
R2961t345 n2962 n346 R=5.238e+00 
R2961t2580 n2962 n2581 R=3.631e+01 
R2963t535 n2964 n536 R=2.901e+01 
R2963t1910 n2964 n1911 R=3.158e+01 
R2963t759 n2964 n760 R=1.170e+01 
R2963t2912 n2964 n2913 R=6.831e+00 
R2965t676 n2966 n677 R=8.529e+00 
R2966t643 n2967 n644 R=7.178e+00 
R2966t2931 n2967 n2932 R=2.617e+00 
R2966t2881 n2967 n2882 R=3.320e+01 
R2967t2378 n2968 n2379 R=4.786e+00 
R2967t2927 n2968 n2928 R=5.506e+01 
R2969t1304 n2970 n1305 R=3.119e+00 
R2971t1389 n2972 n1390 R=1.106e+01 
R2972t34 n2973 n35 R=6.913e+01 
R2972t2789 n2973 n2790 R=1.426e+01 
R2973t1849 n2974 n1850 R=2.019e+00 
R2974t1028 n2975 n1029 R=3.609e+00 
R2975t76 n2976 n77 R=3.877e+00 
R2975t1267 n2976 n1268 R=5.552e+01 
R2975t1242 n2976 n1243 R=6.482e+00 
R2976t1378 n2977 n1379 R=1.895e+00 
R2978t1127 n2979 n1128 R=2.368e+01 
R2979t1807 n2980 n1808 R=2.185e+01 
R2979t815 n2980 n816 R=2.415e+00 
R2979t2788 n2980 n2789 R=2.677e+01 
R2980t1500 n2981 n1501 R=3.374e+00 
R2980t2091 n2981 n1 R=3.095e+00 
R2980t1154 n2981 n1 R=9.673e+00 
R2980t1037 n2981 n1038 R=4.128e+00 
R2981t1404 n2982 n1405 R=5.226e+00 
R2981t177 n2982 n178 R=8.583e+00 
R2982t1118 n2983 n1119 R=1.022e+01 
R2982t2747 n2983 n1 R=1.179e+02 
R2982t1655 n2983 n1656 R=7.170e+00 
R2982t704 n2983 n705 R=3.361e+00 
R2983t1194 n2984 n1195 R=2.031e+01 
R2983t994 n2984 n995 R=8.118e+00 
R2983t1736 n2984 n1737 R=4.553e+00 
R2984t2483 n2985 n2484 R=2.246e+02 
R2985t1024 n2986 n1025 R=9.530e+01 
R2985t1086 n2986 n1087 R=3.629e+00 
R2986t314 n2987 n315 R=3.881e+00 
R2989t1701 n2990 n1702 R=2.213e+00 
R2990t726 n2991 n727 R=2.109e+01 
R2991t2443 n2992 n2444 R=1.074e+01 
R2991t2400 n2992 n2401 R=2.584e+01 
R2993t2507 n2994 n2508 R=1.414e+01 
R2993t267 n2994 n268 R=3.222e+00 
R2994t2787 n2995 n2788 R=3.114e+01 
R2995t2690 n2996 n2691 R=2.428e+00 
R2995t2597 n2996 n2598 R=2.604e+00 
R2996t46 n2997 n47 R=4.831e+01 
R2996t1115 n2997 n1116 R=2.216e+02 
R2997t2194 n2998 n2195 R=6.510e+00 
R2997t2928 n2998 n2929 R=5.405e+00 
R2999t1068 n3000 n1069 R=3.308e+01 
R3000t219 n3001 n220 R=5.447e+00 
R3000t1142 n3001 n1143 R=3.720e+01 
R3000t831 n3001 n832 R=8.586e+00 
R3001t956 n3002 n957 R=3.584e+01 
R3001t2662 n3002 n2663 R=4.435e+00 
R3002t1626 n3003 n1627 R=1.499e+01 
R3002t2781 n3003 n2782 R=7.174e+00 
R3003t806 n3004 n807 R=3.270e+00 
R3003t1224 n3004 n1225 R=5.846e+03 
R3004t493 n3005 n494 R=2.552e+00 
R3005t2020 n3006 n2021 R=5.700e+01 
R3005t12 n3006 n13 R=5.524e+00 
R3006t2357 n3007 n2358 R=5.395e+00 
R3006t1949 n3007 n1950 R=5.838e+00 
R3007t1080 n3008 n1081 R=7.642e+00 
R3007t2505 n3008 n2506 R=7.305e+00 
R3008t1602 n3009 n1603 R=1.115e+01 
R3008t1537 n3009 n1538 R=5.133e+00 
R3010t1446 n3011 n1447 R=7.079e+00 
R3010t659 n3011 n660 R=2.763e+01 
R3010t693 n3011 n694 R=3.239e+00 
R3011t1475 n3012 n1476 R=2.258e+01 
R3011t471 n3012 n472 R=1.856e+01 
R3012t1491 n3013 n1492 R=6.274e+01 
R3013t1636 n3014 n1637 R=3.402e+02 
R3013t2654 n3014 n2655 R=1.079e+01 
R3013t2312 n3014 n2313 R=1.255e+02 
R3013t2812 n3014 n2813 R=6.382e+00 
R3014t1521 n3015 n1522 R=1.137e+01 
R3014t827 n3015 n828 R=2.073e+01 
R3015t431 n3016 n432 R=4.215e+00 
R3016t954 n3017 n955 R=3.051e+00 
R3017t2325 n3018 n2326 R=3.899e+00 
R3017t1099 n3018 n1100 R=4.115e+00 
R3018t956 n3019 n957 R=6.135e+00 
R3018t2364 n3019 n2365 R=6.141e+02 
R3019t2065 n3020 n2066 R=3.938e+00 
R3019t766 n3020 n767 R=5.040e+00 
R3019t1668 n3020 n1669 R=5.239e+00 
R3020t2501 n3021 n2502 R=4.693e+01 
R3020t800 n3021 n801 R=4.424e+00 
R3020t1324 n3021 n1325 R=6.997e+00 
R3021t1131 n3022 n1132 R=6.719e+00 
R3021t1974 n3022 n1975 R=1.548e+02 
R3021t2836 n3022 n2837 R=1.181e+01 
R3022t1743 n3023 n1744 R=2.692e+00 
R3022t394 n3023 n395 R=4.924e+01 
R3023t2335 n3024 n2336 R=5.159e+00 
R3025t2209 n3026 n2210 R=2.640e+01 
R3025t1766 n3026 n1767 R=3.550e+00 
R3025t1638 n3026 n1639 R=1.856e+01 
R3025t2851 n3026 n2852 R=1.368e+01 
R3025t2100 n3026 n2101 R=1.400e+01 
R3026t1435 n3027 n1436 R=4.134e+00 
R3027t1126 n3028 n1127 R=6.613e+01 
R3027t1593 n3028 n1594 R=7.433e+01 
R3027t2052 n3028 n2053 R=2.394e+01 
R3027t2289 n3028 n2290 R=8.659e+00 
R3028t1723 n3029 n1724 R=3.166e+01 
R3028t1978 n3029 n1979 R=1.327e+01 
R3028t2391 n3029 n2392 R=5.122e+00 
R3029t881 n3030 n882 R=6.197e+00 
R3029t373 n3030 n374 R=7.416e+01 
R3030t1501 n3031 n1502 R=2.551e+01 
R3030t1029 n3031 n1030 R=2.516e+01 
R3031t1079 n3032 n1080 R=1.136e+01 
R3032t2421 n3033 n2422 R=1.050e+01 
R3033t1233 n3034 n1234 R=1.273e+01 
R3033t2076 n3034 n2077 R=1.311e+01 
R3033t2491 n3034 n2492 R=5.034e+01 
R3033t2402 n3034 n2403 R=3.475e+01 
R3034t711 n3035 n712 R=1.152e+01 
R3034t2477 n3035 n2478 R=1.914e+01 
R3034t634 n3035 n635 R=8.559e+00 
R3035t2732 n3036 n2733 R=6.234e+00 
R3036t2210 n3037 n2211 R=5.733e+00 
R3036t1158 n3037 n1159 R=6.096e+00 
R3037t1290 n3038 n1291 R=3.022e+00 
R3037t1872 n3038 n1873 R=6.783e+00 
R3038t945 n3039 n946 R=5.481e+00 
R3038t2286 n3039 n2287 R=4.522e+00 
R3038t530 n3039 n531 R=1.529e+01 
R3038t703 n3039 n704 R=7.929e+01 
R3039t1625 n1 n1626 R=7.068e+00 
R3041t577 n3042 n578 R=1.250e+01 
R3041t991 n3042 n992 R=1.937e+01 
R3041t2997 n3042 n2998 R=9.580e+00 
R3042t1662 n3043 n1663 R=9.783e+00 
R3042t353 n3043 n354 R=6.017e+00 
R3043t123 n3044 n124 R=2.294e+01 
R3043t1767 n3044 n1768 R=6.136e+00 
R3044t710 n3045 n711 R=4.153e+00 
R3045t2650 n3046 n2651 R=3.304e+00 
R3045t929 n3046 n930 R=1.214e+01 
R3047t2390 n3048 n2391 R=3.344e+00 
R3048t1783 n3049 n1784 R=1.325e+01 
R3049t738 n3050 n739 R=1.837e+01 
R3049t169 n3050 n170 R=2.421e+00 
R3049t1470 n3050 n1471 R=2.524e+01 
R3050t2135 n3051 n2136 R=1.068e+04 
R3050t1510 n3051 n1511 R=2.568e+01 
R3051t2639 n3052 n2640 R=7.572e+00 
R3052t2455 n3053 n2456 R=2.162e+01 
R3052t212 n3053 n213 R=7.928e+00 
R3053t1125 n3054 n1126 R=1.459e+01 
R3053t2031 n3054 n2032 R=2.471e+00 
R3054t1587 n3055 n1588 R=1.141e+03 
R3055t919 n3056 n920 R=5.013e+00 
R3055t2968 n3056 n2969 R=1.100e+01 
R3056t725 n3057 n726 R=9.645e+00 
R3056t1445 n3057 n1446 R=2.379e+00 
R3057t2113 n3058 n2114 R=2.715e+00 
R3057t1729 n3058 n1730 R=6.252e+00 
R3057t2238 n3058 n2239 R=8.720e+01 
R3058t324 n3059 n325 R=7.942e+00 
R3058t2898 n3059 n2899 R=8.125e+00 
R3058t342 n3059 n343 R=2.137e+01 
R3058t2256 n3059 n2257 R=5.543e+02 
R3058t1884 n3059 n1885 R=4.581e+00 
R3058t422 n3059 n423 R=7.696e+00 
R3059t962 n3060 n963 R=5.200e+00 
R3060t319 n3061 n320 R=1.329e+01 
R3060t1005 n3061 n1006 R=1.138e+01 
R3060t568 n3061 n569 R=3.841e+00 
R3060t388 n3061 n389 R=4.621e+00 
R3062t1452 n3063 n1453 R=3.700e+00 
R3062t196 n3063 n197 R=1.125e+01 
R3062t2033 n3063 n2034 R=1.186e+01 
R3063t448 n3064 n449 R=9.446e+00 
R3064t1183 n3065 n1184 R=1.810e+01 
R3064t2867 n3065 n2868 R=4.130e+00 
R3064t1703 n3065 n1704 R=2.184e+01 
R3065t1892 n3066 n1893 R=8.641e+00 
R3065t1026 n3066 n1027 R=1.604e+01 
R3066t1651 n3067 n1652 R=1.426e+01 
R3066t2799 n3067 n2800 R=4.700e+00 
R3066t1045 n3067 n1046 R=2.888e+02 
R3066t1213 n3067 n1214 R=6.449e+00 
R3066t2712 n3067 n2713 R=1.636e+01 
R3067t427 n3068 n428 R=2.205e+01 
R3067t778 n3068 n779 R=2.287e+00 
R3068t712 n3069 n713 R=3.883e+00 
R3068t2603 n3069 n2604 R=4.533e+00 
R3068t2877 n3069 n2878 R=6.079e+00 
R3069t801 n3070 n802 R=6.459e+01 
R3069t2770 n3070 n2771 R=2.305e+00 
R3070t494 n3071 n495 R=2.593e+00 
R3070t1390 n3071 n1391 R=1.115e+01 
R3071t1993 n3072 n1994 R=3.284e+02 
R3071t1369 n3072 n1370 R=4.682e+01 
R3072t1560 n3073 n1561 R=9.629e+01 
R3072t64 n3073 n65 R=5.225e+00 
R3072t245 n3073 n246 R=4.533e+01 
R3073t1062 n3074 n1063 R=2.208e+01 
R3073t1646 n3074 n1647 R=2.247e+01 
R3073t2547 n3074 n2548 R=2.447e+00 
R3073t1234 n3074 n1235 R=5.734e+01 
R3074t1039 n3075 n1040 R=4.457e+01 
R3074t2678 n3075 n2679 R=2.068e+01 
R3074t2163 n3075 n2164 R=4.133e+01 
R3075t2872 n3076 n2873 R=2.586e+01 
R3076t2392 n3077 n2393 R=3.269e+00 
R3076t104 n3077 n105 R=4.499e+00 
R3077t2228 n3078 n2229 R=2.601e+00 
R3078t1301 n3079 n1302 R=1.682e+01 
R3078t1346 n3079 n1347 R=4.865e+00 
R3078t784 n3079 n785 R=1.043e+01 
R3079t1025 n3080 n1026 R=1.599e+01 
R3079t2419 n3080 n2420 R=1.341e+01 
R3080t2762 n3081 n2763 R=3.668e+01 
R3081t2086 n3082 n2087 R=1.364e+01 
R3082t881 n3083 n882 R=1.998e+01 
R3082t2314 n3083 n2315 R=9.201e+00 
R3083t602 n3084 n603 R=1.199e+01 
R3083t1017 n3084 n1018 R=1.367e+01 
R3083t2808 n3084 n2809 R=7.351e+00 
R3084t2381 n3085 n2382 R=6.296e+00 
R3084t607 n3085 n608 R=4.551e+00 
R3084t2073 n3085 n2074 R=1.329e+02 
R3085t2498 n3086 n2499 R=8.229e+00 
R3085t2259 n3086 n2260 R=1.674e+01 
R3087t921 n3088 n922 R=6.886e+00 
R3089t1495 n3090 n1496 R=2.602e+00 
R3090t2360 n3091 n2361 R=3.546e+02 
R3090t2438 n3091 n2439 R=3.412e+00 
R3090t1631 n3091 n1632 R=2.457e+01 
R3090t98 n3091 n99 R=6.560e+00 
R3090t2546 n3091 n2547 R=4.407e+00 
R3092t608 n3093 n609 R=3.902e+00 
R3093t2163 n3094 n2164 R=1.864e+01 
R3093t2678 n3094 n2679 R=4.624e+01 
R3094t907 n3095 n908 R=7.690e+00 
R3094t2828 n3095 n2829 R=4.052e+00 
R3095t1078 n3096 n1079 R=7.423e+00 
R3095t1685 n3096 n1686 R=4.151e+00 
R3095t1575 n3096 n1576 R=2.010e+01 
R3096t885 n3097 n886 R=2.002e+01 
R3097t42 n1 n43 R=4.667e+00 
R3098t2970 n3099 n2971 R=2.787e+00 
R3098t537 n3099 n538 R=3.839e+01 
R3098t3055 n3099 n3056 R=2.285e+01 
R3099t1978 n3100 n1979 R=2.722e+02 
R3100t2353 n3101 n2354 R=4.717e+00 
R3101t1030 n3102 n1031 R=9.757e+00 
R3102t1047 n3103 n1048 R=1.850e+01 
R3102t348 n3103 n349 R=6.968e+00 
R3102t2795 n3103 n2796 R=2.159e+01 
R3103t1074 n3104 n1075 R=4.158e+00 
R3103t747 n3104 n748 R=4.896e+00 
R3105t866 n3106 n867 R=7.928e+00 
R3105t845 n3106 n846 R=3.360e+01 
R3106t3009 n3107 n3010 R=1.047e+01 
R3107t1174 n3108 n1175 R=2.672e+00 
R3107t1559 n3108 n1560 R=2.176e+02 
R3107t2884 n3108 n2885 R=7.456e+00 
R3108t1456 n3109 n1457 R=1.111e+01 
R3108t1709 n3109 n1710 R=1.079e+01 
R3108t1308 n3109 n1309 R=1.196e+01 
R3108t412 n3109 n413 R=1.567e+02 
R3109t2955 n3110 n2956 R=3.271e+00 
R3110t2534 n3111 n2535 R=8.495e+00 
R3111t3091 n1 n3092 R=8.424e+00 
R3112t2652 n3113 n2653 R=1.507e+01 
R3112t2424 n3113 n2425 R=7.081e+01 
R3113t1751 n3114 n1752 R=3.138e+01 
R3113t249 n3114 n250 R=3.439e+00 
R3115t2183 n3116 n2184 R=5.787e+00 
R3117t2808 n3118 n2809 R=6.566e+00 
R3117t3083 n3118 n3084 R=9.730e+00 
R3117t1267 n3118 n1268 R=4.691e+01 
R3117t76 n3118 n77 R=2.760e+01 
R3117t976 n3118 n977 R=5.678e+00 
R3117t1392 n3118 n1393 R=2.141e+01 
R3118t643 n3119 n644 R=6.797e+00 
R3118t2966 n3119 n2967 R=4.793e+00 
R3119t485 n3120 n486 R=3.891e+00 
R3119t2672 n3120 n2673 R=2.201e+01 
R3119t269 n3120 n270 R=1.054e+02 
R3120t879 n3121 n880 R=3.149e+00 
R3120t2909 n3121 n2910 R=1.173e+01 
R3120t543 n3121 n544 R=1.466e+01 
R3120t418 n3121 n419 R=3.437e+00 
R3120t390 n3121 n391 R=7.680e+01 
R3122t3035 n3123 n3036 R=4.434e+00 
R3123t224 n3124 n225 R=2.757e+01 
R3123t2269 n3124 n2270 R=4.806e+00 
R3123t1402 n3124 n1403 R=1.046e+01 
R3124t66 n3125 n67 R=6.073e+00 
R3124t860 n3125 n861 R=3.097e+01 
R3124t386 n3125 n387 R=5.997e+00 
R3124t2724 n3125 n2725 R=5.549e+00 
R3124t2027 n3125 n2028 R=1.529e+01 
R3125t2324 n3126 n2325 R=1.122e+01 
R3125t2429 n3126 n2430 R=2.063e+01 
R3125t296 n3126 n297 R=3.436e+00 
R3126t2431 n3127 n2432 R=2.251e+01 
R3127t2630 n3128 n2631 R=4.326e+00 
R3128t2172 n3129 n2173 R=1.344e+01 
R3128t1051 n3129 n1052 R=5.304e+01 
R3129t2609 n3130 n2610 R=9.320e+00 
R3130t356 n3131 n357 R=2.556e+00 
R3130t1917 n3131 n1918 R=4.083e+01 
R3130t2485 n3131 n2486 R=5.589e+00 
R3131t2405 n3132 n2406 R=3.765e+00 
R3131t194 n3132 n195 R=6.455e+01 
R3132t2963 n3133 n2964 R=1.452e+01 
R3132t2912 n3133 n2913 R=8.977e+00 
R3133t2561 n3134 n2562 R=9.917e+01 
R3133t1259 n3134 n1260 R=9.687e+00 
R3134t283 n3135 n284 R=3.479e+00 
R3134t1695 n3135 n1696 R=5.925e+00 
R3134t2990 n3135 n2991 R=3.766e+01 
R3135t1797 n3136 n1798 R=3.969e+01 
R3136t604 n3137 n605 R=9.483e+00 
R3137t1911 n3138 n1912 R=2.165e+00 
R3137t37 n3138 n38 R=8.911e+01 
R3138t2435 n3139 n2436 R=1.399e+01 
R3138t1040 n3139 n1041 R=4.479e+00 
R3139t3061 n3140 n3062 R=1.560e+02 
R3140t2313 n3141 n2314 R=1.043e+01 
R3140t1888 n3141 n1889 R=7.821e+00 
R3140t455 n3141 n456 R=1.455e+01 
R3141t929 n3142 n930 R=2.361e+01 
R3141t1986 n3142 n1987 R=3.826e+00 
R3142t2204 n3143 n2205 R=6.606e+00 
R3143t2017 n3144 n2018 R=6.178e+00 
R3143t1428 n3144 n1429 R=5.592e+00 
R3145t3128 n3146 n3129 R=3.114e+00 
R3145t2172 n3146 n2173 R=1.677e+01 
R3146t1041 n3147 n1042 R=1.462e+01 
R3146t2868 n3147 n2869 R=3.923e+00 
R3147t1054 n3148 n1055 R=2.567e+00 
R3148t333 n3149 n334 R=7.380e+00 
R3148t1066 n3149 n1067 R=1.152e+01 
R3149t1113 n3150 n1114 R=5.369e+00 
R3150t480 n3151 n481 R=8.423e+00 
R3150t82 n3151 n83 R=1.202e+01 
R3151t2752 n3152 n2753 R=5.721e+00 
R3152t274 n3153 n275 R=6.682e+00 
R3152t371 n3153 n372 R=1.300e+01 
R3152t2740 n3153 n2741 R=8.863e+01 
R3153t230 n3154 n231 R=7.248e+00 
R3153t204 n3154 n205 R=9.000e+00 
R3155t2976 n3156 n2977 R=3.138e+00 
R3155t1378 n3156 n1379 R=1.081e+01 
R3156t231 n3157 n1 R=8.225e+00 
R3156t2356 n3157 n2357 R=9.366e+00 
R3157t3142 n3158 n3143 R=7.587e+00 
R3158t515 n3159 n516 R=6.422e+00 
R3158t2520 n3159 n2521 R=3.800e+01 
R3158t624 n3159 n625 R=2.505e+00 
R3160t1157 n3161 n1158 R=7.152e+00 
R3160t672 n3161 n673 R=1.683e+02 
R3161t1032 n3162 n1033 R=1.016e+01 
R3162t471 n3163 n472 R=5.413e+01 
R3162t2144 n3163 n2145 R=1.077e+01 
R3163t1672 n3164 n1673 R=6.217e+00 
R3163t2271 n3164 n2272 R=4.413e+00 
R3164t3088 n3165 n3089 R=3.947e+00 
R3164t2681 n3165 n2682 R=2.526e+01 
R3164t360 n3165 n361 R=4.286e+00 
R3164t85 n3165 n86 R=3.000e+01 
R3165t1026 n3166 n1027 R=5.975e+00 
R3165t226 n3166 n227 R=4.359e+00 
R3165t1008 n3166 n1009 R=6.952e+01 
R3167t1356 n3168 n1357 R=2.324e+01 
R3167t690 n3168 n691 R=1.482e+01 
R3169t365 n3170 n366 R=8.503e+00 
R3169t2141 n3170 n2142 R=2.338e+01 
R3170t2115 n3171 n2116 R=1.604e+01 
R3170t2583 n3171 n2584 R=2.092e+01 
R3170t1508 n3171 n1509 R=1.137e+01 
R3171t2614 n3172 n2615 R=3.610e+00 
R3171t1 n3172 n2 R=4.660e+00 
R3172t1507 n3173 n1508 R=4.758e+00 
R3174t2023 n3175 n2024 R=7.122e+00 
R3174t2256 n3175 n2257 R=4.878e+00 
R3174t342 n3175 n343 R=7.739e+00 
R3175t1537 n3176 n1538 R=1.074e+01 
R3175t3008 n3176 n3009 R=7.095e+00 
R3175t1602 n3176 n1603 R=1.492e+02 
R3176t2504 n3177 n2505 R=3.237e+01 
R3177t85 n3178 n86 R=2.581e+00 
R3177t3164 n3178 n3165 R=1.954e+01 
R3177t534 n3178 n535 R=6.629e+01 
R3177t185 n3178 n186 R=7.405e+00 
R3177t360 n3178 n361 R=4.885e+00 
R3178t754 n3179 n755 R=6.869e+00 
R3179t2572 n3180 n2573 R=1.011e+01 
R3179t586 n3180 n587 R=1.051e+01 
R3179t2749 n3180 n2750 R=2.422e+01 
R3180t624 n3181 n625 R=4.658e+00 
R3180t2520 n3181 n2521 R=1.223e+01 
R3181t484 n3182 n485 R=2.126e+01 
R3181t1682 n3182 n1683 R=2.464e+00 
R3181t2237 n3182 n2238 R=2.302e+01 
R3181t161 n3182 n162 R=2.628e+00 
R3181t2960 n3182 n2961 R=2.637e+01 
R3182t248 n3183 n249 R=5.704e+00 
R3182t2736 n3183 n2737 R=4.438e+00 
R3183t2317 n3184 n2318 R=5.061e+01 
R3184t447 n3185 n448 R=8.737e+00 
R3184t1121 n3185 n1122 R=5.366e+00 
R3185t2243 n3186 n2244 R=1.024e+02 
R3186t2058 n3187 n2059 R=4.659e+00 
R3186t2166 n3187 n2167 R=2.754e+01 
R3187t941 n3188 n942 R=1.425e+01 
R3187t1550 n3188 n1551 R=3.028e+00 
R3187t1940 n3188 n1941 R=2.012e+00 
R3187t1025 n3188 n1026 R=2.072e+01 
R3189t300 n3190 n301 R=4.247e+00 
R3189t1435 n3190 n1436 R=3.718e+00 
R3190t2898 n3191 n2899 R=1.396e+01 
R3191t2780 n3192 n2781 R=1.728e+01 
R3192t992 n3193 n993 R=9.626e+00 
R3193t1422 n3194 n1423 R=8.767e+00 
R3194t1162 n3195 n1163 R=9.377e+00 
R3197t2049 n3198 n2050 R=7.814e+00 
R3198t87 n3199 n88 R=1.268e+01 
R3199t1514 n3200 n1515 R=1.561e+02 
R3200t3104 n3201 n3105 R=4.564e+00 
R3200t2312 n3201 n2313 R=7.198e+01 
R3200t3013 n3201 n3014 R=4.949e+00 
R3201t663 n3202 n664 R=8.798e+00 
R3201t1135 n3202 n1136 R=7.606e+00 
R3203t3196 n3204 n3197 R=3.244e+00 
R3203t2369 n3204 n2370 R=6.370e+01 
R3204t227 n3205 n228 R=8.593e+00 
R3204t649 n3205 n650 R=6.125e+00 
R3204t2067 n3205 n2068 R=6.086e+00 
R3205t1534 n3206 n1535 R=1.062e+01 
R3205t561 n3206 n562 R=1.278e+02 
R3206t1994 n3207 n1995 R=1.499e+01 
R3206t1175 n3207 n1176 R=9.971e+01 
R3207t1588 n3208 n1589 R=8.167e+00 
R3207t1007 n3208 n1008 R=6.584e+00 
R3208t1098 n3209 n1099 R=8.456e+01 
R3208t3030 n3209 n3031 R=6.263e+01 
R3208t819 n3209 n820 R=1.314e+01 
R3208t1332 n3209 n1333 R=2.218e+01 
R3209t460 n3210 n461 R=4.965e+00 
R3209t2500 n3210 n2501 R=1.095e+01 
R3210t2220 n3211 n2221 R=1.594e+00 
R3211t1800 n3212 n1801 R=1.795e+01 
R3212t336 n3213 n337 R=3.239e+00 
R3213t2807 n3214 n2808 R=6.455e+00 
R3214t1412 n3215 n1413 R=7.909e+00 
R3214t855 n3215 n856 R=2.115e+01 
R3214t1294 n3215 n1295 R=1.829e+01 
R3214t1221 n3215 n1222 R=2.394e+00 
R3215t1789 n3216 n1790 R=3.025e+00 
R3216t1836 n3217 n1837 R=1.525e+01 
R3216t998 n3217 n999 R=6.127e+00 
R3216t456 n3217 n457 R=1.003e+02 
R3216t1970 n3217 n1971 R=1.233e+01 
R3217t2330 n3218 n2331 R=1.575e+02 
R3218t1323 n3219 n1324 R=5.686e+00 
R3218t2340 n3219 n2341 R=1.423e+02 
R3218t1479 n3219 n1480 R=2.804e+00 
R3218t2295 n3219 n2296 R=3.487e+01 
R3219t54 n3220 n55 R=9.057e+00 
R3219t161 n3220 n162 R=5.962e+01 
R3219t3181 n3220 n3182 R=9.865e+00 
R3219t2237 n3220 n2238 R=2.783e+00 
R3220t737 n3221 n738 R=6.316e+00 
R3220t1725 n3221 n1726 R=3.325e+00 
R3220t404 n3221 n405 R=4.475e+00 
R3221t1128 n3222 n1129 R=1.194e+01 
R3221t390 n3222 n391 R=8.459e+00 
R3221t2521 n3222 n2522 R=1.232e+01 
R3222t1435 n3223 n1436 R=6.714e+00 
R3222t3026 n3223 n3027 R=2.754e+01 
R3224t1092 n3225 n1093 R=3.297e+00 
R3224t1331 n3225 n1332 R=9.047e+00 
R3224t1144 n3225 n1145 R=1.279e+01 
R3225t1924 n3226 n1925 R=3.855e+01 
R3226t56 n3227 n57 R=1.100e+01 
R3226t1964 n3227 n1965 R=6.677e+00 
R3229t1951 n3230 n1952 R=8.664e+00 
R3229t218 n3230 n219 R=1.098e+01 
R3229t2084 n3230 n2085 R=2.504e+01 
R3231t3144 n3232 n3145 R=2.819e+00 
R3232t2598 n3233 n2599 R=3.799e+00 
R3232t1787 n3233 n1788 R=4.543e+01 
R3233t1750 n3234 n1751 R=5.563e+00 
R3233t1441 n3234 n1442 R=5.642e+00 
R3233t1427 n3234 n1428 R=9.805e+00 
R3233t2695 n3234 n2696 R=3.617e+01 
R3235t1366 n3236 n1367 R=1.106e+01 
R3235t1181 n3236 n1182 R=6.035e+01 
R3235t1020 n3236 n1021 R=5.410e+00 
R3235t741 n3236 n742 R=1.488e+01 
R3236t106 n3237 n107 R=2.496e+00 
R3236t1727 n3237 n1 R=1.438e+01 
R3237t3212 n3238 n3213 R=2.752e+01 
R3237t336 n3238 n337 R=4.381e+00 
R3237t702 n3238 n703 R=9.017e+00 
R3238t1553 n3239 n1554 R=3.189e+00 
R3238t286 n3239 n287 R=4.874e+00 
R3239t573 n3240 n574 R=1.639e+01 
R3240t1258 n3241 n1259 R=5.970e+00 
R3240t1716 n3241 n1717 R=6.975e+00 
R3240t2879 n3241 n2880 R=1.336e+01 
R3241t3063 n3242 n3064 R=2.047e+02 
R3242t2155 n3243 n2156 R=1.887e+01 
R3243t431 n3244 n432 R=9.530e+00 
R3243t3015 n3244 n3016 R=4.070e+01 
R3244t1093 n3245 n1094 R=2.804e+01 
R3244t1954 n3245 n1955 R=6.167e+00 
R3244t1484 n3245 n1 R=5.480e+01 
R3245t1665 n3246 n1666 R=2.878e+00 
R3245t3037 n3246 n3038 R=8.690e+00 
R3245t1872 n3246 n1873 R=7.849e+01 
R3247t668 n3248 n669 R=3.242e+01 
R3247t1593 n3248 n1594 R=3.956e+01 
R3247t1490 n3248 n1491 R=8.792e+00 
R3248t1363 n3249 n1364 R=3.440e+00 
R3249t2503 n3250 n2504 R=4.173e+00 
R3249t2195 n3250 n2196 R=2.009e+01 
R3249t1061 n3250 n1062 R=2.510e+01 
R3250t1073 n3251 n1074 R=4.565e+01 
R3250t2404 n3251 n2405 R=3.483e+00 
R3251t1972 n3252 n1973 R=8.950e+00 
R3251t2766 n3252 n2767 R=7.586e+00 
R3252t290 n3253 n291 R=1.050e+01 
R3252t1164 n3253 n1165 R=5.517e+00 
R3252t1340 n3253 n1341 R=5.282e+00 
R3254t3251 n3255 n3252 R=3.718e+01 
R3254t901 n3255 n902 R=3.576e+01 
R3254t750 n3255 n751 R=6.737e+00 
R3254t2568 n3255 n2569 R=3.258e+01 
R3254t2539 n3255 n2540 R=1.591e+01 
R3255t1122 n3256 n1123 R=4.628e+00 
R3255t2977 n3256 n2978 R=2.075e+01 
R3255t1204 n3256 n1205 R=5.758e+00 
R3256t392 n3257 n393 R=2.690e+00 
R3256t883 n3257 n884 R=5.866e+00 
R3256t1815 n3257 n1816 R=1.465e+01 
R3257t1152 n3258 n1153 R=1.146e+01 
R3258t2505 n3259 n2506 R=7.087e+00 
R3259t86 n3260 n87 R=3.792e+00 
R3259t2984 n3260 n2985 R=4.489e+01 
R3260t2604 n3261 n2605 R=6.394e+00 
R3260t1627 n3261 n1628 R=1.997e+01 
R3260t1673 n3261 n1674 R=9.272e+00 
R3261t1512 n3262 n1513 R=4.519e+00 
R3262t3040 n3263 n3041 R=4.637e+00 
R3262t2586 n3263 n2587 R=1.928e+00 
R3263t387 n3264 n388 R=1.009e+01 
R3263t2348 n3264 n2349 R=1.058e+01 
R3263t2611 n3264 n2612 R=6.682e+00 
R3263t1878 n3264 n1879 R=4.265e+00 
R3264t2075 n3265 n2076 R=3.119e+00 
R3264t2140 n3265 n2141 R=4.259e+00 
R3264t2211 n3265 n2212 R=4.236e+01 
R3265t3078 n3266 n3079 R=1.265e+01 
R3265t2917 n3266 n2918 R=7.948e+00 
R3266t2952 n3267 n2953 R=6.574e+00 
R3266t1867 n3267 n1868 R=2.145e+01 
R3267t1416 n3268 n1417 R=1.026e+03 
R3267t1797 n3268 n1798 R=5.506e+00 
R3267t3135 n3268 n3136 R=3.350e+00 
R3269t2051 n3270 n2052 R=2.373e+02 
R3270t1624 n3271 n1625 R=1.630e+01 
R3270t1863 n3271 n1864 R=2.256e+00 
R3270t347 n3271 n348 R=9.510e+01 
R3271t614 n3272 n615 R=1.221e+01 
R3271t1279 n3272 n1280 R=5.459e+00 
R3271t791 n3272 n792 R=3.106e+01 
R3271t2408 n3272 n2409 R=2.963e+00 
R3272t1009 n3273 n1010 R=1.824e+01 
R3272t3050 n3273 n3051 R=6.414e+00 
R3274t1332 n3275 n1333 R=1.938e+01 
R3275t2160 n3276 n2161 R=1.264e+01 
R3275t2088 n3276 n2089 R=3.151e+00 
R3275t105 n3276 n106 R=1.294e+01 
R3276t2019 n3277 n2020 R=9.939e+00 
R3276t1664 n3277 n1665 R=7.632e+00 
R3277t2892 n3278 n2893 R=1.574e+01 
R3279t928 n3280 n929 R=4.908e+01 
R3280t3121 n3281 n3122 R=3.363e+00 
R3281t3231 n3282 n3232 R=7.252e+00 
R3281t3144 n3282 n3145 R=3.797e+01 
R3281t546 n3282 n547 R=2.980e+01 
R3282t1778 n3283 n1779 R=3.686e+00 
R3282t2493 n3283 n2494 R=1.865e+01 
R3282t2968 n3283 n2969 R=1.587e+01 
R3282t937 n3283 n938 R=2.969e+01 
R3283t2846 n3284 n2847 R=2.402e+01 
R3284t1974 n3285 n1975 R=1.236e+01 
R3284t3021 n3285 n3022 R=1.482e+01 
R3284t2172 n3285 n2173 R=1.415e+01 
R3285t1862 n3286 n1863 R=2.965e+00 
R3285t689 n3286 n690 R=3.934e+00 
R3286t605 n3287 n606 R=1.879e+01 
R3286t2596 n3287 n2597 R=6.475e+00 
R3286t2102 n3287 n2103 R=2.732e+01 
R3286t2453 n3287 n2454 R=1.835e+01 
R3287t2651 n3288 n2652 R=4.830e+00 
R3287t1665 n3288 n1666 R=5.604e+00 
R3287t3245 n3288 n3246 R=6.145e+01 
R3288t1611 n3289 n1612 R=1.128e+01 
R3288t2327 n3289 n2328 R=2.517e+00 
R3288t2495 n3289 n2496 R=9.246e+00 
R3290t966 n3291 n967 R=9.760e+00 
R3291t61 n3292 n62 R=4.443e+00 
R3293t1236 n3294 n1237 R=1.146e+01 
R3293t3288 n3294 n3289 R=3.389e+01 
R3293t2495 n3294 n2496 R=5.886e+00 
R3294t2044 n3295 n2045 R=3.348e+00 
R3294t309 n3295 n310 R=9.176e+00 
R3294t1771 n3295 n1772 R=4.417e+00 
R3295t2716 n3296 n2717 R=7.605e+00 
R3295t1860 n3296 n1861 R=1.392e+02 
R3295t1585 n3296 n1586 R=3.390e+00 
R3296t1734 n3297 n1735 R=6.158e+00 
R3297t2844 n3298 n2845 R=5.815e+00 
R3299t931 n3300 n932 R=2.672e+01 
R3299t2758 n3300 n2759 R=7.629e+00 
R3299t2819 n3300 n2820 R=1.657e+01 
R3300t357 n3301 n358 R=1.331e+01 
R3300t1431 n3301 n1432 R=4.788e+00 
R3300t1353 n3301 n1354 R=8.790e+01 
R3301t660 n3302 n661 R=5.629e+00 
R3301t1567 n3302 n1568 R=6.925e+00 
R3301t1056 n3302 n1057 R=4.291e+00 
R3303t3260 n3304 n3261 R=8.745e+00 
R3303t1082 n3304 n1083 R=7.510e+00 
R3304t545 n3305 n546 R=8.386e+00 
R3304t138 n3305 n139 R=3.645e+01 
R3304t2694 n3305 n2695 R=2.769e+00 
R3305t530 n3306 n531 R=5.717e+00 
R3306t2100 n3307 n2101 R=5.843e+00 
R3306t154 n3307 n155 R=3.464e+00 
R3307t863 n3308 n864 R=1.433e+01 
R3307t1130 n3308 n1131 R=1.260e+01 
R3309t2336 n3310 n2337 R=3.163e+00 
R3310t2512 n3311 n2513 R=8.455e+00 
R3310t94 n3311 n95 R=4.543e+00 
R3310t2578 n3311 n2579 R=1.188e+02 
R3310t1243 n3311 n1244 R=6.360e+00 
R3311t1788 n3312 n1789 R=1.042e+01 
R3312t585 n3313 n586 R=2.030e+01 
R3313t2309 n3314 n2310 R=1.725e+01 
R3313t1554 n3314 n1555 R=1.451e+01 
R3314t1438 n3315 n1439 R=8.021e+00 
R3314t1142 n3315 n1143 R=4.505e+00 
R3315t3003 n3316 n3004 R=1.007e+01 
R3316t3205 n3317 n3206 R=2.907e+00 
R3317t675 n3318 n676 R=4.778e+00 
R3317t112 n3318 n113 R=2.178e+02 
R3317t41 n3318 n42 R=4.338e+01 
R3317t714 n3318 n715 R=7.235e+01 
R3318t2504 n3319 n2505 R=5.242e+00 
R3318t519 n3319 n520 R=5.261e+00 
R3319t1362 n3320 n1363 R=6.025e+00 
R3319t2794 n3320 n2795 R=3.410e+00 
R3320t1755 n3321 n1756 R=2.425e+00 
R3321t859 n3322 n860 R=9.539e+00 
R3321t1722 n3322 n1723 R=1.494e+01 
R3321t1503 n3322 n1504 R=6.273e+00 
R3322t1077 n3323 n1078 R=1.100e+01 
R3322t547 n3323 n548 R=1.637e+01 
R3322t1467 n3323 n1468 R=8.280e+00 
R3322t1002 n3323 n1003 R=4.680e+00 
R3323t1565 n3324 n1566 R=5.817e+00 
R3324t112 n3325 n113 R=7.348e+00 
R3325t1552 n3326 n1553 R=2.834e+01 
R3325t398 n3326 n1 R=4.187e+00 
R3325t987 n3326 n988 R=4.430e+01 
R3326t2565 n3327 n2566 R=2.643e+00 
R3326t1425 n3327 n1426 R=8.234e+00 
R3327t1939 n3328 n1940 R=6.126e+01 
R3327t1547 n3328 n1548 R=5.152e+00 
R3328t887 n3329 n888 R=3.998e+00 
R3329t1835 n3330 n1836 R=2.208e+00 
R3330t3143 n3331 n3144 R=1.995e+00 
R3330t268 n3331 n269 R=1.933e+00 
R3331t1171 n3332 n1172 R=1.992e+01 
R3332t1258 n3333 n1259 R=1.024e+01 
R3332t2879 n3333 n2880 R=4.554e+00 
R3332t1622 n3333 n1623 R=1.015e+01 
R3332t124 n3333 n125 R=1.471e+01 
R3333t729 n3334 n730 R=3.331e+00 
R3333t2746 n3334 n2747 R=1.005e+01 
R3333t252 n3334 n253 R=4.121e+00 
R3334t1565 n3335 n1566 R=1.397e+04 
R3334t3323 n3335 n3324 R=1.942e+00 
R3335t2376 n3336 n2377 R=8.958e+00 
R3336t1360 n3337 n1361 R=1.252e+01 
R3336t1480 n3337 n1481 R=1.566e+00 
R3336t2929 n3337 n2930 R=8.876e+00 
R3337t1177 n3338 n1178 R=9.910e+00 
R3337t67 n3338 n68 R=5.120e+00 
R3338t2428 n3339 n2429 R=3.147e+00 
R3338t1880 n3339 n1881 R=2.642e+01 
R3339t1696 n3340 n1697 R=6.640e+00 
R3339t2212 n3340 n2213 R=4.225e+00 
R3340t2814 n3341 n2815 R=1.956e+00 
R3340t2316 n3341 n2317 R=6.878e+01 
R3341t426 n3342 n427 R=2.227e+01 
R3341t1047 n3342 n1048 R=1.144e+01 
R3342t323 n3343 n324 R=2.245e+00 
R3343t350 n3344 n351 R=2.432e+01 
R3343t2045 n3344 n2046 R=2.464e+01 
R3344t1146 n3345 n1147 R=3.890e+00 
R3344t1875 n3345 n1876 R=4.810e+00 
R3344t2261 n3345 n2262 R=1.088e+01 
R3345t1825 n3346 n1826 R=4.974e+00 
R3345t461 n3346 n462 R=6.122e+00 
R3346t1297 n3347 n1298 R=2.265e+01 
R3346t2462 n3347 n2463 R=8.232e+00 
R3346t679 n3347 n680 R=3.375e+00 
R3347t2441 n3348 n2442 R=1.534e+00 
R3347t2478 n3348 n2479 R=1.100e+01 
R3347t334 n3348 n335 R=7.440e+02 
R3347t1166 n3348 n1167 R=9.330e+01 
R3348t2321 n3349 n2322 R=6.455e+00 
R3348t2444 n3349 n2445 R=1.096e+01 
R3349t2245 n3350 n2246 R=9.165e+00 
R3349t645 n3350 n646 R=1.503e+02 
R3349t2667 n3350 n2668 R=1.784e+01 
R3350t1191 n3351 n1192 R=5.800e+00 
R3351t1264 n3352 n1265 R=2.382e+01 
R3353t1881 n3354 n1882 R=4.038e+01 
R3353t1615 n3354 n1616 R=4.800e+01 
R3353t1799 n3354 n1800 R=7.741e+00 
R3353t1368 n3354 n1369 R=1.023e+02 
R3354t513 n3355 n514 R=1.171e+01 
R3354t2137 n3355 n2138 R=4.349e+00 
R3355t1347 n3356 n1348 R=1.387e+01 
R3355t2207 n3356 n2208 R=1.020e+01 
R3356t106 n3357 n107 R=2.436e+00 
R3356t2738 n3357 n2739 R=5.613e+00 
R3356t1727 n3357 n1 R=1.376e+01 
R3357t1832 n3358 n1833 R=1.009e+01 
R3357t313 n3358 n314 R=4.170e+00 
R3358t3137 n3359 n3138 R=8.930e+00 
R3358t37 n3359 n38 R=4.949e+00 
R3358t1402 n3359 n1403 R=5.999e+00 
R3359t2206 n3360 n2207 R=6.334e+00 
R3359t1014 n3360 n1015 R=1.197e+01 
R3360t1055 n3361 n1056 R=7.478e+00 
R3361t2548 n3362 n2549 R=9.043e+00 
R3361t53 n3362 n54 R=1.092e+02 
R3361t1544 n3362 n1545 R=2.325e+00 
R3361t2712 n3362 n2713 R=6.440e+01 
R3362t2249 n3363 n2250 R=3.634e+01 
R3362t2466 n3363 n2467 R=2.947e+00 
R3363t1936 n3364 n1937 R=4.948e+00 
R3364t3087 n3365 n3088 R=1.264e+01 
R3364t982 n3365 n983 R=2.935e+01 
R3364t921 n3365 n922 R=3.018e+00 
R3365t2172 n3366 n2173 R=3.799e+01 
R3365t3284 n3366 n3285 R=6.022e+00 
R3366t1275 n3367 n1276 R=2.057e+01 
R3366t1827 n3367 n1828 R=8.798e+00 
R3367t1824 n3368 n1825 R=1.236e+01 
R3367t2315 n3368 n2316 R=4.076e+01 
R3367t2094 n3368 n2095 R=5.468e+00 
R3368t634 n3369 n635 R=1.406e+02 
R3368t2700 n3369 n2701 R=3.722e+00 
R3369t825 n3370 n826 R=1.285e+01 
R3369t853 n3370 n854 R=4.327e+00 
R3370t422 n3371 n423 R=2.595e+01 
R3370t1884 n3371 n1885 R=3.108e+00 
R3370t2503 n3371 n2504 R=1.088e+01 
R3371t1470 n3372 n1471 R=9.674e+00 
R3371t3278 n3372 n3279 R=3.056e+00 
R3371t16 n3372 n17 R=1.753e+02 
R3372t618 n3373 n619 R=4.743e+00 
R3372t2014 n3373 n2015 R=2.274e+00 
R3373t2210 n3374 n2211 R=4.428e+01 
R3373t3036 n3374 n3037 R=6.078e+00 
R3373t2680 n3374 n2681 R=5.174e+00 
R3374t3276 n3375 n3277 R=5.949e+01 
R3374t2779 n3375 n2780 R=7.965e+01 
R3375t86 n3376 n87 R=1.016e+01 
R3375t3259 n3376 n3260 R=1.718e+01 
R3376t2945 n3377 n2946 R=1.171e+01 
R3376t1256 n3377 n1257 R=2.204e+00 
R3377t1913 n3378 n1914 R=5.637e+00 
R3377t2149 n3378 n2150 R=8.714e+00 
R3378t1730 n3379 n1731 R=5.644e+00 
R3378t794 n3379 n795 R=6.642e+00 
R3379t190 n3380 n191 R=4.410e+00 
R3382t187 n3383 n188 R=2.989e+02 
R3382t2590 n3383 n2591 R=4.820e+00 
R3383t2852 n3384 n2853 R=4.877e+00 
R3383t420 n3384 n421 R=4.828e+00 
R3383t1850 n3384 n1851 R=6.101e+01 
R3384t1175 n3385 n1176 R=3.677e+00 
R3384t2259 n3385 n2260 R=1.217e+01 
R3384t3206 n3385 n3207 R=5.677e+00 
R3385t1923 n3386 n1924 R=8.833e+00 
R3386t204 n3387 n205 R=7.991e+00 
R3386t3153 n3387 n3154 R=7.606e+00 
R3386t478 n3387 n479 R=3.001e+00 
R3388t1956 n3389 n1957 R=1.605e+02 
R3388t221 n3389 n222 R=2.559e+00 
R3389t1639 n1 n1640 R=4.659e+00 
R3390t3251 n3391 n3252 R=1.962e+01 
R3391t1406 n3392 n1407 R=2.417e+01 
R3391t1473 n3392 n1474 R=1.814e+02 
R3392t1686 n3393 n1687 R=6.476e+00 
R3392t1566 n3393 n1567 R=9.989e+00 
R3394t1379 n3395 n1380 R=2.980e+00 
R3394t2576 n3395 n2577 R=3.441e+00 
R3396t1692 n3397 n1693 R=2.100e+01 
R3396t2765 n3397 n2766 R=7.409e+00 
R3396t1775 n3397 n1776 R=1.843e+01 
R3397t2617 n3398 n2618 R=1.156e+01 
R3397t977 n3398 n978 R=9.993e+00 
R3398t886 n3399 n887 R=7.139e+00 
R3399t2542 n3400 n2543 R=1.604e+01 
R3399t2572 n3400 n2573 R=7.716e+00 
R3399t3179 n3400 n3180 R=6.731e+00 
R3399t195 n3400 n196 R=1.566e+01 
R3400t669 n3401 n670 R=2.559e+01 
R3400t2359 n3401 n2360 R=1.802e+01 
R3400t294 n3401 n295 R=1.927e+01 
R3400t1905 n3401 n1906 R=1.188e+01 
R3401t2331 n3402 n2332 R=8.157e+01 
R3401t964 n3402 n965 R=8.140e+01 
R3402t406 n3403 n407 R=8.212e+00 
R3402t91 n3403 n92 R=3.410e+01 
R3402t1883 n3403 n1884 R=4.131e+00 
R3403t1921 n3404 n1922 R=1.158e+01 
R3404t234 n3405 n235 R=8.112e+00 
R3404t1603 n3405 n1604 R=6.904e+00 
R3404t2133 n3405 n2134 R=5.463e+00 
R3405t1782 n3406 n1783 R=4.788e+00 
R3405t3054 n3406 n3055 R=9.710e+00 
R3406t1440 n3407 n1441 R=8.431e+01 
R3406t2583 n3407 n2584 R=1.677e+01 
R3407t599 n3408 n600 R=9.817e+00 
R3407t1254 n3408 n1255 R=4.593e+00 
R3408t1844 n3409 n1845 R=3.001e+00 
R3408t222 n3409 n223 R=4.738e+00 
R3409t1463 n3410 n1464 R=8.495e+00 
R3410t3064 n3411 n3065 R=2.265e+01 
R3410t2867 n3411 n2868 R=5.957e+00 
R3411t1890 n3412 n1891 R=1.568e+01 
R3411t2923 n3412 n2924 R=6.273e+00 
R3411t808 n3412 n809 R=3.598e+00 
R3412t1378 n3413 n1379 R=2.683e+01 
R3413t2049 n3414 n2050 R=9.522e+01 
R3413t1190 n3414 n1191 R=7.672e+01 
R3413t1197 n3414 n1198 R=6.378e+01 
R3413t3197 n3414 n3198 R=1.600e+01 
R3414t939 n3415 n940 R=9.221e+00 
R3414t1230 n3415 n1231 R=1.745e+01 
R3415t1407 n3416 n1408 R=1.817e+01 
R3415t1081 n3416 n1082 R=1.249e+03 
R3416t89 n3417 n90 R=2.690e+02 
R3416t1648 n3417 n1649 R=8.806e+00 
R3416t1096 n3417 n1097 R=5.812e+00 
R3417t3190 n3418 n3191 R=9.007e+00 
R3417t2403 n3418 n2404 R=3.203e+00 
R3418t628 n3419 n629 R=1.360e+00 
R3418t2412 n3419 n2413 R=1.818e+00 
R3418t2461 n3419 n2462 R=1.887e+01 
R3419t469 n3420 n470 R=1.186e+01 
R3419t1594 n3420 n1595 R=9.025e+00 
R3420t1190 n3421 n1191 R=3.699e+00 
R3420t1197 n3421 n1198 R=8.343e+00 
R3421t2600 n3422 n2601 R=7.009e+00 
R3421t1541 n3422 n1542 R=6.732e+00 
R3422t1280 n3423 n1281 R=1.554e+01 
R3422t2593 n3423 n2594 R=9.293e+00 
R3422t2837 n3423 n2838 R=3.115e+00 
R3423t592 n3424 n593 R=7.567e+00 
R3423t2930 n3424 n2931 R=1.137e+01 
R3423t908 n3424 n909 R=9.943e+00 
R3423t838 n3424 n839 R=1.079e+01 
R3424t658 n3425 n659 R=2.115e+01 
R3425t1959 n3426 n1960 R=4.929e+01 
R3425t1001 n3426 n1002 R=1.891e+00 
R3426t3305 n3427 n3306 R=6.400e+01 
R3426t2294 n3427 n2295 R=7.222e+00 
R3427t1857 n3428 n1858 R=5.858e+01 
R3427t945 n3428 n946 R=1.387e+01 
R3428t695 n3429 n696 R=2.724e+00 
R3428t912 n3429 n913 R=3.922e+01 
R3429t891 n3430 n892 R=1.892e+02 
R3429t2882 n3430 n2883 R=1.107e+01 
R3430t284 n3431 n285 R=5.597e+00 
R3430t864 n3431 n865 R=7.110e+00 
R3431t2587 n3432 n2588 R=1.010e+01 
R3432t3260 n3433 n3261 R=1.070e+01 
R3432t3303 n3433 n3304 R=5.008e+00 
R3433t1601 n3434 n1602 R=4.059e+00 
R3434t318 n3435 n319 R=1.406e+01 
R3434t2300 n3435 n2301 R=4.331e+00 
R3434t2623 n3435 n2624 R=1.211e+01 
R3435t2387 n3436 n2388 R=1.724e+01 
R3435t2356 n3436 n2357 R=9.329e+00 
R3435t3156 n3436 n3157 R=4.418e+00 
R3436t2284 n3437 n2285 R=2.825e+01 
R3436t340 n3437 n341 R=1.946e+01 
R3436t1453 n3437 n1454 R=9.243e+00 
R3436t935 n3437 n936 R=8.564e+01 
R3436t2858 n3437 n2859 R=8.190e+00 
R3437t888 n3438 n889 R=1.944e+01 
R3438t2731 n3439 n2732 R=1.390e+01 
R3438t2342 n3439 n2343 R=6.789e+00 
R3438t1342 n3439 n1343 R=4.878e+00 
R3439t2340 n3440 n2341 R=3.560e+01 
R3439t2374 n3440 n2375 R=2.363e+00 
R3439t341 n3440 n342 R=1.479e+01 
R3440t1036 n3441 n1037 R=6.034e+00 
R3440t789 n3441 n790 R=5.442e+02 
R3440t1024 n3441 n1025 R=9.611e+00 
R3441t2630 n3442 n2631 R=9.574e+00 
R3441t3127 n3442 n3128 R=1.125e+01 
R3443t995 n3444 n996 R=1.788e+01 
R3443t29 n3444 n30 R=2.572e+00 
R3443t3166 n3444 n3167 R=6.746e+00 
R3444t1336 n3445 n1337 R=2.303e+01 
R3444t1589 n3445 n1590 R=7.606e+01 
R3444t2303 n3445 n2304 R=2.680e+00 
R3444t2021 n3445 n2022 R=1.887e+01 
R3445t3178 n3446 n3179 R=3.875e+00 
R3445t2805 n3446 n2806 R=4.116e+00 
R3447t1595 n3448 n1596 R=6.928e+00 
R3447t1091 n3448 n1092 R=1.442e+01 
R3448t2648 n3449 n2649 R=1.005e+01 
R3448t1851 n3449 n1852 R=2.610e+01 
R3451t2249 n3452 n2250 R=2.910e+00 
R3451t3362 n3452 n3363 R=4.929e+00 
R3452t932 n3453 n933 R=1.991e+02 
R3454t2287 n3455 n2288 R=5.568e+00 
R3455t3366 n3456 n3367 R=1.582e+02 
R3455t1708 n3456 n1 R=2.289e+01 
R3455t1827 n3456 n1828 R=6.702e+00 
R3456t1872 n3457 n1873 R=4.336e+00 
R3457t536 n3458 n537 R=6.750e+00 
R3457t2951 n3458 n2952 R=6.149e+00 
R3458t564 n3459 n565 R=5.324e+00 
R3458t2717 n3459 n2718 R=4.161e+00 
R3459t1540 n3460 n1541 R=9.195e+00 
R3460t3116 n3461 n3117 R=9.836e+00 
R3461t2788 n3462 n2789 R=4.747e+00 
R3461t432 n3462 n433 R=6.409e+00 
R3461t2440 n3462 n2441 R=1.778e+01 
R3462t93 n3463 n94 R=5.684e+00 
R3463t175 n3464 n176 R=2.850e+00 
R3464t2012 n3465 n2013 R=4.925e+00 
R3465t509 n3466 n510 R=9.266e+01 
R3465t2713 n3466 n2714 R=8.838e+00 
R3465t1683 n3466 n1684 R=1.260e+01 
R3466t3346 n3467 n3347 R=2.561e+01 
R3466t127 n3467 n128 R=7.764e+00 
R3466t679 n3467 n680 R=6.342e+00 
R3467t2466 n3468 n2467 R=5.186e+02 
R3468t1911 n3469 n1912 R=1.032e+01 
R3469t222 n3470 n223 R=1.174e+01 
R3470t1618 n3471 n1619 R=1.574e+00 
R3470t2494 n3471 n2495 R=2.203e+01 
R3470t1105 n3471 n1106 R=6.460e+00 
R3471t2312 n3472 n2313 R=6.807e+01 
R3471t34 n3472 n35 R=8.636e+00 
R3472t3454 n3473 n3455 R=1.800e+02 
R3473t348 n3474 n349 R=7.467e+00 
R3474t214 n3475 n215 R=1.801e+02 
R3474t329 n3475 n330 R=3.501e+00 
R3475t924 n3476 n925 R=6.189e+00 
R3475t2496 n3476 n2497 R=2.589e+01 
R3476t2734 n3477 n2735 R=1.062e+01 
R3477t2728 n3478 n2729 R=8.927e+00 
R3477t312 n3478 n313 R=3.034e+00 
R3478t477 n3479 n478 R=3.599e+00 
R3478t2018 n3479 n2019 R=6.661e+00 
R3479t2628 n3480 n2629 R=6.166e+00 
R3479t1096 n3480 n1097 R=6.188e+00 
R3480t1765 n3481 n1766 R=7.162e+00 
R3480t2167 n3481 n2168 R=2.936e+00 
R3480t1806 n3481 n1807 R=2.605e+01 
R3480t2874 n3481 n2875 R=2.233e+00 
R3481t553 n3482 n554 R=5.660e+00 
R3481t3277 n3482 n3278 R=2.567e+00 
R3482t2836 n3483 n2837 R=3.208e+00 
R3482t1661 n3483 n1662 R=4.389e+00 
R3482t1597 n3483 n1598 R=4.289e+00 
R3483t2741 n3484 n2742 R=1.920e+01 
R3483t1898 n3484 n1899 R=7.357e+00 
R3483t2314 n3484 n2315 R=3.190e+00 
R3484t1400 n3485 n1401 R=1.142e+02 
R3484t661 n3485 n662 R=1.181e+01 
R3484t1976 n3485 n1977 R=2.933e+00 
R3487t63 n3488 n64 R=5.091e+00 
R3487t758 n3488 n759 R=1.868e+01 
R3488t980 n3489 n981 R=4.114e+00 
R3488t1074 n3489 n1075 R=1.904e+01 
R3488t616 n3489 n617 R=3.330e+02 
R3488t2413 n3489 n2414 R=6.704e+00 
R3489t2725 n3490 n2726 R=6.643e+00 
R3489t389 n3490 n390 R=8.584e+00 
R3489t347 n3490 n348 R=3.989e+00 
R3490t7 n3491 n8 R=1.442e+01 
R3490t501 n3491 n502 R=4.564e+00 
R3490t3050 n3491 n3051 R=1.637e+01 
R3491t603 n3492 n604 R=2.276e+00 
R3492t2838 n1 n2839 R=3.893e+00 
R3493t2267 n3494 n2268 R=2.140e+02 
R3493t1516 n3494 n1517 R=3.897e+01 
R3494t1715 n3495 n1716 R=5.862e+00 
R3495t1331 n3496 n1332 R=1.116e+01 
R3495t2077 n3496 n2078 R=9.077e+01 
R3496t1294 n3497 n1295 R=1.359e+01 
R3496t1221 n3497 n1222 R=2.851e+00 
R3497t981 n3498 n982 R=8.848e+01 
R3497t2378 n3498 n2379 R=1.621e+01 
R3497t2749 n3498 n2750 R=4.604e+01 
R3498t138 n3499 n139 R=1.103e+01 
R3498t545 n3499 n546 R=5.579e+01 
R3498t3304 n3499 n3305 R=3.576e+00 
R3499t1693 n3500 n1694 R=4.795e+00 
R3500t222 n3501 n223 R=2.729e+01 
R3500t2273 n3501 n2274 R=1.683e+01 
R3500t2867 n3501 n2868 R=8.163e+01 
R3501t846 n3502 n847 R=2.447e+00 
R3501t2732 n3502 n2733 R=2.220e+01 
R3501t533 n3502 n534 R=4.473e+01 
R3502t3050 n3503 n3051 R=3.458e+00 
R3502t1510 n3503 n1511 R=5.402e+01 
R3503t1584 n3504 n1585 R=3.506e+00 
R3503t1586 n3504 n1587 R=3.288e+01 
R3504t2714 n3505 n2715 R=3.271e+00 
R3504t1901 n3505 n1902 R=7.201e+00 
R3506t1283 n3507 n1284 R=7.157e+00 
R3506t523 n3507 n524 R=8.185e+00 
R3506t2320 n3507 n2321 R=3.402e+00 
R3506t916 n3507 n917 R=1.529e+02 
R3507t1533 n3508 n1534 R=4.947e+00 
R3507t1023 n3508 n1024 R=5.063e+00 
R3508t1326 n3509 n1327 R=3.685e+01 
R3508t1830 n3509 n1831 R=3.643e+00 
R3509t3494 n3510 n3495 R=3.624e+00 
R3509t1715 n3510 n1716 R=1.170e+01 
R3510t591 n3511 n592 R=4.369e+00 
R3510t1156 n3511 n1157 R=9.363e+00 
R3510t3351 n3511 n3352 R=7.162e+00 
R3512t3359 n3513 n3360 R=1.961e+01 
R3513t3448 n3514 n3449 R=3.094e+00 
R3513t1851 n3514 n1852 R=1.051e+01 
R3514t944 n3515 n945 R=1.867e+00 
R3515t320 n3516 n321 R=5.603e+00 
R3515t144 n3516 n145 R=7.348e+00 
R3516t3282 n3517 n3283 R=7.168e+01 
R3516t2493 n3517 n2494 R=3.575e+00 
R3517t621 n3518 n622 R=2.067e+01 
R3517t1984 n3518 n1985 R=3.532e+00 
R3517t2006 n3518 n2007 R=1.412e+01 
R3518t3515 n3519 n3516 R=7.372e+00 
R3519t1415 n3520 n1416 R=1.228e+01 
R3519t204 n3520 n205 R=7.169e+00 
R3520t1595 n3521 n1596 R=7.762e+00 
R3520t3447 n3521 n3448 R=7.070e+00 
R3520t1091 n3521 n1092 R=4.229e+00 
R3520t698 n3521 n699 R=6.528e+00 
R3521t216 n3522 n217 R=4.765e+00 
R3521t2602 n3522 n2603 R=1.443e+01 
R3522t1493 n3523 n1494 R=1.006e+01 
R3523t250 n3524 n251 R=1.322e+01 
R3523t448 n3524 n449 R=6.491e+00 
R3523t1523 n3524 n1524 R=6.567e+00 
R3524t3383 n3525 n3384 R=2.616e+00 
R3524t1850 n3525 n1851 R=2.724e+01 
R3524t246 n3525 n247 R=2.561e+00 
R3525t3163 n3526 n3164 R=1.117e+01 
R3525t2271 n3526 n2272 R=3.225e+00 
R3526t3246 n3527 n3247 R=8.582e+00 
R3527t2664 n3528 n2665 R=6.897e+01 
R3527t96 n3528 n97 R=3.879e+01 
R3527t2796 n3528 n2797 R=4.235e+00 
R3527t155 n3528 n156 R=3.162e+00 
R3528t680 n3529 n681 R=1.418e+01 
R3528t528 n3529 n529 R=7.466e+00 
R3528t70 n3529 n71 R=5.568e+00 
R3528t2054 n3529 n2055 R=1.245e+02 
R3528t105 n3529 n106 R=2.159e+00 
R3528t3275 n3529 n3276 R=4.628e+01 
R3529t1266 n3530 n1267 R=2.968e+01 
R3529t3215 n3530 n3216 R=5.289e+00 
R3529t597 n3530 n598 R=2.398e+01 
R3530t1804 n3531 n1805 R=8.442e+00 
R3531t2220 n3532 n2221 R=4.746e+01 
R3531t570 n3532 n571 R=4.944e+00 
R3532t1966 n3533 n1967 R=6.227e+00 
R3533t2288 n3534 n2289 R=1.395e+01 
R3533t237 n3534 n238 R=4.003e+00 
R3534t818 n3535 n819 R=2.510e+01 
R3534t1339 n3535 n1340 R=2.167e+00 
R3535t370 n3536 n371 R=1.030e+01 
R3535t883 n3536 n884 R=5.407e+00 
R3535t2354 n3536 n2355 R=9.746e+00 
R3536t2154 n3537 n2155 R=1.116e+01 
R3536t560 n3537 n561 R=6.537e+01 
R3537t442 n3538 n443 R=6.853e+00 
R3537t495 n3538 n496 R=1.048e+01 
R3538t2346 n3539 n2347 R=4.852e+00 
R3538t651 n3539 n652 R=1.403e+01 
R3538t1926 n3539 n1927 R=2.147e+02 
R3538t636 n3539 n637 R=1.350e+01 
R3538t436 n3539 n437 R=6.473e+00 
R3539t677 n3540 n678 R=7.068e+00 
R3540t1224 n3541 n1225 R=3.698e+01 
R3540t2108 n3541 n2109 R=3.822e+00 
R3540t433 n3541 n434 R=3.000e+00 
R3540t507 n3541 n508 R=5.462e+00 
R3541t1398 n3542 n1399 R=1.402e+00 
R3541t2893 n3542 n2894 R=3.394e+01 
R3542t2123 n3543 n2124 R=3.510e+00 
R3542t987 n3543 n988 R=1.403e+01 
R3543t86 n3544 n87 R=3.434e+00 
R3544t1263 n3545 n1264 R=8.198e+00 
R3545t17 n3546 n18 R=4.516e+00 
R3545t649 n3546 n650 R=9.899e+00 
R3545t884 n3546 n885 R=1.124e+01 
R3545t1171 n3546 n1172 R=2.781e+01 
R3546t416 n3547 n417 R=3.479e+00 
R3547t1613 n3548 n1614 R=4.818e+00 
R3547t604 n3548 n605 R=1.043e+01 
R3549t3122 n3550 n3123 R=4.178e+00 
R3549t3035 n3550 n3036 R=5.787e+00 
R3549t2732 n3550 n2733 R=6.159e+01 
R3549t1553 n3550 n1554 R=2.555e+00 
R3550t912 n3551 n913 R=8.484e+01 
R3551t1234 n3552 n1235 R=4.776e+00 
R3551t3073 n3552 n3074 R=1.538e+01 
R3552t3 n3553 n4 R=1.173e+02 
R3552t3244 n3553 n3245 R=1.274e+00 
R3552t1484 n3553 n1 R=1.760e+01 
R3552t1383 n3553 n1384 R=1.971e+00 
R3553t279 n3554 n280 R=6.889e+00 
R3553t2354 n3554 n2355 R=4.296e+00 
R3554t1466 n3555 n1467 R=9.594e+00 
R3554t3015 n3555 n3016 R=8.518e+00 
R3555t358 n3556 n359 R=3.285e+00 
R3555t2911 n3556 n2912 R=1.004e+01 
R3556t299 n3557 n300 R=6.982e+01 
R3556t2908 n3557 n2909 R=2.663e+01 
R3556t1956 n3557 n1957 R=2.825e+01 
R3556t221 n3557 n222 R=8.705e+00 
R3556t942 n3557 n943 R=5.634e+00 
R3558t170 n3559 n171 R=3.298e+00 
R3558t1153 n3559 n1154 R=7.820e+00 
R3558t1758 n3559 n1759 R=3.799e+01 
R3558t1414 n3559 n1415 R=2.000e+01 
R3559t3541 n3560 n3542 R=1.747e+00 
R3559t2893 n3560 n2894 R=4.959e+01 
R3560t219 n3561 n220 R=8.551e+00 
R3560t3526 n3561 n3527 R=1.081e+01 
R3560t3000 n3561 n3001 R=4.241e+00 
R3561t1538 n3562 n1539 R=8.413e+00 
R3561t2421 n3562 n2422 R=2.858e+01 
R3562t118 n3563 n119 R=1.082e+01 
R3563t757 n3564 n758 R=2.501e+01 
R3563t900 n3564 n901 R=1.087e+01 
R3563t939 n3564 n940 R=4.289e+01 
R3564t3087 n3565 n3088 R=4.214e+00 
R3565t1628 n3566 n1629 R=3.541e+00 
R3566t1206 n3567 n1207 R=2.192e+01 
R3566t2469 n3567 n2470 R=2.551e+00 
R3566t1662 n3567 n1663 R=5.843e+01 
R3566t2577 n3567 n2578 R=8.652e+00 
R3566t1473 n3567 n1474 R=1.738e+00 
R3567t296 n3568 n297 R=5.496e+00 
R3568t2252 n3569 n2253 R=5.901e+00 
R3569t2385 n3570 n2386 R=1.703e+01 
R3569t457 n3570 n458 R=4.749e+00 
R3570t565 n3571 n566 R=6.726e+00 
R3570t192 n3571 n193 R=3.576e+00 
R3571t1215 n3572 n1216 R=8.620e+00 
R3571t2896 n3572 n2897 R=3.960e+01 
R3573t592 n3574 n593 R=4.754e+00 
R3573t3423 n3574 n3424 R=3.340e+01 
R3573t55 n3574 n56 R=1.117e+01 
R3574t3335 n3575 n3336 R=3.610e+00 
R3574t1684 n3575 n1685 R=4.389e+01 
R3574t2376 n3575 n2377 R=1.000e+01 
R3575t1798 n3576 n1799 R=1.124e+01 
R3576t2482 n3577 n2483 R=5.765e+00 
R3577t811 n3578 n812 R=4.079e+00 
R3578t1961 n3579 n1962 R=9.842e+00 
R3578t1233 n3579 n1234 R=4.672e+00 
R3578t3033 n3579 n3034 R=7.257e+00 
R3579t392 n3580 n393 R=3.827e+01 
R3579t1815 n3580 n1816 R=5.784e+00 
R3579t3256 n3580 n3257 R=1.009e+01 
R3580t1650 n3581 n1651 R=3.961e+00 
R3580t1 n3581 n2 R=5.888e+00 
R3580t3171 n3581 n3172 R=2.896e+01 
R3580t1252 n3581 n1253 R=4.886e+03 
R3581t3071 n3582 n3072 R=5.187e+00 
R3581t597 n3582 n598 R=4.320e+00 
R3582t619 n3583 n620 R=8.420e+00 
R3582t581 n3583 n582 R=3.968e+00 
R3583t1891 n3584 n1892 R=1.087e+01 
R3583t17 n3584 n18 R=7.184e+01 
R3584t1216 n3585 n1217 R=7.646e+00 
R3584t543 n3585 n544 R=8.071e+01 
R3584t354 n3585 n355 R=6.163e+00 
R3585t2600 n3586 n2601 R=6.832e+00 
R3585t569 n3586 n570 R=1.800e+01 
R3586t2647 n3587 n2648 R=3.999e+01 
R3586t2686 n3587 n2687 R=5.716e+00 
R3586t873 n3587 n874 R=8.462e+00 
R3587t1506 n3588 n1507 R=3.158e+01 
R3587t2485 n3588 n2486 R=1.276e+01 
R3587t3130 n3588 n3131 R=5.911e+00 
R3588t2223 n3589 n2224 R=2.729e+00 
R3588t380 n3589 n381 R=8.539e+00 
R3589t263 n3590 n264 R=4.006e+00 
R3589t2534 n3590 n2535 R=1.134e+01 
R3589t1901 n3590 n1902 R=1.933e+01 
R3590t2419 n3591 n2420 R=8.332e+00 
R3590t1367 n3591 n1368 R=1.008e+02 
R3590t3079 n3591 n3080 R=4.869e+00 
R3591t1114 n3592 n1115 R=3.040e+00 
R3591t1108 n3592 n1109 R=1.157e+01 
R3592t529 n3593 n530 R=1.793e+01 
R3592t2711 n3593 n2712 R=2.374e+01 
R3592t242 n3593 n243 R=7.489e+00 
R3593t542 n3594 n543 R=1.713e+01 
R3593t2816 n3594 n2817 R=2.104e+00 
R3593t690 n3594 n691 R=1.755e+00 
R3594t3530 n3595 n3531 R=3.702e+01 
R3594t544 n3595 n545 R=1.373e+01 
R3595t3093 n3596 n3094 R=8.490e+00 
R3595t2298 n3596 n2299 R=1.137e+01 
R3596t2508 n3597 n2509 R=5.806e+00 
R3596t1170 n3597 n1171 R=9.590e+00 
R3597t2988 n3598 n2989 R=7.513e+00 
R3597t300 n3598 n301 R=3.737e+00 
R3598t203 n3599 n204 R=8.161e+01 
R3598t1932 n3599 n1933 R=3.971e+00 
R3598t721 n3599 n722 R=5.827e+00 
R3599t2272 n3600 n2273 R=1.249e+01 
R3600t2818 n3601 n2819 R=5.830e+00 
R3600t2234 n3601 n2235 R=2.824e+01 
R3600t2130 n3601 n2131 R=3.754e+00 
R3600t1570 n3601 n1571 R=5.610e+00 
R3601t1606 n3602 n1607 R=3.994e+00 
R3601t1244 n3602 n1245 R=4.613e+00 
R3601t1000 n3602 n1001 R=1.390e+01 
R3602t1853 n3603 n1854 R=3.785e+00 
R3602t793 n3603 n794 R=3.193e+01 
R3602t459 n3603 n460 R=8.742e+01 
R3602t876 n3603 n877 R=2.909e+01 
R3603t654 n3604 n655 R=1.241e+01 
R3603t2129 n3604 n2130 R=1.020e+01 
R3603t1571 n3604 n1572 R=4.409e+01 
R3604t2033 n3605 n2034 R=4.935e+00 
R3605t2316 n3606 n2317 R=4.160e+01 
R3605t3340 n3606 n3341 R=2.128e+00 
R3605t1123 n3606 n1124 R=1.900e+03 
R3605t1566 n3606 n1567 R=1.330e+01 
R3606t3557 n3607 n3558 R=7.653e+00 
R3606t3009 n3607 n3010 R=3.714e+00 
R3607t1914 n3608 n1915 R=8.166e+00 
R3608t3095 n3609 n3096 R=8.590e+00 
R3608t1078 n3609 n1079 R=5.665e+00 
R3609t291 n3610 n292 R=5.689e+00 
R3609t828 n3610 n829 R=9.890e+00 
R3610t2212 n3611 n2213 R=4.409e+00 
R3610t2566 n3611 n2567 R=2.455e+00 
R3611t399 n3612 n400 R=7.520e+00 
R3611t1136 n3612 n1137 R=6.661e+00 
R3611t1907 n3612 n1908 R=6.582e+00 
R3612t894 n3613 n895 R=2.654e+00 
R3613t827 n3614 n828 R=4.439e+00 
R3614t643 n3615 n644 R=4.843e+00 
R3614t1812 n3615 n1813 R=1.096e+02 
R3614t2881 n3615 n2882 R=9.047e+00 
R3614t2966 n3615 n2967 R=1.476e+01 
R3615t2721 n3616 n2722 R=2.225e+01 
R3615t1747 n3616 n1748 R=6.706e+00 
R3616t388 n3617 n389 R=8.655e+00 
R3616t3060 n3617 n3061 R=4.027e+01 
R3617t3475 n3618 n3476 R=1.981e+00 
R3617t924 n3618 n925 R=8.210e+00 
R3618t3608 n3619 n3609 R=8.737e+00 
R3619t630 n3620 n631 R=3.701e+00 
R3619t1007 n3620 n1008 R=1.742e+01 
R3620t2547 n3621 n2548 R=8.860e+00 
R3620t1646 n3621 n1647 R=8.736e+00 
R3621t697 n3622 n698 R=5.262e+00 
R3622t1755 n3623 n1756 R=3.096e+01 
R3622t3320 n3623 n3321 R=1.742e+01 
R3622t2363 n3623 n2364 R=4.138e+01 
R3622t702 n3623 n703 R=4.740e+00 
R3624t2624 n3625 n2625 R=7.346e+00 
R3625t3613 n3626 n3614 R=2.116e+00 
R3625t827 n3626 n828 R=4.999e+01 
R3626t443 n3627 n444 R=1.532e+01 
R3626t3174 n3627 n3175 R=1.364e+02 
R3627t735 n3628 n736 R=4.401e+01 
R3627t2022 n3628 n2023 R=5.826e+00 
R3628t3512 n3629 n3513 R=8.316e+00 
R3628t3359 n3629 n3360 R=7.970e+00 
R3629t1452 n3630 n1453 R=5.090e+00 
R3629t3062 n3630 n3063 R=1.130e+03 
R3631t2366 n3632 n2367 R=5.873e+00 
R3632t874 n3633 n875 R=8.767e+00 
R3633t2945 n3634 n2946 R=1.027e+01 
R3634t2321 n3635 n2322 R=3.378e+00 
R3634t1812 n3635 n1813 R=2.006e+02 
R3634t3348 n3635 n3349 R=7.012e+00 
R3635t2970 n3636 n2971 R=9.277e+00 
R3635t1569 n3636 n1570 R=9.866e+00 
R3635t837 n3636 n838 R=1.186e+01 
R3636t2637 n3637 n2638 R=3.295e+00 
R3637t3100 n3638 n3101 R=6.153e+00 
R3637t229 n3638 n230 R=1.129e+01 
R3637t2895 n3638 n2896 R=4.427e+01 
R3638t262 n3639 n263 R=2.148e+00 
R3638t2738 n3639 n2739 R=8.127e+00 
R3639t2981 n3640 n2982 R=9.706e+00 
R3639t3068 n3640 n3069 R=2.260e+01 
R3640t634 n3641 n635 R=1.206e+01 
R3640t3034 n3641 n3035 R=4.759e+00 
R3640t3368 n3641 n3369 R=2.061e+00 
R3640t2477 n3641 n2478 R=1.288e+01 
R3641t1687 n3642 n1688 R=7.816e+01 
R3641t3105 n3642 n3106 R=3.170e+00 
R3641t866 n3642 n867 R=3.635e+00 
R3642t2664 n3643 n2665 R=2.877e+00 
R3642t260 n3643 n261 R=3.441e+02 
R3642t890 n3643 n891 R=2.747e+00 
R3642t155 n3643 n156 R=9.448e+00 
R3642t3527 n3643 n3528 R=1.980e+01 
R3643t429 n3644 n430 R=2.653e+00 
R3643t1457 n3644 n1458 R=2.552e+01 
R3643t800 n3644 n801 R=6.000e+00 
R3644t274 n3645 n275 R=2.705e+00 
R3644t409 n3645 n410 R=5.765e+00 
R3644t2365 n3645 n2366 R=8.300e+00 
R3645t291 n3646 n292 R=6.506e+01 
R3645t259 n3646 n260 R=3.733e+00 
R3645t1356 n3646 n1357 R=2.391e+01 
R3646t191 n3647 n192 R=4.252e+00 
R3647t3119 n3648 n3120 R=5.515e+00 
R3647t332 n3648 n333 R=3.547e+00 
R3647t485 n3648 n486 R=8.977e+00 
R3648t2073 n3649 n2074 R=8.587e+01 
R3648t1886 n3649 n1887 R=2.686e+01 
R3649t2015 n3650 n2016 R=3.206e+01 
R3650t2260 n3651 n2261 R=1.033e+02 
R3650t1851 n3651 n1852 R=3.232e+01 
R3650t3513 n3651 n3514 R=2.158e+00 
R3650t739 n3651 n740 R=5.187e+01 
R3651t3234 n3652 n3235 R=5.159e+00 
R3652t2188 n3653 n2189 R=4.690e+01 
R3653t2659 n3654 n2660 R=2.519e+00 
R3653t2706 n3654 n2707 R=6.714e+00 
R3654t870 n3655 n871 R=6.317e+00 
R3654t3327 n3655 n3328 R=9.621e+00 
R3655t1272 n3656 n1273 R=1.907e+01 
R3655t2754 n3656 n2755 R=1.909e+01 
R3655t2163 n3656 n2164 R=4.269e+00 
R3655t674 n3656 n675 R=5.301e+00 
R3658t458 n3659 n459 R=6.599e+00 
R3658t1927 n3659 n1928 R=1.869e+01 
R3658t2558 n3659 n2559 R=5.597e+00 
R3659t2290 n3660 n2291 R=4.038e+00 
R3660t3468 n3661 n3469 R=9.927e+00 
R3661t370 n3662 n371 R=7.243e+01 
R3662t2746 n3663 n2747 R=4.772e+00 
R3662t359 n3663 n360 R=2.913e+00 
R3663t1549 n3664 n1550 R=9.660e+00 
R3663t2957 n3664 n2958 R=6.763e+00 
R3663t567 n3664 n568 R=6.912e+00 
R3663t640 n3664 n641 R=1.411e+01 
R3664t602 n3665 n603 R=2.358e+01 
R3664t3117 n3665 n3118 R=1.212e+01 
R3664t1392 n3665 n1393 R=1.353e+02 
R3664t1591 n3665 n1592 R=8.906e+00 
R3664t1610 n3665 n1611 R=2.939e+01 
R3665t96 n3666 n97 R=8.279e+01 
R3665t2796 n3666 n2797 R=2.529e+00 
R3666t3496 n3667 n3497 R=1.016e+01 
R3666t1294 n3667 n1295 R=3.926e+00 
R3666t2028 n3667 n2029 R=7.038e+00 
R3667t1182 n3668 n1183 R=5.787e+00 
R3668t2946 n3669 n2947 R=2.063e+00 
R3669t3128 n3670 n3129 R=9.550e+00 
R3669t3365 n3670 n3366 R=8.805e+00 
R3670t3516 n3671 n3517 R=3.900e+00 
R3670t680 n3671 n681 R=2.715e+01 
R3670t2393 n3671 n2394 R=7.387e+00 
R3670t2968 n3671 n2969 R=1.229e+01 
R3670t3282 n3671 n3283 R=1.053e+01 
R3671t945 n3672 n946 R=3.804e+01 
R3671t3427 n3672 n3428 R=6.117e+00 
R3672t108 n3673 n109 R=5.157e+00 
R3673t917 n3674 n918 R=3.087e+01 
R3673t789 n3674 n790 R=9.312e+00 
R3674t1652 n3675 n1653 R=1.955e+01 
R3674t2847 n3675 n2848 R=4.101e+00 
R3674t1439 n3675 n1440 R=3.920e+00 
R3674t1337 n3675 n1338 R=9.752e+00 
R3675t109 n3676 n110 R=2.212e+01 
R3676t3228 n3677 n3229 R=4.913e+00 
R3676t1198 n3677 n1199 R=1.285e+01 
R3677t2241 n3678 n2242 R=3.889e+00 
R3677t1329 n3678 n1330 R=1.241e+01 
R3677t2253 n3678 n2254 R=1.089e+01 
R3678t271 n3679 n272 R=3.748e+00 
R3678t730 n3679 n731 R=3.481e+00 
R3678t1374 n3679 n1375 R=3.358e+00 
R3678t1311 n3679 n1312 R=3.877e+01 
R3679t2113 n3680 n2114 R=1.688e+01 
R3680t1463 n3681 n1464 R=5.377e+00 
R3681t1110 n3682 n1111 R=9.052e+01 
R3681t756 n3682 n757 R=4.003e+00 
R3682t2296 n3683 n2297 R=9.265e+00 
R3683t2563 n3684 n2564 R=1.517e+02 
R3683t1185 n3684 n1186 R=5.478e+00 
R3684t3016 n3685 n3017 R=5.556e+00 
R3684t260 n3685 n261 R=1.228e+01 
R3685t2037 n3686 n2038 R=3.848e+00 
R3685t3042 n3686 n3043 R=4.401e+00 
R3686t3007 n3687 n3008 R=1.855e+01 
R3686t1251 n3687 n1252 R=3.737e+00 
R3686t3063 n3687 n3064 R=1.120e+01 
R3687t2197 n3688 n2198 R=4.351e+00 
R3687t3577 n3688 n3578 R=3.519e+00 
R3688t1809 n3689 n1810 R=3.310e+00 
R3688t2465 n3689 n2466 R=5.797e+01 
R3688t2519 n3689 n2520 R=3.442e+00 
R3689t770 n3690 n771 R=8.081e+00 
R3689t1419 n3690 n1420 R=1.023e+01 
R3689t1626 n3690 n1627 R=4.058e+01 
R3690t142 n3691 n143 R=1.223e+01 
R3691t413 n3692 n414 R=1.838e+01 
R3691t1573 n3692 n1574 R=5.596e+00 
R3692t1981 n3693 n1982 R=9.035e+00 
R3692t3136 n3693 n3137 R=1.137e+01 
R3692t604 n3693 n605 R=6.938e+01 
R3692t3547 n3693 n3548 R=4.715e+00 
R3692t1613 n3693 n1614 R=1.008e+01 
R3693t107 n3694 n108 R=7.052e+00 
R3693t2627 n3694 n2628 R=8.736e+00 
R3693t1870 n3694 n1871 R=8.843e+01 
R3694t1010 n3695 n1011 R=3.652e+00 
R3695t494 n3696 n495 R=1.094e+02 
R3695t3070 n3696 n3071 R=5.678e+00 
R3695t778 n3696 n779 R=3.718e+00 
R3695t126 n3696 n127 R=1.575e+02 
R3696t1952 n3697 n1953 R=1.055e+01 
R3696t3387 n3697 n3388 R=5.566e+00 
R3697t2442 n3698 n2443 R=1.107e+01 
R3697t2876 n3698 n2877 R=1.477e+01 
R3698t2992 n3699 n2993 R=3.467e+00 
R3699t804 n3700 n805 R=1.762e+01 
R3699t1253 n3700 n1254 R=3.795e+01 
R3700t2027 n3701 n2028 R=2.962e+01 
R3701t3077 n3702 n3078 R=2.931e+00 
R3703t1032 n3704 n1033 R=5.542e+01 
R3703t1514 n3704 n1515 R=8.354e+00 
R3703t2416 n3704 n2417 R=4.203e+00 
R3704t721 n3705 n722 R=2.867e+01 
R3704t3598 n3705 n3599 R=9.906e+01 
R3705t546 n3706 n547 R=2.166e+00 
R3705t2423 n3706 n2424 R=2.334e+00 
R3705t1225 n3706 n1226 R=1.941e+01 
R3706t3304 n3707 n3305 R=2.073e+01 
R3706t633 n3707 n634 R=1.827e+01 
R3707t3575 n3708 n3576 R=1.160e+01 
R3707t1423 n3708 n1424 R=1.431e+01 
R3708t2977 n3709 n2978 R=4.362e+00 
R3708t2308 n3709 n2309 R=2.811e+00 
R3708t1465 n3709 n1466 R=9.842e+00 
R3708t682 n3709 n683 R=1.914e+01 
R3709t2991 n3710 n2992 R=5.245e+00 
R3709t2443 n3710 n2444 R=6.576e+00 
R3710t3054 n3711 n3055 R=4.503e+00 
R3711t980 n3712 n981 R=4.461e+00 
R3711t993 n3712 n994 R=3.618e+00 
R3711t2413 n3712 n2414 R=3.142e+00 
R3711t3488 n3712 n3489 R=2.933e+01 
R3712t1949 n3713 n1950 R=5.354e+00 
R3713t2599 n3714 n2600 R=1.031e+01 
R3714t3212 n3715 n3213 R=9.965e+00 
R3714t336 n3715 n337 R=1.345e+01 
R3714t2127 n3715 n2128 R=5.411e+01 
R3714t1817 n3715 n1818 R=1.598e+01 
R3714t2186 n3715 n2187 R=2.755e+00 
R3715t1407 n3716 n1408 R=7.230e+01 
R3715t3607 n3716 n3608 R=6.665e+00 
R3715t2383 n3716 n2384 R=2.167e+02 
R3715t1313 n3716 n1314 R=1.006e+02 
R3716t275 n3717 n276 R=7.302e+01 
R3716t1405 n3717 n1406 R=1.374e+01 
R3716t600 n3717 n601 R=2.131e+01 
R3716t1768 n3717 n1769 R=2.302e+00 
R3717t3661 n3718 n3662 R=1.514e+01 
R3717t2944 n3718 n2945 R=6.546e+00 
R3717t2848 n3718 n2849 R=1.217e+01 
R3718t2760 n3719 n2761 R=3.200e+00 
R3719t2513 n3720 n2514 R=7.074e+00 
R3719t3648 n3720 n3649 R=7.592e+00 
R3720t1824 n3721 n1825 R=6.693e+01 
R3720t2315 n3721 n2316 R=5.205e+01 
R3721t2317 n3722 n2318 R=6.666e+00 
R3721t2695 n3722 n2696 R=3.891e+00 
R3722t924 n3723 n925 R=7.426e+00 
R3722t3617 n3723 n3618 R=2.817e+01 
R3722t3186 n3723 n3187 R=4.153e+01 
R3723t1408 n3724 n1409 R=3.638e+00 
R3723t3668 n3724 n3669 R=7.743e+00 
R3723t2946 n3724 n2947 R=5.534e+03 
R3724t1265 n3725 n1266 R=2.049e+01 
R3724t801 n3725 n802 R=3.067e+01 
R3725t658 n3726 n659 R=9.963e+00 
R3725t1790 n3726 n1791 R=1.628e+01 
R3726t3718 n3727 n3719 R=2.311e+02 
R3726t1796 n3727 n1797 R=7.128e+00 
R3726t2337 n3727 n2338 R=4.333e+00 
R3727t1384 n3728 n1385 R=2.754e+01 
R3727t2085 n3728 n2086 R=4.425e+00 
R3728t3166 n3729 n3167 R=6.464e+00 
R3728t3443 n3729 n3444 R=1.268e+01 
R3728t995 n3729 n996 R=3.858e+00 
R3728t461 n3729 n462 R=2.714e+01 
R3729t250 n3730 n251 R=5.189e+00 
R3729t3523 n3730 n3524 R=1.263e+01 
R3729t1523 n3730 n1524 R=4.034e+00 
R3730t2243 n3731 n2244 R=5.060e+00 
R3730t3185 n3731 n3186 R=6.244e+00 
R3730t1026 n3731 n1027 R=1.503e+01 
R3730t3065 n3731 n3066 R=6.747e+00 
R3732t752 n3733 n753 R=3.744e+00 
R3733t1512 n3734 n1513 R=1.144e+02 
R3733t2396 n3734 n2397 R=7.943e+00 
R3733t973 n3734 n974 R=3.123e+01 
R3733t324 n3734 n325 R=1.205e+01 
R3733t3058 n3734 n3059 R=1.221e+01 
R3733t422 n3734 n423 R=7.029e+00 
R3733t1012 n3734 n1013 R=3.117e+01 
R3734t114 n3735 n115 R=1.238e+01 
R3734t346 n3735 n347 R=4.295e+00 
R3734t261 n3735 n262 R=1.008e+01 
R3734t1535 n3735 n1536 R=2.825e+02 
R3734t1817 n3735 n1818 R=9.870e+00 
R3734t918 n3735 n919 R=7.238e+00 
R3735t2067 n3736 n2068 R=3.661e+00 
R3735t771 n3736 n772 R=1.118e+01 
R3736t1157 n3737 n1158 R=2.350e+01 
R3736t3160 n3737 n3161 R=7.339e+00 
R3736t2113 n3737 n2114 R=1.528e+01 
R3737t1637 n3738 n1638 R=2.321e+00 
R3737t1381 n3738 n1382 R=3.586e+01 
R3738t1822 n3739 n1823 R=9.830e+00 
R3738t2710 n3739 n2711 R=4.727e+00 
R3738t1917 n3739 n1918 R=4.012e+00 
R3738t1384 n3739 n1385 R=4.819e+01 
R3739t1671 n3740 n1672 R=5.558e+00 
R3739t3453 n3740 n3454 R=4.613e+00 
R3740t765 n3741 n766 R=1.940e+01 
R3740t140 n3741 n141 R=1.690e+00 
R3740t2493 n3741 n2494 R=3.027e+01 
R3741t1816 n3742 n1817 R=5.123e+00 
R3741t1697 n3742 n1698 R=4.448e+00 
R3741t1220 n3742 n1221 R=4.662e+01 
R3741t559 n3742 n560 R=3.822e+00 
R3741t950 n3742 n951 R=1.858e+01 
R3742t2841 n3743 n2842 R=5.302e+01 
R3742t2144 n3743 n2145 R=4.701e+00 
R3743t1020 n3744 n1021 R=5.814e+00 
R3743t2134 n3744 n2135 R=6.801e+00 
R3743t2559 n3744 n2560 R=4.681e+00 
R3744t626 n3745 n627 R=9.209e+00 
R3744t3574 n3745 n3575 R=4.693e+00 
R3745t2013 n3746 n2014 R=1.436e+01 
R3745t3080 n3746 n3081 R=3.403e+01 
R3745t2762 n3746 n2763 R=1.327e+01 
R3746t1138 n3747 n1139 R=9.300e+01 
R3747t686 n3748 n687 R=1.656e+01 
R3747t745 n3748 n746 R=3.496e+00 
R3747t548 n3748 n549 R=3.712e+00 
R3747t2473 n3748 n2474 R=2.046e+01 
R3748t846 n3749 n847 R=1.212e+01 
R3748t2495 n3749 n2496 R=5.774e+00 
R3748t239 n3749 n240 R=4.946e+00 
R3748t533 n3749 n534 R=1.096e+01 
R3748t3501 n3749 n3502 R=1.016e+01 
R3749t2787 n3750 n2788 R=4.155e+00 
R3750t3012 n3751 n3013 R=3.243e+00 
R3750t1491 n3751 n1492 R=7.326e+00 
R3750t2648 n3751 n2649 R=6.701e+00 
R3751t1718 n3752 n1719 R=7.178e+00 
R3751t2562 n3752 n2563 R=2.144e+01 
R3752t1246 n3753 n1247 R=2.887e+00 
R3752t847 n3753 n848 R=2.337e+00 
R3753t1067 n3754 n1068 R=7.298e+00 
R3754t3172 n3755 n3173 R=1.017e+01 
R3755t1414 n3756 n1415 R=1.096e+01 
R3755t3558 n3756 n3559 R=6.961e+00 
R3756t1699 n3757 n1700 R=9.745e+00 
R3756t2515 n3757 n2516 R=5.007e+00 
R3756t714 n3757 n715 R=2.776e+01 
R3756t41 n3757 n42 R=2.956e+00 
R3757t1069 n3758 n1070 R=2.501e+01 
R3757t1530 n3758 n1531 R=1.814e+01 
R3757t2448 n3758 n2449 R=9.375e+01 
R3757t787 n3758 n788 R=5.588e+00 
R3758t2677 n3759 n2678 R=6.298e+00 
R3758t1575 n3759 n1576 R=6.453e+00 
R3758t3095 n3759 n3096 R=2.333e+01 
R3758t3608 n3759 n3609 R=5.639e+00 
R3759t1825 n3760 n1826 R=4.999e+01 
R3759t3345 n3760 n3346 R=3.722e+00 
R3759t461 n3760 n462 R=1.032e+01 
R3759t475 n3760 n476 R=6.765e+00 
R3759t362 n3760 n363 R=5.299e+00 
R3760t2073 n3761 n2074 R=4.344e+01 
R3760t3648 n3761 n3649 R=1.860e+00 
R3761t2165 n3762 n2166 R=7.134e+00 
R3761t3046 n3762 n3047 R=2.262e+01 
R3762t146 n3763 n147 R=1.133e+01 
R3762t2106 n3763 n2107 R=3.432e+00 
R3762t3175 n3763 n3176 R=1.913e+01 
R3763t1984 n3764 n1985 R=1.851e+00 
R3763t2352 n3764 n2353 R=1.467e+01 
R3763t563 n3764 n564 R=3.294e+00 
R3764t1737 n3765 n1738 R=5.829e+00 
R3765t2718 n3766 n2719 R=5.495e+00 
R3765t556 n3766 n557 R=4.166e+00 
R3766t1459 n3767 n1460 R=2.177e+01 
R3767t1212 n3768 n1213 R=2.754e+01 
R3767t2870 n3768 n2871 R=1.874e+01 
R3767t2142 n3768 n2143 R=1.294e+01 
R3767t1760 n3768 n1761 R=4.448e+00 
R3769t2886 n3770 n2887 R=1.785e+00 
R3769t1745 n3770 n1746 R=3.202e+00 
R3770t1284 n3771 n1285 R=7.382e+01 
R3770t2297 n3771 n2298 R=9.437e+00 
R3770t1880 n3771 n1881 R=1.639e+01 
R3771t2045 n3772 n2046 R=2.241e+01 
R3771t871 n3772 n872 R=1.053e+01 
R3771t2616 n3772 n2617 R=8.797e+00 
R3772t2731 n3773 n2732 R=5.844e+01 
R3773t1973 n3774 n1974 R=6.664e+00 
R3774t3451 n3775 n3452 R=5.137e+00 
R3774t2249 n3775 n2250 R=1.679e+01 
R3774t1672 n3775 n1673 R=7.872e+01 
R3774t3163 n3775 n3164 R=1.067e+01 
R3775t2274 n3776 n2275 R=6.249e+00 
R3775t2230 n3776 n2231 R=3.943e+00 
R3776t3695 n3777 n3696 R=1.428e+01 
R3776t778 n3777 n779 R=6.555e+00 
R3776t3067 n3777 n3068 R=1.160e+02 
R3776t427 n3777 n428 R=6.005e+00 
R3777t332 n3778 n333 R=3.455e+00 
R3777t829 n3778 n830 R=1.267e+02 
R3779t1124 n3780 n1125 R=6.679e+01 
R3779t1174 n3780 n1175 R=1.367e+01 
R3779t3107 n3780 n3108 R=6.194e+00 
R3779t232 n3780 n233 R=6.313e+00 
R3779t1580 n3780 n1581 R=7.437e+01 
R3780t1083 n3781 n1084 R=5.973e+00 
R3780t1791 n3781 n1792 R=1.864e+02 
R3780t1343 n3781 n1344 R=4.441e+00 
R3780t1607 n3781 n1608 R=6.317e+00 
R3781t2884 n3782 n2885 R=1.671e+01 
R3781t1559 n3782 n1560 R=7.029e+00 
R3782t1255 n3783 n1256 R=6.021e+00 
R3783t109 n3784 n110 R=1.307e+01 
R3783t2423 n3784 n2424 R=7.151e+00 
R3783t546 n3784 n547 R=1.436e+01 
R3784t1314 n3785 n1315 R=4.718e+00 
R3784t2967 n3785 n2968 R=1.589e+01 
R3785t737 n3786 n738 R=6.402e+00 
R3785t1725 n3786 n1726 R=1.516e+01 
R3785t82 n3786 n83 R=5.418e+02 
R3785t583 n3786 n584 R=3.612e+01 
R3786t2831 n3787 n2832 R=1.378e+01 
R3786t2326 n3787 n2327 R=1.018e+01 
R3786t337 n3787 n338 R=1.344e+01 
R3786t3493 n3787 n3494 R=5.964e+00 
R3787t743 n3788 n744 R=6.473e+00 
R3787t2615 n3788 n2616 R=3.976e+01 
R3787t198 n3788 n199 R=1.182e+01 
R3788t535 n3789 n536 R=1.249e+02 
R3788t3419 n3789 n3420 R=2.398e+00 
R3788t1594 n3789 n1595 R=2.665e+01 
R3788t2912 n3789 n2913 R=6.590e+00 
R3788t759 n3789 n760 R=2.838e+00 
R3789t376 n3790 n377 R=2.707e+00 
R3789t1920 n3790 n1921 R=2.671e+01 
R3790t2196 n3791 n2197 R=7.522e+00 
R3791t2836 n3792 n2837 R=1.996e+02 
R3791t3482 n3792 n3483 R=1.007e+01 
R3791t1597 n3792 n1598 R=1.134e+01 
R3791t69 n3792 n70 R=6.838e+00 
R3791t194 n3792 n195 R=3.460e+01 
R3791t3131 n3792 n3132 R=9.307e+00 
R3793t1909 n3794 n1910 R=4.338e+00 
R3794t122 n3795 n123 R=8.918e+00 
R3795t1379 n3796 n1380 R=1.890e+00 
R3796t1271 n3797 n1 R=1.854e+01 
R3796t1650 n3797 n1651 R=4.948e+00 
R3797t1572 n3798 n1573 R=4.587e+02 
R3797t1881 n3798 n1882 R=5.327e+00 
R3797t3731 n3798 n3732 R=2.467e+00 
R3798t300 n3799 n301 R=1.604e+01 
R3798t3597 n3799 n3598 R=8.818e+00 
R3798t1642 n3799 n1643 R=9.596e+00 
R3798t328 n3799 n329 R=4.266e+00 
R3798t752 n3799 n753 R=2.593e+01 
R3798t3732 n3799 n3733 R=1.218e+01 
R3798t3189 n3799 n3190 R=8.565e+00 
R3799t3069 n3800 n3070 R=1.140e+01 
R3799t1030 n3800 n1031 R=2.380e+01 
R3799t3724 n3800 n3725 R=4.956e+01 
R3800t2925 n3801 n2926 R=6.236e+00 
R3801t464 n3802 n465 R=3.992e+02 
R3801t1217 n3802 n1218 R=3.101e+00 
R3802t2988 n3803 n2989 R=1.001e+02 
R3802t8 n3803 n9 R=5.183e+00 
R3803t2105 n3804 n2106 R=5.965e+00 
R3803t3175 n3804 n3176 R=4.157e+00 
R3803t3762 n3804 n3763 R=2.399e+01 
R3803t2106 n3804 n2107 R=5.201e+00 
R3804t3511 n3805 n3512 R=9.356e+00 
R3804t1157 n3805 n1158 R=4.136e+00 
R3804t3794 n3805 n3795 R=6.183e+01 
R3805t543 n3806 n544 R=2.522e+01 
R3805t418 n3806 n419 R=1.663e+00 
R3806t2094 n3807 n2095 R=1.129e+01 
R3806t1373 n3807 n1374 R=8.766e+00 
R3807t1850 n3808 n1851 R=8.664e+00 
R3807t2344 n3808 n2345 R=1.237e+01 
R3807t1449 n3808 n1450 R=3.054e+00 
R3808t1955 n3809 n1956 R=9.895e+00 
R3808t1049 n3809 n1050 R=4.965e+00 
R3808t2221 n3809 n2222 R=5.673e+00 
R3809t74 n3810 n75 R=2.999e+01 
R3809t1584 n3810 n1585 R=6.490e+00 
R3809t3503 n3810 n3504 R=9.478e+00 
R3810t1693 n3811 n1694 R=7.485e+01 
R3810t3499 n3811 n3500 R=7.532e+00 
R3811t1450 n3812 n1451 R=3.082e+01 
R3811t1092 n3812 n1093 R=4.771e+00 
R3812t688 n3813 n689 R=4.187e+00 
R3812t813 n3813 n814 R=4.992e+00 
R3813t3619 n3814 n3620 R=5.824e+00 
R3813t3807 n3814 n3808 R=1.972e+01 
R3813t1997 n3814 n1998 R=3.013e+00 
R3814t1204 n3815 n1205 R=3.983e+00 
R3814t1678 n3815 n1679 R=6.256e+00 
R3814t3255 n3815 n3256 R=1.445e+01 
R3815t3761 n3816 n3762 R=1.040e+01 
R3816t2285 n3817 n2286 R=2.333e+00 
R3816t2482 n3817 n2483 R=2.721e+01 
R3816t3576 n3817 n3577 R=2.451e+00 
R3817t2277 n3818 n2278 R=3.220e+00 
R3817t2014 n3818 n2015 R=3.724e+01 
R3818t1139 n3819 n1140 R=6.893e+00 
R3819t2964 n3820 n2965 R=3.519e+00 
R3820t520 n3821 n521 R=1.206e+01 
R3820t566 n3821 n567 R=2.589e+01 
R3821t3075 n3822 n3076 R=2.505e+00 
R3821t3291 n3822 n3292 R=1.745e+00 
R3821t61 n3822 n62 R=2.094e+02 
R3821t91 n3822 n92 R=6.516e+01 
R3822t129 n3823 n130 R=3.181e+00 
R3822t465 n3823 n466 R=6.237e+00 
R3823t2339 n3824 n2340 R=1.099e+01 
R3823t99 n3824 n100 R=3.149e+00 
R3824t1184 n3825 n1185 R=5.135e+02 
R3824t3818 n3825 n3819 R=5.633e+00 
R3824t1307 n3825 n1308 R=4.490e+00 
R3825t2130 n3826 n2131 R=3.873e+00 
R3826t2235 n3827 n2236 R=3.758e+00 
R3826t1907 n3827 n1908 R=1.203e+01 
R3827t748 n3828 n749 R=3.856e+00 
R3828t339 n3829 n340 R=2.552e+01 
R3828t1834 n3829 n1835 R=6.661e+00 
R3828t455 n3829 n456 R=1.296e+01 
R3828t1888 n3829 n1889 R=6.509e+00 
R3829t2334 n3830 n2335 R=7.394e+00 
R3829t1713 n3830 n1714 R=2.135e+00 
R3829t1401 n3830 n1402 R=6.980e+00 
R3829t1968 n3830 n1969 R=7.341e+00 
R3830t464 n3831 n465 R=5.771e+00 
R3830t1819 n3831 n1820 R=5.017e+00 
R3831t701 n3832 n702 R=3.603e+00 
R3832t313 n3833 n314 R=5.571e+00 
R3833t2342 n3834 n2343 R=4.487e+00 
R3834t1900 n3835 n1901 R=7.274e+00 
R3834t2265 n3835 n2266 R=1.204e+01 
R3834t581 n3835 n582 R=6.960e+00 
R3835t1150 n3836 n1151 R=7.735e+00 
R3835t2934 n3836 n2935 R=3.035e+00 
R3835t723 n3836 n724 R=1.075e+02 
R3836t2499 n3837 n2500 R=3.612e+00 
R3836t348 n3837 n349 R=1.317e+01 
R3836t3473 n3837 n3474 R=5.053e+00 
R3837t818 n3838 n819 R=2.805e+00 
R3838t3272 n3839 n3273 R=2.379e+00 
R3838t3050 n3839 n3051 R=1.101e+01 
R3838t3490 n3839 n3491 R=8.665e+00 
R3839t650 n3840 n651 R=1.019e+01 
R3839t2039 n3840 n2040 R=2.095e+01 
R3840t577 n3841 n578 R=4.756e+01 
R3840t1989 n3841 n1990 R=7.227e+00 
R3840t2194 n3841 n2195 R=9.575e+00 
R3840t2997 n3841 n2998 R=1.263e+01 
R3840t3041 n3841 n3042 R=3.938e+00 
R3841t1191 n3842 n1192 R=3.006e+01 
R3841t3350 n3842 n3351 R=3.189e+00 
R3841t2599 n3842 n2600 R=2.117e+01 
R3841t2762 n3842 n2763 R=2.240e+00 
R3841t820 n3842 n821 R=1.064e+02 
R3842t710 n3843 n711 R=3.521e+02 
R3842t3044 n3843 n3045 R=1.671e+01 
R3842t2159 n3843 n2160 R=6.736e+00 
R3843t539 n3844 n540 R=2.741e+00 
R3843t1842 n3844 n1843 R=5.136e+00 
R3844t3030 n3845 n3031 R=1.114e+01 
R3844t1029 n3845 n1030 R=1.808e+00 
R3844t1925 n3845 n1926 R=2.274e+00 
R3845t1908 n3846 n1909 R=7.678e+00 
R3846t852 n3847 n853 R=1.583e+01 
R3846t2613 n3847 n2614 R=9.194e+00 
R3846t2258 n3847 n2259 R=2.345e+01 
R3847t3452 n3848 n3453 R=1.664e+01 
R3848t1131 n3849 n1132 R=3.973e+00 
R3848t2836 n3849 n2837 R=4.755e+00 
R3848t3482 n3849 n3483 R=1.762e+02 
R3848t1661 n3849 n1662 R=1.135e+01 
R3848t3112 n3849 n3113 R=6.076e+00 
R3848t2652 n3849 n2653 R=2.014e+01 
R3849t2683 n3850 n2684 R=1.236e+01 
R3850t740 n3851 n741 R=5.547e+00 
R3850t2008 n3851 n2009 R=8.436e+00 
R3851t2143 n3852 n2144 R=4.162e+00 
R3851t65 n3852 n66 R=5.406e+00 
R3853t3094 n3854 n3095 R=1.279e+01 
R3853t907 n3854 n908 R=2.153e+01 
R3853t3698 n3854 n3699 R=1.190e+01 
R3854t2604 n3855 n2605 R=4.206e+00 
R3854t1931 n3855 n1932 R=8.153e+01 
R3854t2744 n3855 n2745 R=5.042e+00 
R3855t2972 n3856 n2973 R=1.478e+01 
R3855t3466 n3856 n3467 R=2.828e+00 
R3856t467 n3857 n468 R=3.679e+00 
R3856t1198 n3857 n1199 R=1.450e+01 
R3857t1245 n3858 n1246 R=3.501e+00 
R3858t1077 n3859 n1078 R=4.780e+01 
R3858t3322 n3859 n3323 R=2.983e+00 
R3859t3076 n3860 n3077 R=5.416e+00 
R3859t104 n3860 n105 R=5.679e+00 
R3859t1291 n3860 n1292 R=5.936e+00 
R3860t1713 n3861 n1714 R=1.367e+01 
R3860t1814 n3861 n1815 R=2.045e+01 
R3860t2975 n3861 n2976 R=3.588e+02 
R3861t3141 n3862 n3142 R=1.464e+01 
R3861t1574 n3862 n1575 R=4.126e+00 
R3861t835 n3862 n836 R=1.459e+01 
R3863t1327 n3864 n1328 R=4.181e+00 
R3863t2992 n3864 n2993 R=7.428e+01 
R3864t687 n3865 n688 R=4.680e+00 
R3865t896 n3866 n897 R=6.654e+00 
R3865t460 n3866 n461 R=2.475e+02 
R3865t823 n3866 n824 R=6.294e+00 
R3866t2057 n3867 n2058 R=3.657e+00 
R3866t254 n3867 n255 R=2.803e+01 
R3867t1840 n3868 n1841 R=2.293e+01 
R3868t32 n3869 n33 R=1.979e+01 
R3868t3093 n3869 n3094 R=3.988e+02 
R3868t3595 n3869 n3596 R=2.245e+00 
R3869t2872 n3870 n2873 R=1.450e+01 
R3869t2568 n3870 n2569 R=7.757e+00 
R3869t1846 n3870 n1847 R=4.216e+00 
R3870t36 n3871 n37 R=2.323e+01 
R3871t1098 n3872 n1099 R=3.956e+00 
R3871t3208 n3872 n3209 R=7.212e+00 
R3871t3030 n3872 n3031 R=6.645e+00 
R3871t2125 n3872 n2126 R=8.633e+00 
R3872t1539 n3873 n1540 R=4.101e+00 
R3873t121 n3874 n122 R=3.704e+00 
R3873t2784 n3874 n2785 R=9.999e+01 
R3873t2158 n3874 n2159 R=5.626e+00 
R3874t1776 n3875 n1777 R=4.501e+00 
R3874t1925 n3875 n1926 R=4.527e+00 
R3875t1349 n3876 n1350 R=1.313e+01 
R3875t2874 n3876 n2875 R=5.512e+00 
R3875t258 n3876 n259 R=2.047e+00 
R3876t125 n3877 n126 R=6.179e+00 
R3877t2172 n3878 n2173 R=1.210e+01 
R3879t1891 n3880 n1892 R=5.506e+00 
R3879t2557 n3880 n2558 R=1.305e+01 
R3879t2535 n3880 n2536 R=4.228e+01 
R3879t822 n3880 n823 R=5.745e+00 
R3879t17 n3880 n18 R=3.019e+01 
R3879t3583 n3880 n3584 R=4.625e+00 
R3880t1147 n3881 n1148 R=5.218e+00 
R3880t2483 n3881 n2484 R=3.381e+00 
R3881t406 n3882 n407 R=6.516e+00 
R3881t473 n3882 n474 R=4.217e+00 
R3881t1133 n3882 n1134 R=7.200e+00 
R3881t2487 n3882 n2488 R=2.415e+01 
R3882t2833 n3883 n2834 R=1.114e+01 
R3882t3633 n3883 n3634 R=1.589e+01 
R3883t2823 n3884 n2824 R=5.446e+00 
R3883t466 n3884 n467 R=2.605e+02 
R3884t3431 n3885 n3432 R=2.236e+00 
R3884t2386 n3885 n2387 R=4.365e+00 
R3885t1806 n3886 n1807 R=9.213e+00 
R3885t1247 n3886 n1248 R=3.786e+00 
R3886t97 n3887 n98 R=3.441e+00 
R3886t3618 n3887 n3619 R=2.081e+01 
R3888t1046 n3889 n1047 R=1.233e+01 
R3890t2595 n3891 n2596 R=3.240e+00 
R3891t1797 n3892 n1798 R=1.987e+00 
R3891t1519 n3892 n1520 R=1.278e+01 
R3891t631 n3892 n632 R=2.188e+00 
R3892t3396 n3893 n3397 R=1.208e+01 
R3892t43 n3893 n44 R=1.312e+01 
R3892t1524 n3893 n1525 R=3.219e+00 
R3893t2333 n3894 n2334 R=3.108e+00 
R3893t2576 n3894 n2577 R=1.575e+01 
R3894t1211 n3895 n1212 R=4.876e+00 
R3894t1677 n3895 n1678 R=1.957e+01 
R3894t1548 n3895 n1549 R=2.650e+00 
R3895t2331 n3896 n2332 R=7.809e+00 
R3895t108 n3896 n109 R=1.399e+01 
R3895t1836 n3896 n1837 R=2.196e+01 
R3895t964 n3896 n965 R=3.928e+00 
R3896t658 n3897 n659 R=4.703e+00 
R3896t454 n3897 n455 R=2.651e+00 
R3896t3852 n3897 n3853 R=4.492e+01 
R3897t88 n3898 n89 R=1.310e+01 
R3897t1476 n3898 n1477 R=2.280e+02 
R3898t552 n3899 n553 R=4.663e+00 
R3898t2763 n3899 n2764 R=5.685e+01 
R3898t1924 n3899 n1925 R=4.281e+00 
R3898t3225 n3899 n3226 R=3.062e+01 
R3899t3103 n3900 n3104 R=9.615e+00 
R3899t1830 n3900 n1831 R=2.233e+01 
R3899t1077 n3900 n1078 R=2.569e+01 
R3900t60 n3901 n61 R=1.733e+01 
R3900t2258 n3901 n2259 R=2.100e+01 
R3900t3397 n3901 n3398 R=1.000e+01 
R3901t1983 n3902 n1984 R=8.571e+00 
R3901t1487 n3902 n1488 R=3.157e+00 
R3902t1240 n3903 n1241 R=4.040e+00 
R3902t2821 n3903 n2822 R=3.972e+00 
R3903t955 n3904 n956 R=2.109e+01 
R3903t1837 n3904 n1838 R=2.185e+01 
R3904t920 n3905 n921 R=2.074e+01 
R3904t2145 n3905 n2146 R=1.861e+00 
R3905t1960 n3906 n1961 R=2.571e+00 
R3905t2138 n3906 n2139 R=1.739e+01 
R3905t716 n3906 n717 R=1.224e+01 
R3906t464 n3907 n465 R=4.907e+00 
R3906t3830 n3907 n3831 R=1.761e+01 
R3906t2755 n3907 n2756 R=2.237e+01 
R3906t1819 n3907 n1820 R=8.273e+00 
R3907t2478 n3908 n2479 R=7.731e+00 
R3907t3347 n3908 n3348 R=4.557e+00 
R3907t2917 n3908 n2918 R=6.453e+00 
R3908t836 n3909 n837 R=3.544e+00 
R3909t3203 n3910 n3204 R=4.774e+01 
R3910t2273 n3911 n2274 R=3.982e+00 
R3910t851 n3911 n852 R=1.373e+01 
R3911t287 n3912 n288 R=7.472e+00 
R3911t2547 n3912 n2548 R=1.387e+01 
R3911t2178 n3912 n2179 R=1.011e+01 
R3912t1922 n3913 n1923 R=1.288e+01 
R3912t1813 n3913 n1814 R=3.933e+01 
R3913t1707 n3914 n1708 R=4.313e+00 
R3913t3908 n3914 n3909 R=6.189e+00 
R3914t3152 n3915 n3153 R=7.177e+00 
R3915t31 n3916 n32 R=2.534e+01 
R3915t2617 n3916 n2618 R=3.332e+02 
R3915t2098 n3916 n2099 R=7.264e+00 
R3916t698 n3917 n699 R=1.457e+01 
R3916t1091 n3917 n1092 R=1.623e+01 
R3916t497 n3917 n498 R=6.108e+00 
R3916t1847 n3917 n1848 R=4.847e+00 
R3916t1628 n3917 n1629 R=3.543e+01 
R3916t1094 n3917 n1095 R=3.933e+00 
R3917t2941 n3918 n2942 R=5.579e+01 
R3917t1146 n3918 n1147 R=2.777e+00 
R3917t1760 n3918 n1761 R=8.806e+01 
R3917t3767 n3918 n3768 R=1.820e+01 
R3918t542 n3919 n543 R=4.144e+00 
R3919t3514 n3920 n3515 R=2.544e+01 
R3919t1880 n3920 n1881 R=1.237e+01 
R3920t1803 n3921 n1804 R=2.691e+01 
R3920t1716 n3921 n1717 R=9.898e+00 
R3922t1711 n3923 n1712 R=2.911e+00 
R3922t672 n3923 n673 R=2.481e+01 
R3923t3632 n3924 n3633 R=3.097e+00 
R3923t874 n3924 n875 R=5.744e+00 
R3924t2964 n3925 n2965 R=1.085e+01 
R3924t3819 n3925 n3820 R=8.628e+00 
R3924t2522 n3925 n2523 R=2.817e+01 
R3925t2887 n3926 n2888 R=5.645e+00 
R3925t2527 n3926 n2528 R=5.125e+00 
R3925t1511 n3926 n1512 R=4.623e+00 
R3926t3897 n3927 n3898 R=2.363e+00 
R3926t1476 n3927 n1477 R=5.473e+00 
R3927t895 n3928 n896 R=2.128e+00 
R3928t1375 n3929 n1376 R=3.791e+01 
R3928t3656 n3929 n3657 R=6.314e+00 
R3929t710 n3930 n711 R=3.965e+00 
R3929t3842 n3930 n3843 R=8.763e+00 
R3929t2159 n3930 n2160 R=1.003e+01 
R3929t2733 n3930 n2734 R=1.695e+02 
R3930t3443 n3931 n3444 R=3.123e+01 
R3930t29 n3931 n30 R=5.815e+00 
R3930t811 n3931 n812 R=1.694e+01 
R3931t806 n3932 n807 R=1.503e+01 
R3931t756 n3932 n757 R=1.648e+01 
R3931t3681 n3932 n3682 R=1.021e+01 
R3932t401 n3933 n402 R=3.523e+00 
R3932t2719 n3933 n2720 R=7.206e+01 
R3933t1240 n3934 n1241 R=2.707e+01 
R3933t3902 n3934 n3903 R=4.666e+00 
R3934t1582 n3935 n1583 R=2.135e+00 
R3936t2562 n3937 n2563 R=4.491e+00 
R3937t2146 n3938 n2147 R=4.852e+00 
R3937t2218 n3938 n2219 R=1.835e+01 
R3937t2797 n3938 n2798 R=5.405e+00 
R3937t913 n3938 n914 R=9.656e+00 
R3938t1088 n3939 n1089 R=3.959e+00 
R3939t646 n3940 n647 R=4.060e+00 
R3939t1916 n3940 n1917 R=4.357e+00 
R3939t3686 n3940 n3687 R=4.914e+01 
R3939t1251 n3940 n1252 R=6.124e+01 
R3940t1875 n3941 n1876 R=1.322e+02 
R3940t2261 n3941 n2262 R=3.721e+00 
R3941t562 n3942 n563 R=1.427e+01 
R3941t3173 n3942 n3174 R=3.129e+00 
R3942t1783 n3943 n1784 R=3.903e+00 
R3942t165 n3943 n166 R=2.411e+00 
R3943t3900 n3944 n3901 R=2.387e+01 
R3943t60 n3944 n61 R=1.540e+00 
R3943t1353 n3944 n1354 R=4.403e+01 
R3943t920 n3944 n921 R=2.235e+00 
R3944t661 n3945 n662 R=2.181e+01 
R3944t798 n3945 n799 R=4.225e+00 
R3945t3530 n3946 n3531 R=1.058e+01 
R3945t3051 n3946 n3052 R=7.771e+00 
R3945t2639 n3946 n2640 R=1.142e+01 
R3946t2895 n3947 n2896 R=3.210e+00 
R3946t826 n3947 n827 R=6.259e+00 
R3947t2154 n3948 n2155 R=4.654e+00 
R3948t2358 n3949 n2359 R=8.397e+00 
R3948t2764 n3949 n2765 R=5.451e+00 
R3949t3191 n3950 n3192 R=5.031e+00 
R3949t2780 n3950 n2781 R=7.847e+00 
R3949t2844 n3950 n2845 R=5.344e+01 
R3950t612 n3951 n613 R=2.669e+00 
R3952t459 n3953 n460 R=9.412e+02 
R3952t2701 n3953 n2702 R=8.081e+00 
R3952t1649 n3953 n1650 R=5.689e+02 
R3952t788 n3953 n789 R=2.109e+00 
R3952t2231 n3953 n2232 R=8.235e+00 
R3953t3652 n3954 n3653 R=5.414e+00 
R3953t3195 n3954 n3196 R=3.862e+00 
R3954t2659 n3955 n2660 R=2.904e+01 
R3954t3653 n3955 n3654 R=1.470e+01 
R3954t1569 n3955 n1570 R=1.611e+01 
R3954t2706 n3955 n2707 R=2.395e+00 
R3955t2228 n3956 n2229 R=1.990e+01 
R3955t1111 n3956 n1112 R=2.790e+00 
R3956t1811 n3957 n1812 R=4.577e+02 
R3956t1443 n3957 n1444 R=5.203e+01 
R3957t348 n3958 n349 R=4.355e+00 
R3958t132 n3959 n133 R=2.762e+00 
R3959t1328 n3960 n1329 R=6.641e+00 
R3959t2022 n3960 n2023 R=6.251e+00 
R3959t3105 n3960 n3106 R=1.926e+01 
R3959t3641 n3960 n3642 R=3.659e+00 
R3960t198 n3961 n199 R=2.615e+00 
R3961t2268 n3962 n2269 R=9.040e+00 
R3962t965 n3963 n966 R=1.713e+00 
R3963t1454 n3964 n1455 R=9.947e+02 
R3963t1067 n3964 n1068 R=5.432e+00 
R3963t396 n3964 n397 R=6.552e+00 
R3963t293 n3964 n294 R=2.842e+00 
R3964t705 n3965 n706 R=1.950e+02 
R3964t2216 n3965 n2217 R=6.374e+00 
R3965t1130 n3966 n1131 R=5.469e+00 
R3965t2338 n3966 n2339 R=1.084e+01 
R3965t3307 n3966 n3308 R=3.178e+00 
R3965t863 n3966 n864 R=6.773e+00 
R3966t1354 n3967 n1355 R=4.460e+00 
R3966t1420 n3967 n1421 R=3.619e+00 
R3966t1244 n3967 n1245 R=8.747e+01 
R3967t2162 n3968 n2163 R=1.087e+01 
R3967t2160 n3968 n2161 R=3.997e+00 
R3967t3275 n3968 n3276 R=2.691e+01 
R3967t2088 n3968 n2089 R=1.130e+01 
R3969t900 n3970 n901 R=6.946e+00 
R3969t3599 n3970 n3600 R=7.047e+01 
R3970t3274 n3971 n3275 R=7.821e+00 
R3971t720 n3972 n721 R=2.070e+00 
R3971t1549 n3972 n1550 R=4.352e+01 
R3971t567 n3972 n568 R=3.504e+01 
R3971t2957 n3972 n2958 R=7.114e+00 
R3972t2156 n3973 n2157 R=5.825e+00 
R3972t255 n3973 n256 R=5.109e+01 
R3972t2608 n3973 n2609 R=3.786e+00 
R3973t1477 n3974 n1478 R=4.264e+00 
R3973t1001 n3974 n1002 R=2.442e+02 
R3973t3425 n3974 n3426 R=2.008e+01 
R3974t2815 n3975 n2816 R=2.883e+01 
R3975t3915 n3976 n3916 R=1.686e+01 
R3975t31 n3976 n32 R=1.782e+01 
R3975t2613 n3976 n2614 R=2.339e+00 
R3975t3846 n3976 n3847 R=2.720e+01 
R3976t512 n3977 n513 R=4.247e+00 
R3977t538 n3978 n539 R=2.434e+01 
R3978t49 n3979 n50 R=3.186e+01 
R3978t443 n3979 n444 R=1.649e+00 
R3979t1020 n3980 n1021 R=1.808e+01 
R3979t3235 n3980 n3236 R=8.781e+01 
R3980t3175 n3981 n3176 R=9.398e+00 
R3980t1602 n3981 n1603 R=3.550e+00 
R3981t517 n3982 n518 R=4.650e+00 
R3982t3749 n3983 n3750 R=4.455e+00 
R3983t2544 n3984 n2545 R=7.150e+00 
R3983t2781 n3984 n2782 R=6.127e+00 
R3983t1626 n3984 n1627 R=5.396e+01 
R3983t1708 n3984 n1 R=1.312e+01 
R3984t489 n3985 n490 R=1.703e+01 
R3984t2524 n3985 n2525 R=4.933e+01 
R3984t109 n3985 n110 R=3.785e+01 
R3984t3783 n3985 n3784 R=4.461e+00 
R3984t92 n3985 n93 R=1.906e+01 
R3985t773 n3986 n774 R=3.714e+00 
R3985t961 n3986 n962 R=7.551e+00 
R3985t732 n3986 n733 R=6.125e+00 
R3986t140 n3987 n141 R=6.550e+00 
R3987t1761 n3988 n1762 R=1.434e+01 
R3988t2309 n3989 n2310 R=5.805e+00 
R3988t3313 n3989 n3314 R=1.256e+01 
R3988t2032 n3989 n2033 R=4.133e+00 
R3989t3236 n3990 n3237 R=6.395e+00 
R3990t629 n3991 n630 R=1.118e+03 
R3990t1630 n3991 n1631 R=4.725e+00 
R3991t1653 n3992 n1654 R=2.583e+02 
R3991t2537 n3992 n2538 R=6.358e+00 
R3991t2877 n3992 n2878 R=7.837e+00 
R3991t3068 n3992 n3069 R=2.061e+01 
R3991t712 n3992 n713 R=4.968e+01 
R3992t276 n3993 n277 R=6.193e+00 
R3992t1733 n3993 n1734 R=2.918e+01 
R3993t2930 n3994 n2931 R=1.649e+01 
R3993t3423 n3994 n3424 R=4.459e+00 
R3993t3573 n3994 n3574 R=4.733e+00 
R3994t1029 n3995 n1030 R=6.541e+01 
R3994t803 n3995 n804 R=2.947e+00 
R3994t858 n3995 n859 R=1.277e+01 
R3995t3228 n3996 n3229 R=4.455e+01 
R3995t2783 n3996 n2784 R=9.304e+00 
R3997t95 n3998 n96 R=1.228e+01 
R3997t699 n3998 n700 R=5.821e+00 
R3997t2160 n3998 n2161 R=9.690e+00 
R3997t3275 n3998 n3276 R=4.105e+01 
R3998t2802 n3999 n2803 R=7.132e+00 
R3999t2989 n4000 n2990 R=3.819e+00 
R4000t187 n4001 n188 R=3.072e+00 
R4000t2590 n4001 n2591 R=3.237e+00 
R4000t3382 n4001 n3383 R=6.085e+00 
R4001t3453 n4002 n3454 R=3.168e+00 
R4001t726 n4002 n727 R=1.074e+01 
R4001t2825 n4002 n2826 R=9.604e+01 
R4002t2789 n4003 n2790 R=1.731e+01 
R4003t344 n4004 n345 R=3.247e+00 
R4003t176 n4004 n177 R=3.501e+00 
R4004t68 n4005 n69 R=5.003e+00 
R4004t2554 n4005 n2555 R=5.222e+00 
R4004t3493 n4005 n3494 R=9.452e+00 
R4005t2784 n4006 n2785 R=4.945e+00 
R4006t765 n4007 n766 R=4.459e+00 
R4007t87 n4008 n88 R=2.626e+00 
R4007t411 n4008 n412 R=2.021e+01 
R4007t566 n4008 n567 R=4.390e+00 
R4007t3820 n4008 n3821 R=7.051e+00 
R4008t1765 n4009 n1766 R=2.865e+00 
R4008t3843 n4009 n3844 R=6.967e+00 
R4008t1842 n4009 n1843 R=1.220e+01 
R4009t2043 n4010 n2044 R=4.942e+00 
R4009t1270 n4010 n1271 R=2.054e+02 
R4009t268 n4010 n269 R=3.091e+00 
R4010t693 n4011 n694 R=2.567e+00 
R4010t1143 n4011 n1144 R=4.164e+00 
R4010t1023 n4011 n1024 R=1.797e+01 
R4011t1676 n4012 n1677 R=6.295e+00 
R4011t2062 n4012 n2063 R=2.902e+00 
R4011t1252 n4012 n1253 R=1.406e+02 
R4014t874 n4015 n875 R=1.635e+01 
R4015t1077 n4016 n1078 R=2.069e+01 
R4015t3899 n4016 n3900 R=5.097e+00 
R4015t1393 n4016 n1394 R=3.481e+00 
R4015t3508 n4016 n3509 R=6.814e+00 
R4015t1830 n4016 n1831 R=5.219e+00 
R4016t2936 n4017 n2937 R=7.002e+00 
R4016t1873 n4017 n1874 R=4.195e+00 
R4016t1256 n4017 n1257 R=2.233e+01 
R4017t405 n4018 n406 R=8.061e+00 
R4018t3477 n4019 n3478 R=3.712e+00 
R4018t2728 n4019 n2729 R=3.022e+00 
R4019t3755 n4020 n3756 R=7.207e+01 
R4019t696 n4020 n697 R=6.165e+00 
R4019t1414 n4020 n1415 R=3.815e+00 
R4020t2634 n4021 n2635 R=1.894e+01 
R4020t2643 n4021 n2644 R=4.771e+00 
R4020t1186 n4021 n1187 R=1.645e+01 
R4021t402 n4022 n403 R=1.657e+01 
R4021t1439 n4022 n1440 R=1.691e+01 
R4021t1445 n4022 n1446 R=2.047e+01 
R4022t1247 n4023 n1248 R=1.510e+01 
R4022t1304 n4023 n1305 R=6.546e+00 
R4023t1331 n4024 n1332 R=3.160e+01 
R4023t1579 n4024 n1580 R=1.649e+01 
R4026t2776 n4027 n2777 R=7.837e+00 
R4026t1312 n4027 n1313 R=4.981e+00 
R4027t1564 n4028 n1565 R=4.946e+00 
R4028t3228 n4029 n3229 R=7.494e+00 
R4028t3676 n4029 n3677 R=3.921e+01 
R4028t2150 n4029 n2151 R=7.413e+01 
R4028t1198 n4029 n1199 R=4.813e+00 
R4029t1344 n4030 n1345 R=1.707e+02 
R4029t1825 n4030 n1826 R=2.302e+01 
R4029t3345 n4030 n3346 R=3.254e+00 
R4029t461 n4030 n462 R=2.578e+01 
R4029t1483 n4030 n1484 R=1.345e+01 
R4029t2834 n4030 n2835 R=4.772e+00 
R4030t3343 n4031 n3344 R=4.034e+00 
R4031t2457 n4032 n2458 R=5.000e+01 
R4031t2150 n4032 n2151 R=6.507e+00 
R4032t1912 n4033 n1913 R=8.213e+00 
R4033t155 n4034 n156 R=3.629e+01 
R4033t2796 n4034 n2797 R=3.892e+01 
R4033t3665 n4034 n3666 R=1.936e+01 
R4034t1827 n4035 n1828 R=2.274e+01 
R4034t2306 n4035 n2307 R=1.494e+01 
R4034t1419 n4035 n1420 R=1.407e+01 
R4035t3040 n4036 n3041 R=3.878e+00 
R4035t1004 n4036 n1005 R=9.986e+00 
R4035t1306 n4036 n1307 R=6.839e+00 
R4036t3024 n4037 n3025 R=1.145e+01 
R4036t829 n4037 n830 R=5.322e+00 
R4037t978 n4038 n979 R=4.090e+00 
R4038t807 n4039 n808 R=3.844e+01 
R4038t753 n4039 n754 R=3.893e+00 
R4038t1565 n4039 n1566 R=7.633e+00 
R4038t3323 n4039 n3324 R=2.817e+00 
R4040t1000 n4041 n1001 R=1.279e+01 
R4040t3601 n4041 n3602 R=3.352e+01 
R4041t1318 n4042 n1319 R=2.181e+00 
R4041t1621 n4042 n1622 R=9.938e+01 
R4042t3476 n4043 n3477 R=4.913e+00 
R4042t2734 n4043 n2735 R=8.277e+01 
R4043t3454 n4044 n3455 R=1.336e+01 
R4044t498 n4045 n499 R=1.298e+01 
R4044t3986 n4045 n3987 R=4.618e+00 
R4045t3352 n4046 n3353 R=3.027e+00 
R4046t1078 n4047 n1079 R=3.213e+00 
R4046t3095 n4047 n3096 R=1.112e+01 
R4046t1685 n4047 n1686 R=1.400e+01 
R4048t1957 n4049 n1958 R=2.410e+00 
R4048t3059 n4049 n3060 R=2.969e+01 
R4048t962 n4049 n963 R=4.890e+00 
R4049t717 n4050 n718 R=3.965e+00 
R4050t2024 n4051 n2025 R=4.466e+00 
R4050t954 n4051 n955 R=9.812e+00 
R4051t1281 n4052 n1282 R=2.478e+00 
R4051t738 n4052 n739 R=3.326e+01 
R4051t3049 n4052 n3050 R=4.087e+01 
R4052t2814 n4053 n2815 R=2.267e+01 
R4052t3340 n4053 n3341 R=1.222e+01 
R4052t3194 n4053 n3195 R=6.674e+00 
R4052t1123 n4053 n1124 R=2.116e+00 
R4052t3605 n4053 n3606 R=6.753e+00 
R4053t958 n4054 n959 R=4.826e+00 
R4054t44 n4055 n45 R=4.715e+01 
R4054t3352 n4055 n3353 R=1.641e+01 
R4055t816 n4056 n817 R=8.188e+00 
R4055t2381 n4056 n2382 R=3.099e+02 
R4055t607 n4056 n608 R=4.677e+00 
R4057t1456 n4058 n1457 R=2.596e+01 
R4057t3088 n4058 n3089 R=7.263e+00 
R4057t1511 n4058 n1512 R=6.383e+00 
R4058t3823 n4059 n3824 R=1.412e+01 
R4058t2390 n4059 n2391 R=5.611e+01 
R4059t186 n4060 n187 R=6.107e+00 
R4059t990 n4060 n991 R=9.885e+00 
R4059t2071 n4060 n2072 R=1.870e+01 
R4059t2950 n4060 n2951 R=2.265e+02 
R4060t3259 n4061 n3260 R=8.854e+00 
R4060t3052 n4061 n3053 R=7.573e+00 
R4061t1262 n4062 n1263 R=3.143e+01 
R4063t339 n4064 n340 R=2.807e+00 
R4063t1888 n4064 n1889 R=6.969e+00 
R4063t3828 n4064 n3829 R=5.752e+00 
R4064t3411 n4065 n3412 R=1.389e+01 
R4064t808 n4065 n809 R=5.373e+03 
R4065t1207 n4066 n1208 R=2.594e+00 
R4066t486 n4067 n487 R=2.650e+00 
R4066t1465 n4067 n1466 R=1.825e+01 
R4066t1710 n4067 n1711 R=7.926e+01 
R4067t3618 n4068 n3619 R=3.462e+00 
R4067t3608 n4068 n3609 R=1.596e+01 
R4067t1078 n4068 n1079 R=9.892e+00 
R4068t1890 n4069 n1891 R=8.627e+00 
R4068t3411 n4069 n3412 R=7.133e+00 
R4068t4064 n4069 n4065 R=5.207e+00 
R4069t2423 n4070 n2424 R=3.444e+01 
R4070t1411 n4071 n1412 R=4.086e+01 
R4070t3921 n4071 n3922 R=1.562e+01 
R4071t1798 n4072 n1799 R=4.609e+02 
R4071t3380 n4072 n3381 R=5.686e+00 
R4071t799 n4072 n800 R=6.450e+01 
R4072t1495 n4073 n1496 R=1.801e+01 
R4072t1041 n4073 n1042 R=1.031e+01 
R4072t1542 n4073 n1543 R=3.338e+00 
R4073t118 n4074 n119 R=1.088e+02 
R4073t839 n4074 n840 R=1.966e+00 
R4073t1348 n4074 n1349 R=7.153e+00 
R4074t3091 n4075 n3092 R=3.356e+00 
R4075t879 n4076 n880 R=5.818e+00 
R4075t3120 n4076 n3121 R=1.179e+01 
R4076t317 n4077 n318 R=5.095e+01 
R4077t3112 n4078 n3113 R=5.532e+00 
R4077t2424 n4078 n2425 R=1.289e+01 
R4077t549 n4078 n550 R=5.872e+00 
R4078t2809 n4079 n2810 R=4.143e+01 
R4078t3811 n4079 n3812 R=1.144e+01 
R4078t1092 n4079 n1093 R=5.646e+00 
R4078t1331 n4079 n1332 R=4.025e+01 
R4078t4023 n4079 n4024 R=9.128e+00 
R4078t1588 n4079 n1589 R=6.565e+00 
R4079t1076 n4080 n1077 R=4.053e+00 
R4079t2844 n4080 n2845 R=3.323e+00 
R4079t3949 n4080 n3950 R=3.630e+00 
R4080t1842 n4081 n1843 R=5.599e+00 
R4080t1349 n4081 n1350 R=3.959e+00 
R4081t2276 n4082 n2277 R=1.669e+01 
R4081t611 n4082 n612 R=5.833e+00 
R4082t1110 n4083 n1111 R=5.209e+01 
R4082t1648 n4083 n1649 R=1.340e+01 
R4082t1096 n4083 n1097 R=6.605e+00 
R4082t3479 n4083 n3480 R=2.566e+01 
R4083t1958 n4084 n1959 R=4.114e+01 
R4084t596 n4085 n597 R=8.624e+00 
R4084t938 n4085 n939 R=4.178e+01 
R4084t100 n4085 n101 R=4.607e+00 
R4084t1430 n4085 n1431 R=2.941e+00 
R4085t1126 n4086 n1127 R=2.867e+00 
R4085t3027 n4086 n3028 R=4.831e+00 
R4086t1021 n4087 n1022 R=1.099e+01 
R4087t1117 n4088 n1118 R=5.891e+00 
R4088t3677 n4089 n3678 R=1.602e+01 
R4088t2253 n4089 n2254 R=5.405e+01 
R4088t1265 n4089 n1266 R=1.700e+02 
R4088t522 n4089 n523 R=3.425e+00 
R4089t2574 n4090 n2575 R=1.963e+01 
R4090t158 n4091 n159 R=4.906e+00 
R4090t236 n4091 n237 R=6.712e+00 
R4090t1540 n4091 n1541 R=4.750e+01 
R4091t2525 n4092 n2526 R=1.637e+01 
R4091t2860 n4092 n2861 R=4.688e+00 
R4091t2002 n4092 n2003 R=4.477e+00 
R4091t1892 n4092 n1893 R=4.070e+00 
R4092t2591 n4093 n2592 R=9.179e+00 
R4092t2054 n4093 n2055 R=6.278e+00 
R4092t394 n4093 n395 R=4.866e+01 
R4093t1287 n4094 n1288 R=1.905e+01 
R4093t2116 n4094 n2117 R=1.134e+01 
R4093t1317 n4094 n1318 R=1.373e+01 
R4093t892 n4094 n893 R=4.491e+00 
R4094t941 n4095 n942 R=6.303e+00 
R4094t3187 n4095 n3188 R=1.407e+01 
R4094t1025 n4095 n1026 R=5.399e+00 
R4095t2676 n4096 n2677 R=6.701e+00 
R4095t2193 n4096 n2194 R=9.872e+00 
R4096t2938 n4097 n2939 R=4.853e+02 
R4096t1929 n4097 n1930 R=3.221e+00 
R4096t2191 n4097 n2192 R=6.003e+00 
R4096t3973 n4097 n3974 R=3.993e+01 
R4096t1477 n4097 n1478 R=7.741e+00 
R4097t1750 n4098 n1751 R=5.437e+00 
R4097t760 n4098 n761 R=1.434e+01 
R4097t2695 n4098 n2696 R=4.600e+02 
R4097t3233 n4098 n3234 R=5.118e+00 
R4098t425 n4099 n426 R=2.008e+00 
R4099t3450 n4100 n3451 R=4.788e+00 
R4099t307 n4100 n308 R=1.197e+01 
R4100t3623 n4101 n3624 R=4.088e+00 
R4101t2956 n4102 n2957 R=4.696e+00 
R4101t2341 n4102 n2342 R=3.566e+01 
R4102t643 n4103 n644 R=7.034e+00 
R4102t3614 n4103 n3615 R=4.563e+01 
R4102t943 n4103 n944 R=2.358e+01 
R4102t990 n4103 n991 R=8.533e+00 
R4102t4059 n4103 n4060 R=3.080e+00 
R4102t2071 n4103 n2072 R=5.125e+00 
R4103t1270 n4104 n1271 R=6.054e+00 
R4104t2740 n4105 n2741 R=3.172e+00 
R4105t1415 n4106 n1416 R=7.688e+00 
R4105t3519 n4106 n3520 R=4.747e+00 
R4105t204 n4106 n205 R=1.026e+01 
R4106t1351 n4107 n1352 R=5.067e+00 
R4106t3910 n4107 n3911 R=8.533e+00 
R4106t851 n4107 n852 R=5.261e+00 
R4107t2015 n4108 n2016 R=7.192e+00 
R4107t1577 n4108 n1578 R=4.153e+01 
R4107t2560 n4108 n2561 R=3.234e+00 
R4108t459 n4109 n460 R=1.407e+01 
R4108t3602 n4109 n3603 R=7.595e+00 
R4108t793 n4109 n794 R=3.052e+00 
R4108t2036 n4109 n2037 R=2.593e+00 
R4109t468 n4110 n469 R=2.359e+01 
R4109t1132 n4110 n1133 R=2.756e+00 
R4109t1619 n4110 n1620 R=3.438e+01 
R4110t397 n4111 n398 R=2.392e+00 
R4110t2305 n4111 n2306 R=2.821e+01 
R4111t2155 n4112 n2156 R=3.702e+00 
R4111t2440 n4112 n2441 R=4.115e+00 
R4111t3461 n4112 n3462 R=4.139e+00 
R4111t3242 n4112 n3243 R=1.566e+01 
R4112t83 n4113 n84 R=3.936e+00 
R4112t2525 n4113 n2526 R=3.456e+00 
R4112t1288 n4113 n1289 R=5.160e+00 
R4112t2860 n4113 n2861 R=8.858e+00 
R4113t2657 n4114 n2658 R=1.365e+01 
R4113t2545 n4114 n2546 R=3.016e+01 
R4113t219 n4114 n220 R=7.091e+00 
R4114t1144 n4115 n1145 R=2.411e+01 
R4115t3237 n4116 n3238 R=1.297e+01 
R4115t918 n4116 n919 R=1.070e+02 
R4115t336 n4116 n337 R=3.272e+01 
R4116t1440 n4117 n1441 R=4.305e+00 
R4116t1338 n4117 n1339 R=4.785e+01 
R4116t471 n4117 n472 R=7.821e+00 
R4117t1561 n4118 n1562 R=9.292e+00 
R4118t4067 n4119 n4068 R=1.738e+01 
R4119t401 n4120 n402 R=2.589e+02 
R4119t3040 n4120 n3041 R=2.126e+01 
R4119t4035 n4120 n4036 R=1.147e+01 
R4119t1004 n4120 n1005 R=2.887e+00 
R4120t382 n4121 n383 R=1.537e+00 
R4120t3503 n4121 n3504 R=5.223e+00 
R4120t3809 n4121 n3810 R=5.172e+00 
R4121t2819 n4122 n2820 R=4.422e+00 
R4121t1196 n4122 n1197 R=4.807e+00 
R4122t795 n4123 n796 R=4.898e+00 
R4122t1447 n4123 n1448 R=1.216e+01 
R4122t2158 n4123 n2159 R=8.654e+00 
R4123t916 n4124 n917 R=4.670e+00 
R4123t523 n4124 n524 R=1.402e+01 
R4123t2320 n4124 n2321 R=6.037e+00 
R4124t89 n4125 n90 R=4.428e+00 
R4124t154 n4125 n155 R=6.814e+00 
R4124t2100 n4125 n2101 R=4.865e+00 
R4124t1777 n4125 n1778 R=7.190e+00 
R4124t176 n4125 n177 R=4.396e+01 
R4125t1147 n4126 n1148 R=1.149e+02 
R4125t3880 n4126 n3881 R=6.806e+00 
R4126t1605 n4127 n1606 R=6.845e+00 
R4126t334 n4127 n335 R=2.193e+01 
R4126t1166 n4127 n1167 R=1.182e+01 
R4127t583 n4128 n584 R=2.166e+00 
R4127t3785 n4128 n3786 R=9.630e+00 
R4127t82 n4128 n83 R=3.909e+00 
R4127t3150 n4128 n3151 R=2.716e+00 
R4128t1513 n4129 n1514 R=3.259e+00 
R4129t1123 n4130 n1124 R=5.109e+01 
R4129t1566 n4130 n1567 R=1.247e+01 
R4129t925 n4130 n926 R=2.494e+00 
R4129t2372 n4130 n2373 R=3.390e+00 
R4130t383 n4131 n384 R=2.728e+00 
R4130t2532 n4131 n2533 R=6.814e+00 
R4131t4100 n4132 n4101 R=5.365e+00 
R4131t1702 n4132 n1703 R=1.534e+00 
R4132t3742 n4133 n3743 R=9.198e+00 
R4132t2144 n4133 n2145 R=7.827e+00 
R4132t3162 n4133 n3163 R=2.637e+00 
R4133t2681 n4134 n2682 R=2.937e+00 
R4133t3164 n4134 n3165 R=1.940e+02 
R4133t1511 n4134 n1512 R=6.300e+00 
R4133t4057 n4134 n4058 R=8.118e+00 
R4133t3088 n4134 n3089 R=5.281e+00 
R4134t2922 n4135 n2923 R=4.749e+00 
R4134t146 n4135 n147 R=3.869e+01 
R4134t164 n4135 n165 R=7.819e+00 
R4135t1870 n4136 n1871 R=4.578e+00 
R4136t2002 n4137 n2003 R=8.121e+01 
R4136t4091 n4137 n4092 R=1.303e+01 
R4136t1892 n4137 n1893 R=6.494e+01 
R4136t2243 n4137 n2244 R=5.870e+01 
R4136t1485 n4137 n1486 R=3.855e+00 
R4137t921 n4138 n922 R=2.691e+00 
R4137t3087 n4138 n3088 R=2.021e+01 
R4137t1173 n4138 n1174 R=9.672e+00 
R4137t923 n4138 n924 R=2.882e+00 
R4137t3564 n4138 n3565 R=2.072e+01 
R4138t2523 n4139 n2524 R=7.476e+00 
R4138t2418 n4139 n2419 R=9.543e+00 
R4138t102 n4139 n103 R=3.163e+01 
R4138t1466 n4139 n1467 R=5.430e+00 
R4139t2606 n4140 n2607 R=3.329e+00 
R4139t1040 n4140 n1041 R=1.691e+01 
R4140t2318 n4141 n2319 R=3.553e+00 
R4140t1918 n4141 n1919 R=3.363e+00 
R4141t3296 n4142 n3297 R=5.820e+00 
R4141t1734 n4142 n1735 R=2.245e+01 
R4142t536 n4143 n537 R=1.101e+02 
R4142t2724 n4143 n2725 R=6.806e+00 
R4142t2888 n4143 n2889 R=7.480e+00 
R4142t3457 n4143 n3458 R=5.564e+00 
R4143t1247 n4144 n1248 R=4.143e+01 
R4143t3885 n4144 n3886 R=1.334e+02 
R4143t2003 n4144 n2004 R=7.687e+01 
R4143t2969 n4144 n2970 R=4.740e+01 
R4144t410 n4145 n411 R=6.004e+00 
R4144t3581 n4145 n3582 R=9.415e+00 
R4145t1780 n4146 n1781 R=6.667e+00 
R4146t3294 n4147 n3295 R=2.449e+01 
R4146t2044 n4147 n2045 R=5.849e+00 
R4146t1521 n4147 n1522 R=7.111e+00 
R4147t1076 n4148 n1077 R=4.851e+01 
R4147t2575 n4148 n2576 R=8.782e+00 
R4147t3903 n4148 n3904 R=6.272e+00 
R4147t1837 n4148 n1838 R=8.947e+00 
R4147t3949 n4148 n3950 R=1.201e+01 
R4147t4079 n4148 n4080 R=1.744e+01 
R4148t312 n4149 n313 R=5.704e+00 
R4148t3477 n4149 n3478 R=9.420e+00 
R4148t467 n4149 n468 R=1.333e+01 
R4148t3856 n4149 n3857 R=5.608e+00 
R4148t2728 n4149 n2729 R=1.216e+02 
R4149t2965 n4150 n2966 R=4.095e+00 
R4149t676 n4150 n677 R=1.319e+01 
R4149t2158 n4150 n2159 R=1.083e+01 
R4150t1619 n4151 n1620 R=1.206e+01 
R4151t237 n4152 n238 R=3.187e+00 
R4152t1654 n4153 n1655 R=7.543e+00 
R4152t109 n4153 n110 R=3.012e+01 
R4153t2682 n4154 n2683 R=7.824e+00 
R4153t3246 n4154 n3247 R=6.824e+00 
R4154t197 n4155 n198 R=1.809e+00 
R4155t1038 n4156 n1039 R=3.222e+00 
R4155t2545 n4156 n2546 R=9.819e+00 
R4155t4113 n4156 n4114 R=2.434e+01 
R4156t1910 n4157 n1911 R=2.321e+00 
R4156t2963 n4157 n2964 R=1.773e+01 
R4156t1455 n4157 n1456 R=8.026e+01 
R4156t1647 n4157 n1648 R=7.662e+00 
R4157t262 n4158 n263 R=1.609e+02 
R4157t2738 n4158 n2739 R=1.428e+01 
R4158t2807 n4159 n2808 R=7.312e+00 
R4158t3213 n4159 n3214 R=3.335e+00 
R4158t3145 n4159 n3146 R=9.613e+01 
R4158t3502 n4159 n3503 R=2.540e+00 
R4158t1510 n4159 n1511 R=1.671e+01 
R4159t390 n4160 n391 R=1.354e+01 
R4159t418 n4160 n419 R=1.775e+01 
R4159t3805 n4160 n3806 R=1.514e+01 
R4160t3290 n4161 n3291 R=1.769e+01 
R4160t4044 n4161 n4045 R=5.334e+00 
R4161t2048 n4162 n2049 R=6.016e+00 
R4161t2579 n4162 n2580 R=2.335e+00 
R4161t526 n4162 n527 R=1.235e+01 
R4162t3442 n4163 n3443 R=5.678e+00 
R4162t2047 n4163 n2048 R=8.366e+00 
R4162t1812 n4163 n1813 R=1.996e+01 
R4162t3634 n4163 n3635 R=9.825e+00 
R4163t103 n4164 n104 R=1.531e+01 
R4164t2624 n4165 n2625 R=2.770e+01 
R4164t3047 n4165 n3048 R=1.024e+01 
R4164t2255 n4165 n2256 R=6.005e+00 
R4165t2505 n4166 n2506 R=1.056e+02 
R4165t3258 n4166 n3259 R=2.482e+00 
R4165t1172 n4166 n1173 R=6.388e+00 
R4165t2375 n4166 n2376 R=7.087e+00 
R4166t2553 n4167 n2554 R=4.452e+00 
R4166t132 n4167 n133 R=1.504e+01 
R4166t1249 n4167 n1250 R=6.993e+01 
R4167t344 n4168 n345 R=2.850e+00 
R4167t756 n4168 n757 R=9.288e+00 
R4167t4003 n4168 n4004 R=7.853e+00 
R4168t2569 n4169 n2570 R=4.508e+00 
R4168t354 n4169 n355 R=9.007e+00 
R4169t1870 n4170 n1871 R=4.127e+01 
R4169t3693 n4170 n3694 R=2.372e+00 
R4170t3874 n4171 n3875 R=9.205e+00 
R4170t1925 n4171 n1926 R=6.475e+00 
R4170t3844 n4171 n3845 R=1.388e+01 
R4170t3030 n4171 n3031 R=9.412e+00 
R4171t2069 n4172 n2070 R=3.712e+00 
R4171t2137 n4172 n2138 R=9.369e+00 
R4172t363 n4173 n364 R=2.961e+01 
R4173t2464 n4174 n2465 R=3.890e+00 
R4173t2660 n4174 n2661 R=2.061e+01 
R4173t3602 n4174 n3603 R=1.113e+01 
R4174t3886 n4175 n3887 R=2.532e+00 
R4174t3758 n4175 n3759 R=1.839e+01 
R4174t3608 n4175 n3609 R=8.427e+00 
R4174t3618 n4175 n3619 R=6.816e+00 
R4175t1509 n4176 n1510 R=5.851e+00 
R4175t1417 n4176 n1418 R=3.856e+00 
R4176t3155 n4177 n3156 R=2.278e+00 
R4176t1262 n4177 n1263 R=1.187e+01 
R4176t3410 n4177 n3411 R=2.396e+01 
R4176t2867 n4177 n2868 R=4.911e+01 
R4177t397 n4178 n398 R=2.386e+00 
R4177t2728 n4178 n2729 R=4.528e+00 
R4177t2305 n4178 n2306 R=4.151e+01 
R4178t4127 n4179 n4128 R=1.887e+02 
R4178t583 n4179 n584 R=4.367e+00 
R4178t857 n4179 n858 R=1.598e+01 
R4178t1231 n4179 n1232 R=2.465e+01 
R4178t2864 n4179 n2865 R=1.189e+02 
R4179t854 n4180 n855 R=1.030e+01 
R4179t2543 n4180 n2544 R=3.920e+00 
R4180t544 n4181 n545 R=9.357e+00 
R4180t1953 n4181 n1954 R=5.674e+00 
R4181t2210 n4182 n2211 R=8.847e+00 
R4181t502 n4182 n503 R=1.066e+01 
R4181t1729 n4182 n1730 R=8.644e+00 
R4182t3350 n4183 n3351 R=9.029e+00 
R4183t832 n4184 n833 R=7.108e+02 
R4183t2509 n4184 n2510 R=8.301e+00 
R4183t3503 n4184 n3504 R=5.456e+00 
R4183t1586 n4184 n1587 R=2.851e+00 
R4184t1897 n4185 n1898 R=1.876e+01 
R4184t416 n4185 n417 R=1.756e+01 
R4184t3546 n4185 n3547 R=2.414e+00 
R4185t3883 n4186 n3884 R=2.516e+00 
R4186t1956 n4187 n1957 R=1.003e+01 
R4186t3994 n4187 n3995 R=4.866e+01 
R4187t1125 n4188 n1126 R=4.367e+00 
R4187t2316 n4188 n2317 R=5.379e+00 
R4187t2814 n4188 n2815 R=1.114e+01 
R4188t3314 n4189 n3315 R=1.502e+01 
R4189t3156 n1 n3157 R=1.027e+01 
R4189t3435 n1 n3436 R=8.775e+00 
R4189t3232 n1 n3233 R=2.534e+01 
R4190t115 n4191 n116 R=3.541e+00 
R4190t24 n4191 n25 R=3.190e+02 
R4191t2456 n4192 n2457 R=4.061e+00 
R4191t4105 n4192 n4106 R=2.198e+01 
R4191t4185 n4192 n4186 R=3.759e+00 
R4192t613 n4193 n614 R=4.479e+00 
R4192t2389 n4193 n2390 R=1.430e+01 
R4192t247 n4193 n248 R=2.978e+00 
R4192t869 n4193 n870 R=5.291e+01 
R4193t2146 n4194 n2147 R=3.194e+01 
R4193t2218 n4194 n2219 R=1.837e+01 
R4193t2471 n4194 n2472 R=5.835e+00 
R4194t3233 n4195 n3234 R=2.078e+01 
R4194t1441 n4195 n1442 R=5.966e+00 
R4195t1178 n4196 n1179 R=3.880e+01 
R4195t1227 n4196 n1228 R=5.705e+00 
R4196t527 n4197 n528 R=2.218e+00 
R4196t4062 n4197 n4063 R=8.765e+00 
R4197t107 n4198 n108 R=3.112e+01 
R4197t1199 n4198 n1200 R=2.878e+00 
R4197t2812 n4198 n2813 R=1.867e+01 
R4197t4169 n4198 n4170 R=9.246e+00 
R4197t3693 n4198 n3694 R=3.405e+01 
R4198t3116 n4199 n3117 R=3.610e+01 
R4198t3460 n4199 n3461 R=1.702e+01 
R4198t2720 n4199 n2721 R=4.589e+00 
R4199t2224 n4200 n2225 R=3.368e+00 
R4200t336 n4201 n337 R=7.509e+00 
R4200t4115 n4201 n4116 R=5.968e+00 
R4200t918 n4201 n919 R=7.477e+00 
R4200t2127 n4201 n2128 R=3.124e+00 
R4201t32 n4202 n33 R=2.658e+00 
R4201t3868 n4202 n3869 R=3.125e+01 
R4202t3039 n4203 n1 R=1.115e+01 
R4202t1037 n4203 n1038 R=1.822e+01 
R4202t2980 n4203 n2981 R=7.445e+02 
R4202t1500 n4203 n1501 R=5.531e+00 
R4203t2978 n4204 n2979 R=9.519e+00 
R4204t217 n4205 n218 R=4.758e+02 
R4204t933 n4205 n934 R=7.287e+00 
R4204t1442 n4205 n1443 R=2.729e+01 
R4205t363 n4206 n364 R=5.585e+01 
R4206t2632 n4207 n2633 R=3.592e+00 
R4207t453 n4208 n454 R=2.566e+00 
R4207t1908 n4208 n1909 R=4.340e+01 
R4208t4043 n4209 n4044 R=3.140e+00 
R4208t3454 n4209 n3455 R=9.386e+00 
R4209t593 n4210 n594 R=1.627e+01 
R4209t1321 n4210 n1322 R=7.022e+00 
R4210t1082 n4211 n1083 R=3.290e+00 
R4210t2486 n4211 n2487 R=4.666e+00 
R4210t2280 n4211 n2281 R=2.652e+01 
R4211t1522 n4212 n1523 R=8.396e+00 
R4211t1754 n4212 n1755 R=4.594e+00 
R4211t2031 n4212 n2032 R=9.529e+00 
R4212t3269 n4213 n3270 R=3.240e+00 
R4213t3525 n4214 n3526 R=3.667e+01 
R4213t2271 n4214 n2272 R=4.887e+00 
R4214t3709 n4215 n3710 R=3.404e+00 
R4215t888 n4216 n889 R=9.215e+00 
R4215t3321 n4216 n3322 R=6.767e+00 
R4216t3941 n4217 n3942 R=2.194e+02 
R4216t562 n4217 n563 R=8.110e+00 
R4216t3403 n4217 n3404 R=8.447e+00 
R4217t779 n4218 n780 R=5.322e+00 
R4217t2454 n4218 n2455 R=4.528e+00 
R4218t4081 n4219 n4082 R=8.349e+00 
R4218t611 n4219 n612 R=8.499e+00 
R4218t1389 n4219 n1390 R=4.301e+00 
R4219t2902 n4220 n2903 R=1.013e+01 
R4220t1652 n4221 n1653 R=3.725e+00 
R4220t3674 n4221 n3675 R=3.462e+02 
R4221t3755 n4222 n3756 R=8.861e+00 
R4221t3558 n4222 n3559 R=5.048e+00 
R4221t170 n4222 n171 R=1.792e+01 
R4221t2227 n4222 n2228 R=2.564e+01 
R4221t33 n4222 n34 R=1.277e+03 
R4222t3281 n4223 n3282 R=3.011e+00 
R4223t903 n4224 n904 R=1.533e+05 
R4223t2552 n4224 n2553 R=2.491e+00 
R4224t1136 n4225 n1137 R=4.110e+00 
R4224t2476 n4225 n2477 R=6.090e+00 
R4225t205 n4226 n206 R=2.245e+00 
R4226t442 n4227 n443 R=3.114e+01 
R4226t2793 n4227 n2794 R=1.232e+00 
R4227t1403 n4228 n1404 R=3.300e+00 
R4227t1400 n4228 n1401 R=5.884e+00 
R4227t1583 n4228 n1584 R=4.680e+01 
R4228t1863 n4229 n1864 R=1.253e+01 
R4228t2010 n4229 n2011 R=2.192e+00 
R4228t2097 n4229 n2098 R=1.564e+00 
R4229t1436 n4230 n1437 R=2.325e+02 
R4229t3031 n4230 n3032 R=1.005e+01 
R4230t1717 n4231 n1718 R=7.682e+00 
R4230t4207 n4231 n4208 R=4.594e+01 
R4230t1319 n4231 n1320 R=6.980e+00 
R4231t1307 n4232 n1308 R=2.950e+00 
R4232t478 n4233 n479 R=2.648e+02 
R4233t3182 n4234 n3183 R=8.868e+00 
R4233t248 n4234 n249 R=9.909e+00 
R4234t1617 n4235 n1618 R=2.282e+01 
R4234t2661 n4235 n2662 R=8.145e+00 
R4235t3590 n4236 n3591 R=2.274e+01 
R4235t2406 n4236 n2407 R=2.188e+00 
R4235t773 n4236 n774 R=4.081e+01 
R4236t3684 n4237 n3685 R=1.352e+01 
R4236t260 n4237 n261 R=3.727e+00 
R4236t4193 n4237 n4194 R=3.031e+01 
R4237t2670 n4238 n2671 R=9.320e+00 
R4237t957 n4238 n958 R=4.036e+00 
R4237t3264 n4238 n3265 R=1.509e+01 
R4237t2211 n4238 n2212 R=4.219e+00 
R4238t3760 n4239 n3761 R=2.561e+01 
R4238t1600 n4239 n1601 R=6.891e+00 
R4239t3781 n4240 n3782 R=2.111e+01 
R4239t835 n4240 n836 R=4.136e+03 
R4240t2328 n4241 n2329 R=1.109e+01 
R4240t1149 n4241 n1150 R=1.949e+01 
R4240t807 n4241 n808 R=6.417e+00 
R4240t1899 n4241 n1900 R=1.377e+01 
R4241t3710 n4242 n3711 R=7.177e+01 
R4241t3692 n4242 n3693 R=9.477e+01 
R4241t1613 n4242 n1614 R=2.235e+00 
R4243t2772 n4244 n2773 R=8.196e+00 
R4244t2766 n4245 n2767 R=4.456e+00 
R4244t3251 n4245 n3252 R=5.721e+01 
R4244t3390 n4245 n3391 R=2.679e+00 
R4245t751 n4246 n752 R=7.514e+00 
R4245t2691 n4246 n2692 R=3.895e+00 
R4246t3154 n4247 n3155 R=3.704e+00 
R4246t1704 n4247 n1705 R=4.364e+00 
R4247t2882 n4248 n2883 R=2.287e+01 
R4247t1188 n4248 n1189 R=4.825e+00 
R4247t178 n4248 n179 R=1.297e+01 
R4248t1431 n4249 n1432 R=4.616e+01 
R4248t3300 n4249 n3301 R=2.971e+00 
R4248t1353 n4249 n1354 R=3.348e+01 
R4248t1318 n4249 n1319 R=2.857e+01 
R4248t4041 n4249 n4042 R=8.399e+00 
R4249t1261 n4250 n1262 R=1.356e+01 
R4249t3302 n4250 n3303 R=3.827e+00 
R4250t3253 n4251 n3254 R=1.027e+01 
R4250t3441 n4251 n3442 R=4.412e+00 
R4250t3127 n4251 n3128 R=4.364e+00 
R4251t2212 n4252 n2213 R=1.423e+01 
R4251t2566 n4252 n2567 R=3.514e+02 
R4251t2795 n4252 n2796 R=7.811e+00 
R4252t1504 n4253 n1505 R=1.152e+01 
R4252t197 n4253 n198 R=1.868e+02 
R4252t4154 n4253 n4155 R=1.455e+01 
R4253t3032 n4254 n3033 R=9.095e+00 
R4253t3414 n4254 n3415 R=5.508e+00 
R4254t1371 n4255 n1372 R=9.909e+00 
R4254t2761 n4255 n2762 R=1.143e+01 
R4255t1793 n4256 n1794 R=4.305e+02 
R4256t96 n4257 n97 R=2.826e+01 
R4256t1599 n4257 n1600 R=6.287e+00 
R4256t2792 n4257 n2793 R=3.312e+01 
R4256t1763 n4257 n1764 R=8.594e+00 
R4257t1603 n4258 n1604 R=1.154e+01 
R4257t1758 n4258 n1759 R=3.646e+01 
R4257t1079 n4258 n1080 R=2.114e+01 
R4257t696 n4258 n697 R=1.024e+01 
R4258t95 n4259 n96 R=5.347e+00 
R4258t2160 n4259 n2161 R=3.892e+00 
R4258t2703 n4259 n2704 R=3.763e+00 
R4259t1614 n4260 n1615 R=6.369e+00 
R4260t3330 n4261 n3331 R=7.232e+01 
R4260t268 n4261 n269 R=1.266e+01 
R4260t1270 n4261 n1271 R=3.014e+00 
R4260t899 n4261 n900 R=3.484e+00 
R4261t2268 n4262 n2269 R=2.959e+01 
R4261t3961 n4262 n3962 R=3.729e+00 
R4261t3486 n4262 n3487 R=6.201e+00 
R4262t587 n4263 n588 R=2.495e+00 
R4262t100 n4263 n101 R=1.063e+01 
R4263t146 n4264 n147 R=4.614e+00 
R4263t4134 n4264 n4135 R=3.680e+00 
R4263t164 n4264 n165 R=1.537e+01 
R4264t1661 n4265 n1662 R=7.106e+01 
R4264t2513 n4265 n2514 R=4.701e+00 
R4264t438 n4265 n439 R=3.549e+00 
R4264t549 n4265 n550 R=7.271e+00 
R4265t1980 n4266 n1981 R=1.538e+01 
R4265t1716 n4266 n1717 R=5.750e+00 
R4265t3920 n4266 n3921 R=2.796e+01 
R4267t936 n4268 n937 R=7.031e+00 
R4267t1987 n4268 n1988 R=2.506e+01 
R4268t3445 n4269 n3446 R=2.341e+01 
R4269t1459 n4270 n1460 R=4.596e+00 
R4269t3766 n4270 n3767 R=4.334e+00 
R4270t282 n4271 n283 R=1.510e+01 
R4270t1050 n4271 n1051 R=4.016e+00 
R4271t1886 n4272 n1887 R=2.014e+01 
R4271t4195 n4272 n4196 R=5.599e+00 
R4272t3913 n4273 n3914 R=4.661e+00 
R4272t3908 n4273 n3909 R=9.314e+00 
R4272t836 n4273 n837 R=6.265e+01 
R4272t377 n4273 n378 R=2.651e+00 
R4273t3888 n4274 n3889 R=1.562e+01 
R4273t1046 n4274 n1047 R=1.557e+01 
R4275t1216 n4276 n1217 R=1.136e+01 
R4275t955 n4276 n956 R=1.650e+01 
R4275t462 n4276 n463 R=4.795e+00 
R4276t2629 n4277 n2630 R=2.905e+01 
R4276t3901 n4277 n3902 R=5.281e+01 
R4277t1109 n4278 n1110 R=8.789e+00 
R4278t963 n4279 n964 R=6.233e+00 
R4278t1106 n4279 n1107 R=5.835e+00 
R4279t2380 n4280 n2381 R=1.863e+01 
R4280t3203 n4281 n3204 R=3.688e+01 
R4280t3909 n4281 n3910 R=2.631e+00 
R4280t3385 n4281 n3386 R=5.164e+01 
R4280t1923 n4281 n1924 R=5.892e+00 
R4280t885 n4281 n886 R=6.090e+00 
R4281t553 n4282 n554 R=7.201e+00 
R4282t3921 n4283 n3922 R=3.254e+00 
R4282t1411 n4283 n1412 R=6.036e+00 
R4282t4070 n4283 n4071 R=7.176e+00 
R4283t1505 n4284 n1506 R=9.773e+00 
R4283t4065 n4284 n4066 R=6.063e+00 
R4284t2938 n4285 n2939 R=1.122e+01 
R4284t1477 n4285 n1478 R=7.267e+00 
R4284t4070 n4285 n4071 R=1.469e+01 
R4285t1805 n4286 n1806 R=1.817e+01 
R4285t4 n4286 n5 R=2.352e+00 
R4286t426 n4287 n427 R=4.285e+01 
R4287t1250 n4288 n1251 R=7.443e+00 
R4289t2718 n4290 n2719 R=1.040e+01 
R4290t682 n4291 n683 R=4.478e+00 
R4291t815 n4292 n816 R=1.138e+01 
R4291t2788 n4292 n2789 R=2.249e+01 
R4291t2440 n4292 n2441 R=2.670e+00 
R4291t3461 n4292 n3462 R=1.483e+01 
R4292t3817 n4293 n3818 R=1.575e+02 
R4292t2854 n4293 n2855 R=1.365e+01 
R4293t2602 n4294 n2603 R=3.980e+00 
R4294t2051 n4295 n2052 R=5.297e+00 
R4294t3269 n4295 n3270 R=2.881e+00 
R4294t4212 n4295 n4213 R=3.495e+01 
R4295t1788 n4296 n1789 R=4.314e+01 
R4295t156 n4296 n157 R=5.780e+01 
R4296t2805 n4297 n2806 R=5.296e+00 
R4297t2709 n4298 n2710 R=1.551e+01 
R4297t2777 n4298 n2778 R=3.857e+00 
R4297t2942 n4298 n2943 R=1.648e+01 
R4297t2954 n4298 n2955 R=3.681e+00 
R4298t1881 n4299 n1882 R=1.076e+01 
R4298t3797 n4299 n3798 R=1.151e+01 
R4299t2061 n4300 n2062 R=1.343e+01 
R4299t2821 n4300 n2822 R=2.406e+01 
R4299t446 n4300 n447 R=3.316e+00 
R4300t3018 n4301 n3019 R=1.251e+02 
R4300t956 n4301 n957 R=4.859e+00 
R4301t3202 n4302 n3203 R=1.153e+01 
R4301t1186 n4302 n1187 R=7.255e+00 
R4302t1310 n4303 n1311 R=5.381e+00 
R4302t1518 n4303 n1519 R=5.507e+00 
R4302t1465 n4303 n1466 R=1.725e+00 
R4303t2467 n4304 n2468 R=9.110e+01 
R4303t3713 n4304 n3714 R=1.157e+01 
R4303t2599 n4304 n2600 R=6.121e+00 
R4303t2041 n4304 n2042 R=9.227e+00 
R4304t3624 n4305 n3625 R=1.316e+01 
R4304t2624 n4305 n2625 R=3.832e+00 
R4305t2558 n4306 n2559 R=1.255e+01 
R4305t1927 n4306 n1928 R=5.159e+00 
R4305t3658 n4306 n3659 R=5.057e+00 
R4306t1068 n4307 n1069 R=5.072e+00 
R4306t2999 n4307 n3000 R=5.785e+00 
R4306t2556 n4307 n2557 R=3.240e+00 
R4307t545 n4308 n546 R=2.912e+00 
R4307t3498 n4308 n3499 R=1.137e+01 
R4307t697 n4308 n698 R=3.342e+01 
R4307t1986 n4308 n1987 R=3.379e+00 
R4308t3821 n4309 n3822 R=1.774e+03 
R4308t61 n4309 n62 R=1.327e+01 
R4308t3291 n4309 n3292 R=2.766e+00 
R4309t2115 n4310 n2116 R=5.334e+00 
R4310t898 n4311 n899 R=5.412e+01 
R4310t2053 n4311 n2054 R=4.449e+00 
R4311t780 n4312 n781 R=6.024e+00 
R4311t2924 n4312 n2925 R=2.393e+01 
R4312t578 n4313 n579 R=6.640e+01 
R4312t1879 n4313 n1880 R=2.486e+01 
R4312t1781 n4313 n1782 R=3.039e+00 
R4313t2909 n4314 n2910 R=6.410e+00 
R4313t3868 n4314 n3869 R=6.763e+01 
R4314t3717 n4315 n3718 R=2.788e+01 
R4314t279 n4315 n280 R=7.050e+00 
R4314t3553 n4315 n3554 R=4.498e+00 
R4314t1526 n4315 n1527 R=4.963e+01 
R4314t120 n4315 n121 R=2.764e+00 
R4315t561 n4316 n562 R=3.041e+01 
R4315t931 n4316 n932 R=2.830e+00 
R4315t3299 n4316 n3300 R=3.568e+00 
R4316t790 n4317 n791 R=1.680e+01 
R4316t1434 n4317 n1435 R=2.921e+00 
R4317t3507 n4318 n3508 R=9.478e+02 
R4317t538 n4318 n539 R=3.199e+00 
R4317t1143 n4318 n1144 R=3.694e+01 
R4317t1023 n4318 n1024 R=2.457e+02 
R4318t1825 n4319 n1826 R=3.466e+00 
R4318t4029 n4319 n4030 R=2.823e+01 
R4318t1344 n4319 n1345 R=2.315e+00 
R4319t1624 n4320 n1625 R=3.833e+00 
R4320t1580 n4321 n1581 R=4.118e+00 
R4320t2713 n4321 n2714 R=6.889e+00 
R4321t2406 n4322 n2407 R=1.525e+01 
R4321t4235 n4322 n4236 R=8.811e+00 
R4321t3590 n4322 n3591 R=8.807e+01 
R4321t1544 n4322 n1545 R=5.819e+00 
R4321t53 n4322 n54 R=4.265e+00 
R4322t1353 n4323 n1354 R=6.464e+00 
R4322t4248 n4323 n4249 R=2.712e+01 
R4322t1318 n4323 n1319 R=2.418e+00 
R4322t2258 n4323 n2259 R=6.011e+00 
R4322t60 n4323 n61 R=4.689e+00 
R4323t1478 n4324 n1479 R=9.489e+00 
R4323t905 n4324 n906 R=2.435e+00 
R4325t3004 n4326 n3005 R=2.443e+00 
R4325t493 n4326 n494 R=3.188e+02 
R4326t1265 n4327 n1266 R=5.326e+00 
R4326t3724 n4327 n3725 R=4.264e+01 
R4326t1433 n4327 n1434 R=5.426e+00 
R4326t1030 n4327 n1031 R=5.618e+00 
R4326t3799 n4327 n3800 R=4.895e+00 
R4327t898 n4328 n899 R=2.620e+00 
R4327t2053 n4328 n2054 R=1.763e+01 
R4327t4284 n4328 n4285 R=1.864e+01 
R4327t2938 n4328 n2939 R=4.152e+01 
R4327t428 n4328 n429 R=3.478e+00 
R4327t656 n4328 n657 R=1.147e+01 
R4328t2270 n4329 n2271 R=2.728e+00 
R4328t519 n4329 n520 R=9.329e+01 
R4329t1941 n4330 n1942 R=3.945e+00 
R4329t1390 n4330 n1391 R=2.087e+01 
R4329t2418 n4330 n2419 R=1.163e+02 
R4329t322 n4330 n323 R=1.594e+01 
R4331t3091 n1 n3092 R=1.729e+01 
R4331t4074 n1 n4075 R=1.671e+01 
R4332t1145 n4333 n1146 R=2.574e+01 
R4332t3797 n4333 n3798 R=4.872e+00 
R4333t3623 n4334 n3624 R=3.054e+00 
R4334t4123 n4335 n4124 R=3.998e+00 
R4334t523 n4335 n524 R=3.687e+01 
R4335t2958 n4336 n2959 R=7.004e+00 
R4336t404 n4337 n405 R=2.065e+01 
R4336t1725 n4337 n1726 R=2.393e+01 
R4336t3867 n4337 n3868 R=5.940e+00 
R4337t4141 n4338 n4142 R=2.103e+01 
R4337t2807 n4338 n2808 R=7.994e+00 
R4338t3455 n1 n3456 R=6.540e+00 
R4339t2512 n4340 n2513 R=1.377e+01 
R4339t1752 n4340 n1753 R=2.500e+00 
R4340t1500 n4341 n1501 R=7.561e+00 
R4340t2442 n4341 n2443 R=2.155e+01 
R4340t4202 n4341 n4203 R=1.464e+01 
R4340t2614 n4341 n2615 R=1.016e+02 
R4340t2214 n4341 n2215 R=3.332e+00 
R4341t781 n4342 n782 R=9.463e+00 
R4342t3446 n4343 n3447 R=2.878e+00 
R4343t3364 n4344 n3365 R=5.176e+00 
R4343t4314 n4344 n4315 R=9.722e+00 
R4344t228 n4345 n229 R=4.480e+00 
R4344t4138 n4345 n4139 R=4.415e+01 
R4344t1466 n4345 n1467 R=1.653e+02 
R4344t2949 n4345 n2950 R=1.767e+01 
R4345t3449 n4346 n3450 R=4.423e+01 
R4345t1949 n4346 n1950 R=2.559e+01 
R4345t3006 n4346 n3007 R=3.641e+01 
R4345t2357 n4346 n2358 R=3.564e+00 
R4346t429 n4347 n430 R=4.961e+01 
R4346t3643 n4347 n3644 R=6.568e+01 
R4346t2279 n4347 n2280 R=4.078e+00 
R4346t3357 n4347 n3358 R=4.704e+00 
R4346t1832 n4347 n1833 R=3.433e+00 
R4347t3157 n4348 n3158 R=4.429e+00 
R4348t1371 n4349 n1372 R=3.712e+01 
R4348t4267 n4349 n4268 R=1.908e+01 
R4348t936 n4349 n937 R=3.113e+01 
R4348t4254 n4349 n4255 R=7.095e+00 
R4349t3946 n4350 n3947 R=2.460e+00 
R4350t1284 n4351 n1285 R=3.921e+00 
R4350t3770 n4351 n3771 R=3.571e+00 
R4350t683 n4351 n684 R=8.203e+00 
R4351t1075 n4352 n1076 R=4.410e+00 
R4351t3297 n4352 n3298 R=4.683e+00 
R4351t3651 n4352 n3652 R=1.088e+01 
R4352t3094 n4353 n3095 R=1.128e+01 
R4352t3853 n4353 n3854 R=3.172e+00 
R4353t982 n4354 n983 R=6.248e+00 
R4353t3364 n4354 n3365 R=3.096e+01 
R4353t4343 n4354 n4344 R=2.637e+00 
R4353t4314 n4354 n4315 R=5.244e+01 
R4353t120 n4354 n121 R=6.219e+00 
R4353t1823 n4354 n1824 R=8.484e+00 
R4354t3077 n4355 n3078 R=1.494e+01 
R4354t3701 n4355 n3702 R=6.229e+00 
R4354t3776 n4355 n3777 R=1.159e+01 
R4354t3695 n4355 n3696 R=1.169e+02 
R4355t4082 n4356 n4083 R=2.557e+01 
R4356t1063 n4357 n1064 R=7.301e+00 
R4357t907 n4358 n908 R=1.940e+00 
R4357t2802 n4358 n2803 R=3.359e+00 
R4358t1377 n4359 n1378 R=5.395e+00 
R4358t2474 n4359 n2475 R=5.990e+01 
R4358t1969 n4359 n1970 R=2.111e+01 
R4359t3646 n4360 n3647 R=3.991e+00 
R4359t903 n4360 n904 R=2.581e+00 
R4359t4223 n4360 n4224 R=1.289e+01 
R4360t2466 n4361 n2467 R=3.338e+00 
R4360t3467 n4361 n3468 R=4.818e+00 
R4360t2190 n4361 n2191 R=5.138e+01 
R4362t2046 n4363 n1 R=9.732e+00 
R4362t1889 n4363 n1 R=9.423e+00 
R4362t3890 n4363 n3891 R=8.458e+00 
R4362t2595 n4363 n2596 R=6.080e+02 
R4363t1145 n4364 n1146 R=1.592e+01 
R4363t1227 n4364 n1228 R=3.330e+00 
R4363t1233 n4364 n1234 R=5.546e+02 
R4363t331 n4364 n332 R=2.360e+01 
R4364t1726 n4365 n1727 R=1.500e+01 
R4365t3161 n4366 n3162 R=3.019e+00 
R4365t3882 n4366 n3883 R=6.308e+00 
R4366t1462 n4367 n1463 R=1.829e+01 
R4367t1377 n4368 n1378 R=5.423e+00 
R4367t4358 n4368 n4359 R=4.699e+00 
R4367t1969 n4368 n1970 R=7.715e+00 
R4367t2619 n4368 n2620 R=3.213e+00 
R4368t1721 n4369 n1722 R=3.357e+00 
R4369t2258 n4370 n2259 R=2.624e+01 
R4369t3846 n4370 n3847 R=5.759e+00 
R4369t3975 n4370 n3976 R=4.189e+00 
R4370t1205 n4371 n1206 R=2.035e+00 
R4370t1833 n4371 n1834 R=3.790e+00 
R4371t1633 n4372 n1634 R=1.243e+01 
R4371t3146 n4372 n3147 R=1.327e+01 
R4371t2868 n4372 n2869 R=3.212e+00 
R4371t2641 n4372 n2642 R=1.646e+01 
R4372t2310 n4373 n2311 R=1.796e+01 
R4372t4246 n4373 n4247 R=4.187e+00 
R4372t3056 n4373 n3057 R=4.425e+00 
R4373t317 n4374 n318 R=8.560e+00 
R4373t4076 n4374 n4077 R=4.473e+00 
R4374t1649 n4375 n1650 R=5.111e+01 
R4374t1958 n4375 n1959 R=6.319e+00 
R4375t2553 n4376 n2554 R=7.916e+00 
R4375t4166 n4376 n4167 R=1.091e+01 
R4375t132 n4376 n133 R=1.730e+01 
R4375t3958 n4376 n3959 R=6.915e+00 
R4375t2594 n4376 n2595 R=1.488e+01 
R4376t1032 n4377 n1033 R=1.427e+01 
R4376t3161 n4377 n3162 R=5.010e+00 
R4376t1988 n4377 n1989 R=1.082e+01 
R4376t4365 n4377 n4366 R=1.909e+01 
R4377t355 n4378 n356 R=3.345e+00 
R4377t1083 n4378 n1084 R=7.387e+00 
R4377t3780 n4378 n3781 R=3.862e+02 
R4377t4265 n4378 n4266 R=4.475e+01 
R4378t813 n4379 n814 R=8.041e+01 
R4378t1902 n4379 n1903 R=4.071e+00 
R4378t617 n4379 n618 R=7.214e+00 
R4378t3421 n4379 n3422 R=6.268e+00 
R4378t1541 n4379 n1542 R=1.510e+01 
R4378t470 n4379 n471 R=7.131e+00 
R4378t999 n4379 n1000 R=3.912e+01 
R4379t551 n4380 n552 R=1.628e+01 
R4379t2596 n4380 n2597 R=1.475e+01 
R4379t605 n4380 n606 R=4.152e+01 
R4380t229 n4381 n230 R=4.086e+00 
R4380t3637 n4381 n3638 R=8.427e+00 
R4380t3100 n4381 n3101 R=8.388e+00 
R4380t3567 n4381 n3568 R=2.299e+00 
R4381t3145 n4382 n3146 R=3.058e+00 
R4381t4158 n4382 n4159 R=7.458e+00 
R4381t3502 n4382 n3503 R=5.080e+00 
R4382t2281 n4383 n2282 R=7.404e+00 
R4382t257 n4383 n258 R=4.173e+00 
R4382t3694 n4383 n3695 R=1.206e+01 
R4383t298 n4384 n299 R=2.729e+00 
R4383t4103 n4384 n4104 R=3.634e+02 
R4383t902 n4384 n903 R=5.380e+00 
R4384t1122 n4385 n1123 R=7.962e+00 
R4386t1973 n4387 n1974 R=4.910e+01 
R4386t50 n4387 n51 R=1.315e+01 
R4386t2257 n4387 n2258 R=4.718e+00 
R4387t2635 n4388 n2636 R=5.696e+00 
R4387t2880 n4388 n2881 R=5.470e+00 
R4388t628 n4389 n629 R=1.051e+02 
R4388t3418 n4389 n3419 R=4.207e+01 
R4388t2412 n4389 n2413 R=1.280e+01 
R4388t256 n4389 n257 R=2.037e+01 
R4388t3393 n4389 n3394 R=4.115e+00 
R4389t4132 n4390 n4133 R=5.781e+00 
R4389t3742 n4390 n3743 R=1.187e+01 
R4390t2737 n4391 n2738 R=2.214e+01 
R4391t2962 n4392 n2963 R=5.163e+00 
R4392t4389 n4393 n4390 R=9.293e+00 
R4392t708 n4393 n709 R=5.487e+00 
R4393t579 n4394 n580 R=6.618e+01 
R4393t414 n4394 n415 R=1.043e+01 
R4394t610 n4395 n611 R=3.368e+00 
R4394t2744 n4395 n2745 R=6.445e+00 
R4394t141 n4395 n142 R=5.505e+01 
R4395t2566 n4396 n2567 R=1.356e+01 
R4395t3610 n4396 n3611 R=1.472e+01 
R4395t1457 n4396 n1458 R=2.034e+02 
R4395t2883 n4396 n2884 R=3.462e+00 
R4396t4308 n4397 n4309 R=5.357e+00 
R4396t61 n4397 n62 R=6.225e+01 
R4397t1232 n4398 n1233 R=2.198e+01 
R4397t333 n4398 n334 R=5.309e+00 
R4398t1502 n4399 n1503 R=7.633e+00 
R4398t78 n4399 n79 R=7.707e+00 
R4398t256 n4399 n257 R=1.767e+02 
R4399t1293 n4400 n1294 R=1.353e+01 
R4399t472 n4400 n473 R=4.306e+00 
R4399t988 n4400 n989 R=9.729e+00 
R4399t1335 n4400 n1336 R=4.483e+00 
R4400t1457 n4401 n1458 R=4.244e+00 
R4400t4395 n4401 n4396 R=2.033e+00 
R4400t1324 n4401 n1325 R=5.488e+01 
R4401t3056 n4402 n3057 R=2.762e+01 
R4401t4372 n4402 n4373 R=5.706e+00 
R4401t1445 n4402 n1446 R=1.781e+02 
R4401t4021 n4402 n4022 R=6.217e+00 
R4401t3154 n4402 n3155 R=1.348e+01 
R4401t4246 n4402 n4247 R=2.636e+01 
R4402t2162 n4403 n2163 R=7.619e+00 
R4402t2517 n4403 n2518 R=8.682e+00 
R4402t2054 n4403 n2055 R=4.079e+01 
R4402t1293 n4403 n1294 R=4.352e+00 
R4402t2280 n4403 n2281 R=1.109e+01 
R4402t2109 n4403 n2110 R=1.325e+01 
R4403t72 n4404 n73 R=5.757e+00 
R4403t1019 n4404 n1020 R=1.305e+01 
R4404t2522 n4405 n2523 R=1.416e+02 
R4405t1276 n4406 n1277 R=6.527e+00 
R4406t1138 n4407 n1139 R=9.365e+00 
R4407t186 n4408 n187 R=3.960e+00 
R4407t990 n4408 n991 R=1.024e+01 
R4407t4059 n4408 n4060 R=6.441e+00 
R4408t3247 n4409 n3248 R=5.169e+00 
R4408t2742 n4409 n2743 R=2.828e+00 
R4408t1490 n4409 n1491 R=3.512e+00 
R4409t1574 n4410 n1575 R=1.931e+00 
R4409t2758 n4410 n2759 R=4.050e+00 
R4410t2007 n4411 n2008 R=3.825e+01 
R4412t3514 n4413 n3515 R=2.469e+01 
R4412t3942 n4413 n3943 R=3.034e+01 
R4413t2427 n4414 n2428 R=4.457e+00 
R4413t3725 n4414 n3726 R=5.046e+00 
R4414t3312 n4415 n3313 R=3.698e+00 
R4415t2988 n4416 n2989 R=1.996e+00 
R4415t3597 n4416 n3598 R=1.621e+01 
R4415t300 n4416 n301 R=7.779e+01 
R4415t3802 n4416 n3803 R=2.630e+02 
R4416t3620 n4417 n3621 R=1.480e+01 
R4416t1646 n4417 n1647 R=5.413e+00 
R4416t110 n4417 n111 R=4.545e+01 
R4416t3009 n4417 n3010 R=9.567e+00 
R4418t2772 n4419 n2773 R=3.724e+00 
R4418t4243 n4419 n4244 R=1.326e+01 
R4419t2651 n4420 n2652 R=1.474e+01 
R4419t3287 n4420 n3288 R=1.542e+02 
R4419t1665 n4420 n1666 R=3.989e+00 
R4419t192 n4420 n193 R=8.879e+00 
R4419t3570 n4420 n3571 R=2.188e+01 
R4419t565 n4420 n566 R=5.498e+00 
R4420t11 n4421 n12 R=2.274e+01 
R4420t1819 n4421 n1820 R=8.218e+00 
R4420t3830 n4421 n3831 R=3.806e+01 
R4420t304 n4421 n305 R=4.214e+00 
R4420t1015 n4421 n1016 R=7.515e+00 
R4421t900 n4422 n901 R=1.147e+01 
R4421t3969 n4422 n3970 R=4.203e+00 
R4421t757 n4422 n758 R=2.273e+01 
R4421t50 n4422 n51 R=8.419e+00 
R4421t1973 n4422 n1974 R=1.160e+01 
R4421t3773 n4422 n3774 R=6.355e+00 
R4422t3114 n4423 n3115 R=7.109e+00 
R4423t355 n4424 n356 R=5.331e+00 
R4423t2567 n4424 n2568 R=9.593e+00 
R4424t2623 n4425 n2624 R=3.886e+00 
R4424t3434 n4425 n3435 R=4.087e+00 
R4425t4215 n4426 n4216 R=3.481e+01 
R4425t888 n4426 n889 R=3.883e+00 
R4426t2607 n4427 n2608 R=2.665e+01 
R4426t1599 n4427 n1600 R=2.342e+00 
R4427t2066 n4428 n2067 R=5.449e+00 
R4427t1459 n4428 n1460 R=3.536e+00 
R4428t1505 n4429 n1506 R=2.793e+01 
R4428t4283 n4429 n4284 R=5.965e+00 
R4428t4065 n4429 n4066 R=5.133e+00 
R4429t4005 n4430 n4006 R=8.356e+00 
R4429t1619 n4430 n1620 R=7.293e+01 
R4430t3331 n4431 n3332 R=6.085e+01 
R4430t404 n4431 n405 R=3.786e+00 
R4431t3427 n4432 n3428 R=2.860e+00 
R4432t3556 n4433 n3557 R=4.114e+00 
R4432t2908 n4433 n2909 R=4.183e+00 
R4432t2 n4433 n3 R=3.519e+00 
R4433t3772 n4434 n3773 R=6.864e+00 
R4433t2342 n4434 n2343 R=1.253e+02 
R4433t3833 n4434 n3834 R=3.422e+00 
R4434t2281 n4435 n2282 R=2.006e+01 
R4435t3047 n4436 n3048 R=7.483e+00 
R4435t4164 n4436 n4165 R=3.500e+01 
R4435t2255 n4436 n2256 R=4.581e+00 
R4436t1687 n4437 n1688 R=3.268e+00 
R4436t2191 n4437 n2192 R=1.003e+01 
R4437t4393 n4438 n4394 R=3.851e+00 
R4437t1135 n4438 n1136 R=6.299e+00 
R4438t906 n4439 n907 R=1.176e+01 
R4438t2290 n4439 n2291 R=3.222e+01 
R4438t3659 n4439 n3660 R=4.152e+00 
R4438t3585 n4439 n3586 R=9.389e+00 
R4438t569 n4439 n570 R=4.731e+00 
R4439t2782 n4440 n2783 R=3.551e+00 
R4439t741 n4440 n742 R=2.391e+02 
R4439t3413 n4440 n3414 R=2.740e+01 
R4439t1197 n4440 n1198 R=3.466e+00 
R4440t1940 n4441 n1941 R=2.074e+01 
R4440t3187 n4441 n3188 R=3.877e+01 
R4441t3395 n4442 n3396 R=3.327e+01 
R4441t1351 n4442 n1352 R=4.178e+00 
R4441t4106 n4442 n4107 R=1.210e+01 
R4443t1240 n4444 n1241 R=3.977e+02 
R4443t3933 n4444 n3934 R=1.628e+01 
R4443t3734 n4444 n3735 R=1.930e+01 
R4444t630 n4445 n631 R=4.043e+00 
R4444t3619 n4445 n3620 R=1.434e+01 
R4444t3813 n4445 n3814 R=7.204e+00 
R4445t4226 n4446 n4227 R=1.103e+02 
R4445t107 n4446 n108 R=6.960e+00 
R4445t2858 n4446 n2859 R=5.912e+01 
R4445t2793 n4446 n2794 R=1.216e+01 
R4446t1705 n4447 n1706 R=6.051e+01 
R4446t2055 n4447 n2056 R=7.435e+00 
R4447t821 n4448 n822 R=4.211e+00 
R4447t1877 n4448 n1878 R=1.486e+01 
R4447t2804 n4448 n2805 R=4.235e+01 
R4448t1865 n4449 n1866 R=1.026e+01 
R4449t3681 n4450 n3682 R=7.759e+00 
R4449t3931 n4450 n3932 R=4.149e+00 
R4449t806 n4450 n807 R=7.270e+00 
R4450t2761 n4451 n2762 R=2.581e+01 
R4450t834 n4451 n835 R=5.833e+00 
R4451t3968 n4452 n3969 R=1.673e+01 
R4451t3349 n4452 n3350 R=1.459e+01 
R4451t4333 n4452 n4334 R=7.290e+01 
R4451t3623 n4452 n3624 R=5.290e+00 
R4452t1087 n4453 n1088 R=9.628e+00 
R4452t2850 n4453 n1 R=3.138e+01 
R4453t1994 n4454 n1995 R=1.776e+01 
R4453t3206 n4454 n3207 R=9.580e+00 
R4453t3384 n4454 n3385 R=1.422e+02 
R4454t1944 n4455 n1945 R=5.799e+00 
R4454t1919 n4455 n1920 R=1.672e+01 
R4454t2734 n4455 n2735 R=4.293e+00 
R4454t4042 n4455 n4043 R=1.510e+01 
R4455t1994 n4456 n1995 R=2.806e+00 
R4455t4453 n4456 n4454 R=6.581e+00 
R4456t4284 n4457 n4285 R=4.585e+00 
R4456t4327 n4457 n4328 R=1.457e+01 
R4456t898 n4457 n899 R=6.471e+00 
R4457t1704 n4458 n1705 R=4.797e+00 
R4457t4246 n4458 n4247 R=3.334e+01 
R4457t4372 n4458 n4373 R=1.686e+01 
R4457t2310 n4458 n2311 R=2.901e+01 
R4458t545 n4459 n546 R=4.022e+00 
R4458t3304 n4459 n3305 R=4.381e+01 
R4458t1418 n4459 n1419 R=1.149e+01 
R4458t633 n4459 n634 R=5.466e+00 
R4458t3706 n4459 n3707 R=2.600e+00 
R4459t1983 n4460 n1984 R=2.432e+01 
R4459t3901 n4460 n3902 R=6.753e+00 
R4459t4276 n4460 n4277 R=3.464e+00 
R4459t2629 n4460 n2630 R=9.594e+00 
R4459t2935 n4460 n2936 R=7.117e+00 
R4459t2293 n4460 n2294 R=7.168e+00 
R4460t1304 n4461 n1305 R=6.045e+00 
R4460t2969 n4461 n2970 R=8.697e+00 
R4460t4143 n4461 n4144 R=5.734e+00 
R4460t1247 n4461 n1248 R=2.894e+00 
R4460t4022 n4461 n4023 R=1.551e+01 
R4461t116 n4462 n117 R=1.071e+02 
R4461t1134 n4462 n1135 R=7.540e+00 
R4462t2298 n4463 n2299 R=8.394e+00 
R4462t3595 n4463 n3596 R=4.452e+00 
R4462t3093 n4463 n3094 R=4.116e+00 
R4462t2678 n4463 n2679 R=5.119e+00 
R4462t2093 n4463 n2094 R=8.771e+00 
R4463t621 n4464 n622 R=2.170e+01 
R4463t3731 n4464 n3732 R=3.372e+00 
R4463t75 n4464 n76 R=1.132e+01 
R4463t3517 n4464 n3518 R=3.488e+00 
R4464t2714 n4465 n2715 R=1.092e+01 
R4464t1274 n4465 n1275 R=1.118e+01 
R4464t2221 n4465 n2222 R=1.309e+01 
R4465t416 n4466 n417 R=6.600e+00 
R4465t3546 n4466 n3547 R=1.593e+01 
R4466t2611 n4467 n2612 R=4.902e+01 
R4466t1878 n4467 n1879 R=3.073e+00 
R4467t41 n4468 n42 R=4.459e+00 
R4467t1699 n4468 n1700 R=1.727e+01 
R4467t3317 n4468 n3318 R=4.641e+00 
R4468t4312 n4469 n4313 R=5.736e+00 
R4468t2582 n4469 n2583 R=6.568e+00 
R4469t2501 n4470 n2502 R=7.288e+00 
R4469t3149 n4470 n3150 R=1.152e+01 
R4469t1113 n4470 n1114 R=7.625e+00 
R4470t363 n4471 n364 R=8.997e+00 
R4470t4172 n4471 n4173 R=2.118e+00 
R4470t4205 n4471 n4206 R=2.831e+00 
R4471t2265 n4472 n2266 R=1.396e+01 
R4471t2801 n4472 n2802 R=7.636e+00 
R4471t1992 n4472 n1993 R=2.102e+01 
R4471t1749 n4472 n1750 R=3.110e+00 
R4471t3834 n4472 n3835 R=6.437e+00 
R4472t3951 n4473 n1 R=1.368e+01 
R4472t4224 n4473 n4225 R=8.906e+00 
R4472t2476 n4473 n2477 R=2.368e+00 
R4472t987 n4473 n988 R=8.988e+01 
R4472t3325 n4473 n3326 R=9.258e+00 
R4473t454 n4474 n455 R=1.204e+01 
R4473t1352 n4474 n1353 R=3.879e+00 
R4473t133 n4474 n134 R=1.109e+01 
R4473t3852 n4474 n3853 R=7.939e+00 
R4473t3896 n4474 n3897 R=4.028e+01 
R4474t298 n4475 n299 R=2.232e+01 
R4474t899 n4475 n900 R=1.686e+01 
R4474t4260 n4475 n4261 R=3.546e+02 
R4474t1270 n4475 n1271 R=1.647e+01 
R4474t4103 n4475 n4104 R=2.168e+00 
R4474t4383 n4475 n4384 R=2.730e+01 
R4475t2070 n4476 n2071 R=1.141e+01 
R4475t1425 n4476 n1426 R=3.779e+00 
R4475t3326 n4476 n3327 R=4.555e+01 
R4476t1705 n4477 n1706 R=1.280e+01 
R4476t2039 n4477 n2040 R=2.730e+00 
R4476t3839 n4477 n3840 R=2.653e+00 
R4477t189 n4478 n190 R=7.341e+00 
R4477t2674 n4478 n2675 R=6.290e+00 
R4478t1186 n4479 n1187 R=9.259e+00 
R4478t3268 n4479 n3269 R=5.846e+00 
R4479t3188 n4480 n3189 R=5.354e+00 
R4480t2941 n4481 n2942 R=3.923e+00 
R4480t2859 n4481 n2860 R=7.972e+00 
R4481t3504 n4482 n3505 R=5.649e+00 
R4482t1090 n4483 n1091 R=3.904e+01 
R4482t1848 n4483 n1849 R=4.159e+00 
R4482t768 n4483 n769 R=1.162e+01 
R4483t138 n4484 n139 R=1.721e+01 
R4483t2650 n4484 n2651 R=4.073e+00 
R4483t46 n4484 n47 R=5.600e+00 
R4483t849 n4484 n850 R=3.483e+01 
R4484t1438 n4485 n1439 R=6.611e+00 
R4484t2697 n4485 n2698 R=5.531e+00 
R4484t2420 n4485 n2421 R=1.033e+01 
R4484t4188 n4485 n4189 R=4.653e+00 
R4484t3314 n4485 n3315 R=1.637e+01 
R4485t3014 n4486 n3015 R=3.633e+01 
R4485t309 n4486 n310 R=8.009e+00 
R4485t1194 n4486 n1195 R=7.703e+00 
R4485t372 n4486 n373 R=1.176e+01 
R4486t131 n4487 n132 R=1.720e+01 
R4486t1995 n4487 n1996 R=1.399e+01 
R4486t990 n4487 n991 R=8.640e+00 
R4486t4407 n4487 n4408 R=5.306e+00 
R4487t3255 n4488 n3256 R=6.933e+00 
R4487t3814 n4488 n3815 R=1.451e+01 
R4487t4290 n4488 n4291 R=2.991e+00 
R4488t1156 n4489 n1157 R=1.705e+01 
R4488t3510 n4489 n3511 R=4.456e+01 
R4488t3351 n4489 n3352 R=1.051e+01 
R4488t2607 n4489 n2608 R=5.126e+00 
R4489t1296 n4490 n1297 R=3.250e+01 
R4489t4114 n4490 n4115 R=5.008e+01 
R4489t330 n4490 n331 R=6.461e+00 
R4490t612 n4491 n613 R=3.453e+00 
R4490t1668 n4491 n1669 R=2.332e+00 
R4490t3019 n4491 n3020 R=7.662e+00 
R4491t2857 n4492 n2858 R=6.884e+00 
R4491t1809 n4492 n1810 R=5.783e+00 
R4492t2594 n4493 n2595 R=1.193e+01 
R4493t3472 n4494 n3473 R=5.914e+00 
R4493t1459 n4494 n1460 R=1.217e+01 
R4493t2066 n4494 n2067 R=3.055e+00 
R4494t3951 n4495 n1 R=6.140e+00 
R4494t4472 n4495 n4473 R=4.214e+00 
R4494t3325 n4495 n3326 R=5.539e+01 
R4494t398 n4495 n1 R=4.602e+00 
R4495t1206 n4496 n1207 R=3.463e+00 
R4495t2890 n4496 n2891 R=7.141e+00 
R4495t2426 n4496 n2427 R=8.263e+00 
R4495t554 n4496 n555 R=1.206e+01 
R4496t3794 n4497 n3795 R=3.143e+01 
R4496t3804 n4497 n3805 R=6.873e+00 
R4496t1157 n4497 n1158 R=5.489e+00 
R4496t3736 n4497 n3737 R=9.826e+00 
R4497t3109 n4498 n3110 R=4.793e+00 
R4498t2431 n4499 n2432 R=5.179e+01 
R4498t3473 n4499 n3474 R=1.125e+01 
R4498t3836 n4499 n3837 R=3.692e+00 
R4499t3227 n4500 n3228 R=2.915e+00 
R4499t1392 n4500 n1393 R=5.589e+00 
R4499t1591 n4500 n1592 R=5.583e+00 
R4500t2483 n4501 n2484 R=1.028e+02 
R4500t3880 n4501 n3881 R=4.066e+01 
R4500t2984 n4501 n2985 R=3.844e+00 
R4501t538 n4502 n539 R=3.373e+01 
R4501t4317 n4502 n4318 R=7.889e+00 
R4502t3591 n4503 n3592 R=2.402e+02 
R4502t1108 n4503 n1109 R=2.027e+00 
R4503t341 n4504 n342 R=7.654e+00 
R4503t3439 n4504 n3440 R=6.728e+00 
R4503t1775 n4504 n1776 R=1.226e+01 
R4503t201 n4504 n202 R=2.596e+01 
R4504t1552 n4505 n1553 R=6.743e+01 
R4504t2502 n4505 n2503 R=4.234e+00 
R4505t4037 n4506 n4038 R=4.373e+00 
R4505t3992 n4506 n3993 R=3.653e+01 
R4506t1878 n4507 n1879 R=4.137e+00 
R4506t4466 n4507 n4467 R=1.474e+01 
R4506t3263 n4507 n3264 R=2.287e+02 
R4507t3893 n4508 n3894 R=6.442e+00 
R4507t2576 n4508 n2577 R=2.399e+01 
R4507t3394 n4508 n3395 R=2.555e+00 
R4507t1379 n4508 n1380 R=6.664e+01 
R4507t3795 n4508 n3796 R=1.119e+02 
R4508t615 n4509 n616 R=4.328e+00 
R4508t4479 n4509 n4480 R=1.283e+01 
R4509t171 n4510 n172 R=8.410e+00 
R4509t2482 n4510 n2483 R=4.446e+00 
R4510t4134 n4511 n4135 R=1.465e+02 
R4510t164 n4511 n165 R=1.446e+01 
R4510t863 n4511 n864 R=5.961e+01 
R4510t487 n4511 n488 R=2.103e+00 
R4510t2207 n4511 n2208 R=4.230e+02 
R4511t1720 n4512 n1721 R=5.625e+00 
R4511t3636 n4512 n3637 R=4.207e+01 
R4512t1654 n4513 n1655 R=8.283e+00 
R4512t4152 n4513 n4153 R=5.086e+00 
R4513t24 n4514 n25 R=1.742e+00 
R4514t3109 n4515 n3110 R=2.769e+01 
R4514t4497 n4515 n4498 R=1.249e+01 
R4514t2399 n4515 n2400 R=7.866e+01 
R4515t943 n4516 n944 R=4.379e+01 
R4515t1812 n4516 n1813 R=2.967e+01 
R4516t3374 n4517 n3375 R=3.420e+01 
R4516t4225 n4517 n4226 R=2.239e+00 
R4517t3825 n4518 n3826 R=3.982e+00 
R4517t994 n4518 n995 R=5.626e+01 
R4518t401 n4519 n402 R=5.140e+00 
R4518t4119 n4519 n4120 R=2.822e+03 
R4518t2089 n4519 n2090 R=6.863e+00 
R4519t1407 n4520 n1408 R=4.352e+00 
R4519t3415 n4520 n3416 R=2.330e+01 
R4520t765 n4521 n766 R=8.935e+00 
R4520t3740 n4521 n3741 R=4.201e+00 
R4520t2493 n4521 n2494 R=1.025e+01 
R4520t3516 n4521 n3517 R=7.707e+00 
R4520t4006 n4521 n4007 R=1.836e+01 
R4521t1968 n4522 n1969 R=4.563e+00 
R4521t3672 n4522 n3673 R=5.312e+00 
R4522t1268 n4523 n1269 R=4.837e+00 
R4522t1787 n4523 n1788 R=1.865e+01 
R4523t3513 n4524 n3514 R=1.312e+01 
R4523t3448 n4524 n3449 R=7.821e+00 
R4524t160 n4525 n161 R=2.190e+00 
R4524t285 n4525 n286 R=4.848e+00 
R4525t665 n4526 n666 R=4.775e+00 
R4525t1326 n4526 n1327 R=4.259e+00 
R4525t3508 n4526 n3509 R=7.838e+00 
R4526t3401 n4527 n3402 R=2.655e+01 
R4526t1999 n4527 n2000 R=5.355e+00 
R4526t1214 n4527 n1215 R=9.996e+00 
R4526t98 n4527 n99 R=7.505e+00 
R4526t2331 n4527 n2332 R=1.508e+01 
R4527t3508 n4528 n3509 R=6.035e+00 
R4527t4525 n4528 n4526 R=3.846e+00 
R4527t665 n4528 n666 R=7.210e+00 
R4527t325 n4528 n326 R=3.013e+00 
R4528t1079 n4529 n1080 R=1.783e+01 
R4528t64 n4529 n65 R=3.363e+00 
R4528t460 n4529 n461 R=4.308e+01 
R4529t1797 n4530 n1798 R=5.829e+00 
R4529t1579 n4530 n1580 R=5.230e+00 
R4529t3135 n4530 n3136 R=3.259e+00 
R4530t1195 n1 n1196 R=6.274e+00 
R4530t1084 n1 n1085 R=4.668e+01 
R4531t2518 n4532 n2519 R=1.496e+01 
R4531t2205 n4532 n2206 R=5.802e+00 
R4532t2626 n4533 n2627 R=7.524e+00 
R4532t2561 n4533 n2562 R=8.314e+00 
R4532t3133 n4533 n3134 R=8.805e+00 
R4533t2217 n4534 n2218 R=4.472e+00 
R4533t2257 n4534 n2258 R=4.265e+00 
R4534t3449 n4535 n3450 R=3.750e+00 
R4534t1949 n4535 n1950 R=1.472e+01 
R4534t4345 n4535 n4346 R=2.231e+00 
R4535t2260 n4536 n2261 R=4.597e+01 
R4535t1397 n4536 n1398 R=3.434e+00 
R4536t3494 n4537 n3495 R=6.828e+01 
R4536t3509 n4537 n3510 R=6.799e+00 
R4536t4145 n4537 n4146 R=3.616e+00 
R4536t1780 n4537 n1781 R=6.444e+00 
R4537t1064 n4538 n1065 R=3.198e+01 
R4537t1043 n4538 n1044 R=9.177e+00 
R4537t1432 n4538 n1433 R=5.953e+00 
R4538t1532 n4539 n1533 R=1.207e+02 
R4538t2855 n4539 n2856 R=3.179e+01 
R4539t3182 n4540 n3183 R=3.569e+01 
R4539t4233 n4540 n4234 R=3.482e+00 
R4540t4447 n4541 n4448 R=5.279e+00 
R4541t1894 n4542 n1895 R=3.171e+01 
R4541t2729 n4542 n2730 R=8.188e+00 
R4541t357 n4542 n358 R=1.789e+01 
R4542t2744 n4543 n2745 R=5.234e+00 
R4542t3854 n4543 n3855 R=8.267e+00 
R4542t1755 n4543 n1756 R=2.975e+00 
R4542t4394 n4543 n4395 R=1.388e+03 
R4543t1116 n4544 n1117 R=3.866e+00 
R4544t468 n4545 n469 R=2.547e+00 
R4544t507 n4545 n508 R=2.498e+01 
R4544t4109 n4545 n4110 R=2.978e+01 
R4545t3173 n4546 n3174 R=1.638e+00 
R4545t4044 n4546 n4045 R=1.335e+02 
R4545t3986 n4546 n3987 R=8.085e+00 
R4547t167 n4548 n168 R=3.966e+01 
R4547t2753 n4548 n2754 R=5.530e+00 
R4547t3579 n4548 n3580 R=5.492e+00 
R4548t4540 n4549 n4541 R=5.591e+00 
R4548t4447 n4549 n4448 R=1.566e+01 
R4548t2804 n4549 n2805 R=2.787e+00 
R4549t3489 n4550 n3490 R=4.913e+00 
R4550t1094 n4551 n1095 R=8.926e+01 
R4550t1628 n4551 n1629 R=2.328e+01 
R4550t3565 n4551 n3566 R=9.595e+01 
R4550t3959 n4551 n3960 R=2.389e+01 
R4550t2022 n4551 n2023 R=7.878e+00 
R4550t3627 n4551 n3628 R=3.951e+00 
R4551t1905 n4552 n1906 R=5.999e+01 
R4551t294 n4552 n295 R=2.609e+01 
R4552t3512 n4553 n3513 R=4.288e+00 
R4552t3628 n4553 n3629 R=4.043e+01 
R4552t1555 n4553 n1556 R=1.118e+01 
R4553t1182 n4554 n1183 R=2.798e+01 
R4553t3667 n4554 n3668 R=2.230e+00 
R4554t652 n4555 n653 R=6.817e+01 
R4554t673 n4555 n674 R=2.812e+00 
R4554t758 n4555 n759 R=7.450e+00 
R4554t4221 n4555 n4222 R=1.883e+01 
R4554t33 n4555 n34 R=1.906e+00 
R4555t1745 n4556 n1746 R=8.460e+00 
R4556t1292 n4557 n1293 R=9.618e+00 
R4556t1427 n4557 n1428 R=1.586e+02 
R4556t1616 n4557 n1617 R=2.335e+00 
R4557t1959 n4558 n1960 R=9.959e+01 
R4557t3973 n4558 n3974 R=4.162e+00 
R4558t2334 n4559 n2335 R=3.008e+00 
R4558t2388 n4559 n2389 R=5.738e+00 
R4559t2635 n4560 n2636 R=7.415e+00 
R4559t729 n4560 n730 R=2.074e+00 
R4559t359 n4560 n360 R=7.832e+00 
R4560t254 n4561 n255 R=3.873e+00 
R4560t3866 n4561 n3867 R=1.804e+01 
R4560t4162 n4561 n4163 R=1.111e+01 
R4561t546 n4562 n547 R=1.604e+01 
R4561t3705 n4562 n3706 R=1.079e+01 
R4561t1225 n4562 n1226 R=2.854e+00 
R4562t1303 n4563 n1304 R=6.192e+00 
R4562t1299 n4563 n1300 R=2.942e+01 
R4563t4199 n4564 n4200 R=5.499e+00 
R4564t1318 n4565 n1319 R=7.296e+00 
R4564t2258 n4565 n2259 R=9.721e+00 
R4564t4041 n4565 n4042 R=7.597e+00 
R4564t3846 n4565 n3847 R=1.066e+01 
R4565t2968 n4566 n2969 R=1.097e+01 
R4565t3670 n4566 n3671 R=5.371e+00 
R4565t2393 n4566 n2394 R=4.723e+00 
R4566t432 n4567 n433 R=6.225e+02 
R4566t3461 n4567 n3462 R=9.290e+00 
R4566t4111 n4567 n4112 R=1.459e+02 
R4566t3242 n4567 n3243 R=3.109e+00 
R4566t4390 n4567 n4391 R=1.392e+01 
R4567t4222 n4568 n4223 R=1.080e+01 
R4568t3507 n4569 n3508 R=2.746e+00 
R4568t4317 n4569 n4318 R=9.302e+00 
R4568t4501 n4569 n4502 R=4.149e+00 
R4569t1155 n4570 n1156 R=2.638e+00 
R4569t2232 n4570 n2233 R=2.186e+00 
R4570t10 n4571 n11 R=1.604e+01 
R4570t4465 n4571 n4466 R=2.637e+00 
R4571t1098 n4572 n1099 R=2.191e+01 
R4571t3936 n4572 n3937 R=8.763e+00 
R4571t2562 n4572 n2563 R=3.096e+01 
R4571t3751 n4572 n3752 R=1.772e+02 
R4571t1718 n4572 n1719 R=3.282e+00 
R4571t1332 n4572 n1333 R=2.470e+01 
R4571t3208 n4572 n3209 R=4.454e+00 
R4572t3718 n4573 n3719 R=2.602e+00 
R4572t3726 n4573 n3727 R=2.120e+01 
R4572t30 n4573 n31 R=4.178e+00 
R4572t1796 n4573 n1797 R=8.745e+00 
R4573t3433 n4574 n3434 R=8.268e+00 
R4573t991 n4574 n992 R=1.071e+01 
R4574t2295 n4575 n2296 R=2.235e+01 
R4574t43 n4575 n44 R=3.509e+00 
R4575t1835 n4576 n1836 R=2.084e+02 
R4575t3329 n4576 n3330 R=6.994e+00 
R4575t116 n4576 n117 R=1.805e+02 
R4575t2185 n4576 n2186 R=9.904e+00 
R4576t264 n4577 n265 R=1.066e+01 
R4576t2906 n4577 n2907 R=1.058e+01 
R4576t3207 n4577 n3208 R=1.281e+01 
R4577t173 n4578 n174 R=2.999e+01 
R4577t2803 n4578 n2804 R=2.815e+01 
R4577t1093 n4578 n1094 R=9.617e+00 
R4577t627 n4578 n628 R=1.033e+02 
R4578t3193 n4579 n3194 R=4.483e+00 
R4579t4072 n4580 n4073 R=3.491e+01 
R4579t1542 n4580 n1543 R=5.879e+00 
R4579t2365 n4580 n2366 R=4.710e+00 
R4579t2641 n4580 n2642 R=8.494e+00 
R4580t4203 n4581 n4204 R=3.016e+00 
R4581t2329 n4582 n2330 R=5.264e+00 
R4581t917 n4582 n918 R=9.950e+00 
R4582t3543 n4583 n3544 R=2.168e+00 
R4582t4060 n4583 n4061 R=7.103e+01 
R4582t3259 n4583 n3260 R=2.272e+02 
R4582t86 n4583 n87 R=3.437e+01 
R4583t3806 n4584 n3807 R=1.089e+02 
R4583t1373 n4584 n1374 R=2.774e+00 
R4583t2955 n4584 n2956 R=1.637e+01 
R4583t3109 n4584 n3110 R=1.468e+01 
R4584t834 n4585 n835 R=1.731e+02 
R4584t4450 n4585 n4451 R=9.352e+00 
R4584t2175 n4585 n2176 R=3.678e+01 
R4584t1780 n4585 n1781 R=6.773e+00 
R4585t1192 n4586 n1193 R=1.061e+01 
R4585t1630 n4586 n1631 R=5.952e+00 
R4585t629 n4586 n630 R=2.497e+01 
R4586t1774 n4587 n1775 R=7.255e+00 
R4587t2515 n4588 n2516 R=1.541e+02 
R4587t1699 n4588 n1700 R=5.422e+01 
R4587t1310 n4588 n1311 R=1.031e+01 
R4588t2070 n4589 n2071 R=3.230e+01 
R4589t2829 n4590 n2830 R=4.019e+01 
R4589t3723 n4590 n3724 R=1.240e+01 
R4589t2946 n4590 n2947 R=3.830e+00 
R4590t2178 n4591 n2179 R=1.164e+01 
R4590t1813 n4591 n1814 R=1.752e+01 
R4590t3912 n4591 n3913 R=1.197e+01 
R4591t4180 n4592 n4181 R=4.773e+00 
R4591t544 n4592 n545 R=1.222e+01 
R4592t514 n4593 n515 R=1.696e+01 
R4592t1264 n4593 n1265 R=3.149e+01 
R4592t1278 n4593 n1279 R=6.626e+00 
R4592t1461 n4593 n1462 R=1.290e+01 
R4592t2366 n4593 n2367 R=6.819e+00 
R4592t3631 n4593 n3632 R=1.543e+01 
R4593t3040 n4594 n3041 R=1.484e+01 
R4593t2855 n4594 n2856 R=1.208e+01 
R4593t2586 n4594 n2587 R=9.518e+00 
R4593t3262 n4594 n3263 R=1.439e+01 
R4594t3508 n4595 n3509 R=9.548e+00 
R4594t4527 n4595 n4528 R=1.165e+02 
R4594t4015 n4595 n4016 R=4.909e+01 
R4594t1393 n4595 n1394 R=1.752e+01 
R4594t521 n4595 n522 R=7.147e+00 
R4594t325 n4595 n326 R=4.264e+00 
R4595t2483 n4596 n2484 R=4.256e+00 
R4595t2984 n4596 n2985 R=2.455e+00 
R4595t3259 n4596 n3260 R=1.190e+01 
R4595t484 n4596 n485 R=8.327e+00 
R4596t2195 n4597 n2196 R=4.320e+00 
R4596t3249 n4597 n3250 R=7.153e+00 
R4596t2503 n4597 n2504 R=8.958e+00 
R4596t3370 n4597 n3371 R=7.635e+00 
R4597t1146 n4598 n1147 R=4.380e+00 
R4597t3917 n4598 n3918 R=2.219e+01 
R4597t1875 n4598 n1876 R=1.122e+01 
R4597t3344 n4598 n3345 R=2.297e+01 
R4598t3565 n4599 n3566 R=3.336e+01 
R4598t1979 n4599 n1980 R=9.183e+00 
R4598t856 n4599 n857 R=6.008e+00 
R4599t4361 n4600 n4362 R=5.562e+00 
R4599t1672 n4600 n1673 R=5.592e+01 
R4599t2249 n4600 n2250 R=1.347e+01 
R4599t2466 n4600 n2467 R=9.268e+00 
R4599t3889 n4600 n3890 R=1.782e+01 
R4601t1633 n4602 n1634 R=3.980e+00 
R4601t2901 n4602 n2902 R=3.190e+00 
R4602t1734 n4603 n1735 R=8.221e+00 
R4602t3296 n4603 n3297 R=6.791e+00 
R4602t310 n4603 n311 R=4.512e+00 
R4602t1869 n4603 n1870 R=1.524e+01 
R4603t740 n4604 n741 R=1.615e+01 
R4603t3850 n4604 n3851 R=9.408e+00 
R4604t1659 n4605 n1660 R=2.540e+00 
R4605t4097 n4606 n4098 R=1.155e+01 
R4606t2543 n4607 n2544 R=8.011e+01 
R4606t4245 n4607 n4246 R=5.920e+01 
R4606t850 n4607 n851 R=9.508e+00 
R4608t3292 n4609 n3293 R=6.814e+00 
R4609t327 n1 n328 R=3.738e+00 
R4610t2076 n4611 n2077 R=8.128e+00 
R4610t657 n4611 n658 R=3.745e+01 
R4611t903 n4612 n904 R=9.436e+00 
R4611t314 n4612 n315 R=1.220e+01 
R4611t492 n4612 n493 R=3.760e+00 
R4612t3657 n4613 n3658 R=3.336e+00 
R4612t1517 n4613 n1518 R=3.643e+00 
R4613t3643 n4614 n3644 R=2.708e+00 
R4613t4346 n4614 n4347 R=2.625e+01 
R4613t1832 n4614 n1833 R=8.376e+00 
R4613t2370 n4614 n2371 R=1.009e+01 
R4613t800 n4614 n801 R=8.543e+00 
R4614t1256 n4615 n1257 R=3.930e+00 
R4614t4016 n4615 n4017 R=3.528e+00 
R4614t2936 n4615 n2937 R=1.133e+02 
R4615t1027 n4616 n1028 R=2.790e+00 
R4615t1756 n4616 n1757 R=1.018e+01 
R4615t2760 n4616 n2761 R=1.814e+01 
R4616t1271 n4617 n1 R=2.541e+01 
R4616t2046 n4617 n1 R=1.118e+01 
R4616t4362 n4617 n4363 R=6.522e+00 
R4616t3796 n4617 n3797 R=3.821e+00 
R4617t160 n4618 n161 R=8.189e+00 
R4617t3293 n4618 n3294 R=6.185e+00 
R4617t1236 n4618 n1237 R=9.927e+00 
R4618t1180 n4619 n1181 R=6.830e+00 
R4618t117 n4619 n118 R=3.169e+01 
R4618t878 n4619 n879 R=5.815e+00 
R4618t1316 n4619 n1317 R=9.835e+00 
R4618t2400 n4619 n2401 R=9.404e+00 
R4619t4445 n4620 n4446 R=1.412e+01 
R4619t2878 n4620 n2879 R=6.746e+00 
R4619t107 n4620 n108 R=1.001e+02 
R4620t3962 n4621 n3963 R=4.557e+00 
R4621t985 n4622 n986 R=5.661e+00 
R4621t251 n4622 n252 R=3.374e+00 
R4621t2802 n4622 n2803 R=5.052e+00 
R4621t3998 n4622 n3999 R=8.424e+00 
R4622t952 n4623 n953 R=5.087e+00 
R4622t2714 n4623 n2715 R=1.642e+02 
R4622t3504 n4623 n3505 R=7.362e+00 
R4622t1901 n4623 n1902 R=1.844e+01 
R4622t2099 n4623 n2100 R=1.011e+01 
R4623t1491 n4624 n1492 R=1.143e+01 
R4623t1345 n4624 n1346 R=6.568e+00 
R4623t3012 n4624 n3013 R=7.146e+00 
R4624t1659 n4625 n1660 R=5.748e+00 
R4624t579 n4625 n580 R=6.758e+00 
R4625t2591 n4626 n2592 R=5.619e+00 
R4625t4006 n4626 n4007 R=6.738e+00 
R4626t4504 n4627 n4505 R=2.974e+00 
R4626t2502 n4627 n2503 R=9.587e+00 
R4626t2610 n4627 n1 R=3.080e+00 
R4627t2526 n4628 n2527 R=1.751e+00 
R4627t20 n4628 n21 R=8.022e+00 
R4628t1102 n4629 n1103 R=5.677e+00 
R4628t395 n4629 n396 R=1.290e+01 
R4628t895 n4629 n896 R=1.578e+01 
R4629t1364 n4630 n1365 R=3.514e+01 
R4629t2915 n4630 n2916 R=4.012e+00 
R4629t2333 n4630 n2334 R=7.803e+00 
R4630t3945 n4631 n3946 R=1.734e+01 
R4630t2385 n4631 n2386 R=1.812e+01 
R4630t767 n4631 n768 R=7.235e+00 
R4631t1301 n4632 n1302 R=2.216e+00 
R4631t3078 n4632 n3079 R=7.989e+00 
R4631t3265 n4632 n3266 R=3.414e+00 
R4632t1759 n4633 n1760 R=4.831e+00 
R4632t1654 n4633 n1655 R=4.322e+01 
R4632t2886 n4633 n2887 R=6.340e+01 
R4632t3769 n4633 n3770 R=5.531e+01 
R4632t1745 n4633 n1746 R=4.047e+00 
R4632t4555 n4633 n4556 R=4.819e+01 
R4633t1697 n4634 n1698 R=2.622e+00 
R4633t1220 n4634 n1221 R=6.114e+00 
R4634t1890 n4635 n1891 R=6.964e+00 
R4634t4068 n4635 n4069 R=8.302e+00 
R4634t4175 n4635 n4176 R=1.211e+01 
R4635t1165 n4636 n1166 R=1.048e+01 
R4635t1937 n4636 n1938 R=2.497e+01 
R4635t2035 n4636 n2036 R=2.144e+01 
R4635t3385 n4636 n3386 R=1.290e+02 
R4636t4141 n4637 n4142 R=9.032e+00 
R4636t4337 n4637 n4338 R=5.566e+00 
R4636t2807 n4637 n2808 R=5.481e+00 
R4636t3213 n4637 n3214 R=4.513e+01 
R4638t3447 n4639 n3448 R=4.587e+00 
R4638t3806 n4639 n3807 R=2.250e+01 
R4639t4515 n4640 n4516 R=6.540e+01 
R4639t943 n4640 n944 R=9.609e+00 
R4639t4296 n4640 n4297 R=4.614e+00 
R4639t2805 n4640 n2806 R=1.508e+01 
R4640t1847 n4641 n1848 R=2.030e+01 
R4640t1628 n4641 n1629 R=7.988e+00 
R4640t3565 n4641 n3566 R=5.513e+00 
R4640t4598 n4641 n4599 R=9.451e+00 
R4641t1488 n4642 n1489 R=8.250e+00 
R4642t4510 n4643 n4511 R=1.878e+01 
R4642t2207 n4643 n2208 R=2.818e+00 
R4642t3355 n4643 n3356 R=5.111e+00 
R4643t1062 n4644 n1063 R=4.266e+00 
R4644t1761 n4645 n1762 R=8.969e+00 
R4644t2662 n4645 n2663 R=5.933e+01 
R4645t1460 n4646 n1461 R=6.373e+00 
R4645t1520 n4646 n1521 R=3.022e+00 
R4645t2773 n4646 n2774 R=1.249e+01 
R4646t687 n4647 n688 R=3.515e+01 
R4646t2939 n4647 n2940 R=2.347e+00 
R4646t2945 n4647 n2946 R=7.049e+01 
R4647t3202 n4648 n3203 R=1.186e+01 
R4647t4045 n4648 n4046 R=3.792e+01 
R4647t3352 n4648 n3353 R=1.355e+01 
R4647t1715 n4648 n1716 R=2.423e+00 
R4648t447 n4649 n448 R=3.014e+00 
R4648t1321 n4649 n1322 R=3.384e+00 
R4649t382 n4650 n383 R=2.749e+01 
R4649t4120 n4650 n4121 R=1.485e+01 
R4649t4053 n4650 n4054 R=1.316e+01 
R4649t958 n4650 n959 R=5.376e+00 
R4650t2646 n4651 n2647 R=1.895e+01 
R4650t4638 n4651 n4639 R=3.766e+00 
R4650t3806 n4651 n3807 R=2.277e+01 
R4651t621 n4652 n622 R=2.713e+00 
R4651t3517 n4652 n3518 R=4.803e+00 
R4651t2006 n4652 n2007 R=1.586e+01 
R4652t3704 n4653 n3705 R=3.729e+00 
R4652t317 n4653 n318 R=6.286e+00 
R4652t1644 n4653 n1645 R=1.862e+02 
R4653t241 n4654 n242 R=5.129e+00 
R4653t660 n4654 n661 R=5.896e+00 
R4654t2641 n4655 n2642 R=2.483e+01 
R4654t3644 n4655 n3645 R=5.953e+00 
R4654t2365 n4655 n2366 R=4.433e+00 
R4655t4219 n4656 n4220 R=3.982e+00 
R4655t2902 n4656 n2903 R=1.250e+01 
R4655t979 n4656 n980 R=4.622e+00 
R4656t2309 n4657 n2310 R=3.839e+00 
R4656t3988 n4657 n3989 R=1.276e+01 
R4656t2032 n4657 n2033 R=1.031e+01 
R4658t1371 n4659 n1372 R=1.168e+01 
R4658t215 n4659 n216 R=9.196e+00 
R4658t4254 n4659 n4255 R=2.511e+00 
R4659t2607 n4660 n2608 R=5.343e+00 
R4659t4426 n4660 n4427 R=6.540e+00 
R4659t4488 n4660 n4489 R=2.048e+01 
R4659t96 n4660 n97 R=5.518e+00 
R4659t4256 n4660 n4257 R=4.130e+00 
R4659t1599 n4660 n1600 R=3.238e+02 
R4660t2623 n4661 n2624 R=1.464e+00 
R4660t994 n4661 n995 R=1.543e+02 
R4660t4517 n4661 n4518 R=2.548e+00 
R4660t3825 n4661 n3826 R=4.433e+01 
R4661t4299 n4662 n4300 R=1.461e+01 
R4661t1358 n4662 n1359 R=7.155e+01 
R4661t590 n4662 n591 R=7.117e+00 
R4662t1000 n4663 n1001 R=4.440e+00 
R4662t1354 n4663 n1355 R=2.023e+01 
R4662t3601 n4663 n3602 R=2.146e+00 
R4662t1244 n4663 n1245 R=5.934e+01 
R4662t3966 n4663 n3967 R=4.424e+00 
R4663t3970 n4664 n3971 R=5.580e+00 
R4663t3274 n4664 n3275 R=1.784e+01 
R4663t403 n4664 n404 R=1.643e+01 
R4663t1044 n4664 n1045 R=1.001e+01 
R4664t983 n4665 n984 R=2.757e+02 
R4664t2625 n4665 n2626 R=9.677e+00 
R4664t2138 n4665 n2139 R=5.337e+00 
R4664t994 n4665 n995 R=8.493e+00 
R4664t4517 n4665 n4518 R=3.509e+00 
R4664t3825 n4665 n3826 R=1.058e+01 
R4664t2130 n4665 n2131 R=9.824e+01 
R4664t1570 n4665 n1571 R=1.379e+01 
R4665t2001 n4666 n2002 R=4.018e+00 
R4665t996 n4666 n997 R=2.984e+00 
R4666t4042 n1 n4043 R=3.388e+00 
R4667t588 n4668 n589 R=2.685e+00 
R4667t946 n4668 n947 R=4.736e+01 
R4667t2024 n4668 n2025 R=2.659e+01 
R4667t4050 n4668 n4051 R=1.224e+01 
R4668t1406 n4669 n1407 R=3.365e+00 
R4668t3391 n4669 n3392 R=4.983e+00 
R4668t1206 n4669 n1207 R=4.142e+01 
R4668t3566 n4669 n3567 R=3.305e+01 
R4668t1473 n4669 n1474 R=1.754e+00 
R4669t922 n4670 n923 R=2.652e+00 
R4669t392 n4670 n393 R=9.655e+00 
R4669t883 n4670 n884 R=8.265e+00 
R4669t370 n4670 n371 R=4.999e+01 
R4669t3661 n4670 n3662 R=4.002e+00 
R4670t2222 n4671 n2223 R=6.093e+00 
R4670t2864 n4671 n2865 R=1.030e+01 
R4670t4178 n4671 n4179 R=4.729e+00 
R4670t4192 n4671 n4193 R=5.424e+02 
R4670t247 n4671 n248 R=3.734e+00 
R4670t869 n4671 n870 R=8.111e+02 
R4671t2829 n4672 n2830 R=3.126e+00 
R4672t4667 n4673 n4668 R=1.450e+01 
R4672t3381 n4673 n3382 R=3.657e+01 
R4672t946 n4673 n947 R=4.719e+00 
R4673t1831 n4674 n1832 R=8.654e+00 
R4673t950 n4674 n951 R=1.516e+01 
R4673t1688 n4674 n1689 R=4.346e+00 
R4674t35 n4675 n36 R=7.275e+00 
R4674t125 n4675 n126 R=1.346e+01 
R4674t3876 n4675 n3877 R=1.209e+01 
R4674t3424 n4675 n3425 R=6.601e+00 
R4675t3525 n4676 n3526 R=1.271e+01 
R4675t4213 n4676 n4214 R=2.998e+00 
R4676t310 n4677 n311 R=4.941e+00 
R4676t4651 n4677 n4652 R=3.893e+00 
R4676t949 n4677 n950 R=2.111e+01 
R4676t2562 n4677 n2563 R=2.072e+01 
R4677t2817 n4678 n2818 R=2.666e+00 
R4677t3802 n4678 n3803 R=6.778e+00 
R4678t1213 n4679 n1214 R=5.593e+00 
R4678t21 n4679 n22 R=9.727e+00 
R4679t815 n4680 n816 R=2.188e+01 
R4680t129 n4681 n130 R=1.227e+01 
R4680t868 n4681 n869 R=4.674e+01 
R4680t2851 n4681 n2852 R=2.461e+01 
R4680t1638 n4681 n1639 R=3.782e+00 
R4681t983 n4682 n984 R=7.593e+00 
R4681t2507 n4682 n2508 R=7.591e+00 
R4681t1960 n4682 n1961 R=8.574e+00 
R4681t2993 n4682 n2994 R=3.983e+00 
R4682t3307 n4683 n3308 R=3.919e+00 
R4682t1492 n4683 n1493 R=5.222e+00 
R4682t1130 n4683 n1131 R=6.648e+01 
R4683t1895 n4684 n1896 R=2.449e+01 
R4683t3185 n4684 n3186 R=2.746e+00 
R4683t3367 n4684 n3368 R=1.858e+01 
R4684t4380 n4685 n4381 R=4.205e+01 
R4684t3100 n4685 n3101 R=6.609e+00 
R4685t4573 n4686 n4574 R=1.414e+01 
R4685t3433 n4686 n3434 R=6.978e+00 
R4685t1601 n4686 n1602 R=2.898e+01 
R4685t824 n4686 n825 R=1.565e+01 
R4685t367 n4686 n368 R=5.872e+01 
R4686t527 n4687 n528 R=4.644e+00 
R4687t710 n4688 n711 R=1.416e+01 
R4687t3929 n4688 n3930 R=5.796e+00 
R4687t734 n4688 n735 R=7.229e+01 
R4687t150 n4688 n151 R=2.586e+01 
R4688t3694 n4689 n3695 R=4.136e+00 
R4688t3944 n4689 n3945 R=3.499e+00 
R4688t798 n4689 n799 R=1.418e+01 
R4688t500 n4689 n501 R=2.652e+01 
R4689t3122 n4690 n3123 R=1.817e+01 
R4690t1516 n4691 n1517 R=2.282e+01 
R4691t717 n4692 n718 R=7.640e+00 
R4691t1667 n4692 n1668 R=3.451e+00 
R4691t4049 n4692 n4050 R=2.860e+01 
R4692t4411 n4693 n4412 R=8.829e+00 
R4692t3888 n4693 n3889 R=4.341e+00 
R4692t4273 n4693 n4274 R=7.904e+00 
R4693t958 n4694 n959 R=3.741e+00 
R4693t4649 n4694 n4650 R=1.276e+01 
R4693t479 n4694 n480 R=3.917e+00 
R4694t74 n4695 n75 R=3.300e+00 
R4694t4433 n4695 n4434 R=1.185e+01 
R4694t3772 n4695 n3773 R=2.461e+00 
R4695t3721 n4696 n3722 R=1.878e+01 
R4695t2695 n4696 n2696 R=2.773e+01 
R4695t1427 n4696 n1428 R=1.540e+01 
R4695t3099 n4696 n3100 R=3.382e+01 
R4697t1986 n4698 n1987 R=9.109e+00 
R4697t697 n4698 n698 R=7.340e+01 
R4697t3621 n4698 n3622 R=2.611e+00 
R4698t1184 n4699 n1185 R=2.733e+00 
R4698t3824 n4699 n3825 R=9.174e+00 
R4699t3516 n4700 n3517 R=3.192e+01 
R4699t4006 n4700 n4007 R=3.177e+01 
R4699t70 n4700 n71 R=1.953e+01 
R4699t528 n4700 n529 R=3.611e+00 
R4699t680 n4700 n681 R=2.515e+01 
R4699t3670 n4700 n3671 R=7.167e+01 
R4700t3575 n4701 n3576 R=7.478e+00 
R4700t3707 n4701 n3708 R=2.082e+01 
R4700t2398 n4701 n2399 R=5.190e+02 
R4700t502 n4701 n503 R=1.493e+01 
R4701t2008 n4702 n2009 R=4.897e+00 
R4702t2323 n4703 n2324 R=3.433e+01 
R4702t1681 n4703 n1682 R=3.024e+01 
R4702t1969 n4703 n1970 R=8.340e+00 
R4702t2474 n4703 n2475 R=8.381e+00 
R4703t2354 n4704 n2355 R=1.339e+01 
R4703t3535 n4704 n3536 R=1.385e+01 
R4703t1526 n4704 n1527 R=3.255e+00 
R4703t4314 n4704 n4315 R=4.197e+01 
R4703t3553 n4704 n3554 R=2.921e+00 
R4704t2757 n4705 n2758 R=4.936e+00 
R4704t1809 n4705 n1810 R=1.643e+01 
R4704t3688 n4705 n3689 R=1.959e+01 
R4704t2465 n4705 n2466 R=3.325e+00 
R4704t805 n4705 n806 R=5.920e+00 
R4705t1148 n4706 n1149 R=8.278e+00 
R4705t4437 n4706 n4438 R=1.663e+01 
R4706t1137 n4707 n1138 R=1.557e+01 
R4706t3016 n4707 n3017 R=2.830e+00 
R4706t3684 n4707 n3685 R=3.758e+01 
R4707t715 n4708 n716 R=5.118e+00 
R4707t4259 n4708 n4260 R=1.171e+01 
R4708t792 n4709 n793 R=4.097e+00 
R4708t3351 n4709 n3352 R=8.517e+00 
R4708t1264 n4709 n1265 R=3.642e+00 
R4708t1278 n4709 n1279 R=6.075e+00 
R4709t3024 n4710 n3025 R=1.648e+01 
R4709t4036 n4710 n4037 R=6.657e+00 
R4709t205 n4710 n206 R=1.115e+03 
R4709t4225 n4710 n4226 R=3.726e+01 
R4709t4516 n4710 n4517 R=1.190e+02 
R4709t1664 n4710 n1665 R=2.455e+00 
R4709t2019 n4710 n2020 R=8.981e+01 
R4710t886 n4711 n887 R=2.177e+00 
R4710t4047 n4711 n4048 R=4.044e+01 
R4710t1668 n4711 n1669 R=2.236e+01 
R4710t4490 n4711 n4491 R=6.028e+00 
R4710t612 n4711 n613 R=1.093e+01 
R4711t4110 n4712 n4111 R=3.424e+00 
R4711t1198 n4712 n1199 R=3.554e+00 
R4711t2305 n4712 n2306 R=8.538e+00 
R4712t1890 n4713 n1891 R=4.054e+00 
R4712t4634 n4713 n4635 R=3.779e+01 
R4712t1608 n4713 n1609 R=6.255e+00 
R4712t2923 n4713 n2924 R=3.449e+01 
R4713t2023 n4714 n2024 R=3.286e+01 
R4713t1061 n4714 n1062 R=4.932e+01 
R4714t740 n4715 n741 R=3.602e+01 
R4714t1344 n4715 n1345 R=1.060e+01 
R4714t633 n4715 n634 R=1.709e+01 
R4714t3706 n4715 n3707 R=2.619e+00 
R4714t1843 n4715 n1844 R=8.743e+00 
R4714t2834 n4715 n2835 R=3.671e+00 
R4715t4022 n4716 n4023 R=6.074e+00 
R4715t1675 n4716 n1676 R=1.072e+01 
R4716t1908 n4717 n1909 R=6.525e+00 
R4716t4207 n4717 n4208 R=7.289e+00 
R4717t2310 n4718 n2311 R=2.247e+00 
R4717t4457 n4718 n4458 R=3.819e+00 
R4718t746 n4719 n747 R=7.112e+00 
R4718t1218 n4719 n1219 R=5.190e+00 
R4718t1056 n4719 n1057 R=4.068e+00 
R4719t1061 n4720 n1062 R=3.270e+00 
R4719t1643 n4720 n1644 R=1.877e+01 
R4719t1793 n4720 n1794 R=2.878e+01 
R4720t3182 n4721 n3183 R=8.715e+00 
R4720t4539 n4721 n4540 R=5.819e+00 
R4720t2736 n4721 n2737 R=2.650e+01 
R4720t2960 n4721 n2961 R=3.471e+00 
R4721t114 n4722 n115 R=6.327e+00 
R4721t1673 n4722 n1674 R=6.970e+00 
R4721t1627 n4722 n1628 R=7.948e+00 
R4721t1240 n4722 n1241 R=1.968e+01 
R4721t346 n4722 n347 R=7.107e+00 
R4722t2489 n4723 n2490 R=3.022e+00 
R4723t232 n4724 n233 R=2.679e+00 
R4724t2468 n4725 n2469 R=3.631e+01 
R4724t2173 n4725 n2174 R=6.068e+00 
R4725t908 n4726 n909 R=3.640e+00 
R4725t3423 n4726 n3424 R=7.789e+00 
R4725t838 n4726 n839 R=9.333e+00 
R4726t4017 n4727 n4018 R=1.559e+01 
R4726t4083 n4727 n4084 R=9.428e+00 
R4726t2862 n4727 n2863 R=5.763e+00 
R4727t2908 n4728 n2909 R=8.202e+00 
R4728t1602 n4729 n1603 R=1.544e+01 
R4728t2101 n4729 n2102 R=4.199e+00 
R4729t81 n4730 n82 R=1.257e+01 
R4729t2533 n4730 n2534 R=1.691e+01 
R4729t1000 n4730 n1001 R=7.680e+00 
R4729t4040 n4730 n4041 R=3.307e+00 
R4730t991 n4731 n992 R=7.704e+00 
R4730t3041 n4731 n3042 R=3.854e+01 
R4730t2928 n4731 n2929 R=2.334e+01 
R4730t2997 n4731 n2998 R=3.672e+00 
R4731t3487 n4732 n3488 R=6.637e+00 
R4731t758 n4732 n759 R=5.462e+00 
R4732t1507 n4733 n1508 R=3.766e+00 
R4732t3172 n4733 n3173 R=2.033e+01 
R4733t1931 n4734 n1932 R=1.043e+01 
R4733t3854 n4734 n3855 R=4.779e+00 
R4733t4542 n4734 n4543 R=2.315e+01 
R4733t1755 n4734 n1756 R=4.231e+01 
R4733t4115 n4734 n4116 R=4.642e+00 
R4734t1234 n4735 n1235 R=6.343e+00 
R4734t1828 n4735 n1829 R=6.159e+00 
R4734t4234 n4735 n4235 R=5.323e+00 
R4734t1617 n4735 n1618 R=9.340e+00 
R4735t2978 n4736 n2979 R=4.870e+02 
R4735t4203 n4736 n4204 R=6.762e+00 
R4736t2297 n4737 n2298 R=1.826e+01 
R4736t3770 n4737 n3771 R=2.990e+00 
R4736t683 n4737 n684 R=7.513e+00 
R4736t4350 n4737 n4351 R=2.661e+01 
R4737t1734 n4738 n1735 R=2.714e+00 
R4737t4141 n4738 n4142 R=1.563e+02 
R4737t3936 n4738 n3937 R=4.859e+00 
R4738t1059 n4739 n1060 R=1.515e+01 
R4738t601 n4739 n602 R=1.657e+01 
R4738t159 n4739 n160 R=1.986e+00 
R4739t4160 n4740 n4161 R=3.651e+00 
R4739t252 n4740 n253 R=9.478e+01 
R4739t3333 n4740 n3334 R=3.297e+01 
R4739t3290 n4740 n3291 R=1.042e+01 
R4740t2958 n4741 n2959 R=1.023e+01 
R4741t833 n4742 n834 R=7.368e+00 
R4741t2899 n4742 n2900 R=6.414e+00 
R4742t2437 n4743 n2438 R=5.855e+00 
R4743t635 n4744 n636 R=1.790e+01 
R4743t2370 n4744 n2371 R=5.605e+00 
R4743t540 n4744 n541 R=5.683e+00 
R4743t2640 n4744 n2641 R=3.369e+00 
R4744t4074 n4745 n4075 R=9.698e+01 
R4744t172 n4745 n173 R=1.008e+01 
R4744t718 n4745 n719 R=5.776e+01 
R4745t80 n4746 n81 R=5.868e+00 
R4746t1200 n4747 n1201 R=3.451e+00 
R4746t957 n4747 n958 R=2.218e+01 
R4746t4237 n4747 n4238 R=2.677e+01 
R4746t1637 n4747 n1638 R=8.688e+00 
R4747t1228 n4748 n1229 R=1.230e+01 
R4748t4024 n4749 n4025 R=1.460e+01 
R4748t2279 n4749 n2280 R=3.191e+00 
R4748t560 n4749 n561 R=1.254e+01 
R4749t23 n4750 n24 R=8.003e+00 
R4749t1013 n4750 n1014 R=1.423e+01 
R4749t1338 n4750 n1339 R=5.871e+00 
R4750t401 n4751 n402 R=5.364e+00 
R4750t2089 n4751 n2090 R=2.339e+00 
R4750t2719 n4751 n2720 R=4.861e+00 
R4750t3932 n4751 n3933 R=2.733e+01 
R4751t841 n4752 n842 R=1.658e+01 
R4751t2368 n4752 n2369 R=9.269e+00 
R4752t153 n4753 n154 R=1.855e+01 
R4753t1816 n4754 n1817 R=1.200e+01 
R4753t3741 n4754 n3742 R=1.174e+01 
R4754t4277 n4755 n4278 R=3.558e+00 
R4754t1063 n4755 n1064 R=4.997e+00 
R4755t1378 n4756 n1379 R=1.466e+01 
R4755t2976 n4756 n2977 R=7.022e+00 
R4755t3412 n4756 n3413 R=1.139e+01 
R4755t2867 n4756 n2868 R=3.436e+01 
R4755t4176 n4756 n4177 R=6.667e+00 
R4755t3155 n4756 n3156 R=3.742e+01 
R4756t2086 n4757 n2087 R=1.929e+01 
R4756t3081 n4757 n3082 R=6.932e+00 
R4756t3544 n4757 n3545 R=7.173e+01 
R4756t338 n4757 n339 R=4.229e+01 
R4756t1893 n4757 n1894 R=8.315e+00 
R4757t1089 n4758 n1090 R=1.351e+01 
R4757t90 n4758 n91 R=3.850e+01 
R4757t736 n4758 n737 R=6.745e+01 
R4758t4074 n4759 n4075 R=4.304e+01 
R4758t4331 n4759 n1 R=3.866e+00 
R4758t3437 n4759 n3438 R=5.325e+00 
R4759t3927 n4760 n3928 R=4.587e+00 
R4760t4411 n4761 n4412 R=6.494e+00 
R4760t1543 n4761 n1544 R=7.786e+01 
R4760t1348 n4761 n1349 R=2.771e+01 
R4760t4273 n4761 n4274 R=1.917e+01 
R4760t4692 n4761 n4693 R=4.878e+00 
R4761t2371 n4762 n2372 R=4.443e+00 
R4761t1671 n4762 n1672 R=4.570e+01 
R4761t3739 n4762 n3740 R=5.243e+00 
R4761t3453 n4762 n3454 R=2.393e+01 
R4762t2311 n4763 n2312 R=1.786e+01 
R4762t1205 n4763 n1206 R=1.010e+01 
R4763t136 n4764 n137 R=1.630e+01 
R4763t1331 n4764 n1332 R=4.975e+00 
R4763t3495 n4764 n3496 R=4.628e+00 
R4763t2077 n4764 n2078 R=4.818e+00 
R4764t3467 n4765 n3468 R=2.825e+00 
R4764t4360 n4765 n4361 R=1.035e+01 
R4764t2190 n4765 n2191 R=1.242e+01 
R4765t1732 n4766 n1733 R=2.598e+00 
R4766t3014 n4767 n3015 R=2.009e+00 
R4766t4485 n4767 n4486 R=1.978e+01 
R4766t309 n4767 n310 R=1.052e+01 
R4766t2044 n4767 n2045 R=2.823e+00 
R4766t4146 n4767 n4147 R=1.509e+02 
R4766t1521 n4767 n1522 R=1.852e+01 
R4767t4423 n4768 n4424 R=6.198e+01 
R4767t2567 n4768 n2568 R=6.491e+00 
R4768t3632 n4769 n3633 R=3.457e+01 
R4768t3923 n4769 n3924 R=1.458e+01 
R4768t2591 n4769 n2592 R=2.338e+01 
R4768t394 n4769 n395 R=3.858e+00 
R4768t3022 n4769 n3023 R=1.296e+01 
R4769t2425 n4770 n2426 R=2.706e+00 
R4770t4318 n4771 n4319 R=6.676e+00 
R4770t1344 n4771 n1345 R=3.402e+01 
R4770t740 n4771 n741 R=1.396e+02 
R4770t3850 n4771 n3851 R=4.147e+00 
R4770t2008 n4771 n2009 R=1.115e+01 
R4770t4701 n4771 n4702 R=6.203e+00 
R4771t4404 n4772 n4405 R=2.817e+00 
R4771t4504 n4772 n4505 R=1.624e+01 
R4772t3232 n4773 n3233 R=8.749e+00 
R4772t4189 n4773 n1 R=6.978e+01 
R4772t3435 n4773 n3436 R=2.744e+00 
R4773t3699 n4774 n3700 R=5.894e+00 
R4773t550 n4774 n551 R=8.091e+00 
R4773t373 n4774 n374 R=1.724e+01 
R4773t1253 n4774 n1254 R=3.730e+00 
R4774t806 n4775 n807 R=1.378e+01 
R4774t1224 n4775 n1225 R=2.347e+01 
R4774t433 n4775 n434 R=8.398e+00 
R4774t4082 n4775 n4083 R=1.416e+01 
R4774t4355 n4775 n4356 R=3.076e+00 
R4775t2475 n4776 n2476 R=1.115e+01 
R4775t1562 n4776 n1563 R=2.646e+01 
R4776t4590 n4777 n4591 R=1.888e+01 
R4776t4383 n4777 n4384 R=9.305e+01 
R4776t1757 n4777 n1758 R=5.685e+00 
R4777t4583 n4778 n4584 R=4.953e+00 
R4777t4310 n4778 n4311 R=7.427e+01 
R4779t198 n4780 n199 R=1.833e+01 
R4779t3787 n4780 n3788 R=2.084e+00 
R4781t1811 n4782 n1812 R=1.158e+01 
R4781t3956 n4782 n3957 R=2.992e+00 
R4782t4740 n4783 n4741 R=7.477e+00 
R4782t1651 n4783 n1652 R=3.221e+01 
R4783t3780 n4784 n3781 R=1.160e+02 
R4783t4377 n4784 n4378 R=1.942e+00 
R4783t4265 n4784 n4266 R=1.194e+01 
R4783t1980 n4784 n1981 R=5.622e+00 
R4783t1607 n4784 n1608 R=4.160e+00 
R4784t2 n4785 n3 R=1.932e+01 
R4784t4432 n4785 n4433 R=5.834e+02 
R4784t3086 n4785 n3087 R=1.273e+01 
R4784t2782 n4785 n2783 R=1.430e+01 
R4784t2908 n4785 n2909 R=1.881e+02 
R4785t777 n4786 n778 R=2.806e+00 
R4785t1509 n4786 n1510 R=2.217e+03 
R4786t1404 n4787 n1405 R=3.580e+01 
R4787t46 n4788 n47 R=6.966e+00 
R4787t289 n4788 n290 R=3.106e+00 
R4787t2996 n4788 n2997 R=1.077e+01 
R4787t1559 n4788 n1560 R=1.123e+01 
R4787t3781 n4788 n3782 R=1.067e+01 
R4788t444 n4789 n445 R=1.154e+01 
R4788t779 n4789 n780 R=1.355e+01 
R4788t632 n4789 n633 R=9.339e+00 
R4788t508 n4789 n509 R=1.171e+01 
R4788t2454 n4789 n2455 R=4.211e+00 
R4788t4217 n4789 n4218 R=1.535e+01 
R4789t3176 n4790 n3177 R=8.521e+00 
R4789t4537 n4790 n4538 R=4.523e+00 
R4789t2232 n4790 n2233 R=1.948e+01 
R4790t2988 n4791 n2989 R=1.849e+01 
R4790t3802 n4791 n3803 R=7.518e+00 
R4790t4677 n4791 n4678 R=2.302e+01 
R4790t2817 n4791 n2818 R=4.323e+01 
R4791t580 n4792 n581 R=1.513e+01 
R4791t852 n4792 n853 R=5.999e+02 
R4791t1476 n4792 n1477 R=2.759e+00 
R4791t1658 n4792 n1659 R=5.225e+00 
R4791t1239 n4792 n1240 R=3.294e+00 
R4792t573 n4793 n574 R=1.565e+01 
R4792t1612 n4793 n1613 R=3.234e+00 
R4793t3113 n4794 n3114 R=9.125e+00 
R4793t1649 n4794 n1650 R=3.961e+00 
R4793t4374 n4794 n4375 R=1.488e+01 
R4794t1627 n4795 n1628 R=2.527e+00 
R4794t1240 n4795 n1241 R=1.159e+01 
R4795t2941 n4796 n2942 R=3.074e+00 
R4795t3917 n4796 n3918 R=8.780e+00 
R4796t2756 n4797 n2757 R=2.807e+00 
R4797t2977 n4798 n2978 R=5.275e+00 
R4797t3255 n4798 n3256 R=1.123e+01 
R4797t3708 n4798 n3709 R=1.098e+01 
R4797t682 n4798 n683 R=4.165e+00 
R4797t4290 n4798 n4291 R=5.676e+00 
R4797t4487 n4798 n4488 R=9.838e+01 
R4798t4103 n4799 n4104 R=1.930e+00 
R4798t4383 n4799 n4384 R=1.847e+01 
R4798t1270 n4799 n1271 R=4.819e+01 
R4798t902 n4799 n903 R=2.829e+00 
R4799t3273 n4800 n3274 R=1.038e+01 
R4800t1099 n4801 n1100 R=1.536e+01 
R4800t3017 n4801 n3018 R=8.615e+00 
R4800t2325 n4801 n2326 R=1.464e+01 
R4800t3887 n4801 n3888 R=1.422e+01 
R4801t254 n4802 n255 R=1.130e+01 
R4801t4560 n4802 n4561 R=1.186e+01 
R4801t243 n4802 n244 R=7.157e+00 
R4801t2581 n4802 n2582 R=2.120e+02 
R4801t678 n4802 n679 R=3.409e+01 
R4801t3442 n4802 n3443 R=3.275e+00 
R4801t4162 n4802 n4163 R=1.110e+02 
R4802t689 n4803 n690 R=1.364e+01 
R4802t2856 n4803 n2857 R=1.107e+01 
R4802t1222 n4803 n1223 R=1.678e+01 
R4803t4118 n4804 n4119 R=1.387e+01 
R4803t930 n4804 n931 R=4.232e+00 
R4803t2833 n4804 n2834 R=8.371e+00 
R4803t1380 n4804 n1381 R=2.685e+01 
R4804t4451 n4805 n4452 R=1.181e+01 
R4804t3623 n4805 n3624 R=9.253e+00 
R4804t4100 n4805 n4101 R=6.323e+00 
R4805t2841 n4806 n2842 R=1.093e+01 
R4805t3742 n4806 n3743 R=9.086e+00 
R4805t4389 n4806 n4390 R=3.465e+00 
R4805t4392 n4806 n4393 R=1.827e+01 
R4805t3491 n4806 n3492 R=9.886e+00 
R4805t603 n4806 n604 R=3.112e+00 
R4806t985 n4807 n986 R=1.152e+01 
R4806t3444 n4807 n3445 R=1.393e+01 
R4806t1589 n4807 n1590 R=3.685e+00 
R4808t3761 n4809 n3762 R=4.454e+00 
R4808t1180 n4809 n1181 R=2.865e+00 
R4808t3709 n4809 n3710 R=2.956e+01 
R4810t1821 n4811 n1822 R=1.491e+01 
R4810t144 n4811 n145 R=2.900e+00 
R4810t780 n4811 n781 R=1.803e+01 
R4811t423 n4812 n424 R=1.652e+01 
R4812t444 n4813 n445 R=1.904e+01 
R4812t779 n4813 n780 R=5.520e+00 
R4812t1083 n4813 n1084 R=8.110e+00 
R4812t1791 n4813 n1792 R=3.938e+00 
R4813t689 n4814 n690 R=5.116e+00 
R4813t4802 n4814 n4803 R=1.990e+01 
R4813t2856 n4814 n2857 R=2.849e+00 
R4813t708 n4814 n709 R=4.499e+00 
R4814t877 n4815 n878 R=9.079e+00 
R4814t894 n4815 n895 R=1.126e+01 
R4814t3612 n4815 n3613 R=2.329e+01 
R4814t3524 n4815 n3525 R=5.244e+01 
R4815t2693 n4816 n2694 R=6.587e+00 
R4815t4555 n4816 n4556 R=5.614e+00 
R4816t52 n4817 n53 R=9.241e+00 
R4816t823 n4817 n824 R=6.400e+00 
R4817t3292 n4818 n3293 R=7.286e+00 
R4817t4608 n4818 n4609 R=7.409e+00 
R4817t2944 n4818 n2945 R=5.005e+00 
R4818t3084 n4819 n3085 R=6.515e+01 
R4818t1600 n4819 n1601 R=1.557e+03 
R4819t1363 n4820 n1364 R=2.589e+01 
R4819t1587 n4820 n1588 R=3.737e+01 
R4820t86 n4821 n87 R=5.005e+00 
R4820t3543 n4821 n3544 R=1.317e+01 
R4820t3375 n4821 n3376 R=2.468e+00 
R4821t3331 n4822 n3332 R=6.772e+00 
R4821t3867 n4822 n3868 R=4.721e+00 
R4821t4336 n4822 n4337 R=6.568e+00 
R4821t404 n4822 n405 R=4.565e+01 
R4821t4430 n4822 n4431 R=3.577e+00 
R4822t590 n4823 n591 R=9.441e+01 
R4823t4765 n4824 n4766 R=2.747e+00 
R4823t1732 n4824 n1733 R=1.217e+02 
R4823t985 n4824 n986 R=2.647e+01 
R4823t251 n4824 n252 R=4.442e+00 
R4824t3116 n4825 n3117 R=4.194e+00 
R4824t3460 n4825 n3461 R=2.779e+01 
R4824t2068 n4825 n2069 R=4.883e+01 
R4824t1950 n4825 n1951 R=5.670e+00 
R4825t51 n4826 n52 R=2.859e+00 
R4826t4100 n4827 n4101 R=1.535e+02 
R4826t4131 n4827 n4132 R=2.326e+02 
R4826t3623 n4827 n3624 R=2.652e+01 
R4826t4333 n4827 n4334 R=2.684e+01 
R4826t1702 n4827 n1703 R=5.281e+00 
R4827t4427 n4828 n4428 R=6.492e+00 
R4827t1706 n4828 n1707 R=4.555e+00 
R4828t2759 n4829 n2760 R=2.373e+01 
R4828t1685 n4829 n1686 R=2.035e+02 
R4828t1575 n4829 n1576 R=2.274e+00 
R4828t2605 n4829 n2606 R=3.326e+01 
R4829t3471 n4830 n3472 R=1.620e+01 
R4829t1297 n4830 n1298 R=4.315e+00 
R4829t3346 n4830 n3347 R=5.482e+00 
R4829t3466 n4830 n3467 R=9.025e+01 
R4829t34 n4830 n35 R=1.929e+01 
R4830t4584 n4831 n4585 R=4.811e+00 
R4830t3268 n4831 n3269 R=1.257e+01 
R4831t579 n4832 n580 R=3.416e+01 
R4831t4393 n4832 n4394 R=2.344e+00 
R4831t414 n4832 n415 R=5.522e+00 
R4832t948 n4833 n949 R=4.446e+01 
R4832t4632 n4833 n4633 R=1.051e+01 
R4832t4555 n4833 n4556 R=5.445e+00 
R4832t4815 n4833 n4816 R=5.233e+00 
R4832t2693 n4833 n2694 R=1.655e+01 
R4833t1268 n4834 n1269 R=5.568e+00 
R4833t957 n4834 n958 R=2.070e+01 
R4833t351 n4834 n352 R=5.449e+00 
R4833t3232 n4834 n3233 R=7.080e+00 
R4835t1054 n4836 n1055 R=5.978e+00 
R4836t177 n4837 n178 R=2.790e+02 
R4836t2981 n4837 n2982 R=5.654e+00 
R4836t3639 n4837 n3640 R=2.467e+00 
R4836t3068 n4837 n3069 R=9.771e+01 
R4836t2877 n4837 n2878 R=1.639e+00 
R4837t1974 n4838 n1975 R=6.434e+00 
R4837t2845 n4838 n2846 R=8.001e+00 
R4837t2172 n4838 n2173 R=8.736e+01 
R4837t3284 n4838 n3285 R=3.882e+00 
R4838t602 n4839 n603 R=7.335e+00 
R4838t3664 n4839 n3665 R=3.432e+00 
R4838t3117 n4839 n3118 R=7.859e+00 
R4838t3083 n4839 n3084 R=3.743e+00 
R4839t1765 n4840 n1766 R=8.956e+00 
R4839t4008 n4840 n4009 R=1.266e+02 
R4839t1349 n4840 n1350 R=3.112e+01 
R4839t4080 n4840 n4081 R=6.951e+00 
R4839t1842 n4840 n1843 R=6.553e+00 
R4840t2021 n4841 n2022 R=9.309e+00 
R4840t4313 n4841 n4314 R=7.309e+01 
R4840t2909 n4841 n2910 R=2.612e+01 
R4840t1261 n4841 n1262 R=1.984e+02 
R4841t1287 n4842 n1288 R=1.294e+01 
R4841t2365 n4842 n2366 R=1.119e+01 
R4841t409 n4842 n410 R=4.744e+00 
R4842t2606 n4843 n2607 R=3.554e+01 
R4842t3429 n4843 n3430 R=3.568e+00 
R4842t2882 n4843 n2883 R=7.629e+00 
R4843t88 n4844 n89 R=2.903e+00 
R4843t817 n4844 n818 R=5.032e+00 
R4844t4686 n4845 n4687 R=4.588e+00 
R4844t4790 n4845 n4791 R=1.217e+01 
R4845t4289 n4846 n4290 R=2.727e+01 
R4846t812 n4847 n813 R=4.072e+01 
R4847t19 n4848 n20 R=1.401e+01 
R4847t2313 n4848 n2314 R=3.685e+00 
R4847t2824 n4848 n2825 R=1.306e+01 
R4848t1184 n4849 n1185 R=6.805e+00 
R4849t3406 n4850 n3407 R=7.528e+00 
R4850t412 n4851 n413 R=3.737e+00 
R4850t731 n4851 n732 R=5.349e+00 
R4850t3108 n4851 n3109 R=3.129e+00 
R4850t1308 n4851 n1309 R=6.656e+00 
R4851t1685 n4852 n1686 R=8.309e+00 
R4851t4828 n4852 n4829 R=2.181e+00 
R4851t2759 n4852 n2760 R=2.239e+01 
R4852t3023 n4853 n3024 R=1.039e+01 
R4852t2683 n4853 n2684 R=6.442e+00 
R4852t3849 n4853 n3850 R=1.137e+02 
R4853t727 n4854 n728 R=1.135e+02 
R4853t1458 n4854 n1459 R=7.703e+00 
R4853t2771 n4854 n2772 R=2.679e+01 
R4853t2304 n4854 n2305 R=1.020e+01 
R4854t986 n4855 n987 R=1.199e+01 
R4854t4002 n4855 n4003 R=4.119e+01 
R4855t4384 n4856 n4385 R=3.992e+00 
R4855t1404 n4856 n1405 R=8.267e+00 
R4855t4786 n4856 n4787 R=2.846e+00 
R4856t2145 n4857 n2146 R=2.579e+01 
R4856t3904 n4857 n3905 R=4.333e+01 
R4856t476 n4857 n477 R=8.293e+00 
R4856t3596 n4857 n3597 R=1.286e+01 
R4856t2508 n4857 n2509 R=3.514e+02 
R4856t1353 n4857 n1354 R=1.766e+02 
R4856t920 n4857 n921 R=2.440e+00 
R4857t1304 n4858 n1305 R=1.348e+01 
R4857t2969 n4858 n2970 R=1.759e+01 
R4857t2634 n4858 n2635 R=5.960e+00 
R4857t4020 n4858 n4021 R=1.761e+01 
R4857t4022 n4858 n4023 R=6.757e+00 
R4858t1470 n4859 n1471 R=5.356e+02 
R4858t2516 n4859 n2517 R=5.923e+00 
R4858t3450 n4859 n3451 R=2.133e+01 
R4859t3900 n4860 n3901 R=3.436e+00 
R4859t709 n4860 n710 R=1.523e+01 
R4860t3200 n4861 n3201 R=4.645e+02 
R4860t3104 n4861 n3105 R=4.536e+00 
R4860t3557 n4861 n3558 R=5.705e+00 
R4861t4404 n4862 n4405 R=1.986e+00 
R4861t2121 n4862 n2122 R=5.395e+00 
R4861t2522 n4862 n2523 R=1.726e+01 
R4862t4404 n4863 n4405 R=5.958e+00 
R4862t4771 n4863 n4772 R=2.199e+01 
R4862t2522 n4863 n2523 R=8.752e+00 
R4863t3312 n4864 n3313 R=7.042e+00 
R4863t4544 n4864 n4545 R=1.069e+01 
R4863t4005 n4864 n4006 R=6.271e+00 
R4863t4414 n4864 n4415 R=1.470e+01 
R4864t4089 n4865 n4090 R=2.086e+00 
R4864t2574 n4865 n2575 R=1.323e+02 
R4864t2230 n4865 n2231 R=4.614e+01 
R4864t1289 n4865 n1290 R=2.188e+00 
R4864t1681 n4865 n1682 R=9.098e+00 
R4865t2055 n4866 n2056 R=5.605e+01 
R4865t4446 n4866 n4447 R=2.729e+00 
R4865t250 n4866 n251 R=1.164e+01 
R4865t3729 n4866 n3730 R=4.501e+00 
R4865t1705 n4866 n1706 R=1.297e+01 
R4866t2288 n4867 n2289 R=1.173e+01 
R4866t3533 n4867 n3534 R=8.658e+00 
R4866t237 n4867 n238 R=1.521e+02 
R4866t4151 n4867 n4152 R=5.321e+00 
R4866t1138 n4867 n1139 R=1.638e+01 
R4867t3061 n4868 n3062 R=2.438e+01 
R4868t2722 n4869 n2723 R=2.012e+01 
R4868t3667 n4869 n3668 R=5.083e+00 
R4869t2975 n4870 n2976 R=3.025e+00 
R4869t3860 n4870 n3861 R=2.483e+00 
R4870t4642 n4871 n4643 R=2.291e+00 
R4870t4510 n4871 n4511 R=1.915e+01 
R4871t2611 n4872 n2612 R=9.641e+00 
R4872t643 n4873 n644 R=1.768e+02 
R4872t3118 n4873 n3119 R=2.986e+00 
R4872t1785 n4873 n1786 R=6.689e+00 
R4872t2950 n4873 n2951 R=2.376e+01 
R4872t2071 n4873 n2072 R=6.047e+00 
R4873t262 n4874 n263 R=1.894e+00 
R4873t4157 n4874 n4158 R=1.445e+01 
R4874t2429 n4875 n2430 R=1.900e+00 
R4874t1160 n4875 n1161 R=2.597e+00 
R4874t2324 n4875 n2325 R=3.020e+01 
R4875t4457 n4876 n4458 R=1.569e+01 
R4875t4717 n4876 n4718 R=2.577e+02 
R4875t2872 n4876 n2873 R=7.185e+01 
R4875t3869 n4876 n3870 R=3.770e+01 
R4875t1846 n4876 n1847 R=3.070e+00 
R4876t2620 n4877 n2621 R=1.471e+01 
R4876t1719 n4877 n1720 R=8.997e+00 
R4876t3930 n4877 n3931 R=4.434e+00 
R4876t811 n4877 n812 R=5.447e+00 
R4876t3577 n4877 n3578 R=2.568e+01 
R4877t1991 n4878 n1992 R=1.064e+01 
R4877t1033 n4878 n1034 R=3.392e+00 
R4877t4325 n4878 n4326 R=6.763e+01 
R4878t3127 n4879 n3128 R=2.656e+01 
R4878t2630 n4879 n2631 R=3.292e+01 
R4878t1904 n4879 n1905 R=7.917e+00 
R4878t3563 n4879 n3564 R=5.220e+00 
R4879t4074 n4880 n4075 R=5.919e+00 
R4879t4744 n4880 n4745 R=2.899e+00 
R4880t1118 n4881 n1119 R=9.272e+00 
R4881t4698 n4882 n4699 R=5.013e+00 
R4881t1184 n4882 n1185 R=2.883e+01 
R4882t2891 n4883 n2892 R=4.476e+01 
R4882t2324 n4883 n2325 R=1.299e+01 
R4882t862 n4883 n863 R=1.555e+01 
R4883t4873 n4884 n4874 R=6.357e+00 
R4883t4425 n4884 n4426 R=3.102e+00 
R4883t4215 n4884 n4216 R=7.313e+00 
R4884t1994 n4885 n1995 R=4.631e+00 
R4884t3206 n4885 n3207 R=3.591e+00 
R4884t1175 n4885 n1176 R=3.025e+02 
R4885t3412 n4886 n3413 R=3.574e+00 
R4885t3555 n4886 n3556 R=2.980e+00 
R4886t2886 n4887 n2887 R=3.799e+01 
R4886t3769 n4887 n3770 R=4.098e+00 
R4886t1745 n4887 n1746 R=6.216e+01 
R4887t2556 n4888 n2557 R=3.396e+00 
R4887t2897 n4888 n2898 R=1.719e+01 
R4888t2075 n4889 n2076 R=6.381e+00 
R4888t3264 n4889 n3265 R=3.322e+01 
R4888t210 n4889 n211 R=8.947e+00 
R4888t4522 n4889 n4523 R=3.465e+00 
R4889t774 n4890 n775 R=3.325e+00 
R4889t2481 n4890 n2482 R=4.816e+01 
R4890t3847 n4891 n3848 R=4.292e+00 
R4891t2092 n4892 n2093 R=3.777e+00 
R4891t2688 n4892 n2689 R=1.848e+01 
R4891t125 n4892 n126 R=9.486e+00 
R4891t1858 n4892 n1859 R=1.391e+01 
R4892t2758 n4893 n2759 R=2.564e+00 
R4892t3299 n4893 n3300 R=3.602e+00 
R4892t2819 n4893 n2820 R=3.413e+00 
R4893t2494 n4894 n2495 R=8.690e+00 
R4893t79 n4894 n80 R=6.715e+00 
R4894t875 n4895 n876 R=1.698e+01 
R4894t2729 n4895 n2730 R=2.115e+00 
R4894t826 n4895 n827 R=1.337e+01 
R4895t4461 n4896 n4462 R=4.702e+00 
R4895t627 n4896 n628 R=7.406e+00 
R4895t292 n4896 n293 R=5.022e+00 
R4896t378 n4897 n379 R=2.440e+00 
R4896t272 n4897 n273 R=1.698e+01 
R4896t584 n4897 n585 R=2.374e+00 
R4896t1424 n4897 n1425 R=3.059e+01 
R4897t4312 n4898 n4313 R=1.736e+02 
R4897t4468 n4898 n4469 R=4.232e+00 
R4897t1781 n4898 n1782 R=8.881e+01 
R4897t2904 n4898 n2905 R=9.165e+00 
R4897t2582 n4898 n2583 R=1.049e+01 
R4898t1818 n4899 n1819 R=3.051e+00 
R4899t3243 n4900 n3244 R=1.924e+01 
R4899t2716 n4900 n2717 R=1.598e+01 
R4899t1012 n4900 n1013 R=2.408e+00 
R4900t2766 n4901 n2767 R=4.472e+00 
R4900t2539 n4901 n2540 R=3.985e+00 
R4901t2457 n4902 n2458 R=2.570e+00 
R4901t2299 n4902 n2300 R=3.170e+01 
R4901t3047 n4902 n3048 R=1.424e+01 
R4901t4435 n4902 n4436 R=3.384e+00 
R4902t3334 n4903 n3335 R=7.971e+00 
R4903t4270 n4904 n4271 R=7.365e+00 
R4903t4580 n4904 n4581 R=3.401e+01 
R4903t424 n4904 n425 R=1.849e+01 
R4904t3511 n4905 n3512 R=8.599e+00 
R4905t2536 n4906 n2537 R=1.986e+01 
R4905t2717 n4906 n2718 R=8.104e+00 
R4906t2646 n4907 n2647 R=3.932e+00 
R4906t188 n4907 n189 R=8.632e+00 
R4906t656 n4907 n657 R=3.363e+00 
R4907t4047 n4908 n4048 R=7.623e+00 
R4908t3440 n4909 n3441 R=1.004e+01 
R4908t1834 n4909 n1835 R=1.117e+01 
R4908t3417 n4909 n3418 R=3.140e+00 
R4909t1238 n4910 n1239 R=2.119e+00 
R4909t3096 n4910 n3097 R=1.382e+01 
R4909t3048 n4910 n3049 R=6.221e+00 
R4910t1189 n4911 n1190 R=3.998e+00 
R4910t2448 n4911 n2449 R=5.264e+00 
R4910t137 n4911 n138 R=2.234e+01 
R4910t2379 n4911 n2380 R=6.186e+00 
R4911t3604 n4912 n3605 R=7.008e+00 
R4912t4342 n4913 n4343 R=4.641e+01 
R4912t481 n4913 n482 R=5.104e+00 
R4912t1977 n4913 n1978 R=9.157e+00 
R4912t1481 n4913 n1482 R=2.378e+01 
R4912t1849 n4913 n1850 R=3.406e+02 
R4912t2973 n4913 n2974 R=4.528e+00 
R4913t2708 n4914 n2709 R=3.501e+00 
R4913t281 n4914 n282 R=1.696e+01 
R4913t1660 n4914 n1661 R=9.816e+00 
R4915t465 n4916 n466 R=1.106e+01 
R4915t1494 n4916 n1495 R=7.652e+00 
R4916t4453 n4917 n4454 R=1.262e+01 
R4916t4455 n4917 n4456 R=5.526e+00 
R4916t32 n4917 n33 R=5.043e+01 
R4916t4201 n4917 n4202 R=2.985e+01 
R4917t69 n4918 n70 R=1.270e+01 
R4917t4238 n4918 n4239 R=4.241e+00 
R4917t1600 n4918 n1601 R=1.499e+01 
R4918t453 n4919 n454 R=2.381e+01 
R4918t3845 n4919 n3846 R=2.112e+01 
R4918t1908 n4919 n1909 R=1.093e+01 
R4919t1376 n1 n1377 R=5.910e+00 
R4920t4025 n4921 n4026 R=5.435e+00 
R4920t1065 n4921 n1066 R=3.908e+00 
R4921t688 n4922 n689 R=6.932e+00 
R4921t3812 n4922 n3813 R=1.297e+01 
R4922t404 n4923 n405 R=3.397e+01 
R4922t4430 n4923 n4431 R=3.301e+00 
R4923t916 n4924 n917 R=1.966e+01 
R4923t2552 n4924 n2553 R=5.281e+00 
R4923t4223 n4924 n4224 R=1.538e+02 
R4923t4359 n4924 n4360 R=6.550e+00 
R4923t3646 n4924 n3647 R=5.256e+00 
R4923t4334 n4924 n4335 R=3.961e+00 
R4923t4123 n4924 n4124 R=1.679e+01 
R4924t4266 n4925 n4267 R=3.591e+00 
R4925t3904 n4926 n3905 R=4.329e+00 
R4925t920 n4926 n921 R=8.642e+00 
R4925t3943 n4926 n3944 R=8.891e+00 
R4925t3900 n4926 n3901 R=1.341e+01 
R4925t4859 n4926 n4860 R=2.033e+01 
R4926t3477 n4927 n3478 R=8.488e+00 
R4926t4018 n4927 n4019 R=3.690e+00 
R4926t2728 n4927 n2729 R=2.973e+02 
R4926t166 n4927 n167 R=4.575e+00 
R4926t1578 n4927 n1579 R=6.754e+00 
R4926t312 n4927 n313 R=1.825e+01 
R4927t3283 n4928 n3284 R=3.324e+00 
R4927t2846 n4928 n2847 R=1.911e+01 
R4927t295 n4928 n296 R=3.967e+01 
R4928t1080 n4929 n1081 R=2.486e+00 
R4928t1057 n4929 n1058 R=6.758e+00 
R4928t3241 n4929 n3242 R=6.132e+00 
R4928t3063 n4929 n3064 R=3.609e+01 
R4929t59 n4930 n60 R=4.228e+00 
R4929t1405 n4930 n1406 R=3.590e+01 
R4929t463 n4930 n464 R=1.014e+01 
R4929t275 n4930 n276 R=3.919e+00 
R4930t2310 n4931 n2311 R=2.416e+02 
R4930t4717 n4931 n4718 R=1.037e+02 
R4930t2460 n4931 n2461 R=1.193e+01 
R4930t2971 n4931 n2972 R=1.350e+01 
R4931t2566 n4932 n2567 R=5.053e+00 
R4931t4251 n4932 n4252 R=5.078e+00 
R4931t2341 n4932 n2342 R=4.718e+01 
R4931t2883 n4932 n2884 R=1.081e+01 
R4933t790 n4934 n791 R=1.688e+01 
R4933t4316 n4934 n4317 R=6.569e+00 
R4933t4242 n4934 n4243 R=9.139e+00 
R4934t4752 n4935 n4753 R=5.471e+00 
R4935t1463 n4936 n1464 R=5.863e+00 
R4935t2001 n4936 n2002 R=1.770e+01 
R4935t3680 n4936 n3681 R=1.169e+01 
R4935t996 n4936 n997 R=2.244e+01 
R4935t4665 n4936 n4666 R=7.264e+00 
R4936t649 n4937 n650 R=1.167e+01 
R4936t3204 n4937 n3205 R=1.955e+01 
R4936t404 n4937 n405 R=2.103e+01 
R4936t4922 n4937 n4923 R=2.620e+00 
R4937t3385 n4938 n3386 R=7.645e+00 
R4937t1165 n4938 n1166 R=1.836e+02 
R4937t184 n4938 n185 R=1.210e+01 
R4938t2264 n4939 n2265 R=1.831e+01 
R4938t2889 n4939 n2890 R=1.343e+02 
R4938t2998 n4939 n2999 R=9.550e+00 
R4939t2014 n4940 n2015 R=3.173e+00 
R4939t3817 n4940 n3818 R=1.788e+02 
R4939t2112 n4940 n2113 R=1.245e+01 
R4940t2290 n4941 n2291 R=7.225e+00 
R4940t3659 n4941 n3660 R=1.865e+02 
R4940t4378 n4941 n4379 R=6.988e+01 
R4940t617 n4941 n618 R=5.533e+00 
R4941t987 n4942 n988 R=6.254e+01 
R4941t3542 n4942 n3543 R=1.736e+01 
R4941t3847 n4942 n3848 R=7.987e+00 
R4941t3452 n4942 n3453 R=1.298e+01 
R4942t2321 n4943 n2322 R=6.681e+00 
R4942t2805 n4943 n2806 R=3.060e+00 
R4942t4639 n4943 n4640 R=1.426e+01 
R4942t3634 n4943 n3635 R=2.644e+02 
R4943t1535 n4944 n1536 R=4.340e+00 
R4943t2186 n4944 n2187 R=3.313e+00 
R4944t4417 n4945 n4418 R=3.160e+00 
R4945t1675 n4946 n1676 R=1.817e+01 
R4945t655 n4946 n656 R=8.837e-01 
R4946t4794 n4947 n4795 R=1.552e+01 
R4946t1627 n4947 n1628 R=4.656e+00 
R4946t3260 n4947 n3261 R=2.996e+01 
R4946t4600 n4947 n4601 R=3.110e+00 
R4948t973 n4949 n974 R=2.609e+01 
R4948t2403 n4949 n2404 R=3.377e+00 
R4949t2223 n4950 n2224 R=3.591e+00 
R4949t3588 n4950 n3589 R=5.954e+01 
R4949t3864 n4950 n3865 R=4.694e+01 
R4950t2885 n4951 n2886 R=5.827e+00 
R4950t2131 n4951 n2132 R=2.259e+01 
R4951t4231 n4952 n4232 R=3.256e+00 
R4951t4848 n4952 n4849 R=2.148e+01 
R4952t3649 n4953 n3650 R=7.692e+01 
R4952t2644 n4953 n2645 R=3.587e+01 
R4953t3682 n4954 n3683 R=2.750e+01 
R4953t3755 n4954 n3756 R=5.890e+00 
R4953t4221 n4954 n4222 R=8.068e+00 
R4954t78 n4955 n79 R=1.396e+01 
R4954t3393 n4955 n3394 R=6.622e+00 
R4954t4388 n4955 n4389 R=8.012e+00 
R4954t256 n4955 n257 R=3.936e+00 
R4954t4398 n4955 n4399 R=9.581e+00 
R4955t1483 n4956 n1484 R=1.794e+00 
R4955t4029 n4956 n4030 R=7.957e+00 
R4955t1843 n4956 n1844 R=1.801e+01 
R4955t2834 n4956 n2835 R=4.482e+00 
R4956t3596 n4957 n3597 R=1.719e+01 
R4956t4856 n4957 n4857 R=5.248e+00 
R4956t476 n4957 n477 R=5.333e+01 
R4956t3650 n4957 n3651 R=4.138e+01 
R4957t2586 n4958 n2587 R=2.287e+01 
R4957t4593 n4958 n4594 R=7.216e+00 
R4957t2855 n4958 n2856 R=1.088e+02 
R4957t2101 n4958 n2102 R=4.155e+01 
R4957t14 n4958 n15 R=3.452e+00 
R4958t1462 n4959 n1463 R=3.819e+00 
R4958t4366 n4959 n4367 R=6.557e+01 
R4958t2118 n4959 n2119 R=1.024e+01 
R4958t4166 n4959 n4167 R=1.664e+01 
R4958t132 n4959 n133 R=5.805e+00 
R4959t2282 n4960 n2283 R=1.782e+00 
R4959t1972 n4960 n1973 R=8.328e+00 
R4959t2136 n4960 n2137 R=4.784e+00 
R4959t2208 n4960 n2209 R=5.362e+01 
R4960t1347 n4961 n1348 R=8.842e+00 
R4960t3355 n4961 n3356 R=4.954e+00 
R4960t1319 n4961 n1320 R=1.364e+01 
R4961t3218 n4962 n3219 R=2.209e+01 
R4961t2295 n4962 n2296 R=2.775e+01 
R4961t2699 n4962 n2700 R=5.134e+00 
R4961t4440 n4962 n4441 R=3.622e+00 
R4962t2292 n4963 n2293 R=2.436e+00 
R4962t106 n4963 n107 R=5.125e+01 
R4962t3236 n4963 n3237 R=9.749e+01 
R4963t4004 n4964 n4005 R=5.875e+01 
R4963t2554 n4964 n2555 R=3.136e+01 
R4963t119 n4964 n120 R=1.138e+01 
R4963t1151 n4964 n1152 R=9.270e+00 
R4963t3493 n4964 n3494 R=1.317e+01 
R4964t4323 n4965 n4324 R=3.307e+00 
R4964t1478 n4965 n1479 R=5.086e+00 
R4965t1812 n4966 n1813 R=3.036e+02 
R4965t4515 n4966 n4516 R=1.499e+00 
R4965t943 n4966 n944 R=6.556e+00 
R4965t4102 n4966 n4103 R=4.486e+01 
R4965t3614 n4966 n3615 R=2.064e+00 
R4966t3289 n4967 n3290 R=2.857e+00 
R4967t1610 n4968 n1611 R=4.411e+00 
R4967t3664 n4968 n3665 R=4.162e+00 
R4968t3310 n4969 n3311 R=8.267e+00 
R4968t381 n4969 n382 R=3.535e+00 
R4968t2512 n4969 n2513 R=3.652e+00 
R4969t4862 n4970 n4863 R=3.978e+00 
R4969t2522 n4970 n2523 R=5.577e+00 
R4969t3924 n4970 n3925 R=1.496e+01 
R4970t162 n4971 n163 R=1.683e+01 
R4970t1772 n4971 n1773 R=6.166e+00 
R4970t2751 n4971 n2752 R=4.457e+00 
R4970t2679 n4971 n2680 R=4.474e+00 
R4971t3747 n4972 n3748 R=3.467e+01 
R4971t4477 n4972 n4478 R=7.172e+00 
R4971t2674 n4972 n2675 R=7.843e+00 
R4971t2473 n4972 n2474 R=2.068e+00 
R4972t2361 n4973 n2362 R=4.144e+01 
R4972t4532 n4973 n4533 R=4.065e+00 
R4972t2626 n4973 n2627 R=1.311e+01 
R4973t3857 n4974 n3858 R=3.953e+00 
R4973t887 n4974 n888 R=2.533e+01 
R4973t3328 n4974 n3329 R=9.094e+00 
R4974t1381 n4975 n1382 R=1.271e+01 
R4974t1935 n4975 n1936 R=1.893e+01 
R4975t174 n4976 n1 R=4.843e+00 
R4975t1322 n4976 n1 R=1.004e+01 
R4975t3236 n4976 n3237 R=7.967e+00 
R4975t1727 n4976 n1 R=4.905e+00 
R4976t3234 n4977 n3235 R=2.684e+01 
R4976t3651 n4977 n3652 R=4.259e+00 
R4976t1076 n4977 n1077 R=3.687e+00 
R4976t2575 n4977 n2576 R=1.517e+01 
R4977t874 n4978 n875 R=1.995e+01 
R4977t1496 n4978 n1497 R=6.149e+01 
R4977t1845 n4978 n1846 R=2.189e+01 
R4977t3211 n4978 n3212 R=2.192e+01 
R4978t2251 n4979 n2252 R=3.879e+00 
R4978t2785 n4979 n2786 R=3.263e+01 
R4978t4809 n4979 n4810 R=2.631e+00 
R4979t832 n4980 n833 R=1.103e+02 
R4979t2731 n4980 n2732 R=5.844e+01 
R4979t3438 n4980 n3439 R=3.439e+00 
R4980t3539 n4981 n3540 R=2.558e+00 
R4980t677 n4981 n678 R=5.027e+00 
R4981t4104 n4982 n4105 R=1.916e+01 
R4981t2871 n4982 n2872 R=1.031e+01 
R4981t2538 n4982 n2539 R=1.996e+01 
R4981t371 n4982 n372 R=7.124e+00 
R4981t3152 n4982 n3153 R=1.227e+01 
R4981t2740 n4982 n2741 R=3.279e+00 
R4982t1161 n4983 n1162 R=2.856e+02 
R4982t1728 n4983 n1729 R=6.844e+01 
R4982t2356 n4983 n2357 R=4.223e+00 
R4982t2387 n4983 n2388 R=6.774e+00 
R4982t706 n4983 n707 R=3.243e+01 
R4983t1192 n4984 n1193 R=6.767e+00 
R4983t1630 n4984 n1631 R=9.019e+00 
R4983t4585 n4984 n4586 R=6.412e+00 
R4984t1177 n4985 n1178 R=1.170e+01 
R4984t3337 n4985 n3338 R=3.468e+00 
R4985t1720 n4986 n1721 R=1.098e+01 
R4985t2104 n4986 n2105 R=1.695e+01 
R4986t4069 n4987 n4070 R=5.463e+00 
R4986t903 n4987 n904 R=1.192e+01 
R4986t4223 n4987 n4224 R=2.852e+00 
R4987t3347 n4988 n3348 R=2.128e+01 
R4987t2726 n4988 n2727 R=6.569e+00 
R4987t1621 n4988 n1622 R=8.093e+00 
R4987t1166 n4988 n1167 R=6.387e+00 
R4988t1712 n4989 n1713 R=1.383e+01 
R4988t2498 n4989 n2499 R=2.765e+00 
R4989t71 n4990 n72 R=4.796e+00 
R4989t1380 n4990 n1381 R=3.289e+02 
R4989t4803 n4990 n4804 R=3.482e+00 
R4989t4118 n4990 n4119 R=2.691e+00 
R4989t4067 n4990 n4068 R=5.088e+01 
R4990t2756 n4991 n2757 R=9.681e+01 
R4990t4711 n4991 n4712 R=2.578e+01 
R4990t1198 n4991 n1199 R=1.911e+02 
R4990t3676 n4991 n3677 R=9.320e+00 
R4990t1764 n4991 n1765 R=3.925e+00 
R4991t3189 n4992 n3190 R=1.837e+01 
R4991t3798 n4992 n3799 R=2.414e+01 
R4991t3732 n4992 n3733 R=2.619e+00 
R4992t4367 n4993 n4368 R=1.491e+01 
R4992t2619 n4993 n2620 R=5.306e+00 
R4992t1381 n4993 n1382 R=4.444e+01 
R4993t175 n4994 n176 R=6.528e+00 
R4993t3490 n4994 n3491 R=3.127e+01 
R4993t7 n4994 n8 R=5.036e+00 
R4993t751 n4994 n752 R=7.032e+01 
R4994t1216 n4995 n1217 R=1.077e+01 
R4994t3584 n4995 n3585 R=1.613e+01 
R4994t354 n4995 n355 R=3.726e+00 
R4994t3903 n4995 n3904 R=2.680e+01 
R4995t3179 n4996 n3180 R=1.081e+01 
R4995t2749 n4996 n2750 R=2.137e+01 
R4996t2417 n1 n2418 R=1.094e+01 
R4997t4570 n4998 n4571 R=1.599e+01 
R4997t4465 n4998 n4466 R=1.845e+01 
R4998t1997 n4999 n1998 R=1.622e+01 
R4998t3813 n4999 n3814 R=6.903e+01 
R4998t4444 n4999 n4445 R=3.286e+00 
R4999t534 n5000 n535 R=5.015e+00 
R4999t2183 n5000 n2184 R=2.819e+01 
R4999t185 n5000 n186 R=7.390e+00 
R5000t230 n5001 n231 R=5.290e+00 
R5000t2947 n5001 n2948 R=1.564e+01 
R5000t3153 n5001 n3154 R=1.628e+01 
R5001t3726 n5002 n3727 R=9.260e+00 
R5001t2337 n5002 n2338 R=9.077e+00 
R5001t4615 n5002 n4616 R=7.154e+00 
R5001t2760 n5002 n2761 R=5.039e+00 
R5002t3398 n5003 n3399 R=3.708e+01 
R5002t700 n5003 n701 R=6.659e+00 
R5002t2555 n5003 n2556 R=6.420e+00 
R5003t4915 n5004 n4916 R=7.753e+00 
R5003t4203 n5004 n4204 R=1.949e+01 
R5003t4580 n5004 n4581 R=1.096e+01 
R5004t4199 n5005 n4200 R=8.057e+00 
R5004t2215 n5005 n2216 R=1.062e+01 
R5005t107 n5006 n108 R=1.679e+01 
R5005t4619 n5006 n4620 R=2.862e+00 
R5005t1199 n5006 n1200 R=2.783e+00 
R5005t2812 n5006 n2813 R=6.920e+01 
R5005t2878 n5006 n2879 R=1.169e+01 
R5006t3305 n5007 n3306 R=1.848e+01 
R5006t2070 n5007 n2071 R=7.214e+01 
R5006t2643 n5007 n2644 R=4.642e+00 
R5006t1186 n5007 n1187 R=9.635e+00 
R5006t530 n5007 n531 R=4.197e+00 
R5007t2593 n5008 n2594 R=9.870e+00 
R5007t3422 n5008 n3423 R=5.821e+00 
R5008t2346 n5009 n2347 R=1.865e+00 
R5008t3538 n5009 n3539 R=4.517e+01 
R5008t651 n5009 n652 R=2.475e+00 
R5008t1461 n5009 n1462 R=2.926e+01 
R5009t152 n5010 n153 R=3.876e+00 
R5009t1542 n5010 n1543 R=2.635e+01 
R5009t1495 n5010 n1496 R=8.895e+00 
R5009t3089 n5010 n3090 R=7.099e+00 
R5010t2430 n5011 n2431 R=5.624e+00 
R5010t3106 n5011 n3107 R=2.331e+01 
R5010t526 n5011 n527 R=3.750e+01 
R5010t4161 n5011 n4162 R=5.290e+00 
R5010t2048 n5011 n2049 R=2.123e+02 
R5011t3679 n5012 n3680 R=1.005e+01 
R5011t2113 n5012 n2114 R=4.344e+00 
R5011t3736 n5012 n3737 R=1.120e+01 
R5012t222 n5013 n223 R=1.319e+01 
R5012t1844 n5013 n1845 R=4.778e+00 
R5012t3469 n5013 n3470 R=6.709e+00 
R5012t2911 n5013 n2912 R=3.434e+00 
R5012t3412 n5013 n3413 R=3.258e+02 
R5013t1449 n5014 n1450 R=1.905e+01 
R5013t264 n5014 n265 R=3.444e+00 
R5013t4576 n5014 n4577 R=4.483e+00 
R5013t3207 n5014 n3208 R=1.934e+01 
R5013t1007 n5014 n1008 R=3.703e+00 
R5014t1391 n5015 n1392 R=7.936e+00 
R5014t1486 n5015 n1487 R=6.819e+00 
R5014t3599 n5015 n3600 R=3.795e+01 
R5015t1416 n5016 n1417 R=6.011e+00 
R5015t2906 n5016 n2907 R=7.156e+01 
R5016t4365 n5017 n4366 R=2.135e+01 
R5016t4376 n5017 n4377 R=9.122e+00 
R5016t1988 n5017 n1989 R=5.297e+00 
R5017t2146 n5018 n2147 R=1.629e+00 
R5017t4193 n5018 n4194 R=1.678e+01 
R5018t3388 n5019 n3389 R=3.246e+00 
R5018t1956 n5019 n1957 R=1.280e+02 
R5018t4186 n5019 n4187 R=3.051e+00 
R5018t1120 n5019 n1121 R=4.310e+01 
R5019t2919 n5020 n2920 R=7.542e+00 
R5019t115 n5020 n116 R=2.130e+01 
R5020t2990 n5021 n2991 R=7.991e+00 
R5020t1399 n5021 n1400 R=7.879e+01 
R5020t2531 n5021 n2532 R=3.319e+01 
R5020t130 n5021 n131 R=7.050e+00 
R5020t726 n5021 n727 R=4.502e+00 
R5021t4279 n5022 n4280 R=4.713e+00 
R5021t2806 n5022 n2807 R=3.853e+00 
R5022t2386 n5023 n2387 R=7.261e+00 
R5022t3884 n5023 n3885 R=6.569e+00 
R5022t430 n5023 n431 R=4.519e+00 
R5022t1546 n5023 n1547 R=3.945e+01 
R5022t3431 n5023 n3432 R=9.993e+00 
R5023t519 n5024 n520 R=5.175e+00 
R5024t1560 n5025 n1561 R=3.711e+00 
R5024t4019 n5025 n4020 R=1.104e+01 
R5024t3755 n5025 n3756 R=6.367e+00 
R5024t4953 n5025 n4954 R=6.324e+00 
R5024t3682 n5025 n3683 R=1.022e+02 
R5025t111 n5026 n112 R=2.786e+00 
R5026t4871 n5027 n4872 R=3.415e+00 
R5026t3354 n5027 n3355 R=1.789e+01 
R5027t770 n5028 n771 R=5.632e+00 
R5027t2335 n5028 n2336 R=5.432e+01 
R5027t3023 n5028 n3024 R=4.167e+00 
R5027t3689 n5028 n3690 R=7.097e+00 
R5028t784 n5029 n785 R=1.250e+01 
R5028t1602 n5029 n1603 R=1.834e+01 
R5028t3980 n5029 n3981 R=5.971e+00 
R5029t4218 n5030 n4219 R=1.774e+01 
R5029t4081 n5030 n4082 R=4.018e+00 
R5030t3914 n5031 n3915 R=1.035e+01 
R5030t3152 n5031 n3153 R=4.476e+00 
R5030t2740 n5031 n2741 R=5.526e+00 
R5031t1411 n5032 n1412 R=2.755e+00 
R5031t4282 n5032 n4283 R=7.138e+00 
R5031t2880 n5032 n2881 R=5.062e+00 
R5032t2659 n5033 n2660 R=4.154e+01 
R5033t290 n5034 n291 R=7.031e+00 
R5033t1238 n5034 n1239 R=3.380e+00 
R5033t3252 n5034 n3253 R=5.952e+00 
R5033t1340 n5034 n1341 R=1.350e+01 
R5034t118 n5035 n119 R=2.067e+01 
R5034t3515 n5035 n3516 R=1.144e+01 
R5034t144 n5035 n145 R=1.500e+01 
R5034t4810 n5035 n4811 R=3.286e+01 
R5034t1821 n5035 n1822 R=5.421e+00 
R5035t450 n5036 n451 R=4.527e+00 
R5035t3918 n5036 n3919 R=3.036e+01 
R5036t997 n5037 n998 R=3.588e+00 
R5036t80 n5037 n81 R=1.295e+02 
R5037t346 n5038 n347 R=4.536e+00 
R5037t4721 n5038 n4722 R=6.825e+00 
R5037t1240 n5038 n1241 R=6.618e+00 
R5037t4443 n5038 n4444 R=2.471e+00 
R5037t3734 n5038 n3735 R=2.788e+01 
R5038t179 n5039 n180 R=2.565e+00 
R5039t531 n5040 n532 R=9.019e+00 
R5039t2857 n5040 n2858 R=3.567e+01 
R5039t101 n5040 n102 R=1.637e+01 
R5040t1258 n5041 n1259 R=5.854e+00 
R5040t3240 n5041 n3241 R=1.018e+01 
R5040t1506 n5041 n1507 R=9.543e+00 
R5040t124 n5041 n125 R=3.484e+01 
R5041t718 n5042 n719 R=1.635e+01 
R5041t2459 n5042 n2460 R=9.256e+00 
R5041t1248 n5042 n1249 R=2.809e+00 
R5042t2648 n5043 n2649 R=2.621e+01 
R5042t910 n5043 n911 R=1.000e+01 
R5042t1851 n5043 n1852 R=5.860e+00 
R5042t3448 n5043 n3449 R=3.824e+00 
R5043t2162 n5044 n2163 R=1.344e+02 
R5043t2517 n5044 n2518 R=2.335e+00 
R5043t1740 n5044 n1741 R=9.947e+01 
R5043t2088 n5044 n2089 R=7.301e+00 
R5044t4752 n5045 n4753 R=5.675e+00 
R5044t153 n5045 n154 R=4.801e+00 
R5045t1544 n5046 n1545 R=3.004e+02 
R5045t3361 n5046 n3362 R=6.208e+00 
R5045t2712 n5046 n2713 R=4.834e+00 
R5046t1696 n5047 n1697 R=9.851e+00 
R5046t3339 n5047 n3340 R=2.412e+00 
R5047t3450 n5048 n3451 R=7.541e+00 
R5047t4099 n5048 n4100 R=8.826e+03 
R5047t3315 n5048 n3316 R=5.783e+00 
R5048t4157 n5049 n4158 R=6.234e+00 
R5048t3134 n5049 n3135 R=4.399e+00 
R5049t263 n5050 n264 R=7.283e+00 
R5049t3212 n5050 n3213 R=1.557e+01 
R5049t3237 n5050 n3238 R=1.607e+01 
R5049t702 n5050 n703 R=4.745e+00 
R5049t2363 n5050 n2364 R=1.929e+01 
R5050t1387 n5051 n1388 R=1.454e+01 
R5051t698 n5052 n699 R=5.688e+00 
R5051t3974 n5052 n3975 R=2.789e+00 
R5051t1094 n5052 n1095 R=6.607e+00 
R5052t1624 n5053 n1625 R=3.637e+01 
R5052t2854 n5053 n2855 R=1.112e+01 
R5052t4292 n5053 n4293 R=6.129e+00 
R5052t4319 n5053 n4320 R=3.682e+00 
R5053t4843 n5054 n4844 R=5.325e+00 
R5053t14 n5054 n15 R=1.393e+01 
R5053t817 n5054 n818 R=5.586e+00 
R5054t1896 n5055 n1897 R=4.284e+00 
R5054t4056 n5055 n4057 R=1.359e+01 
R5054t25 n5055 n26 R=5.900e+00 
R5055t1333 n5056 n1334 R=4.406e+01 
R5055t1685 n5056 n1686 R=5.859e+02 
R5055t1988 n5056 n1989 R=3.385e+00 
R5055t1032 n5056 n1033 R=6.233e+00 
R5056t3231 n5057 n3232 R=6.103e+00 
R5056t417 n5057 n418 R=1.370e+01 
R5056t3144 n5057 n3145 R=4.599e+01 
R5057t1706 n5058 n1707 R=5.567e+01 
R5057t4827 n5058 n4828 R=1.274e+01 
R5057t4427 n5058 n4428 R=5.955e+01 
R5057t1459 n5058 n1460 R=8.096e+00 
R5057t3766 n5058 n3767 R=1.211e+01 
R5058t744 n5059 n745 R=8.007e+00 
R5058t2631 n5059 n2632 R=8.385e+00 
R5059t1360 n5060 n1361 R=4.304e+00 
R5059t4128 n5060 n4129 R=8.502e+01 
R5060t3599 n5061 n3600 R=2.128e+00 
R5060t3969 n5061 n3970 R=1.996e+01 
R5060t5014 n5061 n5015 R=8.047e+00 
R5060t3773 n5061 n3774 R=1.626e+01 
R5060t4421 n5061 n4422 R=1.283e+01 
R5061t265 n5062 n266 R=6.181e+00 
R5061t1558 n5062 n1559 R=5.646e+00 
R5061t1684 n5062 n1685 R=5.153e+00 
R5062t1955 n5063 n1956 R=3.120e+00 
R5062t1049 n5063 n1050 R=2.415e+01 
R5062t2499 n5063 n2500 R=3.858e+01 
R5062t3836 n5063 n3837 R=1.423e+01 
R5062t4498 n5063 n4499 R=1.182e+01 
R5063t2990 n5064 n2991 R=4.230e+00 
R5063t3134 n5064 n3135 R=5.438e+01 
R5063t283 n5064 n284 R=2.802e+00 
R5064t3870 n5065 n3871 R=2.103e+01 
R5064t2894 n5065 n2895 R=2.119e+01 
R5064t2897 n5065 n2898 R=4.118e+00 
R5064t4887 n5065 n4888 R=4.834e+01 
R5065t2505 n5066 n2506 R=4.430e+00 
R5065t1080 n5066 n1081 R=1.166e+02 
R5065t4928 n5066 n4929 R=1.067e+01 
R5066t421 n5067 n422 R=4.918e+01 
R5066t1219 n5067 n1220 R=4.317e+01 
R5066t616 n5067 n617 R=2.614e+01 
R5067t2703 n5068 n2704 R=1.540e+01 
R5067t4258 n5068 n4259 R=1.352e+01 
R5067t2486 n5068 n2487 R=8.349e+00 
R5067t2160 n5068 n2161 R=1.354e+01 
R5068t1274 n5069 n1275 R=4.871e+00 
R5068t2221 n5069 n2222 R=2.490e+00 
R5068t4101 n5069 n4102 R=1.352e+01 
R5069t4366 n5070 n4367 R=4.764e+00 
R5069t4958 n5070 n4959 R=6.661e+00 
R5069t132 n5070 n133 R=3.888e+00 
R5070t3927 n5071 n3928 R=8.033e+00 
R5070t895 n5071 n896 R=9.134e+00 
R5071t446 n5072 n447 R=1.671e+01 
R5071t4299 n5072 n4300 R=2.328e+01 
R5071t4661 n5072 n4662 R=9.291e+00 
R5071t1800 n5072 n1801 R=9.249e+00 
R5071t1982 n5072 n1983 R=5.461e+01 
R5072t1721 n5073 n1722 R=1.041e+01 
R5072t4368 n5073 n4369 R=6.137e+00 
R5072t1576 n5073 n1577 R=2.478e+01 
R5073t1183 n5074 n1184 R=4.297e+00 
R5073t3239 n5074 n3240 R=3.910e+00 
R5074t3764 n5075 n3765 R=5.477e+00 
R5074t159 n5075 n160 R=2.465e+00 
R5075t541 n5076 n542 R=7.364e+00 
R5075t2573 n5076 n2574 R=5.035e+00 
R5075t859 n5076 n860 R=2.288e+01 
R5075t3321 n5076 n3322 R=9.923e+00 
R5075t1503 n5076 n1504 R=2.948e+00 
R5075t2011 n5076 n2012 R=2.255e+02 
R5076t1769 n5077 n1770 R=1.558e+01 
R5076t3456 n5077 n3457 R=9.525e+01 
R5077t1891 n5078 n1892 R=7.214e+01 
R5077t3270 n5078 n3271 R=3.390e+01 
R5077t2557 n5078 n2558 R=3.700e+00 
R5078t110 n5079 n111 R=5.603e+00 
R5078t4854 n5079 n4855 R=1.024e+01 
R5078t4002 n5079 n4003 R=4.025e+00 
R5079t4090 n5080 n4091 R=1.174e+01 
R5079t1540 n5080 n1541 R=4.648e+00 
R5080t548 n5081 n549 R=1.305e+01 
R5080t2843 n5081 n2844 R=4.952e+01 
R5080t891 n5081 n892 R=6.436e+00 
R5080t2473 n5081 n2474 R=6.220e+00 
R5081t4162 n5082 n4163 R=7.283e+00 
R5081t4560 n5082 n4561 R=3.863e+00 
R5081t3634 n5082 n3635 R=2.986e+02 
R5081t3348 n5082 n3349 R=4.036e+00 
R5081t2057 n5082 n2058 R=1.407e+01 
R5081t3866 n5082 n3867 R=8.412e+00 
R5082t3320 n5083 n3321 R=5.137e+00 
R5082t2081 n5083 n2082 R=1.402e+01 
R5083t305 n5084 n306 R=8.832e+00 
R5083t2449 n5084 n2450 R=2.383e+01 
R5083t1934 n5084 n1935 R=5.598e+00 
R5084t3205 n5085 n3206 R=1.331e+02 
R5084t11 n5085 n12 R=8.688e+00 
R5084t1015 n5085 n1016 R=2.969e+01 
R5084t3987 n5085 n3988 R=4.749e+00 
R5085t3737 n5086 n3738 R=4.226e+00 
R5085t1381 n5086 n1382 R=9.199e+00 
R5085t4992 n5086 n4993 R=4.602e+00 
R5086t3833 n5087 n3834 R=5.611e+00 
R5086t4433 n5087 n4434 R=1.593e+01 
R5087t2585 n5088 n2586 R=3.132e+02 
R5087t965 n5088 n966 R=1.222e+01 
R5088t416 n5089 n417 R=9.532e+01 
R5088t4465 n5089 n4466 R=1.498e+01 
R5088t1057 n5089 n1058 R=3.584e+01 
R5088t1897 n5089 n1898 R=4.265e+01 
R5089t4031 n5090 n4032 R=2.044e+00 
R5089t2150 n5090 n2151 R=1.405e+01 
R5089t3995 n5090 n3996 R=4.139e+00 
R5090t2993 n5091 n2994 R=7.512e+00 
R5090t4681 n5091 n4682 R=7.511e+00 
R5090t267 n5091 n268 R=9.100e+00 
R5090t2371 n5091 n2372 R=2.354e+01 
R5090t4761 n5091 n4762 R=6.719e+00 
R5090t3905 n5091 n3906 R=3.318e+01 
R5090t1960 n5091 n1961 R=4.899e+01 
R5091t3318 n5092 n3319 R=4.655e+00 
R5091t1043 n5092 n1044 R=7.497e+00 
R5091t4537 n5092 n4538 R=8.477e+00 
R5091t4789 n5092 n4790 R=1.116e+01 
R5091t3176 n5092 n3177 R=6.692e+00 
R5091t2504 n5092 n2505 R=1.843e+01 
R5092t4794 n5093 n4795 R=4.415e+00 
R5092t1240 n5093 n1241 R=4.928e+00 
R5092t1034 n5093 n1035 R=2.789e+01 
R5093t2399 n5094 n2400 R=5.868e+00 
R5095t2914 n5096 n2915 R=5.943e+00 
R5095t4696 n5096 n4697 R=8.062e+00 
R5095t606 n5096 n607 R=1.178e+01 
R5096t1951 n5097 n1952 R=4.978e+00 
R5096t3031 n5097 n3032 R=4.793e+00 
R5096t4229 n5097 n4230 R=3.296e+01 
R5097t113 n5098 n114 R=2.940e+00 
R5097t2621 n5098 n2622 R=4.424e+00 
R5098t1739 n5099 n1740 R=5.834e+00 
R5099t329 n5100 n330 R=4.341e+01 
R5099t2284 n5100 n2285 R=5.607e+00 
R5100t847 n5101 n848 R=1.162e+01 
R5100t1715 n5101 n1716 R=9.066e+00 
R5100t3509 n5101 n3510 R=8.283e+00 
R5100t3752 n5101 n3753 R=1.722e+01 
R5101t1298 n5102 n1299 R=6.949e+00 
R5101t788 n5102 n789 R=4.910e+00 
R5101t1649 n5102 n1650 R=4.297e+02 
R5101t4793 n5102 n4794 R=5.700e+00 
R5102t2924 n5103 n2925 R=4.339e+00 
R5102t4311 n5103 n4312 R=6.894e+00 
R5102t1821 n5103 n1822 R=7.258e+00 
R5102t1795 n5103 n1796 R=3.901e+00 
R5103t5059 n5104 n5060 R=3.652e+01 
R5103t1616 n5104 n1617 R=8.968e+00 
R5103t4556 n5104 n4557 R=4.397e+01 
R5103t1292 n5104 n1293 R=1.914e+01 
R5103t4128 n5104 n4129 R=8.269e+00 
R5104t1712 n5105 n1713 R=4.837e+00 
R5104t1349 n5105 n1350 R=1.065e+01 
R5104t4080 n5105 n4081 R=3.284e+01 
R5104t4988 n5105 n4989 R=7.387e+00 
R5105t2045 n5106 n2046 R=2.903e+00 
R5105t3343 n5106 n3344 R=4.711e+00 
R5105t3771 n5106 n3772 R=1.479e+01 
R5107t3114 n5108 n3115 R=4.693e+00 
R5107t4422 n5108 n4423 R=1.723e+01 
R5108t842 n5109 n843 R=3.608e+00 
R5108t3554 n5109 n3555 R=3.615e+01 
R5108t1466 n5109 n1467 R=1.136e+01 
R5108t102 n5109 n103 R=8.917e+00 
R5109t1257 n5110 n1258 R=4.695e+01 
R5109t2910 n5110 n2911 R=1.930e+00 
R5109t3832 n5110 n3833 R=1.760e+00 
R5110t3534 n5111 n3535 R=1.370e+01 
R5110t818 n5111 n819 R=3.948e+02 
R5110t3837 n5111 n3838 R=1.897e+01 
R5110t2546 n5111 n2547 R=3.801e+00 
R5111t3126 n5112 n3127 R=4.282e+00 
R5112t1496 n5113 n1497 R=6.523e+00 
R5112t4977 n5113 n4978 R=3.686e+00 
R5112t4014 n5113 n4015 R=4.791e+01 
R5113t1582 n5114 n1583 R=7.078e+00 
R5113t771 n5114 n772 R=1.455e+01 
R5113t3735 n5114 n3736 R=1.422e+01 
R5113t2067 n5114 n2068 R=1.149e+02 
R5114t1906 n5115 n1907 R=7.741e+00 
R5114t913 n5115 n914 R=8.819e+01 
R5115t2161 n5116 n2162 R=1.702e+00 
R5117t3921 n5118 n3922 R=4.445e+01 
R5117t4070 n5118 n4071 R=6.495e+00 
R5117t4284 n5118 n4285 R=3.869e+01 
R5118t1014 n5119 n1015 R=1.040e+01 
R5118t2666 n5119 n2667 R=2.075e+01 
R5118t511 n5119 n512 R=1.639e+01 
R5118t1241 n5119 n1242 R=1.399e+01 
R5118t557 n5119 n558 R=1.866e+01 
R5119t1416 n5120 n1417 R=1.371e+02 
R5119t3267 n5120 n3268 R=1.952e+00 
R5119t5015 n5120 n5016 R=1.902e+00 
R5120t3486 n5121 n3487 R=3.472e+00 
R5121t2447 n5122 n2448 R=4.182e+00 
R5122t414 n5123 n415 R=5.026e+01 
R5123t955 n5124 n956 R=8.102e+00 
R5123t4275 n5124 n4276 R=2.629e+01 
R5123t809 n5124 n810 R=4.737e+00 
R5123t2521 n5124 n2522 R=2.250e+01 
R5123t1357 n5124 n1358 R=5.019e+00 
R5124t1105 n5125 n1106 R=8.978e+00 
R5124t3377 n5125 n3378 R=1.420e+02 
R5125t3450 n5126 n3451 R=2.799e+01 
R5125t4099 n5126 n4100 R=5.295e+00 
R5125t307 n5126 n308 R=1.503e+01 
R5126t3447 n5127 n3448 R=9.838e+01 
R5126t2094 n5127 n2095 R=8.426e+00 
R5126t3806 n5127 n3807 R=2.986e+00 
R5126t4638 n5127 n4639 R=1.066e+01 
R5127t4269 n5128 n4270 R=2.751e+01 
R5127t3766 n5128 n3767 R=1.564e+01 
R5127t358 n5128 n359 R=3.581e+00 
R5128t4283 n5129 n4284 R=2.424e+00 
R5129t2743 n5130 n2744 R=2.813e+00 
R5130t2970 n5131 n2971 R=1.400e+01 
R5130t2968 n5131 n2969 R=8.236e+00 
R5130t3055 n5131 n3056 R=2.379e+01 
R5130t3098 n5131 n3099 R=1.324e+01 
R5131t2672 n5132 n2673 R=4.593e+00 
R5131t3596 n5132 n3597 R=5.202e+00 
R5131t1170 n5132 n1171 R=6.838e+01 
R5131t269 n5132 n270 R=8.476e+00 
R5131t3119 n5132 n3120 R=5.750e+01 
R5132t178 n5133 n179 R=7.354e+00 
R5132t4781 n5133 n4782 R=3.285e+00 
R5132t1811 n5133 n1812 R=1.106e+01 
R5133t4722 n5134 n4723 R=3.803e+00 
R5133t2489 n5134 n2490 R=6.464e+00 
R5133t2488 n5134 n2489 R=8.332e+00 
R5134t2262 n5135 n2263 R=4.762e+00 
R5134t2602 n5135 n2603 R=2.673e+01 
R5134t356 n5135 n357 R=1.518e+01 
R5134t4293 n5135 n4294 R=6.556e+00 
R5135t4535 n5136 n4536 R=5.342e+01 
R5135t1397 n5136 n1398 R=2.834e+00 
R5135t2813 n5136 n2814 R=1.678e+01 
R5135t476 n5136 n477 R=3.273e+01 
R5136t2733 n5137 n2734 R=3.515e+02 
R5137t1203 n5138 n1204 R=1.848e+01 
R5138t1786 n5139 n1787 R=4.376e+01 
R5138t4628 n5139 n4629 R=5.802e+00 
R5138t1102 n5139 n1103 R=4.510e+00 
R5139t2442 n5140 n2443 R=3.034e+00 
R5139t2935 n5140 n2936 R=8.147e+00 
R5139t2214 n5140 n2215 R=4.302e+00 
R5139t4340 n5140 n4341 R=1.524e+01 
R5140t989 n5141 n990 R=2.033e+00 
R5141t1071 n5142 n1072 R=5.650e+01 
R5141t2927 n5142 n2928 R=5.880e+00 
R5142t2209 n5143 n2210 R=2.059e+01 
R5142t2578 n5143 n2579 R=8.618e+00 
R5142t3025 n5143 n3026 R=1.125e+01 
R5142t1766 n5143 n1767 R=5.908e+01 
R5142t1127 n5143 n1128 R=4.637e+00 
R5142t94 n5143 n95 R=8.123e+00 
R5143t2737 n5144 n2738 R=8.089e+00 
R5143t717 n5144 n718 R=1.125e+01 
R5143t1667 n5144 n1668 R=2.570e+04 
R5143t1106 n5144 n1107 R=1.212e+03 
R5143t4278 n5144 n4279 R=4.570e+00 
R5143t963 n5144 n964 R=2.021e+01 
R5144t1604 n5145 n1605 R=3.653e+00 
R5144t1680 n5145 n1681 R=9.039e+00 
R5144t2114 n5145 n2115 R=1.724e+01 
R5145t4679 n5146 n4680 R=7.210e+00 
R5145t4500 n5146 n4501 R=4.698e+00 
R5146t2705 n5147 n2706 R=1.282e+02 
R5146t4025 n5147 n4026 R=4.152e+00 
R5146t4265 n5147 n4266 R=8.934e+00 
R5147t1182 n5148 n1183 R=1.426e+01 
R5147t2722 n5148 n2723 R=4.424e+00 
R5147t4868 n5148 n4869 R=7.527e+00 
R5147t3667 n5148 n3668 R=5.973e+00 
R5148t1095 n5149 n1096 R=2.905e+00 
R5148t319 n5149 n320 R=9.393e+00 
R5149t2417 n5150 n2418 R=3.588e+00 
R5149t3983 n5150 n3984 R=1.462e+01 
R5149t2544 n5150 n2545 R=1.394e+01 
R5150t371 n5151 n372 R=2.891e+00 
R5150t3152 n5151 n3153 R=3.753e+01 
R5151t3338 n5152 n3339 R=3.256e+00 
R5152t2306 n5153 n2307 R=2.174e+00 
R5152t1827 n5153 n1828 R=1.022e+01 
R5152t4034 n5153 n4035 R=1.104e+02 
R5153t3928 n5154 n3929 R=2.349e+02 
R5153t2673 n5154 n2674 R=5.598e+00 
R5153t2921 n5154 n2922 R=7.242e+00 
R5153t3656 n5154 n3657 R=1.570e+01 
R5154t1991 n5155 n1992 R=3.700e+00 
R5154t4877 n5155 n4878 R=5.374e+00 
R5154t4325 n5155 n4326 R=4.695e+00 
R5155t2612 n5156 n2613 R=1.349e+01 
R5155t2644 n5156 n2645 R=2.860e+00 
R5155t1861 n5156 n1862 R=3.652e+00 
R5156t625 n5157 n626 R=3.983e+00 
R5156t818 n5157 n819 R=2.273e+00 
R5157t2436 n5158 n2437 R=1.532e+01 
R5157t449 n5158 n450 R=5.701e+00 
R5158t1470 n5159 n1471 R=4.873e+00 
R5158t4858 n5159 n4859 R=2.981e+00 
R5159t3431 n5160 n3432 R=4.817e+00 
R5159t2587 n5160 n2588 R=1.151e+01 
R5159t2263 n5160 n2264 R=4.358e+00 
R5159t217 n5160 n218 R=1.019e+02 
R5160t1013 n5161 n1014 R=4.386e+00 
R5160t4749 n5161 n4750 R=6.010e+00 
R5160t4116 n5161 n4117 R=3.036e+00 
R5160t1338 n5161 n1339 R=8.301e+00 
R5161t4204 n5162 n4205 R=2.642e+00 
R5161t217 n5162 n218 R=1.371e+00 
R5161t5159 n5162 n5160 R=1.096e+01 
R5162t642 n5163 n643 R=2.467e+00 
R5162t2082 n5163 n2083 R=8.429e+00 
R5162t1088 n5163 n1089 R=1.568e+01 
R5162t3938 n5163 n3939 R=6.056e+00 
R5162t3082 n5163 n3083 R=6.604e+00 
R5163t761 n5164 n762 R=1.123e+01 
R5163t2840 n5164 n2841 R=2.061e+00 
R5163t1421 n5164 n1422 R=4.500e+00 
R5164t3698 n5165 n3699 R=4.669e+00 
R5164t3853 n5165 n3854 R=6.613e+01 
R5164t907 n5165 n908 R=5.850e+01 
R5164t4357 n5165 n4358 R=3.505e+00 
R5164t2802 n5165 n2803 R=7.395e+01 
R5164t251 n5165 n252 R=5.304e+00 
R5164t4823 n5165 n4824 R=1.504e+02 
R5165t2733 n5166 n2734 R=7.761e+00 
R5165t451 n5166 n452 R=7.821e+00 
R5166t129 n5167 n130 R=4.807e+01 
R5166t3822 n5167 n3823 R=1.055e+01 
R5166t2330 n5167 n2331 R=3.941e+00 
R5167t1168 n5168 n1169 R=5.326e+00 
R5167t2608 n5168 n2609 R=4.789e+01 
R5167t3972 n5168 n3973 R=2.739e+00 
R5167t2156 n5168 n2157 R=1.596e+01 
R5168t4324 n5169 n4325 R=7.275e+00 
R5169t2996 n5170 n2997 R=9.313e+00 
R5169t1965 n5170 n1966 R=4.305e+00 
R5170t294 n5171 n295 R=4.364e+00 
R5170t4551 n5171 n4552 R=7.682e+00 
R5170t2359 n5171 n2360 R=4.564e+01 
R5171t372 n5172 n373 R=4.245e+01 
R5171t4424 n5172 n4425 R=1.311e+01 
R5171t3434 n5172 n3435 R=6.199e+01 
R5171t318 n5172 n319 R=3.091e+00 
R5172t3280 n5173 n3281 R=8.207e+00 
R5172t2093 n5173 n2094 R=4.020e+00 
R5172t2678 n5173 n2679 R=2.962e+01 
R5173t1038 n5174 n1039 R=3.825e+00 
R5173t4155 n5174 n4156 R=1.056e+02 
R5174t598 n5175 n599 R=1.644e+01 
R5174t790 n5175 n791 R=9.878e+00 
R5174t635 n5175 n636 R=1.083e+01 
R5174t1113 n5175 n1114 R=9.323e+00 
R5174t1434 n5175 n1435 R=1.248e+02 
R5175t1524 n5176 n1525 R=9.388e+00 
R5175t3485 n5176 n3486 R=6.416e+00 
R5175t43 n5176 n44 R=1.109e+01 
R5175t3892 n5176 n3893 R=1.752e+01 
R5176t2062 n5177 n2063 R=2.793e+00 
R5176t1676 n5177 n1677 R=3.461e+01 
R5177t1140 n5178 n1141 R=4.155e+01 
R5177t2945 n5178 n2946 R=4.598e+01 
R5177t3376 n5178 n3377 R=3.497e+00 
R5178t2710 n5179 n2711 R=1.383e+00 
R5178t1384 n5179 n1385 R=4.472e+00 
R5178t654 n5179 n655 R=3.821e+00 
R5179t2233 n5180 n2234 R=2.340e+01 
R5179t2757 n5180 n2758 R=3.659e+00 
R5179t4704 n5180 n4705 R=8.352e+00 
R5179t1809 n5180 n1810 R=9.737e+00 
R5180t3504 n5181 n3505 R=9.676e+00 
R5180t4481 n5181 n4482 R=2.693e+00 
R5180t1901 n5181 n1902 R=3.775e+01 
R5181t4881 n5182 n4882 R=9.291e+00 
R5181t128 n5182 n129 R=9.035e+00 
R5181t3818 n5182 n3819 R=1.300e+03 
R5182t1109 n5183 n1110 R=8.723e+01 
R5182t2995 n5183 n2996 R=6.104e+00 
R5182t2690 n5183 n2691 R=5.779e+01 
R5183t1899 n5184 n1900 R=3.161e+00 
R5183t4947 n5184 n4948 R=1.751e+01 
R5184t727 n5185 n728 R=3.085e+00 
R5184t2702 n5185 n2703 R=2.089e+00 
R5184t1458 n5185 n1459 R=6.671e+01 
R5184t4853 n5185 n4854 R=4.186e+00 
R5185t1693 n5186 n1694 R=3.783e+01 
R5185t2332 n5186 n2333 R=1.044e+01 
R5185t2226 n5186 n2227 R=4.384e+00 
R5185t2336 n5186 n2337 R=4.440e+00 
R5186t2421 n5187 n2422 R=6.138e+00 
R5186t3032 n5187 n3033 R=2.463e+00 
R5186t4408 n5187 n4409 R=4.826e+01 
R5186t3247 n5187 n3248 R=6.260e+00 
R5187t2315 n5188 n2316 R=4.189e+00 
R5187t2094 n5188 n2095 R=1.285e+01 
R5188t4962 n5189 n4963 R=1.789e+00 
R5188t3236 n5189 n3237 R=1.285e+01 
R5188t3989 n5189 n3990 R=3.098e+00 
R5189t3935 n5190 n3936 R=2.361e+00 
R5190t978 n5191 n979 R=8.589e+00 
R5190t4505 n5191 n4506 R=7.078e+00 
R5190t4037 n5191 n4038 R=1.489e+01 
R5191t1351 n5192 n1352 R=5.062e+01 
R5191t4106 n5192 n4107 R=3.012e+01 
R5191t25 n5192 n26 R=4.471e+00 
R5193t1487 n5194 n1488 R=1.642e+01 
R5193t3901 n5194 n3902 R=1.382e+02 
R5193t4276 n5194 n4277 R=4.330e+00 
R5194t4303 n5195 n4304 R=4.071e+00 
R5194t3713 n5195 n3714 R=5.869e+00 
R5195t2025 n5196 n2026 R=6.102e+00 
R5195t691 n5196 n692 R=4.052e+00 
R5195t1115 n5196 n1116 R=3.933e+00 
R5195t1150 n5196 n1151 R=2.115e+02 
R5196t3429 n5197 n3430 R=8.185e+00 
R5196t891 n5197 n892 R=4.341e+01 
R5196t2473 n5197 n2474 R=1.145e+01 
R5196t4971 n5197 n4972 R=8.688e+01 
R5196t2674 n5197 n2675 R=4.985e+00 
R5196t1187 n5197 n1188 R=1.277e+01 
R5196t1623 n5197 n1624 R=5.490e+00 
R5197t2035 n5198 n2036 R=3.035e+00 
R5197t4635 n5198 n4636 R=6.434e+00 
R5198t2349 n5199 n2350 R=5.989e+00 
R5198t3996 n5199 n3997 R=7.439e+00 
R5199t2169 n5200 n2170 R=7.165e+00 
R5199t4334 n5200 n4335 R=5.208e+00 
R5199t523 n5200 n524 R=8.327e+00 
R5200t81 n5201 n82 R=2.763e+00 
R5200t311 n5201 n312 R=1.669e+01 
R5200t2180 n5201 n2181 R=1.322e+02 
R5201t1128 n5202 n1129 R=3.319e+01 
R5201t1469 n5202 n1470 R=2.666e+00 
R5202t3069 n5203 n3070 R=4.189e+00 
R5202t801 n5203 n802 R=5.674e+00 
R5202t3724 n5203 n3725 R=8.044e+00 
R5203t2825 n5204 n2826 R=1.548e+01 
R5203t2531 n5204 n2532 R=1.385e+01 
R5203t1730 n5204 n1731 R=4.613e+01 
R5203t794 n5204 n795 R=3.517e+01 
R5203t1784 n5204 n1785 R=3.302e+00 
R5204t2845 n5205 n2846 R=6.124e+00 
R5204t4837 n5205 n4838 R=5.074e+00 
R5204t1615 n5205 n1616 R=5.831e+00 
R5204t2172 n5205 n2173 R=8.385e+00 
R5205t1444 n5206 n1445 R=1.467e+01 
R5205t653 n5206 n654 R=2.498e+00 
R5206t3896 n5207 n3897 R=6.132e+00 
R5206t3852 n5207 n3853 R=9.307e+00 
R5207t182 n5208 n183 R=1.159e+02 
R5207t2705 n5208 n2706 R=6.925e+00 
R5207t5146 n5208 n5147 R=5.547e+00 
R5207t4025 n5208 n4026 R=7.417e+00 
R5208t3343 n5209 n3344 R=1.613e+01 
R5208t4030 n5209 n4031 R=4.665e+00 
R5210t1514 n5211 n1515 R=1.106e+01 
R5210t2416 n5211 n2417 R=7.454e+00 
R5210t1140 n5211 n1141 R=2.982e+01 
R5210t3633 n5211 n3634 R=5.850e+00 
R5211t1554 n5212 n1555 R=3.282e+00 
R5211t3313 n5212 n3314 R=6.784e+00 
R5211t3988 n5212 n3989 R=7.200e+00 
R5212t2527 n5213 n2528 R=7.593e+00 
R5212t1711 n5213 n1712 R=9.704e+00 
R5212t2549 n5213 n2550 R=7.374e+00 
R5213t3542 n5214 n3543 R=4.013e+00 
R5213t4941 n5214 n4942 R=3.414e+00 
R5213t3452 n5214 n3453 R=5.892e+00 
R5214t717 n5215 n718 R=1.322e+01 
R5214t4049 n5215 n4050 R=3.054e+00 
R5214t4390 n5215 n4391 R=3.397e+00 
R5214t2737 n5215 n2738 R=1.951e+01 
R5214t5143 n5215 n5144 R=9.358e+00 
R5215t274 n5216 n275 R=4.401e+00 
R5215t892 n5216 n893 R=9.701e+00 
R5215t3914 n5216 n3915 R=6.608e+00 
R5215t3152 n5216 n3153 R=1.589e+01 
R5216t1955 n5217 n1956 R=2.103e+01 
R5216t3126 n5217 n3127 R=1.721e+02 
R5216t5111 n5217 n5112 R=8.343e+01 
R5216t4464 n5217 n4465 R=4.907e+01 
R5217t250 n5218 n251 R=6.197e+01 
R5217t2055 n5218 n2056 R=4.529e+00 
R5217t3241 n5218 n3242 R=6.710e+00 
R5217t3063 n5218 n3064 R=1.850e+01 
R5217t448 n5218 n449 R=2.342e+00 
R5217t3523 n5218 n3524 R=2.621e+01 
R5218t285 n5219 n286 R=2.787e+01 
R5218t2132 n5219 n2133 R=4.736e+00 
R5218t1611 n5219 n1612 R=2.671e+01 
R5218t4524 n5219 n4525 R=1.774e+01 
R5219t2376 n5220 n2377 R=4.163e+00 
R5220t4273 n5221 n4274 R=3.783e+01 
R5220t5034 n5221 n5035 R=5.943e+00 
R5220t118 n5221 n119 R=3.257e+01 
R5220t4073 n5221 n4074 R=3.538e+00 
R5221t4502 n5222 n4503 R=6.661e+00 
R5221t2383 n5222 n2384 R=6.921e+00 
R5221t3715 n5222 n3716 R=9.113e+00 
R5221t1108 n5222 n1109 R=8.704e+00 
R5222t1913 n5223 n1914 R=3.641e+00 
R5222t3377 n5223 n3378 R=3.522e+01 
R5222t5124 n5223 n5125 R=5.810e+00 
R5222t1105 n5223 n1106 R=1.286e+02 
R5222t3470 n5223 n3471 R=2.411e+01 
R5222t1618 n5223 n1619 R=2.274e+01 
R5223t1145 n5224 n1146 R=2.461e+01 
R5223t4332 n5224 n4333 R=2.533e+00 
R5223t1388 n5224 n1389 R=9.358e+00 
R5223t1572 n5224 n1573 R=2.779e+00 
R5223t3797 n5224 n3798 R=2.425e+01 
R5224t2621 n5225 n2622 R=5.411e+00 
R5224t507 n5225 n508 R=4.392e+01 
R5224t4544 n5225 n4545 R=2.888e+00 
R5225t1403 n5226 n1404 R=7.133e+00 
R5226t1013 n5227 n1014 R=2.926e+00 
R5226t516 n5227 n517 R=2.080e+00 
R5227t1444 n5228 n1445 R=3.894e+00 
R5227t5205 n5228 n5206 R=2.747e+00 
R5228t997 n5229 n998 R=2.015e+00 
R5228t4966 n5229 n4967 R=7.550e+01 
R5229t1750 n5230 n1751 R=1.094e+01 
R5229t4811 n5230 n4812 R=1.017e+01 
R5230t424 n5231 n425 R=9.758e+01 
R5230t4903 n5231 n4904 R=4.058e+00 
R5230t4580 n5231 n4581 R=4.472e+00 
R5230t4203 n5231 n4204 R=2.185e+02 
R5230t4735 n5231 n4736 R=7.404e+00 
R5231t1965 n5232 n1966 R=7.807e+00 
R5231t5169 n5232 n5170 R=1.318e+01 
R5232t2159 n5233 n2160 R=1.490e+01 
R5232t3842 n5233 n3843 R=3.603e+00 
R5232t451 n5233 n452 R=7.308e+01 
R5232t3964 n5233 n3965 R=4.915e+01 
R5233t1483 n5234 n1484 R=2.038e+01 
R5233t4955 n5234 n4956 R=2.740e+01 
R5233t1843 n5234 n1844 R=3.089e+00 
R5233t2689 n5234 n2690 R=4.824e+00 
R5233t691 n5234 n692 R=1.067e+01 
R5234t1740 n5235 n1741 R=5.312e+00 
R5234t2517 n5235 n2518 R=2.572e+00 
R5234t2054 n5235 n2055 R=4.731e+00 
R5234t4402 n5235 n4403 R=1.041e+01 
R5235t1296 n5236 n1297 R=2.723e+00 
R5235t5004 n5236 n5005 R=1.307e+02 
R5235t2215 n5236 n2216 R=9.299e+00 
R5235t330 n5236 n331 R=1.363e+01 
R5236t555 n5237 n556 R=1.064e+01 
R5236t3397 n5237 n3398 R=3.424e+00 
R5237t4552 n5238 n4553 R=4.733e+00 
R5237t1555 n5238 n1556 R=1.013e+01 
R5237t670 n5238 n671 R=1.890e+01 
R5238t3611 n5239 n3612 R=1.981e+01 
R5238t4276 n5239 n4277 R=6.759e+00 
R5238t5193 n5239 n5194 R=5.021e+00 
R5239t3422 n5240 n3423 R=7.216e+02 
R5239t2816 n5240 n2817 R=2.385e+00 
R5239t542 n5240 n543 R=4.836e+01 
R5240t3139 n5241 n3140 R=2.263e+00 
R5240t3061 n5241 n3062 R=1.535e+01 
R5241t1669 n5242 n1670 R=9.872e+01 
R5241t2494 n5242 n2495 R=5.607e+00 
R5241t4893 n5242 n4894 R=5.210e+00 
R5241t4212 n5242 n4213 R=1.866e+01 
R5242t2273 n5243 n2274 R=3.177e+00 
R5242t93 n5243 n94 R=4.383e+01 
R5242t3500 n5243 n3501 R=5.969e+00 
R5243t2980 n1 n2981 R=4.118e+03 
R5245t2164 n5246 n2165 R=3.668e+00 
R5245t2828 n5246 n2829 R=2.017e+01 
R5245t3197 n5246 n3198 R=4.579e+00 
R5245t3413 n5246 n3414 R=2.765e+01 
R5246t1139 n5247 n1140 R=2.778e+02 
R5246t4927 n5247 n4928 R=2.608e+01 
R5246t1350 n5247 n1351 R=3.153e+03 
R5246t3818 n5247 n3819 R=1.069e+01 
R5247t4538 n5248 n4539 R=1.645e+01 
R5247t3040 n5248 n3041 R=3.890e+01 
R5247t4119 n5248 n4120 R=1.839e+01 
R5248t1367 n5249 n1368 R=4.014e+00 
R5248t3590 n5249 n3591 R=3.241e+02 
R5248t1237 n5249 n1238 R=4.060e+00 
R5249t2309 n5250 n2310 R=6.392e+00 
R5249t3313 n5250 n3314 R=8.871e+00 
R5249t3800 n5250 n3801 R=3.157e+01 
R5249t4656 n5250 n4657 R=1.304e+01 
R5250t2505 n5251 n2506 R=2.279e+01 
R5250t3258 n5251 n3259 R=5.386e+00 
R5250t5065 n5251 n5066 R=5.552e+00 
R5250t10 n5251 n11 R=5.533e+00 
R5251t1982 n5252 n1983 R=1.084e+00 
R5251t5071 n5252 n5072 R=1.018e+01 
R5251t988 n5252 n989 R=1.857e+01 
R5252t2521 n5253 n2522 R=2.549e+01 
R5252t1357 n5253 n1358 R=1.562e+00 
R5253t561 n5254 n562 R=1.295e+02 
R5253t2919 n5254 n2920 R=5.461e+00 
R5253t3205 n5254 n3206 R=2.232e+00 
R5253t5084 n5254 n5085 R=5.076e+00 
R5253t11 n5254 n12 R=6.833e+00 
R5254t3699 n5255 n3700 R=2.366e+01 
R5255t1151 n5256 n1152 R=9.705e+00 
R5255t4963 n5256 n4964 R=8.218e+00 
R5255t580 n5256 n581 R=3.366e+01 
R5255t271 n5256 n272 R=7.029e+00 
R5255t119 n5256 n120 R=3.958e+00 
R5256t4083 n5257 n4084 R=1.731e+01 
R5256t4726 n5257 n4727 R=3.948e+01 
R5256t2862 n5257 n2863 R=2.668e+02 
R5256t4947 n5257 n4948 R=6.583e+01 
R5257t2618 n5258 n2619 R=3.629e+00 
R5258t830 n5259 n831 R=2.782e+01 
R5259t277 n5260 n278 R=9.788e+00 
R5259t1538 n5260 n1539 R=2.438e+00 
R5260t620 n5261 n621 R=1.814e+01 
R5260t933 n5261 n934 R=4.125e+00 
R5261t4944 n5262 n4945 R=8.188e+01 
R5262t3970 n5263 n3971 R=1.173e+01 
R5262t26 n5263 n27 R=6.613e+01 
R5262t2409 n5263 n2410 R=3.021e+00 
R5263t2322 n5264 n2323 R=8.265e+00 
R5263t227 n5264 n228 R=2.316e+01 
R5264t907 n5265 n908 R=1.524e+01 
R5264t2802 n5265 n2803 R=1.464e+01 
R5264t3998 n5265 n3999 R=6.136e+00 
R5264t1948 n5265 n1949 R=5.311e+00 
R5264t638 n5265 n639 R=2.241e+01 
R5264t1181 n5265 n1182 R=1.490e+01 
R5265t3909 n5266 n3910 R=1.030e+01 
R5265t3203 n5266 n3204 R=2.110e+00 
R5265t2369 n5266 n2370 R=4.251e+00 
R5266t2664 n5267 n2665 R=3.979e+00 
R5266t96 n5267 n97 R=8.639e+02 
R5266t3527 n5267 n3528 R=3.443e+00 
R5267t5261 n5268 n5262 R=6.574e+01 
R5267t4944 n5268 n4945 R=9.142e+00 
R5268t4567 n5269 n4568 R=3.899e+01 
R5268t4222 n5269 n4223 R=4.204e+00 
R5269t2591 n5270 n2592 R=5.164e+01 
R5269t4625 n5270 n4626 R=4.517e+00 
R5269t4006 n5270 n4007 R=9.224e+00 
R5269t4699 n5270 n4700 R=1.323e+01 
R5269t70 n5270 n71 R=1.165e+01 
R5269t4092 n5270 n4093 R=1.160e+01 
R5270t2414 n5271 n2415 R=4.475e+01 
R5270t1291 n5271 n1292 R=2.124e+01 
R5270t1737 n5271 n1738 R=1.948e+01 
R5270t3363 n5271 n3364 R=3.121e+00 
R5270t1936 n5271 n1937 R=2.608e+01 
R5271t2357 n5272 n2358 R=6.265e+00 
R5271t3006 n5272 n3007 R=6.541e+00 
R5272t407 n5273 n408 R=4.047e+00 
R5272t4311 n5273 n4312 R=2.303e+02 
R5272t2924 n5273 n2925 R=4.677e+00 
R5273t904 n5274 n905 R=9.446e+00 
R5273t2323 n5274 n2324 R=5.463e+01 
R5274t55 n5275 n56 R=1.035e+01 
R5274t613 n5275 n614 R=6.858e+00 
R5274t4192 n5275 n4193 R=1.687e+01 
R5274t4670 n5275 n4671 R=1.760e+01 
R5274t4178 n5275 n4179 R=3.312e+00 
R5274t2102 n5275 n2103 R=2.315e+01 
R5275t4753 n5276 n4754 R=2.819e+00 
R5276t4131 n5277 n4132 R=3.106e+00 
R5276t3522 n5277 n3523 R=1.838e+01 
R5276t4100 n5277 n4101 R=4.598e+00 
R5277t2379 n5278 n2380 R=4.355e+00 
R5277t1689 n5278 n1690 R=1.756e+02 
R5278t1710 n5279 n1711 R=2.028e+01 
R5278t1952 n5279 n1953 R=5.046e+00 
R5278t486 n5279 n487 R=5.722e+00 
R5278t1465 n5279 n1466 R=9.022e+01 
R5278t4302 n5279 n4303 R=1.921e+01 
R5278t3387 n5279 n3388 R=7.265e+00 
R5278t3696 n5279 n3697 R=6.523e+01 
R5279t4255 n5280 n4256 R=1.008e+01 
R5279t2665 n5280 n2666 R=7.289e+00 
R5279t2189 n5280 n2190 R=6.138e+00 
R5280t369 n5281 n370 R=3.986e+00 
R5280t4279 n5281 n4280 R=5.493e+00 
R5280t1561 n5281 n1562 R=1.161e+01 
R5281t2825 n5282 n2826 R=4.585e+01 
R5281t5203 n5282 n5204 R=3.313e+00 
R5281t1784 n5282 n1785 R=5.578e+01 
R5282t2015 n5283 n2016 R=6.067e+01 
R5282t1082 n5283 n1083 R=2.418e+01 
R5282t4210 n5283 n4211 R=9.628e+00 
R5282t1577 n5283 n1578 R=2.154e+00 
R5283t5231 n5284 n5232 R=5.452e+00 
R5283t1559 n5284 n1560 R=4.131e+00 
R5283t1965 n5284 n1966 R=5.360e+00 
R5284t772 n5285 n773 R=1.014e+01 
R5284t385 n5285 n386 R=7.534e+00 
R5285t2180 n5286 n2181 R=1.727e+00 
R5285t5200 n5286 n5201 R=2.522e+02 
R5285t81 n5286 n82 R=7.466e+00 
R5286t3724 n5287 n3725 R=1.046e+01 
R5286t1265 n5287 n1266 R=8.422e+00 
R5286t4088 n5287 n4089 R=4.736e+00 
R5286t2253 n5287 n2254 R=4.751e+00 
R5287t2013 n5288 n2014 R=1.780e+01 
R5287t2307 n5288 n2308 R=4.412e+00 
R5287t3745 n5288 n3746 R=2.089e+00 
R5287t2762 n5288 n2763 R=1.699e+01 
R5287t2866 n5288 n2867 R=6.951e+00 
R5288t2631 n5289 n2632 R=1.871e+01 
R5288t5058 n5289 n5059 R=4.914e+00 
R5288t4098 n5289 n4099 R=4.046e+00 
R5289t1337 n5290 n1338 R=1.060e+01 
R5290t452 n5291 n453 R=3.898e+00 
R5290t2853 n5291 n2854 R=8.923e+00 
R5290t762 n5291 n763 R=3.013e+00 
R5291t3847 n5292 n3848 R=2.039e+01 
R5291t3325 n5292 n3326 R=2.818e+00 
R5291t987 n5292 n988 R=1.069e+01 
R5291t4941 n5292 n4942 R=2.372e+00 
R5293t4324 n5294 n4325 R=3.943e+00 
R5293t3390 n5294 n3391 R=8.116e+00 
R5294t4039 n5295 n4040 R=2.433e+01 
R5294t1810 n5295 n1811 R=8.550e+00 
R5294t1539 n5295 n1540 R=2.228e+01 
R5294t3872 n5295 n3873 R=5.368e+00 
R5295t1183 n5296 n1184 R=1.396e+01 
R5295t5073 n5296 n5074 R=2.258e+00 
R5295t2570 n5296 n2571 R=3.013e+00 
R5295t3239 n5296 n3240 R=1.895e+01 
R5296t1611 n5297 n1612 R=2.159e+00 
R5296t2327 n5297 n2328 R=2.997e+01 
R5296t771 n5297 n772 R=2.369e+01 
R5296t969 n5297 n970 R=9.178e+00 
R5296t2132 n5297 n2133 R=2.332e+01 
R5297t3887 n5298 n3888 R=3.884e+01 
R5297t4800 n5298 n4801 R=6.865e+00 
R5298t1493 n5299 n1494 R=6.324e+00 
R5298t3522 n5299 n3523 R=4.337e+00 
R5298t1563 n5299 n1564 R=8.172e+00 
R5299t4398 n5300 n4399 R=8.985e+00 
R5299t256 n5300 n257 R=4.272e+00 
R5300t4406 n5301 n4407 R=3.263e+00 
R5300t1138 n5301 n1139 R=8.565e+00 
R5301t2856 n5302 n2857 R=4.188e+00 
R5302t2410 n5303 n2411 R=3.240e+00 
R5302t1410 n5303 n1411 R=6.970e+01 
R5302t253 n5303 n254 R=4.851e+00 
R5303t1721 n5304 n1722 R=4.078e+01 
R5303t4368 n5304 n4369 R=6.029e+00 
R5303t2942 n5304 n2943 R=5.495e+00 
R5304t205 n5305 n206 R=1.360e+01 
R5304t2893 n5305 n2894 R=3.502e+01 
R5304t3777 n5305 n3778 R=2.550e+00 
R5305t1939 n5306 n1940 R=2.550e+00 
R5305t3327 n5306 n3328 R=1.831e+01 
R5305t3654 n5306 n3655 R=1.529e+00 
R5306t2373 n5307 n2374 R=2.265e+00 
R5306t2081 n5307 n2082 R=1.060e+01 
R5306t2363 n5307 n2364 R=3.476e+01 
R5306t263 n5307 n264 R=2.456e+01 
R5307t915 n5308 n916 R=1.011e+01 
R5307t1254 n5308 n1255 R=3.536e+00 
R5307t917 n5308 n918 R=1.388e+01 
R5308t2752 n5309 n2753 R=2.394e+01 
R5308t585 n5309 n586 R=3.455e+00 
R5308t1355 n5309 n1356 R=5.466e+00 
R5309t4244 n5310 n4245 R=4.274e+00 
R5309t2766 n5310 n2767 R=1.031e+03 
R5310t4849 n5311 n4850 R=6.280e+00 
R5310t3406 n5311 n3407 R=1.145e+01 
R5310t2583 n5311 n2584 R=4.615e+00 
R5310t2115 n5311 n2116 R=3.262e+00 
R5311t1070 n5312 n1071 R=4.281e+00 
R5311t537 n5312 n538 R=1.511e+01 
R5311t1634 n5312 n1635 R=2.480e+01 
R5311t865 n5312 n866 R=3.819e+00 
R5312t4675 n5313 n4676 R=1.031e+02 
R5312t3636 n5313 n3637 R=1.102e+01 
R5313t3751 n5314 n3752 R=8.229e+00 
R5314t2334 n5315 n2335 R=7.220e+00 
R5314t3671 n5315 n3672 R=5.783e+00 
R5314t4558 n5315 n4559 R=7.754e+01 
R5315t2963 n5316 n2964 R=3.404e+00 
R5315t1455 n5316 n1456 R=7.398e+00 
R5315t4156 n5316 n4157 R=2.803e+01 
R5316t470 n5317 n471 R=2.793e+01 
R5316t5038 n5317 n5039 R=5.110e+00 
R5316t179 n5317 n180 R=1.066e+02 
R5316t3715 n5317 n3716 R=2.008e+01 
R5316t2383 n5317 n2384 R=2.189e+00 
R5317t2970 n5318 n2971 R=4.941e+02 
R5317t532 n5318 n533 R=7.479e+00 
R5317t1569 n5318 n1570 R=1.418e+01 
R5317t3635 n5318 n3636 R=2.323e+00 
R5318t529 n5319 n530 R=1.488e+01 
R5318t2051 n5319 n2052 R=7.207e+00 
R5318t4011 n5319 n4012 R=2.373e+01 
R5318t2062 n5319 n2063 R=6.007e+00 
R5318t5176 n5319 n5177 R=6.561e+00 
R5318t242 n5319 n243 R=2.413e+01 
R5319t2513 n5320 n2514 R=1.664e+01 
R5319t4264 n5320 n4265 R=8.187e+00 
R5319t3719 n5320 n3720 R=2.133e+00 
R5319t438 n5320 n439 R=4.036e+01 
R5320t3612 n5321 n3613 R=2.607e+00 
R5320t65 n5321 n66 R=2.655e+01 
R5320t3851 n5321 n3852 R=6.234e+00 
R5321t183 n5322 n184 R=8.571e+00 
R5321t1235 n5322 n1236 R=2.930e+00 
R5322t2323 n5323 n2324 R=6.313e+00 
R5322t5273 n5323 n5274 R=2.578e+00 
R5322t2474 n5323 n2475 R=1.162e+02 
R5322t4702 n5323 n4703 R=2.736e+00 
R5323t2117 n5324 n2118 R=1.357e+01 
R5323t664 n5324 n665 R=2.900e+00 
R5324t3026 n5325 n3027 R=1.208e+01 
R5324t4848 n5325 n4849 R=7.357e+00 
R5325t3106 n5326 n3107 R=4.245e+00 
R5326t1824 n5327 n1825 R=4.897e+00 
R5326t3720 n5327 n3721 R=7.032e+00 
R5326t4683 n5327 n4684 R=4.305e+01 
R5326t3367 n5327 n3368 R=1.052e+02 
R5327t2826 n5328 n2827 R=6.016e+01 
R5327t2083 n5328 n2084 R=4.506e+00 
R5327t3109 n5328 n3110 R=1.492e+01 
R5327t4310 n5328 n4311 R=1.391e+01 
R5328t2239 n5329 n2240 R=4.434e+00 
R5328t2366 n5329 n2367 R=5.855e+02 
R5328t2920 n5329 n2921 R=9.627e+00 
R5328t3631 n5329 n3632 R=6.510e+00 
R5329t187 n5330 n188 R=1.497e+01 
R5329t3382 n5330 n3383 R=1.976e+00 
R5329t4924 n5330 n4925 R=1.010e+01 
R5330t1787 n5331 n1788 R=2.903e+01 
R5330t3232 n5331 n3233 R=4.071e+00 
R5330t4189 n5331 n1 R=3.297e+00 
R5331t2431 n5332 n2432 R=3.128e+00 
R5332t2854 n5333 n2855 R=7.732e+00 
R5333t21 n5334 n22 R=2.284e+00 
R5333t4678 n5334 n4679 R=5.665e+00 
R5333t2699 n5334 n2700 R=1.700e+00 
R5333t2295 n5334 n2296 R=3.379e+01 
R5334t2634 n5335 n2635 R=3.166e+00 
R5334t4020 n5335 n4021 R=5.638e+00 
R5334t1186 n5335 n1187 R=7.854e+00 
R5334t4478 n5335 n4479 R=4.531e+00 
R5335t1747 n5336 n1748 R=7.243e+00 
R5335t3615 n5336 n3616 R=4.757e+00 
R5336t1712 n5337 n1713 R=9.480e+00 
R5336t5104 n5337 n5105 R=4.508e+00 
R5336t1349 n5337 n1350 R=6.626e+00 
R5336t258 n5337 n259 R=1.486e+01 
R5337t1325 n5338 n1326 R=3.584e+00 
R5337t2078 n5338 n2079 R=2.257e+01 
R5337t1915 n5338 n1916 R=2.285e+01 
R5338t2919 n5339 n2920 R=6.075e+00 
R5338t5253 n5339 n5254 R=2.690e+01 
R5338t11 n5339 n12 R=1.494e+02 
R5338t115 n5339 n116 R=1.593e+01 
R5338t5019 n5339 n5020 R=3.092e+00 
R5339t4086 n5340 n4087 R=5.721e+01 
R5339t4983 n5340 n4984 R=2.462e+01 
R5340t640 n5341 n641 R=4.937e+00 
R5340t1571 n5341 n1572 R=4.976e+00 
R5340t3603 n5341 n3604 R=8.111e+00 
R5341t2501 n5342 n2502 R=1.477e+01 
R5341t3020 n5342 n3021 R=2.601e+00 
R5341t1113 n5342 n1114 R=3.040e+01 
R5341t4469 n5342 n4470 R=3.702e+00 
R5342t3815 n5343 n3816 R=6.181e+00 
R5342t5290 n5343 n5291 R=4.047e+01 
R5342t762 n5343 n763 R=9.341e+00 
R5342t436 n5343 n437 R=7.554e+00 
R5343t588 n5344 n589 R=1.089e+01 
R5343t2490 n5344 n2491 R=1.118e+01 
R5344t1937 n5345 n1938 R=2.762e+00 
R5344t193 n5345 n194 R=1.195e+02 
R5345t1552 n5346 n1553 R=1.346e+01 
R5345t4504 n5346 n4505 R=2.339e+00 
R5345t4771 n5346 n4772 R=9.553e+00 
R5346t3802 n5347 n3803 R=1.127e+01 
R5346t4677 n5347 n4678 R=3.711e+00 
R5346t8 n5347 n9 R=2.343e+01 
R5347t180 n5348 n181 R=1.685e+01 
R5347t4027 n5348 n4028 R=3.387e+00 
R5347t1564 n5348 n1565 R=1.739e+01 
R5348t1563 n5349 n1564 R=5.691e+00 
R5348t4868 n5349 n4869 R=2.830e+01 
R5349t5315 n5350 n5316 R=5.115e+00 
R5349t1455 n5350 n1456 R=9.432e+00 
R5349t4274 n5350 n4275 R=1.898e+01 
R5350t4497 n5351 n4498 R=3.870e+02 
R5350t4514 n5351 n4515 R=2.478e+00 
R5352t4759 n5353 n4760 R=1.109e+01 
R5352t2792 n5353 n2793 R=2.502e+01 
R5353t1621 n5354 n1622 R=6.837e+00 
R5353t4041 n5354 n4042 R=2.751e+01 
R5353t4564 n5354 n4565 R=2.384e+00 
R5353t3846 n5354 n3847 R=5.635e+00 
R5354t1436 n5355 n1437 R=1.097e+01 
R5354t4229 n5355 n4230 R=1.343e+01 
R5355t2642 n5356 n2643 R=3.235e+00 
R5355t7 n5356 n8 R=1.839e+01 
R5355t4993 n5356 n4994 R=7.880e+00 
R5355t5023 n5356 n5024 R=3.729e+01 
R5356t1948 n5357 n1949 R=2.441e+00 
R5356t3998 n5357 n3999 R=1.102e+01 
R5356t5264 n5357 n5265 R=3.094e+01 
R5357t2787 n5358 n2788 R=4.100e+00 
R5357t2994 n5358 n2995 R=4.780e+00 
R5357t3059 n5358 n3060 R=1.534e+01 
R5357t962 n5358 n963 R=1.071e+01 
R5358t2643 n5359 n2644 R=1.136e+01 
R5358t4020 n5359 n4021 R=4.845e+00 
R5358t1675 n5359 n1676 R=8.410e+00 
R5359t3405 n5360 n3406 R=6.165e+00 
R5359t3054 n5360 n3055 R=4.792e+01 
R5359t3572 n5360 n3573 R=2.058e+01 
R5360t3924 n5361 n3925 R=4.016e+00 
R5360t2522 n5361 n2523 R=8.605e+00 
R5361t1492 n5362 n1493 R=2.678e+01 
R5362t3086 n5363 n3087 R=3.725e+00 
R5362t741 n5363 n742 R=1.054e+02 
R5362t3814 n5363 n3815 R=3.952e+01 
R5362t1204 n5363 n1205 R=2.173e+01 
R5363t3565 n5364 n3566 R=8.544e+00 
R5363t4550 n5364 n4551 R=3.454e+00 
R5363t3959 n5364 n3960 R=2.005e+01 
R5363t1979 n5364 n1980 R=1.700e+01 
R5364t3575 n5365 n3576 R=6.008e+01 
R5364t3707 n5365 n3708 R=2.118e+00 
R5364t2926 n5365 n2927 R=6.474e+00 
R5364t2093 n5365 n2094 R=6.773e+01 
R5364t1423 n5365 n1424 R=1.377e+01 
R5365t4822 n5366 n4823 R=3.096e+00 
R5365t4397 n5366 n4398 R=3.834e+01 
R5365t1232 n5366 n1233 R=3.012e+00 
R5366t1695 n5367 n1696 R=9.106e+00 
R5366t1041 n5367 n1042 R=8.112e+00 
R5368t971 n5369 n972 R=6.515e+00 
R5368t2552 n5369 n2553 R=7.828e+01 
R5368t4223 n5369 n4224 R=1.072e+01 
R5368t4986 n5369 n4987 R=8.962e+00 
R5369t1364 n5370 n1365 R=1.632e+00 
R5369t2915 n5370 n2916 R=2.575e+01 
R5370t2051 n5371 n2052 R=6.033e+00 
R5370t2595 n5371 n2596 R=2.886e+00 
R5370t1252 n5371 n1253 R=1.337e+01 
R5370t4011 n5371 n4012 R=1.065e+01 
R5370t5318 n5371 n5319 R=6.133e+00 
R5371t2114 n5372 n2115 R=3.960e+00 
R5372t4149 n5373 n4150 R=2.521e+01 
R5372t4150 n5373 n4151 R=1.370e+02 
R5372t3873 n5373 n3874 R=4.999e+00 
R5372t2158 n5373 n2159 R=7.053e+00 
R5373t2131 n5374 n2132 R=2.964e+00 
R5373t3978 n5374 n3979 R=1.141e+01 
R5374t1836 n5375 n1837 R=5.889e+00 
R5374t3895 n5375 n3896 R=7.735e+00 
R5374t998 n5375 n999 R=3.098e+01 
R5374t76 n5375 n77 R=3.308e+01 
R5374t2975 n5375 n2976 R=1.515e+01 
R5374t4869 n5375 n4870 R=3.828e+00 
R5374t3860 n5375 n3861 R=2.499e+01 
R5374t3672 n5375 n3673 R=4.142e+01 
R5374t108 n5375 n109 R=8.891e+00 
R5375t696 n5376 n697 R=9.737e+00 
R5375t1079 n5376 n1080 R=2.735e+00 
R5375t4019 n5376 n4020 R=6.365e+01 
R5375t64 n5376 n65 R=6.554e+00 
R5375t4528 n5376 n4529 R=1.462e+01 
R5377t214 n5378 n215 R=6.320e+00 
R5377t3537 n5378 n3538 R=5.105e+00 
R5377t3474 n5378 n3475 R=5.255e+00 
R5378t5261 n5379 n5262 R=4.040e+00 
R5379t3715 n5380 n3716 R=1.825e+00 
R5379t5316 n5380 n5317 R=5.011e+01 
R5379t1313 n5380 n1314 R=1.252e+01 
R5379t236 n5380 n237 R=5.492e+00 
R5379t179 n5380 n180 R=5.139e+00 
R5380t3689 n5381 n3690 R=3.588e+00 
R5380t3002 n5381 n3003 R=2.313e+00 
R5380t1626 n5381 n1627 R=8.361e+00 
R5381t882 n5382 n883 R=2.345e+01 
R5381t4696 n5382 n4697 R=2.195e+01 
R5381t2034 n5382 n2035 R=7.637e+00 
R5382t2994 n5383 n2995 R=1.221e+01 
R5382t2563 n5383 n2564 R=9.593e+00 
R5383t3188 n5384 n3189 R=1.663e+01 
R5383t3452 n5384 n3453 R=3.826e+00 
R5383t4479 n5384 n4480 R=3.946e+00 
R5384t2213 n5385 n2214 R=9.936e+00 
R5384t339 n5385 n340 R=4.597e+01 
R5384t4063 n5385 n4064 R=1.197e+01 
R5385t1243 n5386 n1244 R=2.482e+01 
R5385t748 n5386 n749 R=5.509e+00 
R5385t3550 n5386 n3551 R=1.092e+01 
R5386t1261 n5387 n1262 R=3.612e+00 
R5386t4249 n5387 n4250 R=3.804e+00 
R5387t3348 n5388 n3349 R=6.092e+00 
R5387t1018 n5388 n1019 R=1.510e+01 
R5387t2057 n5388 n2058 R=4.147e+00 
R5387t5081 n5388 n5082 R=3.205e+01 
R5388t826 n5389 n827 R=6.368e+01 
R5388t3946 n5389 n3947 R=1.558e+01 
R5388t2508 n5389 n2509 R=1.019e+01 
R5388t2278 n5389 n2279 R=2.158e+00 
R5388t4349 n5389 n4350 R=3.669e+00 
R5389t3196 n5390 n3197 R=9.934e+00 
R5389t3203 n5390 n3204 R=6.851e+00 
R5389t4280 n5390 n4281 R=3.382e+01 
R5389t885 n5390 n886 R=4.205e+00 
R5390t3720 n5391 n3721 R=4.551e+00 
R5390t646 n5391 n647 R=1.031e+01 
R5390t1644 n5391 n1645 R=4.142e+00 
R5391t1228 n5392 n1229 R=7.763e+00 
R5391t2465 n5392 n2466 R=7.962e+00 
R5391t3688 n5392 n3689 R=5.681e+00 
R5391t2519 n5392 n2520 R=1.996e+01 
R5392t2208 n5393 n2209 R=2.025e+01 
R5392t2622 n5393 n2623 R=4.697e+00 
R5393t3767 n5394 n3768 R=4.144e+00 
R5393t3917 n5394 n3918 R=3.916e+02 
R5394t1005 n5395 n1006 R=3.437e+00 
R5394t3379 n5395 n3380 R=1.550e+01 
R5394t1885 n5395 n1886 R=1.136e+02 
R5395t943 n5396 n944 R=1.179e+02 
R5395t4639 n5396 n4640 R=1.543e+01 
R5395t4296 n5396 n4297 R=2.087e+00 
R5395t2805 n5396 n2806 R=9.277e+00 
R5395t3445 n5396 n3446 R=5.710e+01 
R5395t4268 n5396 n4269 R=2.733e+01 
R5396t4385 n5397 n1 R=7.583e+00 
R5396t210 n5397 n211 R=1.433e+01 
R5397t2994 n5398 n2995 R=4.852e+00 
R5397t5382 n5398 n5383 R=1.882e+01 
R5397t3059 n5398 n3060 R=3.789e+00 
R5397t5357 n5398 n5358 R=1.335e+01 
R5398t497 n5399 n498 R=2.472e+01 
R5399t423 n5400 n424 R=4.499e+00 
R5399t1360 n5400 n1361 R=1.073e+01 
R5399t65 n5400 n66 R=1.720e+02 
R5399t2929 n5400 n2930 R=6.460e+00 
R5399t3336 n5400 n3337 R=2.568e+00 
R5400t1039 n5401 n1040 R=8.092e+00 
R5400t3074 n5401 n3075 R=1.268e+00 
R5400t2163 n5401 n2164 R=2.604e+01 
R5400t3655 n5401 n3656 R=5.625e+00 
R5400t674 n5401 n675 R=5.309e+00 
R5401t2298 n5402 n2299 R=5.451e+00 
R5401t3595 n5402 n3596 R=2.610e+01 
R5401t3868 n5402 n3869 R=2.053e+01 
R5402t5360 n5403 n5361 R=2.351e+01 
R5402t3924 n5403 n3925 R=4.531e+00 
R5402t3819 n5403 n3820 R=1.864e+01 
R5402t4104 n5403 n4105 R=1.930e+01 
R5403t74 n5404 n75 R=1.641e+01 
R5403t841 n5404 n842 R=1.057e+02 
R5403t3809 n5404 n3810 R=5.114e+00 
R5404t4253 n5405 n4254 R=1.913e+02 
R5404t3563 n5405 n3564 R=2.058e+00 
R5404t939 n5405 n940 R=2.490e+00 
R5404t3414 n5405 n3415 R=8.422e+00 
R5405t371 n5406 n372 R=1.068e+01 
R5405t2538 n5406 n2539 R=4.269e+02 
R5405t5150 n5406 n5151 R=1.767e+01 
R5405t2901 n5406 n2902 R=4.373e+00 
R5406t1801 n5407 n1802 R=9.983e+00 
R5406t2768 n5407 n2769 R=8.567e+00 
R5406t1631 n5407 n1632 R=5.187e+00 
R5406t1214 n5407 n1215 R=2.841e+01 
R5407t605 n5408 n606 R=7.526e+00 
R5407t4379 n5408 n4380 R=2.448e+00 
R5407t2297 n5408 n2298 R=1.746e+02 
R5407t4736 n5408 n4737 R=2.004e+00 
R5407t683 n5408 n684 R=6.413e+01 
R5407t551 n5408 n552 R=1.475e+01 
R5408t1952 n5409 n1953 R=1.832e+01 
R5408t4013 n5409 n4014 R=1.042e+01 
R5408t326 n5409 n327 R=2.131e+00 
R5409t1333 n5410 n1334 R=4.372e+00 
R5409t5055 n5410 n5056 R=4.805e+00 
R5409t2759 n5410 n2760 R=6.157e+00 
R5409t4851 n5410 n4852 R=3.017e+00 
R5409t1685 n5410 n1686 R=5.199e+01 
R5410t5169 n5411 n5170 R=2.067e+01 
R5410t1965 n5411 n1966 R=7.734e+00 
R5410t4723 n5411 n4724 R=9.256e+00 
R5410t5106 n5411 n5107 R=6.343e+00 
R5411t2646 n5412 n2647 R=2.925e+00 
R5411t4650 n5412 n4651 R=6.978e+01 
R5411t3806 n5412 n3807 R=3.071e+00 
R5411t4583 n5412 n4584 R=5.727e+01 
R5411t656 n5412 n657 R=1.094e+02 
R5411t4906 n5412 n4907 R=1.713e+01 
R5412t408 n5413 n409 R=1.606e+02 
R5412t3888 n5413 n3889 R=2.339e+01 
R5413t2215 n5414 n2216 R=1.821e+01 
R5413t5004 n5414 n5005 R=3.724e+00 
R5413t4199 n5414 n4200 R=9.937e+00 
R5413t2224 n5414 n2225 R=9.185e+01 
R5414t139 n5415 n140 R=3.263e+00 
R5414t1747 n5415 n1748 R=1.293e+01 
R5414t3974 n5415 n3975 R=4.996e+01 
R5414t2815 n5415 n2816 R=4.194e+00 
R5415t3145 n5416 n3146 R=9.583e+00 
R5415t4381 n5416 n4382 R=4.968e+00 
R5416t3633 n5417 n3634 R=3.449e+00 
R5416t3882 n5417 n3883 R=7.648e+00 
R5417t2013 n5418 n2014 R=4.883e+00 
R5417t3745 n5418 n3746 R=2.791e+00 
R5417t3080 n5418 n3081 R=2.348e+00 
R5418t2634 n5419 n2635 R=7.618e+00 
R5418t4857 n5419 n4858 R=1.824e+01 
R5418t4143 n5419 n4144 R=6.970e+01 
R5418t834 n5419 n835 R=6.536e+00 
R5418t1874 n5419 n1875 R=7.896e+00 
R5419t3935 n5420 n3936 R=1.114e+01 
R5419t5189 n5420 n5190 R=1.962e+01 
R5419t2857 n5420 n2858 R=1.262e+01 
R5420t1636 n5421 n1637 R=3.903e+01 
R5420t3013 n5421 n3014 R=2.286e+00 
R5420t2812 n5421 n2813 R=1.033e+01 
R5420t5005 n5421 n5006 R=1.309e+01 
R5420t2878 n5421 n2879 R=2.534e+00 
R5421t3082 n5422 n3083 R=5.440e+00 
R5421t5162 n5422 n5163 R=2.577e+01 
R5421t3938 n5422 n3939 R=4.178e+00 
R5421t1088 n5422 n1089 R=7.321e+00 
R5422t1372 n5423 n1373 R=1.125e+01 
R5422t2954 n5423 n2955 R=5.221e+00 
R5422t3129 n5423 n3130 R=4.834e+00 
R5423t1369 n5424 n1370 R=9.130e+00 
R5423t1993 n5424 n1994 R=5.581e+00 
R5423t2612 n5424 n2613 R=8.786e+00 
R5423t1365 n5424 n1366 R=8.713e+02 
R5424t2137 n5425 n2138 R=1.784e+01 
R5424t3354 n5425 n3355 R=1.303e+01 
R5424t5026 n5425 n5027 R=2.136e+00 
R5425t939 n5426 n940 R=4.798e+00 
R5425t1230 n5426 n1231 R=5.052e+00 
R5426t2462 n5427 n2463 R=3.932e+00 
R5428t3414 n5429 n3415 R=4.136e+01 
R5428t4253 n5429 n4254 R=6.962e+00 
R5428t3032 n5429 n3033 R=3.333e+00 
R5429t2394 n5430 n2395 R=1.192e+01 
R5430t2240 n5431 n2241 R=1.277e+01 
R5430t694 n5431 n695 R=2.902e+00 
R5430t2105 n5431 n2106 R=5.661e+00 
R5431t1803 n5432 n1804 R=6.127e+00 
R5431t3920 n5432 n3921 R=3.740e+00 
R5431t1716 n5432 n1717 R=8.890e+01 
R5431t3240 n5432 n3241 R=4.428e+00 
R5431t5040 n5432 n5041 R=7.144e+00 
R5432t3933 n5433 n3934 R=4.232e+00 
R5432t4443 n5433 n4444 R=5.061e+00 
R5432t3981 n5433 n3982 R=5.844e+00 
R5433t2889 n5434 n2890 R=2.179e+00 
R5433t4938 n5434 n4939 R=6.233e+00 
R5434t2273 n5435 n2274 R=1.390e+01 
R5434t3910 n5435 n3911 R=4.394e+00 
R5434t851 n5435 n852 R=2.259e+01 
R5434t3500 n5435 n3501 R=6.110e+00 
R5435t2941 n5436 n2942 R=1.772e+01 
R5435t4480 n5436 n4481 R=3.124e+01 
R5435t2859 n5436 n2860 R=2.842e+00 
R5435t4795 n5436 n4796 R=8.548e+00 
R5436t1366 n5437 n1367 R=1.208e+01 
R5436t5245 n5437 n5246 R=1.413e+01 
R5436t3413 n5437 n3414 R=2.344e+00 
R5436t4439 n5437 n4440 R=3.895e+00 
R5436t741 n5437 n742 R=1.358e+02 
R5437t40 n5438 n41 R=1.139e+01 
R5437t1688 n5438 n1689 R=2.817e+00 
R5438t1268 n5439 n1269 R=4.119e+00 
R5438t4522 n5439 n4523 R=8.510e+00 
R5438t1787 n5439 n1788 R=2.191e+01 
R5438t2598 n5439 n2599 R=1.845e+00 
R5438t3232 n5439 n3233 R=5.206e+01 
R5438t4833 n5439 n4834 R=1.307e+01 
R5439t1135 n5440 n1136 R=5.063e+00 
R5441t111 n5442 n112 R=1.903e+00 
R5441t5025 n5442 n5026 R=2.092e+01 
R5442t2747 n5443 n1 R=2.663e+01 
R5442t2982 n5443 n2983 R=4.872e+00 
R5442t704 n5443 n705 R=7.329e+00 
R5442t1212 n5443 n1213 R=6.294e+00 
R5442t3767 n5443 n3768 R=6.438e+01 
R5443t1089 n5444 n1090 R=8.001e+00 
R5443t4757 n5444 n4758 R=3.666e+00 
R5443t736 n5444 n737 R=2.561e+01 
R5443t2920 n5444 n2921 R=1.794e+01 
R5444t1024 n5445 n1025 R=1.161e+01 
R5444t2985 n5445 n2986 R=2.269e+00 
R5444t1036 n5445 n1037 R=1.172e+02 
R5444t2199 n5445 n2200 R=4.525e+01 
R5444t19 n5445 n20 R=7.522e+00 
R5445t3933 n5446 n3934 R=4.295e+00 
R5445t2593 n5446 n2594 R=2.847e+01 
R5445t5007 n5446 n5008 R=3.583e+00 
R5445t3981 n5446 n3982 R=2.021e+01 
R5445t5432 n5446 n5433 R=1.739e+01 
R5446t1362 n5447 n1363 R=1.308e+01 
R5446t2790 n5447 n2791 R=8.778e+00 
R5446t2636 n5447 n2637 R=5.670e+00 
R5447t2684 n5448 n2685 R=7.293e+00 
R5447t915 n5448 n916 R=2.134e+01 
R5447t4950 n5448 n4951 R=3.417e+01 
R5448t2097 n5449 n2098 R=2.200e+01 
R5448t893 n5449 n894 R=4.161e+00 
R5448t2010 n5449 n2011 R=1.536e+01 
R5448t4228 n5449 n4229 R=1.827e+01 
R5449t1116 n5450 n1117 R=1.169e+01 
R5449t4543 n5450 n4544 R=1.074e+01 
R5449t2896 n5450 n2897 R=5.322e+00 
R5450t782 n5451 n783 R=6.083e+01 
R5450t4914 n5451 n4915 R=5.419e+00 
R5451t848 n5452 n849 R=1.507e+01 
R5451t1769 n5452 n1770 R=6.041e+00 
R5451t4718 n5452 n4719 R=2.191e+01 
R5451t1056 n5452 n1057 R=1.445e+01 
R5451t3301 n5452 n3302 R=5.370e+01 
R5451t2287 n5452 n2288 R=2.198e+01 
R5452t4151 n5453 n4152 R=2.037e+00 
R5452t2585 n5453 n2586 R=3.182e+00 
R5452t4866 n5453 n4867 R=1.940e+01 
R5453t5041 n5454 n5042 R=8.111e+01 
R5453t3142 n5454 n3143 R=1.433e+01 
R5453t1220 n5454 n1221 R=7.393e+00 
R5453t2080 n5454 n2081 R=6.550e+00 
R5453t1248 n5454 n1249 R=5.171e+00 
R5454t3298 n5455 n3299 R=2.730e+00 
R5454t5324 n5455 n5325 R=1.631e+01 
R5454t4848 n5455 n4849 R=1.217e+01 
R5454t1184 n5455 n1185 R=5.681e+00 
R5454t4881 n5455 n4882 R=1.800e+01 
R5455t262 n5456 n263 R=7.154e+00 
R5455t4873 n5456 n4874 R=6.898e+01 
R5455t3638 n5456 n3639 R=1.068e+01 
R5455t4425 n5456 n4426 R=2.388e+01 
R5455t4883 n5456 n4884 R=7.434e+00 
R5456t3172 n5457 n3173 R=1.859e+01 
R5456t2711 n5457 n2712 R=3.998e+00 
R5456t3592 n5457 n3593 R=1.889e+01 
R5456t3782 n5457 n3783 R=1.139e+01 
R5456t4732 n5457 n4733 R=2.072e+01 
R5457t1859 n5458 n1860 R=1.477e+01 
R5457t4239 n5458 n4240 R=5.752e+00 
R5457t835 n5458 n836 R=3.885e+00 
R5457t135 n5458 n136 R=3.600e+00 
R5458t2843 n5459 n2844 R=3.713e+00 
R5459t3548 n5460 n3549 R=2.884e+00 
R5459t5019 n5460 n5020 R=3.746e+01 
R5460t815 n5461 n816 R=8.707e+00 
R5460t4679 n5461 n4680 R=4.495e+00 
R5461t3387 n5462 n3388 R=1.387e+01 
R5461t3696 n5462 n3697 R=4.687e+00 
R5461t2069 n5462 n2070 R=2.707e+02 
R5461t4171 n5462 n4172 R=6.217e+00 
R5461t2137 n5462 n2138 R=2.154e+01 
R5462t4452 n1 n4453 R=2.030e+00 
R5463t5309 n5464 n5310 R=1.167e+01 
R5463t2766 n5464 n2767 R=4.498e+00 
R5463t4900 n5464 n4901 R=2.408e+01 
R5463t4012 n5464 n4013 R=4.148e+00 
R5464t5173 n5465 n5174 R=3.262e+00 
R5464t4155 n5465 n4156 R=8.810e+01 
R5464t3314 n5465 n3315 R=4.294e+00 
R5464t4188 n5465 n4189 R=6.841e+00 
R5465t2083 n5466 n2084 R=2.771e+00 
R5465t5327 n5466 n5328 R=1.764e+01 
R5465t2399 n5466 n2400 R=1.013e+01 
R5466t699 n5467 n700 R=1.398e+01 
R5466t2913 n5467 n2914 R=3.033e+02 
R5466t532 n5467 n533 R=2.340e+01 
R5466t3997 n5467 n3998 R=4.177e+00 
R5467t766 n5468 n767 R=2.906e+00 
R5467t1579 n5468 n1580 R=1.908e+01 
R5467t2065 n5468 n2066 R=1.705e+02 
R5467t3495 n5468 n3496 R=1.291e+01 
R5467t4023 n5468 n4024 R=1.707e+01 
R5468t447 n5469 n448 R=5.418e+00 
R5468t4648 n5469 n4649 R=1.647e+01 
R5468t1321 n5469 n1322 R=2.554e+01 
R5468t4209 n5469 n4210 R=4.252e+00 
R5469t4482 n5470 n4483 R=1.479e+00 
R5469t1090 n5470 n1091 R=2.951e+01 
R5470t2675 n5471 n2676 R=5.409e+00 
R5470t3465 n5471 n3466 R=2.151e+01 
R5470t2713 n5471 n2714 R=5.720e+00 
R5470t5106 n5471 n5107 R=3.711e+03 
R5470t775 n5471 n776 R=1.642e+01 
R5471t408 n5472 n409 R=1.054e+02 
R5471t5412 n5472 n5413 R=2.872e+00 
R5471t3888 n5472 n3889 R=5.420e+00 
R5471t1046 n5472 n1047 R=7.178e+01 
R5472t89 n5473 n90 R=2.992e+00 
R5472t3416 n5473 n3417 R=7.713e+00 
R5472t1648 n5473 n1649 R=8.066e+00 
R5472t1110 n5473 n1111 R=1.957e+01 
R5473t1859 n5474 n1860 R=3.512e+00 
R5473t5457 n5474 n5458 R=2.179e+01 
R5473t4239 n5474 n4240 R=3.161e+00 
R5474t4226 n5475 n4227 R=1.243e+00 
R5474t4445 n5475 n4446 R=1.484e+01 
R5474t442 n5475 n443 R=6.791e+01 
R5475t3872 n5476 n3873 R=6.266e+00 
R5475t1539 n5476 n1540 R=1.227e+01 
R5475t662 n5476 n663 R=6.520e+01 
R5476t992 n5477 n993 R=4.060e+01 
R5476t3192 n5477 n3193 R=2.519e+00 
R5476t5387 n5477 n5388 R=3.366e+01 
R5477t515 n5478 n516 R=8.748e+00 
R5477t3823 n5478 n3824 R=1.057e+01 
R5477t4058 n5478 n4059 R=2.380e+00 
R5478t1095 n5479 n1096 R=2.641e+01 
R5478t4407 n5479 n4408 R=3.655e+01 
R5478t4486 n5479 n4487 R=6.949e+00 
R5479t5422 n5480 n5423 R=1.079e+02 
R5479t2954 n5480 n2955 R=7.710e+00 
R5479t4297 n5480 n4298 R=9.266e+00 
R5479t2942 n5480 n2943 R=1.373e+01 
R5479t5303 n5480 n5304 R=2.098e+01 
R5480t4300 n5481 n4301 R=8.648e+00 
R5480t1072 n5481 n1073 R=1.165e+01 
R5480t3018 n5481 n3019 R=5.689e+00 
R5481t922 n5482 n923 R=1.784e+01 
R5481t4669 n5482 n4670 R=3.278e+01 
R5481t5423 n5482 n5424 R=3.968e+00 
R5481t3661 n5482 n3662 R=2.085e+01 
R5482t3316 n5483 n3317 R=1.543e+01 
R5483t1670 n5484 n1671 R=2.513e+01 
R5483t2247 n5484 n2248 R=4.764e+00 
R5483t2871 n5484 n2872 R=8.329e+00 
R5483t1084 n5484 n1085 R=5.502e+00 
R5483t2506 n5484 n2507 R=1.460e+01 
R5484t3367 n5485 n3368 R=4.239e+00 
R5484t4683 n5485 n4684 R=7.183e+00 
R5484t3185 n5485 n3186 R=9.880e+03 
R5485t4267 n5486 n4268 R=7.398e+00 
R5485t4762 n5486 n4763 R=4.037e+01 
R5486t322 n5487 n323 R=6.531e+00 
R5486t4329 n5487 n4330 R=3.155e+00 
R5487t5137 n5488 n5138 R=2.964e+00 
R5488t4461 n5489 n4462 R=1.192e+01 
R5488t1087 n5489 n1088 R=5.168e+00 
R5488t1134 n5489 n1135 R=3.702e+00 
R5489t459 n5490 n460 R=5.166e+00 
R5489t3602 n5490 n3603 R=8.913e+00 
R5489t4173 n5490 n4174 R=3.234e+00 
R5489t2660 n5490 n2661 R=2.598e+01 
R5490t4362 n5491 n4363 R=4.013e+00 
R5490t4616 n5491 n4617 R=7.560e+00 
R5490t3796 n5491 n3797 R=1.810e+01 
R5490t1650 n5491 n1651 R=1.240e+02 
R5491t305 n5492 n306 R=7.396e+00 
R5491t5083 n5492 n5084 R=4.049e+00 
R5491t570 n5492 n571 R=4.488e+00 
R5491t3531 n5492 n3532 R=6.218e+00 
R5492t4082 n5493 n4083 R=7.264e+00 
R5492t3479 n5493 n3480 R=1.322e+01 
R5492t2628 n5493 n2629 R=3.081e+00 
R5493t5300 n5494 n5301 R=5.617e+00 
R5493t1531 n5494 n1532 R=9.230e+00 
R5493t1609 n5494 n1610 R=2.645e+00 
R5494t3571 n5495 n3572 R=1.035e+01 
R5494t3289 n5495 n3290 R=4.827e+00 
R5495t4511 n5496 n4512 R=2.588e+00 
R5495t2637 n5496 n2638 R=3.174e+00 
R5495t3636 n5496 n3637 R=2.634e+01 
R5496t26 n5497 n27 R=7.611e+00 
R5496t819 n5497 n820 R=2.638e+00 
R5496t5262 n5497 n5263 R=3.894e+01 
R5496t3970 n5497 n3971 R=3.799e+00 
R5496t3208 n5497 n3209 R=1.550e+01 
R5497t456 n5498 n457 R=4.022e+01 
R5497t3569 n5498 n3570 R=3.144e+00 
R5497t457 n5498 n458 R=1.405e+01 
R5497t58 n5498 n59 R=9.702e+01 
R5498t4907 n5499 n4908 R=5.228e+00 
R5498t4047 n5499 n4048 R=9.395e+00 
R5498t4128 n5499 n4129 R=4.926e+01 
R5499t3213 n5500 n3214 R=2.054e+00 
R5499t4158 n5500 n4159 R=2.519e+02 
R5499t3145 n5500 n3146 R=4.590e+01 
R5499t2172 n5500 n2173 R=1.128e+01 
R5499t3877 n5500 n3878 R=1.835e+00 
R5500t3221 n5501 n3222 R=1.024e+01 
R5500t4184 n5501 n4185 R=2.343e+01 
R5500t3546 n5501 n3547 R=3.596e+01 
R5501t1319 n5502 n1320 R=3.125e+01 
R5501t4087 n5502 n4088 R=2.548e+00 
R5502t1841 n5503 n1842 R=2.434e+01 
R5502t774 n5503 n775 R=9.889e+00 
R5502t4889 n5503 n4890 R=5.772e+00 
R5502t2481 n5503 n2482 R=1.634e+01 
R5503t1037 n1 n1038 R=1.719e+00 
R5503t4202 n1 n4203 R=1.384e+01 
R5504t2720 n5505 n2721 R=6.082e+00 
R5504t4198 n5505 n4199 R=8.462e+00 
R5504t329 n5505 n330 R=8.534e+00 
R5504t3474 n5505 n3475 R=1.096e+01 
R5504t214 n5505 n215 R=3.031e+02 
R5506t2881 n5507 n2882 R=4.409e+00 
R5506t2936 n5507 n2937 R=5.717e+00 
R5506t3614 n5507 n3615 R=6.997e+00 
R5507t3581 n5508 n3582 R=7.067e+00 
R5507t3071 n5508 n3072 R=4.456e+00 
R5507t1369 n5508 n1370 R=4.267e+00 
R5508t2322 n5509 n2323 R=3.128e+01 
R5508t5263 n5509 n5264 R=2.871e+00 
R5508t518 n5509 n519 R=1.989e+01 
R5508t1762 n5509 n1763 R=1.561e+01 
R5509t1099 n5510 n1100 R=8.924e+00 
R5509t3017 n5510 n3018 R=7.340e+00 
R5510t3159 n5511 n3160 R=7.899e+00 
R5510t368 n5511 n369 R=4.632e+00 
R5511t3062 n5512 n3063 R=2.598e+00 
R5511t3629 n5512 n3630 R=9.650e+00 
R5512t2463 n5513 n2464 R=7.411e+00 
R5512t4633 n5513 n4634 R=6.196e+01 
R5512t1697 n5513 n1698 R=2.355e+00 
R5512t3741 n5513 n3742 R=6.739e+02 
R5512t4753 n5513 n4754 R=3.106e+01 
R5512t5275 n5513 n5276 R=9.516e+01 
R5513t1068 n5514 n1069 R=4.901e+02 
R5513t2556 n5514 n2557 R=1.049e+01 
R5513t4887 n5514 n4888 R=9.623e+00 
R5513t5064 n5514 n5065 R=4.294e+00 
R5513t3870 n5514 n3871 R=4.012e+00 
R5514t3393 n5515 n3394 R=2.924e+00 
R5514t4585 n5515 n4586 R=3.842e+00 
R5514t2875 n5515 n2876 R=1.625e+01 
R5515t2783 n5516 n2784 R=1.586e+01 
R5515t3995 n5516 n3996 R=1.298e+01 
R5515t5089 n5516 n5090 R=7.639e+02 
R5515t4031 n5516 n4032 R=1.775e+01 
R5515t2255 n5516 n2256 R=6.930e+00 
R5515t4164 n5516 n4165 R=1.246e+01 
R5515t2624 n5516 n2625 R=5.005e+00 
R5515t4304 n5516 n4305 R=3.149e+01 
R5516t152 n5517 n153 R=6.726e+00 
R5516t5009 n5517 n5010 R=8.223e+00 
R5516t1542 n5517 n1543 R=3.936e+00 
R5516t4579 n5517 n4580 R=1.037e+02 
R5517t4563 n5518 n4564 R=1.598e+01 
R5517t2065 n5518 n2066 R=4.567e+00 
R5517t5467 n5518 n5468 R=8.936e+00 
R5517t3495 n5518 n3496 R=7.410e+00 
R5518t5097 n5519 n5098 R=1.165e+01 
R5518t113 n5519 n114 R=1.343e+01 
R5518t1355 n5519 n1356 R=7.864e+00 
R5518t585 n5519 n586 R=6.275e+00 
R5519t4312 n5520 n4313 R=3.870e+00 
R5519t4468 n5520 n4469 R=7.293e+00 
R5519t578 n5520 n579 R=1.913e+02 
R5519t4503 n5520 n4504 R=3.771e+01 
R5519t341 n5520 n342 R=6.095e+00 
R5519t2582 n5520 n2583 R=9.011e+00 
R5520t2658 n5521 n2659 R=1.112e+01 
R5520t1714 n5521 n1715 R=3.885e+00 
R5520t4903 n5521 n4904 R=5.330e+00 
R5521t500 n5522 n501 R=3.915e+00 
R5521t1829 n5522 n1830 R=1.420e+01 
R5521t2119 n5522 n2120 R=9.201e+01 
R5522t2914 n5523 n2915 R=5.046e+00 
R5522t382 n5523 n383 R=5.554e+00 
R5522t606 n5523 n607 R=6.065e+00 
R5523t1376 n1 n1377 R=3.530e+00 
R5524t2958 n5525 n2959 R=8.568e+00 
R5524t4335 n5525 n4336 R=4.036e+00 
R5525t410 n5526 n411 R=3.272e+00 
R5525t4144 n5526 n4145 R=2.641e+01 
R5525t4952 n5526 n4953 R=1.790e+02 
R5526t4007 n5527 n4008 R=1.168e+01 
R5526t3820 n5527 n3821 R=3.900e+00 
R5527t733 n5528 n734 R=7.311e+00 
R5527t2007 n5528 n2008 R=2.305e+01 
R5527t3458 n5528 n3459 R=3.691e+00 
R5527t564 n5528 n565 R=8.008e+00 
R5527t6 n5528 n7 R=1.818e+01 
R5527t799 n5528 n800 R=2.055e+01 
R5527t2016 n5528 n2017 R=4.508e+00 
R5528t4328 n5529 n4329 R=1.222e+01 
R5528t1043 n5529 n1044 R=2.877e+00 
R5528t5091 n5529 n5092 R=9.158e+01 
R5528t3318 n5529 n3319 R=4.910e+01 
R5528t519 n5529 n520 R=3.645e+00 
R5529t1213 n5530 n1214 R=1.140e+01 
R5529t2712 n5530 n2713 R=6.444e+00 
R5529t5045 n5530 n5046 R=7.327e+00 
R5529t2699 n5530 n2700 R=7.392e+00 
R5529t5333 n5530 n5334 R=4.480e+01 
R5529t4678 n5530 n4679 R=2.437e+01 
R5530t4240 n5531 n4241 R=3.231e+01 
R5530t807 n5531 n808 R=2.992e+00 
R5530t4947 n5531 n4948 R=3.731e+01 
R5531t4104 n5532 n4105 R=9.803e+01 
R5531t4981 n5532 n4982 R=6.220e+00 
R5531t2871 n5532 n2872 R=1.652e+01 
R5531t2247 n5532 n2248 R=4.543e+00 
R5531t3819 n5532 n3820 R=5.954e+00 
R5531t5402 n5532 n5403 R=5.929e+00 
R5532t722 n5533 n723 R=3.032e+00 
R5532t4796 n5533 n4797 R=2.357e+01 
R5533t2367 n5534 n2368 R=4.441e+00 
R5533t676 n5534 n677 R=6.877e+00 
R5534t3081 n5535 n3082 R=4.746e+00 
R5534t2086 n5535 n2087 R=8.747e+00 
R5535t970 n5536 n971 R=5.185e+00 
R5535t2455 n5536 n2456 R=8.607e+00 
R5536t1341 n5537 n1342 R=4.663e+01 
R5536t2864 n5537 n2865 R=4.765e+00 
R5536t1231 n5537 n1232 R=5.909e+00 
R5536t5121 n5537 n5122 R=8.189e+00 
R5537t852 n5538 n853 R=2.557e+00 
R5537t3846 n5538 n3847 R=2.244e+02 
R5537t2613 n5538 n2614 R=7.355e+00 
R5537t31 n5538 n32 R=5.650e+00 
R5537t589 n5538 n590 R=5.599e+00 
R5538t667 n5539 n668 R=1.045e+01 
R5539t667 n5540 n668 R=3.185e+00 
R5539t1220 n5540 n1221 R=1.422e+02 
R5539t3142 n5540 n3143 R=1.020e+01 
R5539t5453 n5540 n5454 R=3.093e+00 
R5540t2217 n5541 n2218 R=2.088e+01 
R5540t2940 n5541 n2941 R=7.727e+00 
R5540t663 n5541 n664 R=6.314e+00 
R5540t984 n5541 n985 R=8.770e+00 
R5540t4533 n5541 n4534 R=5.664e+00 
R5541t2832 n5542 n2833 R=6.591e+00 
R5541t3507 n5542 n3508 R=1.696e+01 
R5541t4568 n5542 n4569 R=5.758e+00 
R5541t4501 n5542 n4502 R=9.552e+00 
R5542t2165 n5543 n2166 R=3.699e+00 
R5542t782 n5543 n783 R=1.496e+01 
R5542t5450 n5543 n5451 R=1.711e+01 
R5542t4808 n5543 n4809 R=1.057e+01 
R5542t3761 n5543 n3762 R=1.300e+01 
R5543t3012 n5544 n3013 R=5.289e+00 
R5543t1277 n5544 n1278 R=3.753e+01 
R5543t4341 n5544 n4342 R=9.242e+00 
R5544t3968 n5545 n3969 R=1.247e+01 
R5544t4804 n5545 n4805 R=1.092e+02 
R5544t2152 n5545 n2153 R=3.769e+00 
R5544t3578 n5545 n3579 R=1.181e+03 
R5544t3033 n5545 n3034 R=3.035e+01 
R5545t3253 n5546 n3254 R=6.691e+00 
R5545t757 n5546 n758 R=3.528e+00 
R5545t3127 n5546 n3128 R=1.428e+01 
R5545t4250 n5546 n4251 R=8.418e+00 
R5546t3714 n5547 n3715 R=1.134e+01 
R5547t687 n5548 n688 R=2.105e+01 
R5547t4646 n5548 n4647 R=2.064e+00 
R5548t888 n5549 n889 R=8.230e+00 
R5549t1760 n5550 n1761 R=7.343e+01 
R5549t1962 n5550 n1963 R=2.202e+00 
R5549t2142 n5550 n2143 R=2.668e+00 
R5550t447 n5551 n448 R=2.189e+01 
R5550t3184 n5551 n3185 R=2.317e+00 
R5550t1121 n5551 n1122 R=3.242e+01 
R5550t4648 n5551 n4649 R=5.991e+01 
R5551t4508 n5552 n4509 R=3.954e+00 
R5551t3049 n5552 n3050 R=6.132e+00 
R5552t606 n5553 n607 R=3.081e+00 
R5552t2437 n5553 n2438 R=1.058e+01 
R5552t4742 n5553 n4743 R=6.381e+00 
R5552t382 n5553 n383 R=5.085e+00 
R5554t1941 n5555 n1942 R=5.879e+00 
R5554t2228 n5555 n2229 R=4.731e+01 
R5554t3077 n5555 n3078 R=1.937e+01 
R5555t1319 n5556 n1320 R=1.036e+01 
R5555t5501 n5556 n5502 R=5.211e+00 
R5555t4960 n5556 n4961 R=3.388e+00 
R5555t1117 n5556 n1118 R=8.566e+00 
R5555t4087 n5556 n4088 R=1.935e+01 
R5556t3348 n5557 n3349 R=1.621e+01 
R5556t5387 n5557 n5388 R=6.643e+01 
R5556t1018 n5557 n1019 R=2.842e+00 
R5556t2444 n5557 n2445 R=5.130e+00 
R5557t4879 n5558 n4880 R=7.499e+00 
R5557t4744 n5558 n4745 R=1.959e+01 
R5557t718 n5558 n719 R=3.865e+00 
R5557t1248 n5558 n1249 R=6.529e+01 
R5557t2080 n5558 n2081 R=6.596e+00 
R5557t327 n5558 n328 R=3.728e+01 
R5558t4104 n5559 n4105 R=4.850e+00 
R5558t1281 n5559 n1282 R=8.101e+00 
R5559t4434 n5560 n4435 R=5.146e+00 
R5559t5521 n5560 n5522 R=2.807e+00 
R5559t2119 n5560 n2120 R=6.078e+00 
R5560t3298 n5561 n3299 R=1.810e+01 
R5560t5454 n5561 n5455 R=1.485e+01 
R5560t3222 n5561 n3223 R=1.135e+01 
R5560t3026 n5561 n3027 R=4.448e+00 
R5560t5324 n5561 n5325 R=5.254e+00 
R5561t2672 n5562 n2673 R=6.516e+00 
R5561t1851 n5562 n1852 R=3.385e+00 
R5562t3271 n5563 n3272 R=3.805e+00 
R5562t614 n5563 n615 R=4.513e+00 
R5563t4261 n5564 n4262 R=3.372e+00 
R5563t3486 n5564 n3487 R=5.896e+01 
R5563t5120 n5564 n5121 R=5.792e+00 
R5564t15 n5565 n16 R=2.530e+00 
R5564t2264 n5565 n2265 R=5.453e+00 
R5564t4938 n5565 n4939 R=5.342e+00 
R5564t2231 n5565 n2232 R=9.119e+01 
R5564t1975 n5565 n1976 R=3.081e+02 
R5565t5151 n5566 n5152 R=7.157e+00 
R5566t310 n5567 n311 R=7.849e+00 
R5566t1472 n5567 n1473 R=3.303e+00 
R5566t1869 n5567 n1870 R=1.299e+01 
R5566t4602 n5567 n4603 R=4.204e+01 
R5567t4745 n5568 n4746 R=7.210e+00 
R5567t945 n5568 n946 R=5.680e+00 
R5567t2059 n5568 n2060 R=1.145e+01 
R5568t1112 n5569 n1113 R=2.805e+00 
R5568t1168 n5569 n1169 R=1.883e+01 
R5568t2458 n5569 n2459 R=1.743e+01 
R5568t5482 n5569 n5483 R=4.866e+00 
R5569t3782 n5570 n3783 R=5.072e+00 
R5569t3592 n5570 n3593 R=6.322e+00 
R5569t5456 n5570 n5457 R=7.392e+00 
R5571t1701 n5572 n1702 R=3.607e+00 
R5571t2989 n5572 n2990 R=1.453e+01 
R5571t2947 n5572 n2948 R=5.436e+00 
R5572t4932 n5573 n4933 R=1.537e+01 
R5572t4032 n5573 n4033 R=6.606e+00 
R5572t1389 n5573 n1390 R=2.341e+02 
R5572t4218 n5573 n4219 R=2.118e+01 
R5573t1167 n5574 n1168 R=3.320e+00 
R5574t2754 n5575 n2755 R=1.530e+01 
R5574t4607 n5575 n4608 R=3.434e+01 
R5575t4826 n5576 n4827 R=7.025e+00 
R5575t2732 n5576 n2733 R=6.072e+00 
R5575t1553 n5576 n1554 R=1.247e+01 
R5576t3445 n5577 n3446 R=4.372e+00 
R5576t4268 n5577 n4269 R=8.037e+00 
R5576t3178 n5577 n3179 R=1.184e+01 
R5577t3200 n5578 n3201 R=1.474e+01 
R5577t4860 n5578 n4861 R=7.921e+00 
R5577t2654 n5578 n2655 R=1.681e+01 
R5578t4997 n5579 n4998 R=4.617e+00 
R5578t4570 n5579 n4571 R=6.689e+00 
R5579t2374 n5580 n2375 R=4.552e+00 
R5579t1479 n5580 n1480 R=2.745e+01 
R5580t1926 n5581 n1927 R=1.020e+01 
R5580t1396 n5581 n1397 R=1.656e+01 
R5580t636 n5581 n637 R=1.056e+01 
R5580t3538 n5581 n3539 R=8.232e+00 
R5581t3101 n5582 n3102 R=9.670e+00 
R5581t5138 n5582 n5139 R=6.323e+01 
R5581t4628 n5582 n4629 R=5.891e+00 
R5581t395 n5582 n396 R=2.987e+01 
R5581t1011 n5582 n1012 R=2.525e+00 
R5582t4397 n5583 n4398 R=8.372e+00 
R5582t3651 n5583 n3652 R=1.210e+01 
R5582t4351 n5583 n4352 R=1.726e+01 
R5582t1075 n5583 n1076 R=5.379e+00 
R5582t333 n5583 n334 R=1.729e+01 
R5583t2340 n5584 n2341 R=2.041e+01 
R5583t341 n5584 n342 R=6.669e+00 
R5583t3439 n5584 n3440 R=3.501e+00 
R5584t5035 n5585 n5036 R=1.431e+01 
R5584t3918 n5585 n3919 R=1.330e+02 
R5584t542 n5585 n543 R=2.085e+01 
R5584t690 n5585 n691 R=2.293e+00 
R5584t1356 n5585 n1357 R=5.328e+00 
R5585t3265 n5586 n3266 R=9.707e+00 
R5585t3078 n5586 n3079 R=2.335e+01 
R5585t1346 n5586 n1347 R=3.991e+00 
R5585t2922 n5586 n2923 R=1.914e+01 
R5586t648 n5587 n649 R=3.506e+00 
R5586t272 n5587 n273 R=4.366e+00 
R5587t5192 n5588 n5193 R=2.023e+00 
R5587t4950 n5588 n4951 R=1.049e+01 
R5587t2131 n5588 n2132 R=9.870e+00 
R5588t1545 n5589 n1546 R=4.239e+00 
R5588t2823 n5589 n2824 R=1.801e+01 
R5588t2948 n5589 n2949 R=2.589e+01 
R5588t339 n5589 n340 R=9.271e+00 
R5588t5384 n5589 n5385 R=8.777e+00 
R5589t5361 n5590 n5362 R=5.668e+00 
R5589t4551 n5590 n4552 R=3.080e+00 
R5589t5170 n5590 n5171 R=1.522e+01 
R5590t1928 n5591 n1929 R=2.911e+00 
R5590t337 n5591 n338 R=3.237e+00 
R5591t175 n5592 n176 R=1.738e+01 
R5591t3463 n5592 n3464 R=8.603e+00 
R5591t4993 n5592 n4994 R=1.231e+01 
R5591t3490 n5592 n3491 R=1.196e+01 
R5591t501 n5592 n502 R=1.036e+01 
R5591t1051 n5592 n1052 R=5.003e+00 
R5592t4053 n5593 n4054 R=1.025e+01 
R5592t5498 n5593 n5499 R=3.537e+00 
R5593t3218 n5594 n3219 R=1.643e+01 
R5593t4961 n5594 n4962 R=6.120e+00 
R5594t1800 n5595 n1801 R=4.226e+01 
R5594t3211 n5595 n3212 R=2.881e+00 
R5595t1310 n5596 n1311 R=2.049e+00 
R5595t4302 n5596 n4303 R=2.715e+01 
R5595t1518 n5596 n1519 R=3.817e+00 
R5596t1423 n5597 n1424 R=3.491e+00 
R5596t3707 n5597 n3708 R=3.152e+00 
R5597t2174 n5598 n2175 R=3.926e+00 
R5597t255 n5598 n256 R=1.723e+01 
R5598t807 n5599 n808 R=3.827e+01 
R5598t4038 n5599 n4039 R=6.136e+01 
R5598t5530 n5599 n5531 R=1.056e+01 
R5598t3334 n5599 n3335 R=8.972e+01 
R5598t3323 n5599 n3324 R=6.594e+00 
R5599t3171 n5600 n3172 R=1.749e+01 
R5599t3580 n5600 n3581 R=2.580e+00 
R5599t1252 n5600 n1253 R=1.600e+01 
R5600t2258 n5601 n2259 R=4.699e+00 
R5600t3900 n5601 n3901 R=8.319e+00 
R5600t4369 n5601 n4370 R=1.753e+01 
R5600t555 n5601 n556 R=1.091e+01 
R5600t5236 n5601 n5237 R=1.092e+01 
R5600t3397 n5601 n3398 R=1.242e+01 
R5601t451 n5602 n452 R=7.736e+00 
R5601t5232 n5602 n5233 R=4.345e+00 
R5602t3796 n1 n3797 R=1.748e+01 
R5603t225 n5604 n226 R=1.057e+01 
R5603t4765 n5604 n4766 R=1.712e+01 
R5603t1732 n5604 n1733 R=7.111e+00 
R5604t2319 n5605 n2320 R=4.687e+00 
R5605t3188 n5606 n3189 R=4.183e+01 
R5605t5383 n5606 n5384 R=9.333e+01 
R5605t3452 n5606 n3453 R=5.711e+00 
R5605t3847 n5606 n3848 R=8.440e+00 
R5605t4890 n5606 n4891 R=6.375e+00 
R5606t2218 n5607 n2219 R=6.226e+00 
R5606t4193 n5607 n4194 R=1.487e+01 
R5606t2797 n5607 n2798 R=8.760e+00 
R5606t787 n5607 n788 R=3.220e+01 
R5606t2471 n5607 n2472 R=6.003e+00 
R5607t3062 n5608 n3063 R=1.667e+01 
R5607t2033 n5608 n2034 R=1.594e+01 
R5607t1962 n5608 n1963 R=4.905e+00 
R5607t1746 n5608 n1747 R=2.556e+00 
R5608t812 n5609 n813 R=4.595e+01 
R5608t3279 n5609 n3280 R=2.326e+00 
R5609t94 n5610 n95 R=1.617e+01 
R5609t5142 n5610 n5143 R=1.020e+01 
R5609t2978 n5610 n2979 R=9.513e+00 
R5609t1127 n5610 n1128 R=4.412e+00 
R5610t1916 n5611 n1917 R=3.584e+00 
R5610t3939 n5611 n3940 R=3.296e+01 
R5610t646 n5611 n647 R=1.211e+02 
R5610t5390 n5611 n5391 R=2.419e+01 
R5611t4076 n5612 n4077 R=4.686e+00 
R5611t4373 n5612 n4374 R=3.231e+00 
R5612t4182 n5613 n4183 R=4.242e+00 
R5613t4480 n5614 n4481 R=1.484e+01 
R5613t1779 n5614 n1 R=4.010e+00 
R5613t2727 n5614 n2728 R=6.488e+00 
R5614t355 n5615 n356 R=7.213e+01 
R5614t4423 n5615 n4424 R=4.856e+00 
R5614t1083 n5615 n1084 R=3.740e+00 
R5614t4377 n5615 n4378 R=8.895e+00 
R5615t2931 n5616 n2932 R=5.197e+00 
R5615t2881 n5616 n2882 R=5.844e+00 
R5615t5506 n5616 n5507 R=3.081e+01 
R5615t2936 n5616 n2937 R=6.355e+00 
R5616t2312 n5617 n2313 R=4.986e+00 
R5616t3200 n5617 n3201 R=6.716e+00 
R5616t5078 n5617 n5079 R=1.123e+02 
R5616t110 n5617 n111 R=3.564e+01 
R5616t3104 n5617 n3105 R=3.401e+00 
R5617t3128 n5618 n3129 R=1.144e+01 
R5617t3669 n5618 n3670 R=8.484e+00 
R5617t2172 n5618 n2173 R=3.287e+00 
R5617t3365 n5618 n3366 R=3.263e+00 
R5618t606 n5619 n607 R=1.112e+01 
R5618t2437 n5619 n2438 R=8.204e+00 
R5618t2743 n5619 n2744 R=3.509e+02 
R5618t5129 n5619 n5130 R=5.255e+00 
R5618t4696 n5619 n4697 R=4.683e+02 
R5618t5095 n5619 n5096 R=6.439e+00 
R5620t3976 n5621 n3977 R=3.427e+00 
R5620t2974 n5621 n2975 R=1.234e+02 
R5620t4288 n5621 n4289 R=2.471e+01 
R5621t812 n5622 n813 R=2.501e+01 
R5621t4846 n5622 n4847 R=4.497e+00 
R5622t1536 n5623 n1537 R=2.702e+00 
R5622t4645 n5623 n4646 R=9.064e+01 
R5622t1520 n5623 n1521 R=7.839e+00 
R5622t2184 n5623 n2185 R=1.528e+01 
R5623t617 n5624 n618 R=2.297e+01 
R5623t4940 n5624 n4941 R=4.978e+00 
R5623t2290 n5624 n2291 R=1.132e+02 
R5623t4422 n5624 n4423 R=8.296e+00 
R5624t4258 n5625 n4259 R=2.417e+01 
R5624t95 n5625 n96 R=3.138e+00 
R5624t1789 n5625 n1790 R=1.202e+01 
R5625t4492 n5626 n4493 R=1.916e+01 
R5625t2594 n5626 n2595 R=4.632e+00 
R5626t2201 n5627 n2202 R=7.465e+00 
R5627t3875 n5628 n3876 R=8.019e+01 
R5627t1247 n5628 n1248 R=7.112e+00 
R5627t4022 n5628 n4023 R=6.558e+01 
R5627t4715 n5628 n4716 R=3.558e+00 
R5627t258 n5628 n259 R=3.411e+01 
R5628t3964 n5629 n3965 R=2.629e+01 
R5628t5232 n5629 n5233 R=6.776e+00 
R5628t3842 n5629 n3843 R=1.509e+01 
R5628t3044 n5629 n3045 R=3.833e+00 
R5629t1194 n5630 n1195 R=6.062e+00 
R5629t2983 n5630 n2984 R=1.264e+01 
R5629t1736 n5630 n1737 R=6.742e+00 
R5630t1205 n5631 n1206 R=2.285e+02 
R5630t4370 n5631 n4371 R=1.207e+01 
R5631t490 n5632 n491 R=1.579e+00 
R5631t1040 n5632 n1041 R=1.958e+01 
R5632t500 n5633 n501 R=3.784e+00 
R5632t4688 n5633 n4689 R=3.327e+00 
R5632t3694 n5633 n3695 R=1.327e+02 
R5632t4382 n5633 n4383 R=8.361e+00 
R5633t5292 n5634 n5293 R=1.274e+01 
R5633t5419 n5634 n5420 R=1.358e+01 
R5634t178 n5635 n179 R=1.179e+01 
R5634t5132 n5635 n5133 R=6.516e+00 
R5634t4781 n5635 n4782 R=2.011e+01 
R5634t5371 n5635 n5372 R=2.677e+00 
R5634t2114 n5635 n2115 R=3.612e+01 
R5634t5144 n5635 n5145 R=1.673e+01 
R5635t4914 n5636 n4915 R=2.064e+02 
R5635t4214 n5636 n4215 R=5.047e+00 
R5635t3709 n5636 n3710 R=1.429e+01 
R5635t2443 n5636 n2444 R=4.903e+00 
R5636t3768 n5637 n3769 R=3.710e+00 
R5636t1202 n5637 n1203 R=4.563e+00 
R5638t1059 n5639 n1060 R=8.976e+01 
R5638t4383 n5639 n4384 R=6.150e+00 
R5638t4776 n5639 n4777 R=3.290e+00 
R5640t5408 n5641 n5409 R=6.171e+01 
R5641t2741 n5642 n2742 R=8.332e+00 
R5641t5421 n5642 n5422 R=3.085e+01 
R5641t1088 n5642 n1089 R=2.907e+01 
R5641t1409 n5642 n1410 R=4.228e+00 
R5642t4384 n5643 n4385 R=6.985e+00 
R5642t2977 n5643 n2978 R=2.788e+00 
R5642t3255 n5643 n3256 R=2.813e+03 
R5642t1122 n5643 n1123 R=6.495e+00 
R5643t4212 n5644 n4213 R=2.716e+00 
R5643t5241 n5644 n5242 R=1.263e+01 
R5643t4893 n5644 n4894 R=1.294e+01 
R5644t2671 n5645 n2672 R=2.141e+00 
R5644t811 n5645 n812 R=1.230e+01 
R5644t3577 n5645 n3578 R=5.807e+01 
R5644t3687 n5645 n3688 R=9.321e+00 
R5644t2197 n5645 n2198 R=4.329e+00 
R5645t497 n5646 n498 R=3.358e+00 
R5645t1091 n5646 n1092 R=9.645e+00 
R5645t3447 n5646 n3448 R=1.323e+03 
R5645t4638 n5646 n4639 R=7.399e+00 
R5645t4650 n5646 n4651 R=5.838e+00 
R5646t1915 n5647 n1916 R=1.211e+01 
R5647t52 n5648 n53 R=1.477e+01 
R5647t4816 n5648 n4817 R=1.594e+01 
R5647t3682 n5648 n3683 R=5.922e+00 
R5647t2296 n5648 n2297 R=5.936e+00 
R5647t823 n5648 n824 R=5.816e+00 
R5648t2384 n5649 n2385 R=8.458e+00 
R5648t2783 n5649 n2784 R=1.001e+01 
R5648t2932 n5649 n2933 R=5.818e+00 
R5648t769 n5649 n770 R=2.184e+01 
R5648t1683 n5649 n1684 R=7.759e+00 
R5649t49 n5650 n50 R=9.271e+00 
R5649t3978 n5650 n3979 R=7.010e+00 
R5649t5373 n5650 n5374 R=2.980e+00 
R5650t3172 n5651 n3173 R=8.232e+00 
R5650t1507 n5651 n1508 R=2.894e+00 
R5650t1580 n5651 n1581 R=7.336e+01 
R5651t63 n5652 n64 R=1.937e+01 
R5651t3487 n5652 n3488 R=3.491e+00 
R5651t2750 n5652 n2751 R=2.841e+00 
R5651t4731 n5652 n4732 R=9.452e+00 
R5652t235 n5653 n236 R=3.273e+00 
R5652t2673 n5653 n2674 R=4.138e+00 
R5653t2182 n5654 n2183 R=3.521e+00 
R5653t2235 n5654 n2236 R=7.000e+00 
R5653t3826 n5654 n3827 R=4.039e+01 
R5653t1907 n5654 n1908 R=3.123e+00 
R5653t399 n5654 n400 R=1.796e+01 
R5653t2584 n5654 n2585 R=1.138e+01 
R5654t739 n5655 n740 R=4.825e+00 
R5654t1474 n5655 n1475 R=7.247e+00 
R5655t3821 n5656 n3822 R=2.204e+01 
R5655t1704 n5656 n1705 R=2.342e+01 
R5655t4246 n5656 n4247 R=1.895e+01 
R5655t3154 n5656 n3155 R=1.251e+01 
R5656t1188 n5657 n1189 R=8.106e+00 
R5656t1187 n5657 n1188 R=9.609e+00 
R5656t1320 n5657 n1321 R=5.493e+00 
R5657t3114 n5658 n3115 R=3.725e+00 
R5657t3420 n5658 n3421 R=1.194e+02 
R5658t3204 n5659 n3205 R=1.001e+01 
R5658t227 n5659 n228 R=1.764e+01 
R5658t1762 n5659 n1763 R=4.496e+00 
R5659t2312 n5660 n2313 R=8.363e+00 
R5659t2812 n5660 n2813 R=5.312e+00 
R5660t2846 n5661 n2847 R=3.563e+01 
R5660t2528 n5661 n2529 R=5.619e+00 
R5660t671 n5661 n672 R=1.929e+01 
R5660t2487 n5661 n2488 R=1.244e+01 
R5661t3611 n5662 n3612 R=1.490e+01 
R5661t5238 n5662 n5239 R=6.500e+01 
R5661t1907 n5662 n1908 R=3.375e+00 
R5661t3826 n5662 n3827 R=3.516e+01 
R5661t5193 n5662 n5194 R=5.292e+00 
R5662t4523 n5663 n4524 R=5.230e+00 
R5662t1345 n5663 n1346 R=2.867e+00 
R5663t2872 n5664 n2873 R=2.953e+00 
R5663t4875 n5664 n4876 R=6.256e+00 
R5663t3075 n5664 n3076 R=2.407e+00 
R5664t574 n5665 n575 R=1.053e+01 
R5664t4024 n5665 n4025 R=2.237e+01 
R5665t5332 n5666 n5333 R=1.913e+01 
R5665t618 n5666 n619 R=6.689e+01 
R5666t4775 n5667 n4776 R=4.741e+00 
R5667t49 n5668 n50 R=7.737e+00 
R5667t934 n5668 n935 R=1.460e+01 
R5667t2665 n5668 n2666 R=3.215e+00 
R5668t1299 n5669 n1300 R=6.310e+00 
R5668t2219 n5669 n2220 R=1.595e+01 
R5668t1516 n5669 n1517 R=1.494e+01 
R5668t4690 n5669 n4691 R=9.530e+00 
R5669t2549 n5670 n2550 R=1.352e+01 
R5669t5212 n5670 n5213 R=1.971e+01 
R5669t2680 n5670 n2681 R=1.078e+02 
R5669t672 n5670 n673 R=7.998e+00 
R5670t1993 n5671 n1994 R=7.946e+00 
R5670t2612 n5671 n2613 R=1.092e+01 
R5670t2644 n5671 n2645 R=5.981e+00 
R5670t3071 n5671 n3072 R=3.796e+00 
R5671t5367 n5672 n5368 R=1.432e+01 
R5671t2906 n5672 n2907 R=2.061e+01 
R5671t2126 n5672 n2127 R=3.702e+00 
R5671t2344 n5672 n2345 R=2.780e+01 
R5671t246 n5672 n247 R=1.319e+01 
R5672t4584 n5673 n4585 R=5.531e+00 
R5672t4830 n5673 n4831 R=4.756e+00 
R5672t834 n5673 n835 R=2.785e+01 
R5672t1874 n5673 n1875 R=7.331e+00 
R5672t3268 n5673 n3269 R=1.815e+01 
R5673t3870 n5674 n3871 R=3.685e+00 
R5673t36 n5674 n37 R=3.084e+00 
R5674t2018 n5675 n2019 R=2.097e+01 
R5674t1660 n5675 n1661 R=4.064e+00 
R5674t4913 n5675 n4914 R=6.956e+00 
R5674t281 n5675 n282 R=9.045e+00 
R5674t477 n5675 n478 R=2.895e+00 
R5675t1236 n5676 n1237 R=5.648e+00 
R5675t1611 n5676 n1612 R=5.179e+01 
R5675t3288 n5676 n3289 R=3.197e+00 
R5675t3293 n5676 n3294 R=6.353e+00 
R5676t1622 n5677 n1623 R=9.074e+00 
R5676t3332 n5677 n3333 R=7.788e+00 
R5676t571 n5677 n572 R=1.964e+01 
R5677t586 n5678 n587 R=6.474e+00 
R5677t3179 n5678 n3180 R=7.831e+00 
R5677t981 n5678 n982 R=4.081e+00 
R5677t3497 n5678 n3498 R=9.393e+01 
R5678t2789 n5679 n2790 R=1.163e+01 
R5678t2972 n5679 n2973 R=2.722e+00 
R5678t2475 n5679 n2476 R=5.864e+00 
R5679t3421 n5680 n3422 R=7.150e+00 
R5679t3659 n5680 n3660 R=8.472e+00 
R5679t4940 n5680 n4941 R=2.598e+00 
R5679t4378 n5680 n4379 R=2.662e+01 
R5680t5534 n5681 n5535 R=1.313e+01 
R5680t3081 n5681 n3082 R=8.785e+00 
R5680t84 n5681 n85 R=5.517e+00 
R5681t1073 n5682 n1074 R=1.116e+01 
R5681t4688 n5682 n4689 R=4.164e+01 
R5681t3944 n5682 n3945 R=1.874e+00 
R5681t661 n5682 n662 R=1.384e+02 
R5682t5678 n5683 n5679 R=6.918e+00 
R5682t2475 n5683 n2476 R=1.238e+01 
R5682t644 n5683 n645 R=1.554e+01 
R5682t1129 n5683 n1130 R=1.396e+01 
R5682t2254 n5683 n2255 R=4.645e+00 
R5683t26 n5684 n27 R=5.941e+00 
R5683t803 n5684 n804 R=6.942e+00 
R5683t1501 n5684 n1502 R=1.729e+01 
R5684t4107 n5685 n4108 R=9.391e+00 
R5684t4144 n5685 n4145 R=1.810e+01 
R5684t410 n5685 n411 R=5.113e+00 
R5685t3994 n5686 n3995 R=1.405e+02 
R5685t858 n5686 n859 R=1.917e+00 
R5686t4866 n5687 n4867 R=1.533e+01 
R5686t5452 n5687 n5453 R=8.814e+00 
R5686t1138 n5687 n1139 R=1.174e+01 
R5686t3746 n5687 n3747 R=5.514e+00 
R5686t2842 n5687 n2843 R=4.941e+00 
R5686t2585 n5687 n2586 R=2.684e+01 
R5687t5597 n5688 n5598 R=2.573e+01 
R5688t421 n5689 n422 R=8.857e+00 
R5688t5066 n5689 n5067 R=5.903e+00 
R5688t1219 n5689 n1220 R=1.150e+01 
R5688t3660 n5689 n3661 R=5.836e+00 
R5689t2337 n5690 n2338 R=8.522e+00 
R5689t5001 n5690 n5002 R=9.137e+00 
R5689t4615 n5690 n4616 R=8.601e+00 
R5689t469 n5690 n470 R=6.149e+00 
R5690t260 n5691 n261 R=2.158e+00 
R5690t3642 n5691 n3643 R=5.317e+01 
R5690t890 n5691 n891 R=4.184e+00 
R5691t4511 n5692 n4512 R=1.375e+02 
R5691t4675 n5692 n4676 R=2.840e+00 
R5691t5312 n5692 n5313 R=2.995e+00 
R5691t3636 n5692 n3637 R=5.745e+00 
R5692t882 n5693 n883 R=5.708e+00 
R5692t5095 n5693 n5096 R=4.800e+00 
R5692t4696 n5693 n4697 R=2.144e+01 
R5692t5381 n5693 n5382 R=5.958e+00 
R5693t4345 n5694 n4346 R=4.247e+01 
R5693t3449 n5694 n3450 R=8.737e+00 
R5693t576 n5694 n577 R=1.870e+01 
R5693t747 n5694 n748 R=8.441e+00 
R5694t2353 n5695 n2354 R=1.178e+01 
R5694t4295 n5695 n4296 R=2.706e+00 
R5694t1788 n5695 n1789 R=1.528e+01 
R5694t2905 n5695 n2906 R=8.882e+00 
R5695t2360 n5696 n2361 R=6.679e+01 
R5695t1990 n5696 n1991 R=2.310e+00 
R5695t2839 n5696 n2840 R=9.252e+00 
R5695t1339 n5696 n1340 R=9.583e+01 
R5695t3534 n5696 n3535 R=5.557e+00 
R5696t5010 n5697 n5011 R=2.383e+01 
R5696t2430 n5697 n2431 R=2.895e+01 
R5696t2268 n5697 n2269 R=6.300e+00 
R5696t2048 n5697 n2049 R=3.246e+00 
R5697t2166 n5698 n2167 R=3.464e+00 
R5697t3186 n5698 n3187 R=2.621e+03 
R5697t2058 n5698 n2059 R=2.626e+00 
R5698t386 n5699 n387 R=3.748e+01 
R5698t4142 n5699 n4143 R=6.483e+00 
R5698t1953 n5699 n1954 R=4.958e+00 
R5699t1450 n5700 n1451 R=1.590e+01 
R5699t4967 n5700 n4968 R=1.459e+01 
R5700t3609 n5701 n3610 R=8.428e+00 
R5700t828 n5701 n829 R=7.346e+00 
R5701t2458 n5702 n2459 R=6.013e+00 
R5701t2771 n5702 n2772 R=2.178e+01 
R5701t1196 n5702 n1197 R=8.642e+00 
R5701t5482 n5702 n5483 R=9.536e+00 
R5701t5568 n5702 n5569 R=7.985e+00 
R5702t640 n5703 n641 R=9.494e+00 
R5702t3663 n5703 n3664 R=4.830e+00 
R5702t567 n5703 n568 R=2.591e+01 
R5702t1571 n5703 n1572 R=6.079e+00 
R5702t5340 n5703 n5341 R=3.666e+01 
R5703t871 n5704 n872 R=1.599e+01 
R5703t3771 n5704 n3772 R=6.716e+00 
R5703t4917 n5704 n4918 R=9.477e+00 
R5703t69 n5704 n70 R=3.701e+00 
R5704t1540 n5705 n1541 R=1.116e+01 
R5704t2518 n5705 n2519 R=3.507e+00 
R5705t782 n5706 n783 R=5.456e+00 
R5705t5450 n5706 n5451 R=2.454e+00 
R5705t4914 n5706 n4915 R=3.231e+01 
R5706t5665 n5707 n5666 R=2.655e+01 
R5706t4292 n5707 n4293 R=8.702e+00 
R5706t2854 n5707 n2855 R=3.792e+00 
R5706t5332 n5707 n5333 R=1.505e+01 
R5707t3789 n1 n3790 R=3.588e+00 
R5707t1920 n1 n1921 R=1.368e+01 
R5708t4074 n5709 n4075 R=2.041e+01 
R5708t4879 n5709 n4880 R=4.823e+01 
R5709t2023 n5710 n2024 R=4.931e+00 
R5709t3174 n5710 n3175 R=1.254e+01 
R5709t3626 n5710 n3627 R=7.506e+00 
R5710t1109 n5711 n1110 R=9.028e+01 
R5710t5182 n5711 n5183 R=2.132e+00 
R5710t303 n5711 n304 R=2.501e+00 
R5711t4934 n5712 n4935 R=3.986e+00 
R5712t2343 n5713 n2344 R=7.176e+00 
R5712t1795 n5713 n1796 R=2.514e+01 
R5712t1821 n5713 n1822 R=5.033e+00 
R5712t5034 n5713 n5035 R=9.218e+00 
R5712t5220 n5713 n5221 R=1.210e+01 
R5712t4273 n5713 n4274 R=2.316e+01 
R5713t2057 n5714 n2058 R=1.146e+01 
R5713t3866 n5714 n3867 R=1.015e+01 
R5713t66 n5714 n67 R=2.847e+01 
R5713t860 n5714 n861 R=2.252e+01 
R5713t2433 n5714 n2434 R=5.979e+00 
R5713t254 n5714 n255 R=8.013e+00 
R5714t3197 n5715 n3198 R=1.265e+01 
R5714t2205 n5715 n2206 R=1.692e+02 
R5714t2225 n5715 n2226 R=8.583e+00 
R5715t3778 n5716 n3779 R=6.223e+00 
R5715t746 n5716 n747 R=2.001e+01 
R5716t828 n5717 n829 R=7.753e+00 
R5716t3609 n5717 n3610 R=8.072e+00 
R5716t291 n5717 n292 R=1.366e+01 
R5716t3645 n5717 n3646 R=7.753e+00 
R5716t259 n5717 n260 R=6.001e+00 
R5717t1858 n5718 n1859 R=3.003e+00 
R5717t125 n5718 n126 R=7.424e+00 
R5717t4674 n5718 n4675 R=8.862e+00 
R5717t35 n5718 n36 R=6.175e+00 
R5718t3296 n5719 n3297 R=2.278e+01 
R5718t4141 n5719 n4142 R=1.827e+01 
R5718t4636 n5719 n4637 R=3.276e+00 
R5718t3213 n5719 n3214 R=1.324e+01 
R5718t5499 n5719 n5500 R=3.609e+01 
R5718t1869 n5719 n1870 R=2.176e+01 
R5719t386 n5720 n387 R=3.216e+00 
R5719t5698 n5720 n5699 R=2.439e+01 
R5719t1953 n5720 n1954 R=6.126e+00 
R5720t3849 n5721 n3850 R=2.184e+01 
R5720t1068 n5721 n1069 R=9.840e+00 
R5720t2999 n5721 n3000 R=1.776e+01 
R5721t4170 n5722 n4171 R=2.000e+00 
R5721t2125 n5722 n2126 R=3.508e+00 
R5721t3871 n5722 n3872 R=1.837e+01 
R5721t3030 n5722 n3031 R=1.634e+01 
R5722t1282 n5723 n1283 R=1.478e+03 
R5722t793 n5723 n794 R=1.337e+01 
R5722t2036 n5723 n2037 R=6.826e+01 
R5722t2701 n5723 n2702 R=1.081e+01 
R5722t1649 n5723 n1650 R=9.107e+00 
R5722t4374 n5723 n4375 R=4.195e+00 
R5722t1958 n5723 n1959 R=1.802e+01 
R5723t1987 n5724 n1988 R=4.015e+00 
R5723t4267 n5724 n4268 R=5.175e+00 
R5724t3863 n5725 n3864 R=7.212e+00 
R5724t3853 n5725 n3854 R=7.917e+00 
R5724t3698 n5725 n3699 R=3.988e+00 
R5724t2992 n5725 n2993 R=1.809e+01 
R5725t1972 n5726 n1973 R=1.257e+01 
R5725t3251 n5726 n3252 R=1.636e+01 
R5725t128 n5726 n129 R=3.566e+00 
R5725t5181 n5726 n5182 R=1.601e+01 
R5726t3466 n5727 n3467 R=9.226e+00 
R5726t4829 n5727 n4830 R=2.809e+00 
R5726t3855 n5727 n3856 R=1.628e+01 
R5727t62 n5728 n63 R=2.198e+00 
R5727t2681 n5728 n2682 R=9.649e+00 
R5727t1711 n5728 n1712 R=9.027e+00 
R5728t1360 n5729 n1361 R=8.009e+02 
R5728t5059 n5729 n5060 R=5.543e+00 
R5728t1480 n5729 n1481 R=1.077e+01 
R5728t2811 n5729 n2812 R=4.436e+00 
R5729t4844 n5730 n4845 R=5.743e+00 
R5729t4790 n5730 n4791 R=4.718e+00 
R5729t2988 n5730 n2989 R=2.478e+00 
R5730t2113 n5731 n2114 R=1.996e+01 
R5730t3057 n5731 n3058 R=1.511e+01 
R5730t3736 n5731 n3737 R=1.212e+01 
R5730t3160 n5731 n3161 R=4.028e+00 
R5730t672 n5731 n673 R=8.294e+00 
R5730t2680 n5731 n2681 R=7.409e+00 
R5731t1894 n5732 n1895 R=3.943e+00 
R5731t4541 n5732 n4542 R=5.204e+01 
R5731t1431 n5732 n1432 R=8.244e+00 
R5731t357 n5732 n358 R=3.215e+00 
R5732t5099 n5733 n5100 R=6.928e+00 
R5732t3630 n5733 n3631 R=4.890e+00 
R5733t3015 n5734 n3016 R=7.065e+00 
R5733t3554 n5734 n3555 R=5.449e+00 
R5733t5108 n5734 n5109 R=8.274e+00 
R5733t842 n5734 n843 R=5.881e+00 
R5734t782 n5735 n783 R=1.077e+01 
R5734t5705 n5735 n5706 R=3.178e+00 
R5734t512 n5735 n513 R=9.185e+00 
R5734t3976 n5735 n3977 R=1.128e+01 
R5734t5620 n5735 n5621 R=1.860e+01 
R5734t4914 n5735 n4915 R=1.480e+01 
R5735t5709 n5736 n5710 R=8.483e+00 
R5735t1003 n5736 n1004 R=4.137e+00 
R5735t443 n5736 n444 R=2.528e+00 
R5735t3626 n5736 n3627 R=8.634e+00 
R5736t4952 n5737 n4953 R=2.014e+01 
R5737t2260 n5738 n2261 R=2.867e+01 
R5737t2813 n5738 n2814 R=4.254e+00 
R5737t476 n5738 n477 R=7.424e+00 
R5737t4956 n5738 n4957 R=3.305e+00 
R5737t3650 n5738 n3651 R=5.010e+00 
R5738t1630 n5739 n1631 R=6.722e+00 
R5738t3990 n5739 n3991 R=4.544e+00 
R5739t191 n5740 n192 R=3.029e+00 
R5739t2192 n5740 n2193 R=7.708e+00 
R5739t1753 n5740 n1754 R=4.165e+00 
R5740t1930 n5741 n1931 R=3.650e+00 
R5740t302 n5741 n303 R=3.337e+01 
R5741t1342 n5742 n1343 R=1.668e+01 
R5742t832 n5743 n833 R=1.677e+01 
R5742t2509 n5743 n2510 R=3.420e+01 
R5742t2540 n5743 n2541 R=5.881e+00 
R5743t536 n5744 n537 R=3.154e+00 
R5744t3982 n5745 n3983 R=2.592e+00 
R5745t4040 n5746 n4041 R=1.588e+03 
R5745t5284 n5746 n5285 R=1.367e+01 
R5745t772 n5746 n773 R=3.972e+00 
R5745t194 n5746 n195 R=6.591e+02 
R5746t1829 n5747 n1830 R=6.000e+00 
R5746t5521 n5747 n5522 R=6.297e+00 
R5746t1583 n5747 n1584 R=8.041e+00 
R5746t2751 n5747 n2752 R=7.983e+00 
R5746t2679 n5747 n2680 R=6.303e+01 
R5746t2128 n5747 n2129 R=7.484e+00 
R5746t2119 n5747 n2120 R=8.689e+01 
R5747t5428 n5748 n5429 R=3.312e+01 
R5747t3518 n5748 n3519 R=7.420e+00 
R5747t1230 n5748 n1231 R=1.104e+02 
R5748t5227 n5749 n5228 R=2.871e+01 
R5748t1444 n5749 n1445 R=1.191e+01 
R5748t2454 n5749 n2455 R=9.790e+00 
R5748t508 n5749 n509 R=4.014e+00 
R5749t2165 n5750 n2166 R=1.265e+01 
R5749t5630 n5750 n5631 R=3.390e+00 
R5749t452 n5750 n453 R=7.825e+01 
R5749t3046 n5750 n3047 R=4.677e+00 
R5750t56 n5751 n57 R=1.119e+01 
R5750t3226 n5751 n3227 R=9.609e+00 
R5750t1964 n5751 n1965 R=8.785e+00 
R5750t474 n5751 n475 R=2.022e+01 
R5750t2103 n5751 n2104 R=6.884e+00 
R5750t1482 n5751 n1483 R=5.736e+00 
R5751t1741 n5752 n1742 R=2.147e+00 
R5751t1072 n5752 n1073 R=6.922e+00 
R5751t5480 n5752 n5481 R=2.205e+01 
R5752t868 n5753 n869 R=4.940e+00 
R5752t909 n5753 n910 R=1.287e+01 
R5752t4680 n5753 n4681 R=1.549e+01 
R5752t1638 n5753 n1639 R=4.960e+00 
R5752t1766 n5753 n1767 R=9.210e+00 
R5753t1022 n5754 n1023 R=4.855e+00 
R5753t3370 n5754 n3371 R=4.856e+00 
R5753t422 n5754 n423 R=6.618e+00 
R5754t2180 n5755 n2181 R=1.770e+00 
R5755t4842 n5756 n4843 R=4.335e+00 
R5755t2435 n5756 n2436 R=4.146e+00 
R5756t5169 n5757 n5170 R=1.316e+01 
R5756t1150 n5757 n1151 R=3.674e+00 
R5756t3835 n5757 n3836 R=7.793e+01 
R5756t2934 n5757 n2935 R=2.853e+01 
R5756t134 n5757 n135 R=2.786e+02 
R5757t2115 n5758 n2116 R=2.336e+01 
R5757t3170 n5758 n3171 R=2.895e+00 
R5758t1703 n5759 n1704 R=4.786e+00 
R5758t3064 n5759 n3065 R=3.764e+00 
R5758t851 n5759 n852 R=8.862e+00 
R5758t5434 n5759 n5435 R=3.429e+00 
R5758t3500 n5759 n3501 R=2.710e+01 
R5758t2867 n5759 n2868 R=9.529e+01 
R5759t3682 n5760 n3683 R=1.050e+01 
R5759t4953 n5760 n4954 R=5.763e+00 
R5759t5647 n5760 n5648 R=1.027e+01 
R5759t52 n5760 n53 R=3.984e+00 
R5759t758 n5760 n759 R=1.234e+01 
R5759t4554 n5760 n4555 R=4.806e+01 
R5759t4221 n5760 n4222 R=5.095e+00 
R5760t1926 n5761 n1927 R=3.189e+00 
R5760t5580 n5761 n5581 R=3.765e+00 
R5760t328 n5761 n329 R=2.822e+00 
R5761t1709 n5762 n1710 R=2.716e+00 
R5761t3108 n5762 n3109 R=1.795e+01 
R5761t412 n5762 n413 R=5.260e+02 
R5761t641 n5762 n642 R=1.095e+01 
R5761t85 n5762 n86 R=1.087e+01 
R5762t2208 n5763 n2209 R=7.677e+00 
R5762t5392 n5763 n5393 R=5.822e+00 
R5762t901 n5763 n902 R=4.816e+00 
R5763t2056 n5764 n2057 R=1.454e+01 
R5763t1749 n5764 n1750 R=3.051e+02 
R5764t293 n5765 n294 R=3.288e+00 
R5764t2739 n5765 n2740 R=3.737e+01 
R5765t466 n5766 n467 R=2.175e+01 
R5765t521 n5766 n522 R=2.893e+00 
R5765t4594 n5766 n4595 R=8.226e+00 
R5765t1393 n5766 n1394 R=1.781e+01 
R5766t3529 n5767 n3530 R=1.419e+01 
R5766t2913 n5767 n2914 R=3.943e+01 
R5767t1692 n5768 n1693 R=4.273e+00 
R5767t3396 n5768 n3397 R=4.259e+01 
R5767t3892 n5768 n3893 R=7.763e+00 
R5767t1524 n5768 n1525 R=5.076e+00 
R5768t1852 n5769 n1853 R=2.643e+01 
R5768t5711 n5769 n5712 R=1.320e+01 
R5768t4934 n5769 n4935 R=4.664e+00 
R5768t4752 n5769 n4753 R=5.988e+01 
R5768t5044 n5769 n5045 R=1.931e+01 
R5769t190 n5770 n191 R=8.520e+00 
R5769t3379 n5770 n3380 R=1.105e+01 
R5770t734 n5771 n735 R=2.175e+00 
R5770t4687 n5771 n4688 R=4.505e+00 
R5770t1690 n5771 n1691 R=1.259e+01 
R5770t1790 n5771 n1791 R=2.065e+01 
R5771t4562 n5772 n4563 R=4.716e+00 
R5771t1299 n5772 n1300 R=6.649e+00 
R5771t2219 n5772 n2220 R=2.449e+00 
R5772t1266 n5773 n1267 R=3.699e+00 
R5772t3529 n5773 n3530 R=5.281e+00 
R5772t5766 n5773 n5767 R=3.361e+00 
R5773t1958 n5774 n1959 R=1.651e+01 
R5773t4374 n5774 n4375 R=4.239e+00 
R5774t5135 n5775 n5136 R=4.740e+00 
R5774t4535 n5775 n4536 R=1.156e+01 
R5774t558 n5775 n559 R=9.516e+00 
R5775t4062 n5776 n4063 R=7.319e+00 
R5776t3754 n5777 n3755 R=7.543e+00 
R5776t3194 n5777 n3195 R=3.829e+00 
R5777t825 n5778 n826 R=4.529e+01 
R5777t853 n5778 n854 R=6.099e+00 
R5777t1656 n5778 n1657 R=2.111e+01 
R5778t1789 n5779 n1790 R=5.445e+01 
R5778t3215 n5779 n3216 R=6.498e+00 
R5778t3529 n5779 n3530 R=2.132e+01 
R5778t5766 n5779 n5767 R=7.680e+00 
R5778t2913 n5779 n2914 R=4.596e+00 
R5778t5624 n5779 n5625 R=5.118e+00 
R5779t4055 n5780 n4056 R=2.814e+01 
R5779t816 n5780 n817 R=3.873e+00 
R5780t4160 n5781 n4161 R=3.454e+00 
R5780t3290 n5781 n3291 R=2.324e+01 
R5781t925 n5782 n926 R=1.323e+01 
R5782t5267 n5783 n5268 R=2.803e+00 
R5782t4944 n5783 n4945 R=9.663e+00 
R5782t4417 n5783 n4418 R=8.941e+00 
R5783t832 n5784 n833 R=3.194e+00 
R5783t4979 n5784 n4980 R=7.374e+00 
R5783t5742 n5784 n5743 R=1.042e+01 
R5784t5510 n5785 n5511 R=1.599e+00 
R5784t3624 n5785 n3625 R=1.130e+01 
R5785t1473 n5786 n1474 R=2.387e+01 
R5785t2577 n5786 n2578 R=3.076e+00 
R5785t3391 n5786 n3392 R=7.754e+00 
R5785t3113 n5786 n3114 R=4.418e+00 
R5785t1751 n5786 n1752 R=5.557e+01 
R5786t3977 n5787 n3978 R=2.941e+00 
R5786t2412 n5787 n2413 R=6.968e+01 
R5786t3418 n5787 n3419 R=1.559e+01 
R5786t2461 n5787 n2462 R=1.176e+01 
R5786t538 n5787 n539 R=5.286e+00 
R5787t3308 n5788 n1 R=3.596e+01 
R5787t1787 n5788 n1788 R=3.527e+00 
R5787t4522 n5788 n4523 R=1.741e+02 
R5787t5396 n5788 n5397 R=1.109e+01 
R5787t4385 n5788 n1 R=6.311e+02 
R5788t1098 n5789 n1099 R=2.029e+01 
R5788t5553 n5789 n5554 R=5.570e+00 
R5788t4737 n5789 n4738 R=1.418e+01 
R5788t3936 n5789 n3937 R=3.671e+00 
R5788t4571 n5789 n4572 R=7.941e+00 
R5789t2196 n5790 n2197 R=6.145e+00 
R5789t3790 n5790 n3791 R=8.792e+00 
R5789t1489 n5790 n1490 R=2.722e+01 
R5789t1430 n5790 n1431 R=7.562e+00 
R5790t381 n5791 n382 R=3.551e+00 
R5790t5136 n5791 n5137 R=1.057e+01 
R5790t2266 n5791 n2267 R=2.000e+01 
R5791t4104 n5792 n4105 R=6.001e+01 
R5791t5558 n5792 n5559 R=5.043e+00 
R5791t2740 n5792 n2741 R=1.664e+01 
R5791t5030 n5792 n5031 R=1.715e+01 
R5792t3504 n5793 n3505 R=1.116e+02 
R5792t4481 n5793 n4482 R=1.926e+00 
R5792t2714 n5793 n2715 R=1.465e+01 
R5792t4464 n5793 n4465 R=1.681e+02 
R5792t1274 n5793 n1275 R=1.867e+00 
R5792t5180 n5793 n5181 R=9.330e+01 
R5793t101 n5794 n102 R=1.095e+01 
R5793t1550 n5794 n1551 R=4.653e+00 
R5793t5593 n5794 n5594 R=3.394e+00 
R5793t4961 n5794 n4962 R=1.464e+01 
R5793t4440 n5794 n4441 R=4.086e+01 
R5793t3187 n5794 n3188 R=5.393e+01 
R5794t5494 n5795 n5495 R=4.498e+00 
R5794t3571 n5795 n3572 R=5.342e+00 
R5795t876 n5796 n877 R=3.599e+00 
R5795t3602 n5796 n3603 R=2.555e+01 
R5795t4173 n5796 n4174 R=7.780e+00 
R5795t2464 n5796 n2465 R=6.935e+00 
R5796t978 n5797 n979 R=3.358e+00 
R5796t1487 n5797 n1488 R=9.245e+00 
R5796t2124 n5797 n2125 R=3.129e+00 
R5797t3488 n5798 n3489 R=2.538e+01 
R5797t616 n5798 n617 R=7.371e+00 
R5797t974 n5798 n975 R=3.966e+01 
R5797t576 n5798 n577 R=9.176e+00 
R5798t2766 n5799 n2767 R=4.115e+01 
R5798t3251 n5799 n3252 R=6.947e+00 
R5798t3254 n5799 n3255 R=2.900e+00 
R5798t2539 n5799 n2540 R=3.261e+01 
R5798t4900 n5799 n4901 R=3.030e+00 
R5799t5630 n5800 n5631 R=3.869e+00 
R5799t5749 n5800 n5750 R=7.281e+01 
R5799t1205 n5800 n1206 R=9.211e+00 
R5799t940 n5800 n941 R=7.446e+00 
R5799t452 n5800 n453 R=4.211e+00 
R5800t323 n5801 n324 R=4.812e+00 
R5800t2734 n5801 n2735 R=4.186e+00 
R5801t5415 n5802 n5416 R=1.000e+01 
R5801t501 n5802 n502 R=3.878e+00 
R5801t3490 n5802 n3491 R=9.602e+00 
R5801t3050 n5802 n3051 R=6.162e+01 
R5801t3502 n5802 n3503 R=1.102e+01 
R5801t4381 n5802 n4382 R=1.003e+01 
R5802t695 n5803 n696 R=7.429e+00 
R5802t1576 n5803 n1577 R=9.031e+01 
R5802t2609 n5803 n2610 R=4.684e+00 
R5802t3129 n5803 n3130 R=2.101e+01 
R5803t2328 n5804 n2329 R=8.391e+00 
R5803t4240 n5804 n4241 R=2.582e+00 
R5803t1899 n5804 n1900 R=5.687e+01 
R5804t3116 n5805 n3117 R=4.002e+01 
R5804t272 n5805 n273 R=5.523e+01 
R5804t5586 n5805 n5587 R=2.296e+01 
R5804t648 n5805 n649 R=4.172e+01 
R5804t1906 n5805 n1907 R=3.711e+00 
R5805t1679 n5806 n1680 R=4.885e+02 
R5805t1619 n5806 n1620 R=9.643e+00 
R5805t2367 n5806 n2368 R=5.250e+02 
R5806t1951 n5807 n1952 R=8.599e+00 
R5806t5096 n5807 n5097 R=2.017e+01 
R5806t3229 n5807 n3230 R=2.835e+01 
R5806t2084 n5807 n2085 R=1.057e+01 
R5806t3031 n5807 n3032 R=5.115e+00 
R5807t4022 n5808 n4023 R=8.864e+00 
R5807t4715 n5808 n4716 R=1.397e+01 
R5807t4857 n5808 n4858 R=6.440e+00 
R5807t4020 n5808 n4021 R=1.385e+01 
R5807t5358 n5808 n5359 R=2.291e+01 
R5807t1675 n5808 n1676 R=2.803e+00 
R5808t1185 n5809 n1186 R=2.133e+01 
R5808t3683 n5809 n3684 R=5.815e+00 
R5808t4809 n5809 n4810 R=3.294e+01 
R5808t4978 n5809 n4979 R=1.558e+01 
R5809t5332 n5810 n5333 R=4.541e+01 
R5809t2369 n5810 n2370 R=1.276e+01 
R5810t1959 n5811 n1960 R=1.235e+01 
R5810t4557 n5811 n4558 R=6.481e+00 
R5810t3973 n5811 n3974 R=7.044e+00 
R5810t3425 n5811 n3426 R=2.152e+00 
R5811t4548 n5812 n4549 R=5.491e+00 
R5811t2804 n5812 n2805 R=2.075e+01 
R5811t2452 n5812 n2453 R=8.211e+00 
R5811t67 n5812 n68 R=1.464e+01 
R5811t3337 n5812 n3338 R=1.139e+01 
R5811t4984 n5812 n4985 R=9.430e+00 
R5812t1803 n5813 n1804 R=1.466e+01 
R5813t2300 n5814 n2301 R=5.172e+00 
R5813t4660 n5814 n4661 R=5.454e+02 
R5813t2623 n5814 n2624 R=5.834e+00 
R5813t3434 n5814 n3435 R=5.805e+00 
R5814t2041 n5815 n2042 R=4.912e+00 
R5814t73 n5815 n74 R=3.840e+00 
R5815t4643 n5816 n4644 R=4.471e+00 
R5815t1062 n5816 n1063 R=4.432e+01 
R5815t986 n5816 n987 R=2.856e+01 
R5815t4854 n5816 n4855 R=2.626e+00 
R5815t4002 n5816 n4003 R=1.775e+01 
R5816t381 n5817 n382 R=2.088e+01 
R5816t157 n5817 n158 R=7.521e+00 
R5816t5136 n5817 n5137 R=4.212e+00 
R5816t5790 n5817 n5791 R=4.756e+00 
R5817t1922 n5818 n1923 R=9.567e+00 
R5817t601 n5818 n602 R=1.149e+01 
R5817t2564 n5818 n2565 R=3.224e+00 
R5818t44 n5819 n45 R=2.461e+00 
R5818t1450 n5819 n1451 R=8.201e+01 
R5818t2809 n5819 n2810 R=1.616e+01 
R5819t3720 n5820 n3721 R=9.394e+01 
R5819t5326 n5820 n5327 R=2.693e+00 
R5819t4683 n5820 n4684 R=4.477e+00 
R5820t62 n5821 n63 R=6.247e+00 
R5820t2529 n5821 n2530 R=1.047e+01 
R5820t5727 n5821 n5728 R=5.248e+02 
R5820t1711 n5821 n1712 R=2.842e+01 
R5820t3922 n5821 n3923 R=1.410e+01 
R5821t3193 n5822 n3194 R=6.370e+00 
R5821t2099 n5822 n2100 R=1.312e+02 
R5822t4067 n5823 n4068 R=7.089e+00 
R5822t4118 n5823 n4119 R=2.787e+00 
R5822t1078 n5823 n1079 R=1.703e+01 
R5822t4046 n5823 n4047 R=5.301e+01 
R5822t930 n5823 n931 R=1.389e+01 
R5822t4803 n5823 n4804 R=2.883e+01 
R5823t3332 n5824 n3333 R=7.404e+00 
R5823t5676 n5824 n5677 R=4.745e+00 
R5823t571 n5824 n572 R=8.023e+01 
R5823t208 n5824 n209 R=5.837e+00 
R5823t124 n5824 n125 R=5.395e+00 
R5824t3437 n5825 n3438 R=4.088e+00 
R5824t888 n5825 n889 R=1.467e+01 
R5824t4425 n5825 n4426 R=8.457e+00 
R5825t2414 n5826 n2415 R=5.362e+00 
R5825t5270 n5826 n5271 R=4.517e+00 
R5825t1291 n5826 n1292 R=6.320e+00 
R5826t3588 n5827 n3589 R=9.688e+00 
R5826t2965 n5827 n2966 R=3.069e+00 
R5826t2380 n5827 n2381 R=8.857e+00 
R5826t240 n5827 n241 R=1.806e+02 
R5826t380 n5827 n381 R=4.380e+00 
R5827t1371 n5828 n1372 R=1.211e+02 
R5827t4658 n5828 n4659 R=3.983e+00 
R5827t215 n5828 n216 R=2.643e+00 
R5828t3781 n5829 n3782 R=1.110e+01 
R5828t4239 n5829 n4240 R=2.937e+00 
R5829t4605 n5830 n4606 R=3.966e+01 
R5829t3449 n5830 n3450 R=1.170e+01 
R5830t1017 n5831 n1018 R=3.028e+00 
R5830t3083 n5831 n3084 R=1.913e+01 
R5831t2092 n5832 n2093 R=2.568e+00 
R5831t2688 n5832 n2689 R=1.351e+01 
R5831t3398 n5832 n3399 R=2.892e+00 
R5831t5002 n5832 n5003 R=1.159e+01 
R5831t1858 n5832 n1859 R=7.566e+02 
R5832t2899 n5833 n2900 R=5.644e+00 
R5832t5277 n5833 n5278 R=4.313e+00 
R5833t38 n5834 n39 R=3.629e+00 
R5833t2733 n5834 n2734 R=9.043e+00 
R5833t3929 n5834 n3930 R=5.374e+01 
R5833t4687 n5834 n4688 R=4.717e+02 
R5833t734 n5834 n735 R=2.642e+00 
R5834t4745 n5835 n4746 R=2.635e+00 
R5834t2059 n5835 n2060 R=7.487e+00 
R5834t5567 n5835 n5568 R=7.783e+00 
R5835t3710 n5836 n3711 R=9.466e+00 
R5835t4241 n5836 n4242 R=1.893e+00 
R5836t4513 n5837 n4514 R=9.715e+01 
R5836t4211 n5837 n4212 R=8.638e+00 
R5836t1522 n5837 n1523 R=2.696e+00 
R5836t1859 n5837 n1860 R=1.874e+01 
R5836t5457 n5837 n5458 R=3.085e+03 
R5836t24 n5837 n25 R=4.175e+01 
R5837t2748 n5838 n2749 R=3.369e+00 
R5837t2637 n5838 n2638 R=4.300e+00 
R5837t5495 n5838 n5496 R=1.153e+01 
R5838t1786 n5839 n1787 R=5.114e+00 
R5838t5138 n5839 n5139 R=7.171e+00 
R5838t1102 n5839 n1103 R=2.907e+01 
R5838t895 n5839 n896 R=6.809e+01 
R5838t5070 n5839 n5071 R=5.606e+00 
R5839t1976 n5840 n1977 R=4.411e+00 
R5839t661 n5840 n662 R=8.185e+01 
R5840t3359 n5841 n3360 R=6.432e+00 
R5840t3512 n5841 n3513 R=2.779e+00 
R5841t1142 n5842 n1143 R=3.452e+00 
R5841t1773 n5842 n1774 R=1.226e+01 
R5841t3000 n5842 n3001 R=1.586e+01 
R5841t831 n5842 n832 R=2.075e+01 
R5841t1367 n5842 n1368 R=3.624e+01 
R5841t1237 n5842 n1238 R=5.246e+01 
R5842t1659 n5843 n1660 R=9.870e+00 
R5842t4604 n5843 n4605 R=1.343e+01 
R5842t579 n5843 n580 R=8.091e+00 
R5842t4624 n5843 n4625 R=1.050e+01 
R5843t1805 n5844 n1806 R=1.734e+01 
R5844t4607 n5845 n4608 R=1.587e+00 
R5844t524 n5845 n525 R=1.456e+01 
R5845t2475 n5846 n2476 R=1.982e+01 
R5845t1635 n5846 n1636 R=7.896e+00 
R5845t439 n5846 n440 R=6.210e+01 
R5845t2009 n5846 n2010 R=3.101e+00 
R5845t1562 n5846 n1563 R=1.920e+02 
R5845t4775 n5846 n4776 R=4.696e+00 
R5846t4867 n5847 n4868 R=6.378e+00 
R5846t914 n5847 n915 R=3.649e+00 
R5847t5665 n5848 n5666 R=1.286e+01 
R5847t618 n5848 n619 R=1.064e+01 
R5847t1412 n5848 n1413 R=1.865e+01 
R5847t3214 n5848 n3215 R=3.208e+01 
R5847t1221 n5848 n1222 R=5.450e+00 
R5848t1171 n5849 n1172 R=5.154e+01 
R5848t3331 n5849 n3332 R=1.287e+01 
R5848t4936 n5849 n4937 R=5.689e+01 
R5848t649 n5849 n650 R=7.441e+00 
R5849t1159 n5850 n1160 R=2.090e+02 
R5849t1488 n5850 n1489 R=7.118e+00 
R5849t196 n5850 n197 R=9.497e+00 
R5849t3576 n5850 n3577 R=8.419e+00 
R5849t2775 n5850 n2776 R=1.105e+01 
R5850t2992 n5851 n2993 R=3.973e+01 
R5850t3698 n5851 n3699 R=1.165e+01 
R5850t4823 n5851 n4824 R=3.182e+00 
R5850t5164 n5851 n5165 R=6.154e+00 
R5851t628 n5852 n629 R=2.221e+00 
R5851t195 n5852 n196 R=1.536e+01 
R5851t2461 n5852 n2462 R=6.896e+00 
R5852t5312 n5853 n5313 R=7.296e+00 
R5853t310 n5854 n311 R=8.775e+00 
R5853t4676 n5854 n4677 R=5.113e+00 
R5853t2562 n5854 n2563 R=4.651e+00 
R5853t3936 n5854 n3937 R=1.287e+01 
R5853t4737 n5854 n4738 R=6.130e+01 
R5853t1734 n5854 n1735 R=1.463e+01 
R5854t1079 n5855 n1080 R=6.561e+00 
R5854t4257 n5855 n4258 R=3.103e+00 
R5854t3031 n5855 n3032 R=2.240e+01 
R5854t4229 n5855 n4230 R=2.157e+00 
R5855t1765 n5856 n1766 R=3.131e+01 
R5855t3480 n5856 n3481 R=1.907e+01 
R5855t4839 n5856 n4840 R=5.228e+00 
R5855t1349 n5856 n1350 R=5.069e+00 
R5855t3875 n5856 n3876 R=1.969e+01 
R5855t2874 n5856 n2875 R=4.808e+00 
R5856t4467 n5857 n4468 R=8.807e+00 
R5856t112 n5857 n113 R=3.773e+00 
R5856t3317 n5857 n3318 R=1.305e+01 
R5857t608 n5858 n609 R=3.585e+01 
R5857t142 n5858 n143 R=1.908e+01 
R5857t3092 n5858 n3093 R=3.507e+00 
R5858t4053 n5859 n4054 R=7.450e+00 
R5858t5592 n5859 n5593 R=4.863e+00 
R5858t5498 n5859 n5499 R=3.482e+01 
R5858t4907 n5859 n4908 R=1.924e+01 
R5858t4693 n5859 n4694 R=6.781e+01 
R5858t958 n5859 n959 R=1.914e+01 
R5859t4512 n5860 n4513 R=4.087e+00 
R5860t2940 n5861 n2941 R=8.739e+00 
R5860t5439 n5861 n5440 R=2.618e+01 
R5860t4386 n5861 n4387 R=3.533e+01 
R5861t675 n5862 n676 R=2.634e+01 
R5861t1340 n5862 n1341 R=1.331e+01 
R5861t3324 n5862 n3325 R=1.706e+01 
R5861t112 n5862 n113 R=5.593e+00 
R5861t3317 n5862 n3318 R=3.770e+00 
R5862t2290 n5863 n2291 R=3.292e+00 
R5862t5623 n5863 n5624 R=1.889e+01 
R5862t906 n5863 n907 R=1.504e+01 
R5862t5657 n5863 n5658 R=7.527e+00 
R5862t3114 n5863 n3115 R=8.562e+00 
R5862t4422 n5863 n4423 R=8.527e+00 
R5863t5295 n5864 n5296 R=7.825e+02 
R5863t1183 n5864 n1184 R=5.410e+00 
R5863t3064 n5864 n3065 R=6.217e+00 
R5863t3410 n5864 n3411 R=6.561e+00 
R5864t4026 n5865 n4027 R=9.526e+00 
R5864t1312 n5865 n1313 R=2.636e+01 
R5864t220 n5865 n221 R=1.023e+01 
R5864t2761 n5865 n2762 R=1.290e+02 
R5864t1882 n5865 n1883 R=1.046e+01 
R5864t5775 n5865 n5776 R=4.185e+00 
R5865t103 n5866 n104 R=9.994e+00 
R5865t3714 n5866 n3715 R=5.403e+02 
R5865t5546 n5866 n5547 R=3.235e+00 
R5866t639 n5867 n640 R=1.885e+01 
R5866t354 n5867 n355 R=1.150e+01 
R5866t4168 n5867 n4169 R=3.476e+00 
R5867t1098 n5868 n1099 R=2.330e+00 
R5867t5788 n5868 n5789 R=6.822e+00 
R5867t5553 n5868 n5554 R=5.248e+00 
R5869t4852 n5870 n4853 R=4.808e+00 
R5869t5673 n5870 n5674 R=2.197e+00 
R5869t5720 n5870 n5721 R=2.531e+01 
R5869t3849 n5870 n3850 R=3.020e+00 
R5870t143 n5871 n144 R=2.427e+01 
R5871t3282 n5872 n3283 R=1.661e+03 
R5871t3055 n5872 n3056 R=3.403e+00 
R5871t2968 n5872 n2969 R=3.596e+00 
R5872t423 n5873 n424 R=5.904e+01 
R5872t4811 n5873 n4812 R=2.706e+00 
R5872t4194 n5873 n4195 R=1.126e+01 
R5873t1540 n5874 n1541 R=3.633e+00 
R5873t5704 n5874 n5705 R=1.442e+01 
R5873t3459 n5874 n3460 R=1.016e+01 
R5873t2518 n5874 n2519 R=6.362e+00 
R5874t459 n5875 n460 R=6.123e+00 
R5874t3952 n5875 n3953 R=2.457e+00 
R5874t2231 n5875 n2232 R=1.335e+01 
R5874t1975 n5875 n1976 R=3.812e+00 
R5875t2835 n5876 n2836 R=2.168e+00 
R5875t5700 n5876 n5701 R=2.763e+01 
R5876t2015 n5877 n2016 R=6.510e+00 
R5876t3649 n5877 n3650 R=2.989e+00 
R5876t4952 n5877 n4953 R=2.440e+01 
R5877t5639 n5878 n5640 R=1.804e+01 
R5877t3727 n5878 n3728 R=3.597e+00 
R5878t2470 n5879 n2471 R=5.738e+00 
R5878t1124 n5879 n1125 R=2.948e+00 
R5878t3779 n5879 n3780 R=3.435e+01 
R5879t1109 n5880 n1110 R=3.458e+00 
R5879t5182 n5880 n5183 R=1.625e+01 
R5879t4277 n5880 n4278 R=3.256e+01 
R5880t2601 n5881 n2602 R=4.463e+01 
R5880t3295 n5881 n3296 R=4.392e+01 
R5881t1624 n5882 n1625 R=5.594e+00 
R5881t5244 n5882 n5245 R=2.101e+00 
R5881t3583 n5882 n3584 R=1.074e+01 
R5882t219 n5883 n220 R=8.782e+00 
R5882t3560 n5883 n3561 R=8.920e+00 
R5882t2657 n5883 n2658 R=5.568e+00 
R5882t2682 n5883 n2683 R=1.711e+01 
R5882t4153 n5883 n4154 R=5.723e+01 
R5882t3246 n5883 n3247 R=3.784e+00 
R5882t3526 n5883 n3527 R=1.052e+01 
R5883t1252 n5884 n1253 R=7.002e+01 
R5883t2139 n5884 n2140 R=9.079e+00 
R5884t1924 n5885 n1925 R=1.538e+01 
R5884t3898 n5885 n3899 R=4.230e+00 
R5884t2763 n5885 n2764 R=4.552e+00 
R5884t1222 n5885 n1223 R=5.180e+00 
R5885t1315 n5886 n1316 R=2.614e+00 
R5885t2487 n5886 n2488 R=1.041e+01 
R5885t3881 n5886 n3882 R=2.377e+01 
R5886t324 n5887 n325 R=8.342e+00 
R5886t3058 n5887 n3059 R=2.796e+01 
R5886t2898 n5887 n2899 R=2.537e+00 
R5886t3190 n5887 n3191 R=3.758e+00 
R5887t5757 n5888 n5758 R=8.578e+00 
R5887t3239 n5888 n3240 R=9.783e+00 
R5888t5116 n5889 n5117 R=5.109e+00 
R5888t5257 n5889 n5258 R=1.690e+01 
R5889t1618 n5890 n1619 R=4.343e+01 
R5889t1669 n5890 n1670 R=8.761e+01 
R5889t5222 n5890 n5223 R=4.505e+00 
R5889t3592 n5890 n3593 R=7.402e+00 
R5890t2049 n5891 n2050 R=2.281e+00 
R5890t3197 n5891 n3198 R=6.442e+00 
R5890t3413 n5891 n3414 R=2.088e+00 
R5891t2120 n5892 n2121 R=5.498e+00 
R5892t1480 n5893 n1481 R=2.868e+00 
R5892t631 n5893 n632 R=1.028e+01 
R5892t2811 n5893 n2812 R=1.808e+01 
R5892t5728 n5893 n5729 R=6.168e+00 
R5893t3746 n5894 n3747 R=5.864e+00 
R5893t2669 n5894 n2670 R=5.596e+00 
R5894t407 n5895 n408 R=8.745e+00 
R5894t2924 n5895 n2925 R=3.378e+00 
R5894t1795 n5895 n1796 R=1.720e+01 
R5894t1173 n5895 n1174 R=1.170e+01 
R5894t4137 n5895 n4138 R=1.380e+01 
R5894t923 n5895 n924 R=1.401e+01 
R5895t1593 n5896 n1594 R=4.514e+00 
R5895t3027 n5896 n3028 R=3.017e+00 
R5895t4691 n5896 n4692 R=1.306e+01 
R5895t1667 n5896 n1668 R=8.139e+00 
R5896t5761 n5897 n5762 R=2.694e+01 
R5896t641 n5897 n642 R=1.045e+01 
R5896t754 n5897 n755 R=3.901e+00 
R5896t1035 n5897 n1036 R=3.873e+00 
R5897t1301 n5898 n1302 R=2.239e+01 
R5897t88 n5898 n89 R=1.018e+01 
R5897t817 n5898 n818 R=1.034e+02 
R5897t2101 n5898 n2102 R=4.255e+01 
R5898t4759 n5899 n4760 R=3.289e+00 
R5898t5352 n5899 n5353 R=2.116e+00 
R5898t3927 n5899 n3928 R=3.505e+01 
R5898t5070 n5899 n5071 R=1.040e+01 
R5899t1899 n5900 n1900 R=1.246e+01 
R5899t5183 n5900 n5184 R=2.888e+00 
R5899t2201 n5900 n2202 R=1.052e+01 
R5899t5626 n5900 n5627 R=1.781e+02 
R5899t5256 n5900 n5257 R=8.692e+01 
R5899t4947 n5900 n4948 R=6.782e+00 
R5900t5261 n5901 n5262 R=1.654e+01 
R5900t3287 n5901 n3288 R=2.370e+01 
R5900t3245 n5901 n3246 R=3.672e+00 
R5901t5176 n5902 n5177 R=5.295e+00 
R5901t1162 n5902 n1163 R=6.546e+00 
R5902t2221 n5903 n2222 R=1.159e+02 
R5902t2795 n5903 n2796 R=2.235e+02 
R5902t2499 n5903 n2500 R=3.137e+00 
R5902t1049 n5903 n1050 R=3.443e+00 
R5903t2590 n5904 n2591 R=4.556e+01 
R5903t3382 n5904 n3383 R=9.504e+00 
R5903t5329 n5904 n5330 R=1.826e+01 
R5903t1387 n5904 n1388 R=5.063e+00 
R5903t5050 n5904 n5051 R=5.822e+00 
R5905t5367 n5906 n5368 R=8.361e+00 
R5905t877 n5906 n878 R=1.348e+01 
R5905t4814 n5906 n4815 R=5.653e+00 
R5906t368 n5907 n369 R=5.610e+00 
R5906t5510 n5907 n5511 R=5.909e+02 
R5906t2325 n5907 n2326 R=3.747e+01 
R5906t3180 n5907 n3181 R=4.294e+01 
R5906t3159 n5907 n3160 R=3.291e+00 
R5907t812 n5908 n813 R=2.227e+01 
R5907t5608 n5908 n5609 R=2.520e+00 
R5907t498 n5908 n499 R=2.226e+01 
R5907t2655 n5908 n2656 R=5.040e+00 
R5908t819 n5909 n820 R=7.621e+00 
R5908t3208 n5909 n3209 R=8.022e+00 
R5908t3030 n5909 n3031 R=4.465e+00 
R5909t4758 n1 n4759 R=4.657e+00 
R5911t1077 n5912 n1078 R=9.861e+00 
R5911t3858 n5912 n3859 R=2.301e+00 
R5912t906 n5913 n907 R=7.182e+00 
R5912t2225 n5913 n2226 R=3.065e+00 
R5912t569 n5913 n570 R=3.153e+00 
R5913t16 n5914 n17 R=1.157e+01 
R5913t1072 n5914 n1073 R=7.930e+00 
R5913t1855 n5914 n1856 R=5.953e+00 
R5913t5751 n5914 n5752 R=4.129e+00 
R5914t3971 n5915 n3972 R=3.073e+00 
R5914t567 n5915 n568 R=9.055e+00 
R5914t3248 n5915 n3249 R=5.898e+00 
R5915t4094 n5916 n4095 R=1.348e+02 
R5915t5039 n5916 n5040 R=4.639e+00 
R5915t2719 n5916 n2720 R=1.381e+01 
R5916t5437 n5917 n5438 R=5.611e+00 
R5916t1688 n5917 n1689 R=6.007e+01 
R5916t4673 n5917 n4674 R=1.051e+01 
R5916t1660 n5917 n1661 R=4.310e+00 
R5916t4913 n5917 n4914 R=1.159e+01 
R5917t691 n5918 n692 R=5.396e+00 
R5917t2689 n5918 n2690 R=3.869e+00 
R5918t1345 n5919 n1346 R=5.071e+01 
R5918t5662 n5919 n5663 R=2.192e+01 
R5918t4523 n5919 n4524 R=5.796e+00 
R5918t3513 n5919 n3514 R=2.200e+01 
R5918t3650 n5919 n3651 R=3.066e+02 
R5918t739 n5919 n740 R=4.944e+00 
R5918t5654 n5919 n5655 R=5.940e+00 
R5919t3542 n5920 n3543 R=9.702e+00 
R5919t932 n5920 n933 R=4.299e+00 
R5919t3452 n5920 n3453 R=5.125e+01 
R5919t5213 n5920 n5214 R=7.245e+00 
R5920t2526 n5921 n2527 R=4.938e+01 
R5920t4627 n5921 n4628 R=1.167e+01 
R5920t20 n5921 n21 R=6.425e+00 
R5920t306 n5921 n307 R=1.156e+02 
R5920t2026 n5921 n2027 R=5.572e+00 
R5921t1034 n5922 n1035 R=1.269e+01 
R5921t4210 n5922 n4211 R=1.988e+02 
R5921t1082 n5922 n1083 R=3.291e+01 
R5922t1783 n5923 n1784 R=1.130e+01 
R5922t3048 n5923 n3049 R=4.821e+00 
R5922t4909 n5923 n4910 R=9.930e+00 
R5922t1238 n5923 n1239 R=2.501e+02 
R5922t290 n5923 n291 R=8.226e+00 
R5922t308 n5923 n309 R=3.410e+01 
R5922t165 n5923 n166 R=3.595e+01 
R5922t3942 n5923 n3943 R=2.792e+01 
R5923t970 n5924 n971 R=4.962e+00 
R5923t5843 n5924 n5844 R=4.919e+00 
R5923t1805 n5924 n1806 R=2.930e+02 
R5924t2814 n5925 n2815 R=4.192e+00 
R5924t4187 n5925 n4188 R=1.423e+01 
R5924t4052 n5925 n4053 R=1.010e+01 
R5924t3194 n5925 n3195 R=4.260e+00 
R5925t2683 n5926 n2684 R=3.228e+01 
R5925t166 n5926 n167 R=1.044e+01 
R5925t1578 n5926 n1579 R=5.001e+00 
R5925t2484 n5926 n2485 R=7.907e+00 
R5926t5386 n5927 n5387 R=1.310e+01 
R5926t4249 n5927 n4250 R=1.717e+01 
R5926t3584 n5927 n3585 R=5.951e+00 
R5927t4269 n5928 n4270 R=1.769e+00 
R5927t1459 n5928 n1460 R=3.760e+01 
R5928t2027 n5929 n2028 R=9.164e+00 
R5928t3700 n5929 n3701 R=1.233e+01 
R5929t1229 n5930 n1230 R=1.230e+01 
R5929t1983 n5930 n1984 R=4.621e+00 
R5929t3901 n5930 n3902 R=1.533e+01 
R5930t4337 n5931 n4338 R=4.760e+00 
R5930t2807 n5931 n2808 R=2.002e+01 
R5930t1510 n5931 n1511 R=8.194e+00 
R5930t572 n5931 n573 R=2.803e+00 
R5931t1792 n5932 n1793 R=3.601e+03 
R5931t1444 n5932 n1445 R=2.991e+00 
R5931t2937 n5932 n2938 R=1.047e+01 
R5932t1920 n1 n1921 R=7.145e+00 
R5932t701 n1 n702 R=1.409e+02 
R5932t3831 n1 n3832 R=3.802e+00 
R5933t951 n5934 n952 R=4.117e+00 
R5934t2343 n5935 n2344 R=6.567e+00 
R5934t5712 n5935 n5713 R=9.279e+00 
R5934t1046 n5935 n1047 R=4.929e+00 
R5934t4273 n5935 n4274 R=5.324e+00 
R5935t2001 n5936 n2002 R=4.956e+00 
R5935t2003 n5936 n2004 R=2.760e+00 
R5935t4665 n5936 n4666 R=8.210e+02 
R5936t3282 n5937 n3283 R=2.499e+00 
R5936t5871 n5937 n5872 R=4.550e+00 
R5936t937 n5937 n938 R=2.490e+01 
R5936t919 n5937 n920 R=1.857e+01 
R5936t3055 n5937 n3056 R=5.652e+01 
R5937t5927 n5938 n5928 R=2.871e+00 
R5937t1459 n5938 n1460 R=8.912e+01 
R5937t4493 n5938 n4494 R=4.237e+01 
R5937t3469 n5938 n3470 R=1.146e+01 
R5938t2817 n5939 n2818 R=5.067e+00 
R5938t4677 n5939 n4678 R=1.624e+01 
R5939t2765 n5940 n2766 R=5.022e+00 
R5939t2168 n5940 n2169 R=4.875e+00 
R5940t4949 n5941 n4950 R=1.037e+01 
R5940t4095 n5941 n4096 R=5.756e+00 
R5941t574 n5942 n575 R=5.168e+00 
R5941t1257 n5942 n1258 R=1.797e+01 
R5941t313 n5942 n314 R=6.061e+01 
R5942t3292 n5943 n3293 R=3.247e+00 
R5942t4608 n5943 n4609 R=7.103e+00 
R5942t2179 n5943 n2180 R=3.275e+00 
R5942t1674 n5943 n1675 R=2.270e+01 
R5942t2659 n5943 n2660 R=7.855e+00 
R5943t978 n5944 n979 R=7.548e+00 
R5943t5190 n5944 n5191 R=4.470e+00 
R5943t5796 n5944 n5797 R=1.260e+01 
R5944t379 n5945 n380 R=1.268e+01 
R5944t5532 n5945 n5533 R=3.277e+01 
R5944t4796 n5945 n4797 R=2.767e+00 
R5944t5124 n5945 n5125 R=6.992e+01 
R5945t875 n5946 n876 R=6.772e+00 
R5945t2729 n5946 n2730 R=1.145e+01 
R5945t5427 n5946 n5428 R=2.950e+01 
R5946t3115 n5947 n3116 R=4.634e+00 
R5946t66 n5947 n67 R=4.680e+00 
R5947t2698 n5948 n2699 R=6.345e+00 
R5947t2842 n5948 n2843 R=2.700e+02 
R5948t1831 n5949 n1832 R=2.555e+00 
R5948t4634 n5949 n4635 R=1.035e+01 
R5948t4712 n5949 n4713 R=2.420e+00 
R5949t1946 n5950 n1947 R=2.984e+01 
R5949t2769 n5950 n2770 R=4.731e+00 
R5950t4822 n5951 n4823 R=2.282e+01 
R5950t5365 n5951 n5366 R=8.717e+00 
R5950t1232 n5951 n1233 R=2.556e+01 
R5950t3167 n5951 n3168 R=4.128e+00 
R5950t690 n5951 n691 R=4.568e+01 
R5950t3593 n5951 n3594 R=7.627e+00 
R5950t2816 n5951 n2817 R=1.978e+01 
R5951t4597 n5952 n4598 R=2.750e+00 
R5951t2727 n5952 n2728 R=6.796e+02 
R5952t3267 n5953 n3268 R=6.129e+01 
R5952t5119 n5953 n5120 R=9.244e+00 
R5952t5015 n5953 n5016 R=2.652e+01 
R5952t4023 n5953 n4024 R=4.880e+00 
R5952t1579 n5953 n1580 R=4.286e+02 
R5952t4529 n5953 n4530 R=1.298e+01 
R5952t3135 n5953 n3136 R=5.507e+00 
R5953t4512 n5954 n4513 R=2.250e+01 
R5953t4152 n5954 n4153 R=2.350e+01 
R5953t109 n5954 n110 R=7.099e+00 
R5953t3675 n5954 n3676 R=3.747e+00 
R5954t4384 n5955 n4385 R=1.090e+01 
R5954t1122 n5955 n1123 R=9.101e+00 
R5955t4509 n5956 n4510 R=6.052e+00 
R5955t2775 n5956 n2776 R=6.638e+01 
R5956t420 n5957 n421 R=7.370e+00 
R5956t1478 n5957 n1479 R=1.458e+01 
R5956t4323 n5957 n4324 R=1.849e+02 
R5956t905 n5957 n906 R=5.400e+00 
R5957t1032 n5958 n1033 R=8.577e+00 
R5957t3703 n5958 n3704 R=3.691e+00 
R5957t5055 n5958 n5056 R=4.962e+00 
R5957t1333 n5958 n1334 R=4.211e+01 
R5958t1669 n5959 n1670 R=4.832e+00 
R5958t5889 n5959 n5890 R=3.318e+00 
R5958t3592 n5959 n3593 R=2.150e+01 
R5959t5619 n5960 n5620 R=2.583e+00 
R5959t84 n5960 n85 R=3.647e+00 
R5960t61 n5961 n62 R=4.297e+00 
R5960t4396 n5961 n4397 R=1.034e+01 
R5960t5885 n5961 n5886 R=2.505e+01 
R5961t973 n5962 n974 R=2.356e+01 
R5961t4948 n5962 n4949 R=6.975e+00 
R5961t2396 n5962 n2397 R=8.785e+00 
R5962t4127 n5963 n4128 R=8.309e+01 
R5962t4178 n5963 n4179 R=3.888e+01 
R5962t3150 n5963 n3151 R=4.015e+00 
R5962t480 n5963 n481 R=4.093e+00 
R5962t551 n5963 n552 R=1.859e+01 
R5962t2596 n5963 n2597 R=1.263e+01 
R5962t2102 n5963 n2103 R=2.744e+00 
R5962t5274 n5963 n5275 R=1.655e+01 
R5963t1755 n5964 n1756 R=4.137e+00 
R5963t4733 n5964 n4734 R=3.689e+01 
R5963t4115 n5964 n4116 R=5.050e+00 
R5963t3237 n5964 n3238 R=4.158e+00 
R5963t702 n5964 n703 R=1.859e+01 
R5963t3622 n5964 n3623 R=1.116e+01 
R5964t725 n5965 n726 R=5.817e+00 
R5964t1445 n5965 n1446 R=3.913e+00 
R5965t4732 n5966 n4733 R=3.841e+00 
R5965t3782 n5966 n3783 R=3.280e+00 
R5965t5456 n5966 n5457 R=7.099e+00 
R5966t1203 n5967 n1204 R=1.040e+01 
R5966t5137 n5967 n5138 R=5.083e+00 
R5966t5487 n5967 n5488 R=4.741e+01 
R5967t2178 n5968 n2179 R=1.611e+01 
R5967t3551 n5968 n3552 R=4.724e+00 
R5967t1813 n5968 n1814 R=2.865e+00 
R5967t4590 n5968 n4591 R=5.858e+00 
R5968t2550 n5969 n2551 R=2.722e+00 
R5968t213 n5969 n214 R=1.947e+00 
R5968t677 n5969 n678 R=2.784e+01 
R5969t1603 n5970 n1604 R=7.252e+00 
R5969t4257 n5970 n4258 R=5.635e+00 
R5969t3404 n5970 n3405 R=5.858e+00 
R5969t1436 n5970 n1437 R=2.391e+01 
R5969t4229 n5970 n4230 R=1.752e+01 
R5969t5854 n5970 n5855 R=1.011e+01 
R5970t3192 n5971 n3193 R=2.929e+00 
R5970t1370 n5971 n1371 R=1.302e+01 
R5970t992 n5971 n993 R=4.298e+00 
R5971t2060 n5972 n2061 R=1.979e+01 
R5971t3289 n5972 n3290 R=3.240e+01 
R5971t4966 n5972 n4967 R=6.083e+00 
R5972t4248 n5973 n4249 R=2.269e+01 
R5972t4126 n5973 n4127 R=1.612e+01 
R5972t1166 n5973 n1167 R=6.195e+00 
R5973t812 n5974 n813 R=7.239e+00 
R5973t928 n5974 n929 R=8.374e+00 
R5973t4846 n5974 n4847 R=4.801e+00 
R5974t1336 n5975 n1337 R=3.283e+01 
R5974t5603 n5975 n5604 R=2.206e+01 
R5974t225 n5975 n226 R=2.719e+00 
R5974t1261 n5975 n1262 R=4.758e+00 
R5974t4840 n5975 n4841 R=2.869e+02 
R5975t4251 n5976 n4252 R=6.283e+00 
R5975t5068 n5976 n5069 R=7.134e+00 
R5975t4101 n5976 n4102 R=2.876e+00 
R5975t2341 n5976 n2342 R=4.724e+01 
R5975t4931 n5976 n4932 R=6.418e+00 
R5976t964 n5977 n965 R=1.016e+01 
R5976t3401 n5977 n3402 R=8.672e+00 
R5976t5743 n5977 n5744 R=5.375e+00 
R5977t4588 n5978 n4589 R=2.546e+00 
R5978t1358 n5979 n1359 R=3.755e+00 
R5978t2837 n5979 n2838 R=1.162e+01 
R5979t2060 n5980 n2061 R=5.082e+00 
R5979t5971 n5980 n5972 R=1.374e+01 
R5979t3679 n5980 n3680 R=1.461e+01 
R5979t122 n5980 n123 R=8.440e+01 
R5980t654 n5981 n655 R=5.388e+00 
R5980t2129 n5981 n2130 R=1.761e+01 
R5980t1384 n5981 n1385 R=1.376e+01 
R5980t3727 n5981 n3728 R=3.216e+00 
R5980t5877 n5981 n5878 R=1.712e+01 
R5981t4411 n5982 n4412 R=4.484e+01 
R5981t4692 n5982 n4693 R=1.071e+01 
R5981t3888 n5982 n3889 R=7.388e+00 
R5981t5412 n5982 n5413 R=6.762e+00 
R5981t865 n5982 n866 R=1.887e+01 
R5982t2382 n5983 n2383 R=2.412e+00 
R5982t2831 n5983 n2832 R=3.450e+00 
R5983t4412 n5984 n4413 R=4.606e+00 
R5983t308 n5984 n309 R=1.575e+01 
R5984t1814 n5985 n1815 R=1.652e+00 
R5984t3860 n5985 n3861 R=9.907e+00 
R5984t2975 n5985 n2976 R=4.169e+01 
R5984t1242 n5985 n1243 R=3.184e+00 
R5985t553 n5986 n554 R=4.506e+00 
R5986t2351 n5987 n2352 R=3.169e+00 
R5986t938 n5987 n939 R=1.639e+01 
R5986t3381 n5987 n3382 R=4.104e+00 
R5987t1900 n5988 n1901 R=8.507e+00 
R5987t3834 n5988 n3835 R=7.219e+00 
R5987t581 n5988 n582 R=2.547e+01 
R5987t3582 n5988 n3583 R=1.261e+01 
R5988t2921 n5989 n2922 R=6.571e+00 
R5988t5153 n5989 n5154 R=9.485e+00 
R5989t1686 n5990 n1687 R=5.645e+00 
R5989t2031 n5990 n2032 R=2.200e+02 
R5989t3053 n5990 n3054 R=4.954e+00 
R5989t2316 n5990 n2317 R=1.077e+01 
R5989t3605 n5990 n3606 R=1.225e+01 
R5990t3131 n5991 n3132 R=2.428e+00 
R5990t194 n5991 n195 R=1.225e+01 
R5990t385 n5991 n386 R=5.492e+00 
R5990t2615 n5991 n2616 R=1.117e+01 
R5991t5639 n5992 n5640 R=3.000e+00 
R5991t5877 n5992 n5878 R=3.769e+00 
R5992t2825 n5993 n2826 R=4.563e+00 
R5992t5281 n5993 n5282 R=6.997e+00 
R5993t4375 n5994 n4376 R=4.798e+00 
R5993t1260 n5994 n1261 R=8.684e+00 
R5994t2008 n5995 n2009 R=6.852e+00 
R5994t5631 n5995 n5632 R=1.331e+01 
R5994t1040 n5995 n1041 R=8.781e+00 
R5994t4139 n5995 n4140 R=1.857e+01 
R5995t4724 n5996 n4725 R=4.562e+01 
R5996t2180 n5997 n2181 R=2.118e+01 
R5996t5754 n5997 n5755 R=2.017e+00 
R5997t1087 n5998 n1088 R=1.090e+02 
R5997t4452 n5998 n4453 R=2.520e+00 
R5997t2838 n5998 n2839 R=1.923e+02 
R5998t2632 n5999 n2633 R=2.867e+01 
R5998t2861 n5999 n2862 R=9.287e+00 
R5998t3559 n5999 n3560 R=5.910e+01 
R5998t4206 n5999 n4207 R=5.575e+00 
R5999t3459 n6000 n3460 R=3.645e+00 
R5999t1540 n6000 n1541 R=2.323e+01 
R5999t4090 n6000 n4091 R=2.777e+00 
R5999t236 n6000 n237 R=8.422e+00 
R6000t2928 n6001 n2929 R=3.321e+00 
R6000t4730 n6001 n4731 R=8.817e+00 
R6000t5933 n6001 n5934 R=1.593e+01 
R6001t3932 n6002 n3933 R=1.896e+02 
R6001t3079 n6002 n3080 R=1.261e+01 
R6001t3590 n6002 n3591 R=8.852e+00 
R6001t5248 n6002 n5249 R=4.136e+00 
R6002t2595 n6003 n2596 R=1.041e+01 
R6003t4461 n6004 n4462 R=1.571e+01 
R6003t4895 n6004 n4896 R=9.871e+00 
R6003t627 n6004 n628 R=1.830e+01 
R6003t2497 n6004 n2498 R=4.431e+00 
R6003t2827 n6004 n2828 R=1.985e+01 
R6003t1087 n6004 n1088 R=1.993e+01 
R6003t5488 n6004 n5489 R=5.101e+00 
R6004t956 n6005 n957 R=4.421e+00 
R6004t3001 n6005 n3002 R=7.479e+00 
R6004t3018 n6005 n3019 R=8.026e+00 
R6005t2322 n6006 n2323 R=3.850e+00 
R6005t364 n6006 n365 R=2.294e+01 
R6005t2535 n6006 n2536 R=3.362e+00 
R6005t3879 n6006 n3880 R=2.269e+01 
R6005t822 n6006 n823 R=4.095e+00 
R6006t719 n6007 n720 R=3.373e+01 
R6006t1223 n6007 n1224 R=4.926e+00 
R6007t177 n6008 n178 R=3.122e+00 
R6007t2981 n6008 n2982 R=5.150e+01 
R6007t1404 n6008 n1405 R=1.068e+01 
R6007t4786 n6008 n4787 R=3.128e+00 
R6008t1560 n6009 n1561 R=2.985e+00 
R6008t5024 n6009 n5025 R=2.765e+01 
R6008t3682 n6009 n3683 R=2.743e+00 
R6008t2296 n6009 n2297 R=1.441e+01 
R6008t245 n6009 n246 R=1.835e+01 
R6009t4017 n6010 n4018 R=3.946e+00 
R6009t405 n6010 n406 R=5.866e+01 
R6009t2668 n6010 n2669 R=3.760e+00 
R6009t1206 n6010 n1207 R=5.421e+00 
R6009t1406 n6010 n1407 R=1.018e+01 
R6010t1466 n6011 n1467 R=7.327e+02 
R6010t3554 n6011 n3555 R=2.833e+00 
R6010t1515 n6011 n1516 R=2.534e+01 
R6010t2949 n6011 n2950 R=1.154e+01 
R6011t426 n6012 n427 R=5.195e+00 
R6011t3957 n6012 n3958 R=9.629e+00 
R6011t1047 n6012 n1048 R=6.691e+00 
R6011t3341 n6012 n3342 R=8.970e+01 
R6012t4074 n6013 n4075 R=7.613e+00 
R6012t4744 n6013 n4745 R=7.205e+00 
R6012t3437 n6013 n3438 R=7.879e+00 
R6012t4758 n6013 n4759 R=6.600e+00 
R6013t2726 n6014 n2727 R=4.289e+00 
R6013t352 n6014 n353 R=3.953e+00 
R6013t4987 n6014 n4988 R=5.598e+01 
R6014t3945 n6015 n3946 R=2.376e+00 
R6014t4630 n6015 n4631 R=6.500e+01 
R6014t2385 n6015 n2386 R=4.258e+00 
R6014t2639 n6015 n2640 R=4.309e+01 
R6015t757 n6016 n758 R=3.472e+00 
R6015t5545 n6016 n5546 R=2.243e+01 
R6015t3563 n6016 n3564 R=1.464e+01 
R6015t4878 n6016 n4879 R=2.239e+00 
R6015t3127 n6016 n3128 R=2.126e+01 
R6016t3412 n6017 n3413 R=5.173e+00 
R6016t5012 n6017 n5013 R=3.025e+01 
R6016t2911 n6017 n2912 R=3.265e+00 
R6016t3555 n6017 n3556 R=1.401e+02 
R6016t4885 n6017 n4886 R=8.168e+00 
R6017t2252 n6018 n2253 R=4.039e+00 
R6017t3774 n6018 n3775 R=7.414e+00 
R6018t1284 n6019 n1285 R=3.940e+01 
R6018t4350 n6019 n4351 R=5.840e+00 
R6018t683 n6019 n684 R=9.667e+00 
R6018t1840 n6019 n1841 R=7.953e+00 
R6018t3867 n6019 n3868 R=3.245e+00 
R6019t3283 n6020 n3284 R=8.771e+00 
R6019t3402 n6020 n3403 R=2.494e+02 
R6019t5392 n6020 n5393 R=9.725e+00 
R6019t2622 n6020 n2623 R=1.008e+02 
R6020t5509 n6021 n5510 R=5.009e+00 
R6020t3835 n6021 n3836 R=3.420e+01 
R6020t2934 n6021 n2935 R=5.319e+00 
R6020t2325 n6021 n2326 R=7.799e+00 
R6020t3017 n6021 n3018 R=2.955e+01 
R6021t5685 n6022 n5686 R=4.119e+00 
R6021t4186 n6022 n4187 R=5.860e+00 
R6021t3994 n6022 n3995 R=6.805e+00 
R6022t4540 n6023 n4541 R=2.767e+01 
R6022t708 n6023 n709 R=2.384e+01 
R6022t4392 n6023 n4393 R=6.406e+00 
R6023t2728 n6024 n2729 R=5.178e+00 
R6023t4177 n6024 n4178 R=3.249e+01 
R6023t4926 n6024 n4927 R=1.497e+01 
R6023t166 n6024 n167 R=2.357e+01 
R6023t2683 n6024 n2684 R=1.148e+01 
R6023t3849 n6024 n3850 R=7.590e+00 
R6024t410 n6025 n411 R=8.324e+00 
R6024t5876 n6025 n5877 R=7.440e+00 
R6024t4952 n6025 n4953 R=7.530e+00 
R6024t5525 n6025 n5526 R=3.954e+00 
R6025t1673 n6026 n1674 R=5.255e+00 
R6025t114 n6026 n115 R=2.986e+01 
R6025t47 n6026 n48 R=3.252e+00 
R6026t2248 n6027 n2249 R=6.298e+00 
R6026t3753 n6027 n3754 R=1.641e+01 
R6026t2484 n6027 n2485 R=9.292e+00 
R6026t5925 n6027 n5926 R=1.490e+01 
R6027t4840 n6028 n4841 R=7.777e+00 
R6027t4313 n6028 n4314 R=1.834e+00 
R6027t3868 n6028 n3869 R=2.078e+02 
R6027t5401 n6028 n5402 R=5.972e+00 
R6028t3 n6029 n4 R=2.020e+00 
R6028t3552 n6029 n3553 R=3.661e+01 
R6028t4470 n6029 n4471 R=5.394e+01 
R6028t4172 n6029 n4173 R=5.190e+00 
R6029t575 n6030 n576 R=2.903e+01 
R6029t2276 n6030 n2277 R=3.138e+00 
R6029t4130 n6030 n4131 R=5.104e+00 
R6030t1725 n6031 n1726 R=1.328e+01 
R6030t4336 n6031 n4337 R=2.174e+00 
R6030t1700 n6031 n1701 R=1.744e+00 
R6030t1840 n6031 n1841 R=2.735e+01 
R6030t3867 n6031 n3868 R=1.386e+02 
R6031t1132 n6032 n1133 R=4.596e+00 
R6031t3479 n6032 n3480 R=7.968e+00 
R6031t1096 n6032 n1097 R=9.160e+00 
R6031t3416 n6032 n3417 R=1.156e+01 
R6031t1619 n6032 n1620 R=3.295e+01 
R6031t4109 n6032 n4110 R=1.111e+01 
R6032t2609 n6033 n2610 R=4.445e+00 
R6032t3129 n6033 n3130 R=5.916e+00 
R6032t5422 n6033 n5423 R=3.121e+01 
R6032t5479 n6033 n5480 R=8.733e+00 
R6033t1737 n6034 n1738 R=8.040e+00 
R6033t2564 n6034 n2565 R=1.416e+01 
R6034t1954 n6035 n1955 R=1.082e+01 
R6034t1093 n6035 n1094 R=2.051e+01 
R6034t4577 n6035 n4578 R=1.530e+01 
R6035t3610 n6036 n3611 R=8.227e+00 
R6035t4395 n6036 n4396 R=3.284e+01 
R6035t4400 n6036 n4401 R=1.095e+01 
R6035t3339 n6036 n3340 R=6.388e+00 
R6035t2212 n6036 n2213 R=1.031e+01 
R6036t1401 n6037 n1402 R=2.922e+00 
R6036t1968 n6037 n1969 R=3.486e+01 
R6036t4521 n6037 n4522 R=6.654e+00 
R6036t3672 n6037 n3673 R=5.322e+00 
R6036t5374 n6037 n5375 R=7.402e+01 
R6036t3860 n6037 n3861 R=5.304e+00 
R6036t1713 n6037 n1714 R=4.736e+01 
R6037t3287 n6038 n3288 R=7.644e+00 
R6037t5900 n6038 n5901 R=1.369e+01 
R6037t5378 n6038 n5379 R=1.070e+01 
R6037t5261 n6038 n5262 R=6.389e+00 
R6038t3966 n6039 n3967 R=5.418e+00 
R6038t1420 n6039 n1421 R=9.497e+00 
R6039t485 n6040 n486 R=1.450e+01 
R6039t829 n6040 n830 R=3.959e+01 
R6039t5042 n6040 n5043 R=3.021e+01 
R6039t910 n6040 n911 R=3.990e+00 
R6040t1151 n6041 n1152 R=4.472e+00 
R6040t4963 n6041 n4964 R=4.646e+02 
R6040t3493 n6041 n3494 R=9.606e+00 
R6040t3786 n6041 n3787 R=6.542e+00 
R6040t337 n6041 n338 R=1.107e+01 
R6040t5590 n6041 n5591 R=4.270e+00 
R6040t1928 n6041 n1929 R=6.123e+01 
R6042t4726 n6043 n4727 R=1.062e+02 
R6042t5773 n6043 n5774 R=2.642e+01 
R6042t1958 n6043 n1959 R=7.245e+00 
R6042t4083 n6043 n4084 R=2.485e+00 
R6043t461 n6044 n462 R=9.456e+01 
R6043t1483 n6044 n1484 R=2.326e+00 
R6044t2392 n6045 n2393 R=1.044e+01 
R6044t1936 n6045 n1937 R=3.228e+00 
R6044t2653 n6045 n2654 R=1.349e+01 
R6045t401 n6046 n402 R=5.556e+00 
R6045t4119 n6046 n4120 R=3.778e+00 
R6045t2420 n6046 n2421 R=3.418e+00 
R6045t3932 n6046 n3933 R=2.128e+01 
R6046t3400 n6047 n3401 R=3.326e+00 
R6046t669 n6047 n670 R=7.283e+00 
R6046t2106 n6047 n2107 R=1.226e+01 
R6046t3762 n6047 n3763 R=1.386e+01 
R6047t363 n6048 n364 R=6.731e+00 
R6047t4172 n6048 n4173 R=5.707e+00 
R6047t1655 n6048 n1656 R=1.792e+01 
R6047t2982 n6048 n2983 R=3.050e+01 
R6047t704 n6048 n705 R=1.133e+01 
R6047t1212 n6048 n1213 R=1.974e+02 
R6048t656 n6049 n657 R=8.937e+01 
R6048t2053 n6049 n2054 R=5.332e+00 
R6048t5411 n6049 n5412 R=4.537e+00 
R6048t4583 n6049 n4584 R=7.411e+00 
R6048t4777 n6049 n4778 R=2.731e+00 
R6048t4310 n6049 n4311 R=4.563e+01 
R6049t1379 n6050 n1380 R=5.993e+00 
R6049t3795 n6050 n3796 R=2.391e+01 
R6049t2017 n6050 n2018 R=3.568e+00 
R6049t2213 n6050 n2214 R=1.314e+02 
R6049t1053 n6050 n1054 R=1.734e+01 
R6049t2576 n6050 n2577 R=2.142e+01 
R6049t3394 n6050 n3395 R=5.243e+02 
R6050t3012 n6051 n3013 R=2.331e+02 
R6050t4623 n6051 n4624 R=3.656e+00 
R6050t1345 n6051 n1346 R=8.078e+01 
R6050t4341 n6051 n4342 R=3.021e+00 
R6050t5543 n6051 n5544 R=9.948e+00 
R6051t5408 n6052 n5409 R=3.473e+00 
R6051t4013 n6052 n4014 R=2.225e+00 
R6052t1028 n6053 n1029 R=5.229e+00 
R6052t2974 n6053 n2975 R=4.686e+00 
R6052t5620 n6053 n5621 R=3.615e+00 
R6053t5814 n6054 n5815 R=9.232e+00 
R6053t2041 n6054 n2042 R=4.480e+00 
R6053t4281 n6054 n4282 R=3.795e+00 
R6053t553 n6054 n554 R=3.206e+01 
R6053t3481 n6054 n3482 R=4.502e+00 
R6054t5361 n6055 n5362 R=1.033e+01 
R6054t5589 n6055 n5590 R=7.888e+00 
R6055t5000 n6056 n5001 R=5.108e+00 
R6055t3153 n6056 n3154 R=6.135e+00 
R6055t3386 n6056 n3387 R=2.702e+01 
R6055t1517 n6056 n1518 R=7.865e+01 
R6055t4612 n6056 n4613 R=5.810e+00 
R6056t4187 n6057 n4188 R=2.077e+00 
R6056t3172 n6057 n3173 R=8.757e+00 
R6056t3754 n6057 n3755 R=2.898e+00 
R6056t5776 n6057 n5777 R=3.879e+01 
R6056t3194 n6057 n3195 R=5.754e+01 
R6056t5924 n6057 n5925 R=1.270e+01 
R6057t3704 n6058 n3705 R=5.667e+00 
R6057t1211 n6058 n1212 R=7.453e+01 
R6057t1677 n6058 n1678 R=5.562e+00 
R6057t317 n6058 n318 R=7.489e+00 
R6057t4652 n6058 n4653 R=7.390e+00 
R6058t2563 n6059 n2564 R=4.338e+01 
R6058t5382 n6059 n5383 R=1.049e+01 
R6058t5397 n6059 n5398 R=3.749e+00 
R6058t3059 n6059 n3060 R=5.298e+01 
R6058t3683 n6059 n3684 R=1.326e+01 
R6059t3313 n6060 n3314 R=1.551e+01 
R6059t662 n6060 n663 R=6.695e+00 
R6059t3800 n6060 n3801 R=1.000e+02 
R6059t5249 n6060 n5250 R=2.758e+00 
R6060t3151 n6061 n3152 R=6.146e+00 
R6060t4841 n6061 n4842 R=4.202e+00 
R6061t2008 n6062 n2009 R=6.234e+01 
R6061t3850 n6062 n3851 R=8.085e+00 
R6061t4603 n6062 n4604 R=3.772e+00 
R6062t5206 n6063 n5207 R=6.403e+00 
R6062t3852 n6063 n3853 R=7.269e+00 
R6062t469 n6063 n470 R=1.355e+01 
R6062t1594 n6063 n1595 R=2.226e+01 
R6063t1238 n6064 n1239 R=4.815e+00 
R6063t4909 n6064 n4910 R=4.943e+01 
R6063t3096 n6064 n3097 R=2.455e+01 
R6063t3324 n6064 n3325 R=8.647e+00 
R6063t5861 n6064 n5862 R=4.693e+00 
R6063t1340 n6064 n1341 R=7.866e+00 
R6063t5033 n6064 n5034 R=1.736e+01 
R6064t347 n6065 n348 R=9.053e+00 
R6064t3270 n6065 n3271 R=3.908e+00 
R6064t2557 n6065 n2558 R=2.691e+02 
R6064t5077 n6065 n5078 R=4.630e+00 
R6065t152 n6066 n153 R=1.669e+01 
R6065t5009 n6066 n5010 R=6.028e+01 
R6065t3151 n6066 n3152 R=1.164e+01 
R6065t2752 n6066 n2753 R=6.292e+00 
R6065t794 n6066 n795 R=1.792e+01 
R6065t3378 n6066 n3379 R=5.508e+00 
R6066t2459 n6067 n2460 R=5.161e+01 
R6066t5041 n6067 n5042 R=2.068e+00 
R6066t3157 n6067 n3158 R=8.332e+00 
R6066t3142 n6067 n3143 R=8.259e+00 
R6066t5453 n6067 n5454 R=4.787e+01 
R6067t1028 n6068 n1029 R=6.489e+01 
R6067t2974 n6068 n2975 R=2.105e+00 
R6067t1596 n6068 n1597 R=3.853e+00 
R6067t4288 n6068 n4289 R=6.321e+00 
R6067t5620 n6068 n5621 R=4.816e+01 
R6068t4592 n6069 n4593 R=9.170e+00 
R6068t3631 n6069 n3632 R=5.872e+00 
R6069t2494 n6070 n2495 R=5.090e+00 
R6069t3470 n6070 n3471 R=1.668e+01 
R6069t2556 n6070 n2557 R=1.463e+02 
R6069t4887 n6070 n4888 R=3.774e+01 
R6070t173 n6071 n174 R=1.706e+01 
R6070t4577 n6071 n4578 R=2.546e+00 
R6070t627 n6071 n628 R=3.294e+00 
R6070t292 n6071 n293 R=6.748e+00 
R6071t2141 n6072 n2142 R=5.149e+00 
R6071t3169 n6072 n3170 R=4.037e+00 
R6071t365 n6072 n366 R=7.408e+00 
R6071t2422 n6072 n2423 R=3.639e+00 
R6072t1266 n6073 n1267 R=3.748e+01 
R6072t3529 n6073 n3530 R=8.358e+00 
R6072t597 n6073 n598 R=2.432e+00 
R6073t4799 n6074 n4800 R=5.305e+00 
R6074t4222 n6075 n4223 R=6.635e+01 
R6074t4567 n6075 n4568 R=5.800e+00 
R6074t5056 n6075 n5057 R=1.024e+01 
R6074t3231 n6075 n3232 R=4.351e+00 
R6074t3281 n6075 n3282 R=3.307e+01 
R6075t479 n6076 n480 R=4.707e+00 
R6075t4693 n6076 n4694 R=8.736e+01 
R6075t5858 n6076 n5859 R=2.824e+00 
R6075t4907 n6076 n4908 R=4.337e+01 
R6075t2688 n6076 n2689 R=1.385e+01 
R6076t5073 n6077 n5074 R=3.668e+01 
R6076t3395 n6077 n3396 R=1.939e+00 
R6076t5887 n6077 n5888 R=1.861e+01 
R6077t1712 n6078 n1713 R=5.877e+00 
R6077t4607 n6078 n4608 R=6.419e+01 
R6077t2498 n6078 n2499 R=1.684e+01 
R6077t4988 n6078 n4989 R=5.013e+00 
R6078t2200 n6079 n2201 R=1.433e+01 
R6078t2903 n6079 n2904 R=3.233e+00 
R6078t4985 n6079 n4986 R=1.551e+01 
R6079t880 n6080 n881 R=4.572e+00 
R6079t2385 n6080 n2386 R=1.958e+01 
R6079t3569 n6080 n3570 R=2.350e+00 
R6080t2157 n6081 n2158 R=6.972e+01 
R6080t3381 n6081 n3382 R=1.261e+01 
R6080t4672 n6081 n4673 R=3.851e+00 
R6080t946 n6081 n947 R=1.913e+01 
R6081t20 n6082 n21 R=5.804e+00 
R6081t4627 n6082 n4628 R=7.903e+00 
R6081t963 n6082 n964 R=1.363e+01 
R6082t3331 n6083 n3332 R=5.070e+01 
R6082t5344 n6083 n5345 R=2.664e+03 
R6082t1171 n6083 n1172 R=6.575e+00 
R6083t2197 n6084 n2198 R=5.043e+00 
R6083t3687 n6084 n3688 R=1.000e+01 
R6083t3577 n6084 n3578 R=4.276e+01 
R6084t4932 n6085 n4933 R=1.658e+01 
R6084t5029 n6085 n5030 R=1.315e+01 
R6085t96 n6086 n97 R=2.663e+00 
R6085t3665 n6086 n3666 R=7.123e+01 
R6085t4659 n6086 n4660 R=8.953e+01 
R6085t4488 n6086 n4489 R=8.773e+00 
R6085t1264 n6086 n1265 R=3.006e+02 
R6086t555 n6087 n556 R=2.747e+00 
R6087t3337 n6088 n3338 R=8.645e+00 
R6087t67 n6088 n68 R=4.813e+00 
R6087t59 n6088 n60 R=7.900e+00 
R6087t4929 n6088 n4930 R=1.206e+01 
R6087t463 n6088 n464 R=3.260e+00 
R6088t4422 n6089 n4423 R=3.638e+00 
R6088t5623 n6089 n5624 R=3.494e+01 
R6088t5107 n6089 n5108 R=6.557e+00 
R6088t2064 n6089 n2065 R=5.002e+00 
R6089t3199 n6090 n3200 R=5.041e+00 
R6089t4591 n6090 n4592 R=3.496e+00 
R6090t3168 n6091 n1 R=4.391e+00 
R6091t183 n6092 n184 R=1.581e+01 
R6091t5321 n6092 n5322 R=1.443e+01 
R6091t1235 n6092 n1236 R=6.021e+00 
R6091t2778 n6092 n2779 R=6.865e+00 
R6092t216 n6093 n217 R=1.578e+01 
R6092t3521 n6093 n3522 R=3.185e+00 
R6092t1384 n6093 n1385 R=1.983e+01 
R6092t3738 n6093 n3739 R=9.952e+00 
R6092t1917 n6093 n1918 R=2.862e+02 
R6093t2895 n6094 n2896 R=1.341e+02 
R6093t3946 n6094 n3947 R=5.462e+02 
R6093t229 n6094 n230 R=5.393e+00 
R6093t5388 n6094 n5389 R=5.897e+00 
R6093t4349 n6094 n4350 R=3.672e+00 
R6094t922 n6095 n923 R=2.846e+00 
R6094t5481 n6095 n5482 R=4.055e+00 
R6094t392 n6095 n393 R=2.785e+01 
R6094t1365 n6095 n1366 R=4.726e+00 
R6094t5423 n6095 n5424 R=1.466e+01 
R6095t846 n6096 n847 R=4.966e+00 
R6095t2495 n6096 n2496 R=9.094e+00 
R6095t3748 n6096 n3749 R=2.013e+01 
R6096t1153 n6097 n1154 R=3.336e+00 
R6096t1865 n6097 n1866 R=1.301e+01 
R6096t4448 n6097 n4449 R=6.392e+00 
R6096t170 n6097 n171 R=3.039e+01 
R6097t5877 n6098 n5878 R=4.594e+02 
R6097t4557 n6098 n4558 R=8.161e+00 
R6097t2085 n6098 n2086 R=2.642e+00 
R6097t3727 n6098 n3728 R=2.855e+01 
R6098t217 n6099 n218 R=4.236e+01 
R6098t2401 n6099 n2402 R=2.293e+00 
R6099t4479 n6100 n4480 R=3.470e+01 
R6099t5383 n6100 n5384 R=3.081e+00 
R6099t3452 n6100 n3453 R=2.082e+01 
R6099t932 n6100 n933 R=1.912e+00 
R6100t3471 n6101 n3472 R=1.940e+01 
R6100t5888 n6101 n5889 R=1.078e+01 
R6100t1297 n6101 n1298 R=3.596e+00 
R6100t4829 n6101 n4830 R=4.831e+01 
R6101t653 n6102 n654 R=5.145e+01 
R6101t1805 n6102 n1806 R=8.582e+00 
R6101t4285 n6102 n4286 R=2.041e+00 
R6102t1176 n6103 n1177 R=6.715e+00 
R6102t881 n6103 n882 R=8.082e+00 
R6102t3029 n6103 n3030 R=7.603e+00 
R6103t2498 n6104 n2499 R=5.406e+00 
R6103t2169 n6104 n2170 R=1.317e+01 
R6103t523 n6104 n524 R=1.656e+02 
R6103t3506 n6104 n3507 R=1.206e+01 
R6103t3085 n6104 n3086 R=3.301e+01 
R6104t4779 n6105 n4780 R=3.065e+01 
R6104t3787 n6105 n3788 R=3.860e+00 
R6104t2615 n6105 n2616 R=2.701e+00 
R6104t5990 n6105 n5991 R=2.254e+01 
R6105t23 n6106 n24 R=9.060e+00 
R6105t3491 n6106 n3492 R=1.238e+01 
R6105t603 n6106 n604 R=5.067e+00 
R6105t4805 n6106 n4806 R=3.110e+01 
R6105t2841 n6106 n2842 R=7.171e+00 
R6106t2248 n6107 n2249 R=2.298e+01 
R6106t3753 n6107 n3754 R=4.118e+00 
R6106t6026 n6107 n6027 R=1.792e+01 
R6107t1883 n6108 n1884 R=3.197e+01 
R6107t3402 n6108 n3403 R=2.122e+02 
R6107t901 n6108 n902 R=2.799e+01 
R6107t5762 n6108 n5763 R=6.501e+00 
R6107t5392 n6108 n5393 R=5.022e+00 
R6107t6019 n6108 n6020 R=1.949e+01 
R6108t5332 n6109 n5333 R=2.238e+01 
R6108t2369 n6109 n2370 R=1.916e+01 
R6108t3666 n6109 n3667 R=2.864e+01 
R6109t2448 n6110 n2449 R=3.714e+00 
R6109t3757 n6110 n3758 R=6.566e+00 
R6109t4910 n6110 n4911 R=6.954e+00 
R6109t137 n6110 n138 R=1.557e+01 
R6109t1069 n6110 n1070 R=6.096e+00 
R6110t3604 n6111 n3605 R=2.988e+01 
R6110t4911 n6111 n4912 R=8.708e+00 
R6111t991 n6112 n992 R=2.511e+01 
R6111t4231 n6112 n4232 R=8.733e+00 
R6111t1307 n6112 n1308 R=2.512e+02 
R6112t1252 n6113 n1253 R=8.099e+00 
R6112t5599 n6113 n5600 R=1.542e+01 
R6112t2244 n6113 n2245 R=5.088e+00 
R6112t1943 n6113 n1944 R=9.819e+00 
R6113t4198 n6114 n4199 R=2.375e+00 
R6113t5804 n6114 n5805 R=6.829e+00 
R6113t3116 n6114 n3117 R=3.071e+00 
R6114t2842 n6115 n2843 R=2.483e+00 
R6114t2585 n6115 n2586 R=2.088e+01 
R6115t4939 n6116 n4940 R=2.017e+01 
R6115t3991 n6116 n3992 R=4.524e+01 
R6115t2112 n6116 n2113 R=1.869e+01 
R6116t1699 n6117 n1700 R=5.171e+00 
R6116t4587 n6117 n4588 R=5.179e+00 
R6116t2028 n6117 n2029 R=6.812e+00 
R6116t1518 n6117 n1519 R=3.190e+01 
R6116t5595 n6117 n5596 R=8.680e+00 
R6116t1310 n6117 n1311 R=1.477e+02 
R6117t3200 n6118 n3201 R=3.760e+00 
R6117t5577 n6118 n5578 R=3.274e+00 
R6117t3013 n6118 n3014 R=3.843e+00 
R6117t2654 n6118 n2655 R=4.085e+01 
R6118t4141 n6119 n4142 R=2.616e+00 
R6118t4337 n6119 n4338 R=1.500e+01 
R6118t5553 n6119 n5554 R=3.603e+00 
R6118t5788 n6119 n5789 R=4.914e+02 
R6118t4737 n6119 n4738 R=7.602e+00 
R6119t1195 n1 n1196 R=6.451e+00 
R6119t2901 n1 n2902 R=1.064e+01 
R6120t885 n6121 n886 R=7.243e+00 
R6120t3096 n6121 n3097 R=5.087e+00 
R6120t3464 n6121 n3465 R=5.941e+00 
R6120t2012 n6121 n2013 R=5.347e+00 
R6121t4144 n6122 n4145 R=2.047e+01 
R6121t5684 n6122 n5685 R=4.329e+00 
R6121t3529 n6122 n3530 R=1.616e+01 
R6121t597 n6122 n598 R=4.549e+00 
R6121t3581 n6122 n3582 R=3.467e+01 
R6122t5562 n6123 n5563 R=1.738e+02 
R6122t3271 n6123 n3272 R=2.821e+01 
R6122t2408 n6123 n2409 R=3.809e+01 
R6122t2148 n6123 n2149 R=3.598e+00 
R6122t6083 n6123 n6084 R=4.285e+00 
R6123t4417 n6124 n4418 R=3.008e+00 
R6123t4944 n6124 n4945 R=2.120e+01 
R6123t1745 n6124 n1746 R=6.556e+00 
R6123t4555 n6124 n4556 R=5.806e+00 
R6123t647 n6124 n648 R=8.532e+01 
R6124t4950 n6125 n4951 R=5.487e+00 
R6124t5587 n6125 n5588 R=1.303e+01 
R6124t2885 n6125 n2886 R=5.030e+00 
R6124t5192 n6125 n5193 R=1.995e+01 
R6125t5562 n6126 n5563 R=5.384e+01 
R6125t614 n6126 n615 R=1.436e+01 
R6125t1208 n6126 n1209 R=1.175e+01 
R6125t2339 n6126 n2340 R=8.403e+00 
R6125t2520 n6126 n2521 R=5.430e+00 
R6126t1457 n6127 n1458 R=5.112e+00 
R6126t560 n6127 n561 R=8.670e+00 
R6126t429 n6127 n430 R=7.591e+00 
R6127t3625 n6128 n3626 R=9.530e+00 
R6127t3691 n6128 n3692 R=1.950e+01 
R6127t1573 n6128 n1574 R=6.025e+00 
R6127t369 n6128 n370 R=2.837e+01 
R6127t1945 n6128 n1946 R=2.304e+01 
R6128t2013 n6129 n2014 R=2.166e+01 
R6128t5417 n6129 n5418 R=2.698e+01 
R6128t163 n6129 n164 R=5.956e+00 
R6128t2916 n6129 n2917 R=1.744e+01 
R6128t2721 n6129 n2722 R=5.685e+00 
R6129t68 n6130 n69 R=5.622e+00 
R6129t4004 n6130 n4005 R=1.231e+02 
R6129t4690 n6130 n4691 R=5.443e+00 
R6129t1516 n6130 n1517 R=2.022e+00 
R6129t3493 n6130 n3494 R=2.932e+01 
R6130t2707 n6131 n2708 R=2.177e+01 
R6130t1095 n6131 n1096 R=4.764e+00 
R6130t605 n6131 n606 R=3.650e+00 
R6130t2297 n6131 n2298 R=8.472e+00 
R6131t2789 n6132 n2790 R=1.646e+01 
R6131t4002 n6132 n4003 R=1.225e+01 
R6131t5078 n6132 n5079 R=3.835e+00 
R6131t5616 n6132 n5617 R=1.315e+01 
R6131t2312 n6132 n2313 R=3.737e+00 
R6132t1798 n6133 n1799 R=2.845e+01 
R6132t3444 n6133 n3445 R=4.804e+00 
R6132t1589 n6133 n1590 R=6.506e+00 
R6132t2016 n6133 n2017 R=1.270e+01 
R6132t5527 n6133 n5528 R=3.308e+02 
R6132t799 n6133 n800 R=9.749e+01 
R6133t375 n6134 n376 R=4.938e+00 
R6133t686 n6134 n687 R=2.511e+00 
R6134t1471 n6135 n1472 R=4.967e+00 
R6134t1770 n6135 n1771 R=3.404e+00 
R6134t5201 n6135 n5202 R=2.791e+01 
R6135t3518 n6136 n3519 R=3.017e+01 
R6135t3561 n6136 n3562 R=4.771e+00 
R6135t320 n6136 n321 R=4.551e+00 
R6135t3515 n6136 n3516 R=9.010e+00 
R6136t2029 n6137 n2030 R=9.077e+00 
R6136t2798 n6137 n2799 R=1.456e+01 
R6136t5722 n6137 n5723 R=7.819e+00 
R6136t1958 n6137 n1959 R=4.510e+00 
R6137t826 n6138 n827 R=1.022e+01 
R6137t1353 n6138 n1354 R=5.165e+00 
R6137t3300 n6138 n3301 R=5.087e+00 
R6138t2634 n6139 n2635 R=7.717e+00 
R6138t5334 n6139 n5335 R=4.479e+02 
R6138t1874 n6139 n1875 R=3.061e+00 
R6138t5672 n6139 n5673 R=1.286e+01 
R6138t3268 n6139 n3269 R=4.779e+00 
R6138t4478 n6139 n4479 R=1.393e+01 
R6139t1737 n6140 n1738 R=3.300e+01 
R6139t3764 n6140 n3765 R=8.112e+00 
R6139t5074 n6140 n5075 R=3.891e+00 
R6139t6033 n6140 n6034 R=8.206e+00 
R6140t3061 n6141 n3062 R=3.744e+00 
R6140t3766 n6141 n3767 R=1.162e+01 
R6140t5240 n6141 n5241 R=2.829e+01 
R6142t1412 n6143 n1413 R=3.357e+01 
R6142t5847 n6143 n5848 R=7.122e+00 
R6142t1653 n6143 n1654 R=1.254e+01 
R6143t3718 n6144 n3719 R=7.041e+00 
R6143t3726 n6144 n3727 R=7.128e+00 
R6143t5001 n6144 n5002 R=9.908e+00 
R6143t2760 n6144 n2761 R=1.067e+01 
R6144t1871 n6145 n1872 R=6.444e+00 
R6144t600 n6145 n601 R=1.100e+01 
R6145t3456 n6146 n3457 R=3.082e+00 
R6145t5076 n6146 n5077 R=1.603e+00 
R6145t1769 n6146 n1770 R=6.748e+00 
R6146t4801 n6147 n4802 R=2.829e+01 
R6146t678 n6147 n679 R=2.984e+00 
R6146t1140 n6147 n1141 R=1.714e+00 
R6147t4876 n6148 n4877 R=1.063e+01 
R6147t2918 n6148 n2919 R=5.620e+00 
R6147t2114 n6148 n2115 R=1.925e+02 
R6147t5371 n6148 n5372 R=2.194e+01 
R6147t1719 n6148 n1720 R=7.625e+00 
R6148t464 n6149 n465 R=9.571e+01 
R6148t3801 n6149 n3802 R=3.807e+00 
R6149t2388 n6150 n2389 R=7.028e+00 
R6149t818 n6150 n819 R=5.935e+00 
R6150t5039 n6151 n5040 R=1.808e+01 
R6150t5179 n6151 n5180 R=2.301e+01 
R6150t2233 n6151 n2234 R=2.115e+03 
R6150t5915 n6151 n5916 R=1.384e+01 
R6151t1243 n6152 n1244 R=5.671e+00 
R6151t5385 n6152 n5386 R=4.752e+00 
R6151t2209 n6152 n2210 R=8.047e+00 
R6151t3550 n6152 n3551 R=3.923e+00 
R6152t1456 n6153 n1457 R=2.983e+00 
R6152t1709 n6153 n1710 R=3.531e+00 
R6153t5273 n6154 n5274 R=6.368e+01 
R6153t904 n6154 n905 R=1.609e+01 
R6153t116 n6154 n117 R=2.954e+00 
R6153t4575 n6154 n4576 R=7.355e+00 
R6154t530 n6155 n531 R=4.099e+01 
R6154t3038 n6155 n3039 R=9.418e+00 
R6154t703 n6155 n704 R=2.069e+00 
R6155t3241 n6156 n3242 R=9.677e+00 
R6155t1897 n6156 n1898 R=1.417e+01 
R6156t3349 n6157 n3350 R=4.538e+01 
R6156t533 n6157 n534 R=1.326e+02 
R6156t239 n6157 n240 R=3.460e+00 
R6156t2245 n6157 n2246 R=2.422e+00 
R6157t1121 n6158 n1122 R=1.432e+01 
R6157t3184 n6158 n3185 R=6.049e+00 
R6157t447 n6158 n448 R=7.725e+00 
R6157t2250 n6158 n2251 R=5.239e+00 
R6158t4879 n6159 n4880 R=1.052e+01 
R6158t5557 n6159 n5558 R=3.818e+00 
R6158t327 n6159 n328 R=1.182e+01 
R6158t5708 n6159 n5709 R=5.102e+00 
R6159t590 n6160 n591 R=5.932e+00 
R6159t4397 n6160 n4398 R=2.632e+01 
R6160t205 n6161 n206 R=2.504e+00 
R6160t5304 n6161 n5305 R=3.356e+01 
R6160t4709 n6161 n4710 R=1.906e+01 
R6160t4036 n6161 n4037 R=4.877e+00 
R6160t829 n6161 n830 R=6.425e+00 
R6160t3777 n6161 n3778 R=8.894e+00 
R6161t552 n6162 n553 R=5.277e+00 
R6161t3225 n6162 n3226 R=1.286e+01 
R6161t3898 n6162 n3899 R=7.916e+00 
R6162t5314 n6163 n5315 R=5.095e+00 
R6162t4558 n6163 n4559 R=2.302e+00 
R6162t2388 n6163 n2389 R=3.002e+01 
R6163t784 n6164 n785 R=9.385e+00 
R6163t5028 n6164 n5029 R=5.577e+00 
R6163t1602 n6164 n1603 R=6.754e+00 
R6163t4728 n6164 n4729 R=7.723e+00 
R6164t151 n6165 n152 R=8.675e+00 
R6164t2323 n6165 n2324 R=1.341e+01 
R6165t1140 n6166 n1141 R=2.308e+00 
R6165t5177 n6166 n5178 R=4.581e+00 
R6165t5210 n6166 n5211 R=6.387e+01 
R6165t3633 n6166 n3634 R=4.351e+00 
R6165t2945 n6166 n2946 R=8.090e+00 
R6166t3417 n6167 n3418 R=6.633e+01 
R6166t4908 n6167 n4909 R=2.961e+01 
R6166t2403 n6167 n2404 R=1.401e+01 
R6166t1933 n6167 n1934 R=6.976e+00 
R6166t1834 n6167 n1835 R=4.902e+00 
R6167t4364 n6168 n4365 R=4.846e+00 
R6167t1527 n6168 n1528 R=2.804e+00 
R6168t1702 n6169 n1703 R=1.081e+02 
R6168t4131 n6169 n4132 R=1.323e+02 
R6168t1169 n6169 n1170 R=1.588e+02 
R6168t2698 n6169 n2699 R=5.548e+00 
R6168t5947 n6169 n5948 R=5.966e+01 
R6168t3522 n6169 n3523 R=9.698e+00 
R6168t5276 n6169 n5277 R=3.326e+00 
R6169t2682 n6170 n2683 R=3.755e+00 
R6169t2626 n6170 n2627 R=9.595e+00 
R6169t4972 n6170 n4973 R=2.398e+00 
R6169t2361 n6170 n2362 R=2.784e+01 
R6170t3380 n6171 n3381 R=1.331e+02 
R6170t1410 n6171 n1411 R=7.752e+00 
R6171t3556 n6172 n3557 R=1.998e+01 
R6171t4432 n6172 n4433 R=2.157e+01 
R6171t1404 n6172 n1405 R=1.124e+01 
R6171t4855 n6172 n4856 R=7.457e+00 
R6171t4384 n6172 n4385 R=2.771e+01 
R6171t5954 n6172 n5955 R=5.260e+00 
R6172t650 n6173 n651 R=3.402e+01 
R6172t5610 n6173 n5611 R=2.914e+01 
R6172t3704 n6173 n3705 R=1.898e+00 
R6172t721 n6173 n722 R=9.590e+00 
R6173t491 n6174 n492 R=3.876e+00 
R6173t3702 n6174 n3703 R=4.077e+00 
R6174t5613 n1 n5614 R=3.028e+02 
R6175t911 n6176 n912 R=6.965e+00 
R6175t30 n6176 n31 R=4.239e+00 
R6175t1796 n6176 n1797 R=2.632e+01 
R6176t3014 n6177 n3015 R=1.122e+01 
R6176t4485 n6177 n4486 R=1.564e+01 
R6176t413 n6177 n414 R=2.265e+00 
R6176t3691 n6177 n3692 R=7.045e+01 
R6176t827 n6177 n828 R=5.810e+00 
R6177t5486 n6178 n5487 R=6.345e+00 
R6177t4138 n6178 n4139 R=4.153e+00 
R6177t2418 n6178 n2419 R=4.166e+00 
R6177t4329 n6178 n4330 R=2.009e+01 
R6178t4802 n6179 n4803 R=3.700e+00 
R6178t689 n6179 n690 R=2.022e+01 
R6178t3285 n6179 n3286 R=1.277e+01 
R6178t1862 n6179 n1863 R=1.564e+01 
R6178t338 n6179 n339 R=3.971e+00 
R6178t1209 n6179 n1210 R=2.027e+01 
R6179t694 n6180 n695 R=1.960e+01 
R6179t525 n6180 n526 R=2.599e+00 
R6180t1596 n6181 n1597 R=5.679e+01 
R6180t6067 n6181 n6068 R=2.706e+01 
R6180t1028 n6181 n1029 R=7.867e+00 
R6181t1320 n6182 n1321 R=4.025e+00 
R6181t1898 n6182 n1899 R=8.941e+01 
R6181t5641 n6182 n5642 R=5.749e+01 
R6182t1790 n6183 n1791 R=4.085e+00 
R6182t5770 n6183 n5771 R=3.694e+01 
R6183t1897 n6184 n1898 R=2.391e+00 
R6183t5088 n6184 n5089 R=3.788e+00 
R6183t6155 n6184 n6156 R=5.963e+00 
R6183t3241 n6184 n3242 R=2.878e+01 
R6184t3426 n6185 n3427 R=3.439e+00 
R6184t2294 n6185 n2295 R=3.679e+00 
R6185t5359 n6186 n5360 R=3.124e+00 
R6185t3054 n6186 n3055 R=8.732e+00 
R6185t5702 n6186 n5703 R=2.866e+01 
R6185t1571 n6186 n1572 R=8.635e+00 
R6186t1854 n6187 n1855 R=4.528e+01 
R6186t2467 n6187 n2468 R=4.401e+00 
R6186t4303 n6187 n4304 R=5.600e+01 
R6186t2041 n6187 n2042 R=3.388e+00 
R6187t126 n6188 n127 R=2.875e+00 
R6187t2488 n6188 n2489 R=2.867e+01 
R6187t3695 n6188 n3696 R=1.038e+01 
R6187t494 n6188 n495 R=1.133e+01 
R6188t4262 n6189 n4263 R=9.064e+00 
R6188t4769 n6189 n4770 R=7.400e+00 
R6189t4144 n6190 n4145 R=3.206e+00 
R6189t6121 n6190 n6122 R=7.991e+00 
R6189t3581 n6190 n3582 R=4.514e+00 
R6190t663 n6191 n664 R=4.246e+00 
R6190t248 n6191 n249 R=4.096e+00 
R6190t984 n6191 n985 R=2.212e+01 
R6190t5540 n6191 n5541 R=3.019e+01 
R6191t2198 n6192 n1 R=4.737e+00 
R6192t4914 n6193 n4915 R=4.303e+00 
R6192t5635 n6193 n5636 R=5.596e+00 
R6192t1028 n6193 n1029 R=3.668e+01 
R6192t6052 n6193 n6053 R=4.727e+00 
R6192t5620 n6193 n5621 R=4.192e+01 
R6192t5734 n6193 n5735 R=1.404e+01 
R6193t2707 n6194 n2708 R=1.840e+00 
R6193t6130 n6194 n6131 R=2.530e+01 
R6193t131 n6194 n132 R=4.604e+00 
R6194t1868 n6195 n1869 R=5.448e+00 
R6195t3573 n6196 n3574 R=3.105e+00 
R6195t3993 n6196 n3994 R=9.958e+00 
R6195t2930 n6196 n2931 R=1.111e+01 
R6196t3421 n6197 n3422 R=1.052e+01 
R6196t5679 n6197 n5680 R=5.674e+00 
R6196t3659 n6197 n3660 R=8.106e+00 
R6196t4438 n6197 n4439 R=1.067e+01 
R6196t3585 n6197 n3586 R=2.495e+01 
R6196t2600 n6197 n2601 R=4.599e+00 
R6197t226 n6198 n227 R=2.008e+01 
R6197t3165 n6198 n3166 R=2.198e+01 
R6197t4154 n6198 n4155 R=5.104e+00 
R6197t4252 n6198 n4253 R=3.475e+01 
R6198t3450 n6199 n3451 R=7.401e+00 
R6198t5125 n6199 n5126 R=6.733e+00 
R6198t4858 n6199 n4859 R=2.581e+01 
R6198t5158 n6199 n5159 R=6.309e+00 
R6199t232 n6200 n233 R=3.088e+00 
R6199t1580 n6200 n1581 R=1.247e+01 
R6199t4320 n6200 n4321 R=3.647e+00 
R6199t2713 n6200 n2714 R=8.219e+00 
R6200t3568 n6201 n3569 R=2.803e+00 
R6200t3878 n6201 n3879 R=2.047e+00 
R6200t6017 n6201 n6018 R=5.857e+00 
R6200t2252 n6201 n2253 R=1.108e+02 
R6201t2626 n6202 n2627 R=2.283e+01 
R6201t2657 n6202 n2658 R=3.847e+01 
R6201t6179 n6202 n6180 R=4.903e+00 
R6202t3132 n6203 n3133 R=7.420e+00 
R6202t2963 n6203 n2964 R=1.546e+01 
R6202t5315 n6203 n5316 R=9.775e+00 
R6202t5349 n6203 n5350 R=7.073e+00 
R6203t2040 n6204 n2041 R=1.690e+01 
R6203t3948 n6204 n3949 R=6.972e+01 
R6203t2358 n6204 n2359 R=1.148e+01 
R6204t5219 n6205 n5220 R=6.353e+00 
R6204t5441 n6205 n5442 R=1.387e+01 
R6204t111 n6205 n112 R=1.230e+02 
R6205t886 n6206 n887 R=7.483e+00 
R6205t2820 n6206 n2821 R=1.231e+00 
R6205t3398 n6206 n3399 R=3.387e+00 
R6205t5831 n6206 n5832 R=3.266e+01 
R6205t2688 n6206 n2689 R=6.301e+01 
R6206t5219 n6207 n5220 R=3.497e+00 
R6206t4291 n6207 n4292 R=9.013e+00 
R6207t235 n6208 n236 R=5.810e+00 
R6207t2748 n6208 n2749 R=2.132e+01 
R6207t5837 n6208 n5838 R=8.960e+00 
R6208t5729 n6209 n5730 R=9.237e+00 
R6208t1642 n6209 n1643 R=3.886e+00 
R6208t3798 n6209 n3799 R=1.992e+01 
R6208t3597 n6209 n3598 R=5.514e+00 
R6208t2988 n6209 n2989 R=4.203e+01 
R6209t415 n6210 n416 R=4.850e+00 
R6209t1908 n6210 n1909 R=8.435e+00 
R6209t3845 n6210 n3846 R=2.619e+00 
R6210t5323 n6211 n5324 R=4.289e+00 
R6210t3807 n6211 n3808 R=1.675e+01 
R6211t208 n6212 n209 R=5.555e+00 
R6211t1460 n6212 n1461 R=4.628e+00 
R6211t2773 n6212 n2774 R=1.464e+01 
R6212t1685 n6213 n1686 R=8.689e+00 
R6212t4046 n6213 n4047 R=4.521e+00 
R6212t1988 n6213 n1989 R=9.587e+00 
R6212t5016 n6213 n5017 R=9.733e+00 
R6213t63 n6214 n64 R=7.287e+01 
R6213t3487 n6214 n3488 R=5.022e+00 
R6213t2690 n6214 n2691 R=7.492e+00 
R6213t5182 n6214 n5183 R=1.771e+01 
R6213t5710 n6214 n5711 R=1.061e+01 
R6213t303 n6214 n304 R=6.587e+00 
R6213t13 n6214 n14 R=1.248e+01 
R6213t758 n6214 n759 R=4.930e+01 
R6214t1793 n6215 n1794 R=7.222e+00 
R6214t4719 n6215 n4720 R=6.407e+00 
R6215t2546 n6216 n2547 R=4.851e+00 
R6215t3090 n6216 n3091 R=8.837e+00 
R6215t2360 n6216 n2361 R=6.467e+00 
R6216t1540 n6217 n1541 R=3.154e+01 
R6216t3918 n6217 n3919 R=2.832e+00 
R6216t5035 n6217 n5036 R=1.126e+01 
R6216t450 n6217 n451 R=4.105e+00 
R6217t92 n6218 n93 R=6.407e+01 
R6217t3984 n6218 n3985 R=2.078e+01 
R6217t3783 n6218 n3784 R=2.306e+00 
R6218t265 n6219 n266 R=5.493e+00 
R6218t5145 n6219 n5146 R=5.386e+00 
R6218t4679 n6219 n4680 R=2.186e+02 
R6219t3238 n6220 n3239 R=2.608e+00 
R6219t286 n6220 n287 R=1.728e+01 
R6219t2574 n6220 n2575 R=4.867e+00 
R6219t2230 n6220 n2231 R=2.188e+01 
R6220t3264 n6221 n3265 R=1.119e+01 
R6220t4888 n6221 n4889 R=1.060e+01 
R6220t4237 n6221 n4238 R=7.359e+00 
R6220t957 n6221 n958 R=5.453e+00 
R6220t4833 n6221 n4834 R=7.481e+01 
R6220t1268 n6221 n1269 R=7.687e+00 
R6220t4522 n6221 n4523 R=1.082e+01 
R6221t1733 n6222 n1734 R=4.644e+02 
R6221t4835 n6222 n4836 R=3.503e+01 
R6222t2193 n6223 n2194 R=8.448e+01 
R6222t1873 n6223 n1874 R=5.614e+00 
R6223t1963 n6224 n1964 R=1.019e+02 
R6223t646 n6224 n647 R=1.460e+01 
R6223t437 n6224 n438 R=4.231e+00 
R6223t948 n6224 n949 R=1.083e+01 
R6224t873 n6225 n874 R=2.745e+00 
R6224t1989 n6225 n1990 R=5.404e+00 
R6224t2432 n6225 n2433 R=1.940e+01 
R6225t1336 n6226 n1337 R=1.547e+00 
R6225t3444 n6226 n3445 R=1.856e+01 
R6225t4806 n6226 n4807 R=1.064e+01 
R6225t5603 n6226 n5604 R=3.037e+02 
R6225t5974 n6226 n5975 R=6.086e+00 
R6226t1723 n6227 n1724 R=5.728e+00 
R6226t2692 n6227 n2693 R=7.512e+00 
R6226t2391 n6227 n2392 R=7.789e+01 
R6227t1155 n6228 n1156 R=4.748e+00 
R6227t4569 n6228 n4570 R=6.813e+00 
R6227t2962 n6228 n2963 R=9.780e+00 
R6227t2232 n6228 n2233 R=1.882e+01 
R6228t2618 n6229 n2619 R=4.538e+02 
R6228t5292 n6229 n5293 R=5.010e+00 
R6229t4114 n6230 n4115 R=4.659e+01 
R6229t1610 n6230 n1611 R=8.766e+00 
R6229t1591 n6230 n1592 R=7.755e+01 
R6229t4499 n6230 n4500 R=7.425e+00 
R6229t3227 n6230 n3228 R=2.307e+01 
R6230t1100 n6231 n1101 R=5.831e+00 
R6230t1938 n6231 n1939 R=3.262e+00 
R6230t914 n6231 n915 R=7.248e+00 
R6231t4074 n6232 n4075 R=1.356e+01 
R6231t5708 n6232 n5709 R=5.430e+00 
R6231t3091 n6232 n3092 R=6.093e+01 
R6232t1063 n6233 n1064 R=4.907e+00 
R6232t4356 n6233 n4357 R=6.339e+00 
R6233t590 n6234 n591 R=3.241e+00 
R6233t4822 n6234 n4823 R=2.060e+01 
R6233t5365 n6234 n5366 R=5.231e+00 
R6233t4397 n6234 n4398 R=3.965e+00 
R6233t6159 n6234 n6160 R=1.693e+01 
R6234t3587 n6235 n3588 R=5.216e+00 
R6234t3130 n6235 n3131 R=2.180e+01 
R6234t356 n6235 n357 R=1.310e+01 
R6235t4050 n6236 n4051 R=4.900e+00 
R6235t4667 n6236 n4668 R=2.750e+01 
R6236t4882 n6237 n4883 R=1.303e+01 
R6236t862 n6237 n863 R=3.770e+00 
R6237t1286 n6238 n1287 R=2.397e+00 
R6237t2128 n6238 n2129 R=4.628e+01 
R6237t2119 n6238 n2120 R=4.514e+01 
R6237t4769 n6238 n4770 R=5.549e+00 
R6237t6188 n6238 n6189 R=4.871e+00 
R6238t460 n6239 n461 R=5.718e+01 
R6238t3865 n6239 n3866 R=1.148e+01 
R6238t1330 n6239 n1331 R=5.938e+00 
R6238t1279 n6239 n1280 R=1.417e+01 
R6238t2500 n6239 n2501 R=1.264e+01 
R6238t3209 n6239 n3210 R=2.603e+00 
R6239t138 n6240 n139 R=8.086e+00 
R6239t3498 n6240 n3499 R=4.209e+00 
R6239t929 n6240 n930 R=1.095e+01 
R6239t1986 n6240 n1987 R=8.185e+00 
R6239t4307 n6240 n4308 R=7.195e+00 
R6240t4898 n6241 n4899 R=5.607e+00 
R6240t84 n6241 n85 R=4.138e+00 
R6240t5680 n6241 n5681 R=1.118e+02 
R6241t5063 n6242 n5064 R=1.117e+01 
R6241t3089 n6242 n3090 R=1.493e+01 
R6241t1495 n6242 n1496 R=4.171e+01 
R6241t4072 n6242 n4073 R=2.425e+01 
R6241t1695 n6242 n1696 R=7.677e+01 
R6241t283 n6242 n284 R=6.137e+00 
R6242t310 n6243 n311 R=9.042e+00 
R6242t5566 n6243 n5567 R=2.683e+00 
R6242t1472 n6243 n1473 R=1.510e+01 
R6242t1615 n6243 n1616 R=2.872e+01 
R6242t3353 n6243 n3354 R=1.130e+01 
R6242t4676 n6243 n4677 R=1.796e+03 
R6243t829 n6244 n830 R=9.417e+00 
R6243t4036 n6244 n4037 R=9.131e+00 
R6243t6039 n6244 n6040 R=4.343e+00 
R6243t3024 n6244 n3025 R=3.894e+00 
R6244t1243 n6245 n1244 R=1.049e+01 
R6244t5385 n6245 n5386 R=5.090e+00 
R6244t3310 n6245 n3311 R=3.413e+02 
R6244t3827 n6245 n3828 R=9.830e+00 
R6244t748 n6245 n749 R=1.194e+01 
R6245t3343 n6246 n3344 R=2.791e+01 
R6245t4030 n6246 n4031 R=3.275e+00 
R6245t1244 n6246 n1245 R=4.599e+00 
R6245t634 n6246 n635 R=5.222e+00 
R6246t282 n6247 n283 R=3.069e+00 
R6246t2156 n6247 n2157 R=7.888e+00 
R6246t297 n6247 n298 R=2.651e+00 
R6246t255 n6247 n256 R=3.372e+01 
R6246t3972 n6247 n3973 R=1.400e+01 
R6247t2949 n6248 n2950 R=1.301e+01 
R6247t4344 n6248 n4345 R=1.830e+00 
R6247t5337 n6248 n5338 R=6.788e+00 
R6248t3979 n6249 n3980 R=2.509e+00 
R6248t1020 n6249 n1021 R=3.421e+01 
R6248t5640 n6249 n5641 R=6.771e+01 
R6249t5779 n6250 n5780 R=4.223e+00 
R6249t981 n6250 n982 R=2.549e+00 
R6249t816 n6250 n817 R=6.603e+00 
R6250t4962 n6251 n4963 R=1.145e+01 
R6250t5188 n6251 n5189 R=1.790e+01 
R6250t3989 n6251 n3990 R=1.323e+01 
R6250t1633 n6251 n1634 R=2.400e+01 
R6250t3146 n6251 n3147 R=2.636e+01 
R6251t689 n6252 n690 R=5.392e+00 
R6251t3285 n6252 n3286 R=2.395e+01 
R6251t4813 n6252 n4814 R=1.874e+01 
R6251t708 n6252 n709 R=1.287e+01 
R6251t4392 n6252 n4393 R=5.905e+00 
R6251t4805 n6252 n4806 R=4.872e+02 
R6251t3491 n6252 n3492 R=2.814e+01 
R6252t1559 n6253 n1560 R=6.143e+00 
R6252t5283 n6253 n5284 R=2.227e+01 
R6252t3107 n6253 n3108 R=2.578e+00 
R6252t3779 n6253 n3780 R=4.816e+01 
R6252t232 n6253 n233 R=3.119e+01 
R6252t4723 n6253 n4724 R=7.125e+00 
R6252t5410 n6253 n5411 R=1.010e+01 
R6252t1965 n6253 n1966 R=8.514e+00 
R6253t731 n6254 n732 R=2.500e+01 
R6253t840 n6254 n841 R=4.169e+00 
R6253t1164 n6254 n1165 R=2.261e+01 
R6253t412 n6254 n413 R=4.636e+00 
R6254t3238 n6255 n3239 R=5.670e+01 
R6254t6219 n6255 n6220 R=5.230e+00 
R6254t1553 n6255 n1554 R=1.651e+01 
R6254t5575 n6255 n5576 R=2.664e+01 
R6254t4826 n6255 n4827 R=5.083e+00 
R6254t2230 n6255 n2231 R=2.978e+01 
R6255t5921 n6256 n5922 R=8.145e+00 
R6255t4210 n6256 n4211 R=7.803e+00 
R6255t2280 n6256 n2281 R=4.065e+00 
R6256t4635 n6257 n4636 R=2.599e+01 
R6256t1165 n6257 n1166 R=4.236e+00 
R6256t4937 n6257 n4938 R=3.860e+01 
R6256t3385 n6257 n3386 R=2.046e+00 
R6257t2043 n6258 n2044 R=5.459e+00 
R6257t902 n6258 n903 R=3.681e+00 
R6257t4383 n6258 n4384 R=3.973e+01 
R6257t4776 n6258 n4777 R=1.759e+01 
R6257t1757 n6258 n1758 R=3.371e+00 
R6258t2187 n6259 n2188 R=8.029e+00 
R6258t2474 n6259 n2475 R=6.296e+00 
R6258t5322 n6259 n5323 R=6.708e+01 
R6258t5273 n6259 n5274 R=4.838e+00 
R6258t6153 n6259 n6154 R=4.315e+00 
R6259t325 n6260 n326 R=9.137e+00 
R6259t4594 n6260 n4595 R=8.020e+01 
R6259t5961 n6260 n5962 R=1.163e+01 
R6260t122 n6261 n123 R=4.960e+00 
R6260t5979 n6261 n5980 R=5.945e+00 
R6260t3679 n6261 n3680 R=3.668e+00 
R6260t5011 n6261 n5012 R=3.032e+02 
R6261t1405 n6262 n1406 R=1.120e+01 
R6261t59 n6262 n60 R=6.418e+00 
R6261t2452 n6262 n2453 R=3.254e+00 
R6262t870 n6263 n871 R=7.068e+01 
R6262t1879 n6263 n1880 R=1.043e+01 
R6263t1314 n6264 n1315 R=1.573e+01 
R6263t1529 n6264 n1530 R=6.449e+00 
R6263t3784 n6264 n3785 R=1.641e+01 
R6263t981 n6264 n982 R=7.085e+00 
R6264t1866 n6265 n1867 R=6.701e+00 
R6264t4281 n6265 n4282 R=7.643e+01 
R6264t5985 n6265 n5986 R=3.319e+01 
R6265t5926 n6266 n5927 R=8.104e+00 
R6265t5386 n6266 n5387 R=4.473e+00 
R6265t1261 n6266 n1262 R=2.290e+01 
R6266t1856 n6267 n1857 R=2.504e+00 
R6266t2759 n6267 n2760 R=6.009e+01 
R6266t1647 n6267 n1648 R=1.497e+01 
R6268t5140 n6269 n5141 R=3.385e+00 
R6269t1455 n6270 n1456 R=1.202e+01 
R6269t1856 n6270 n1857 R=6.934e+00 
R6269t1647 n6270 n1648 R=1.308e+01 
R6270t407 n6271 n408 R=1.221e+01 
R6270t5272 n6271 n5273 R=3.787e+00 
R6270t780 n6271 n781 R=8.217e+00 
R6270t4311 n6271 n4312 R=6.857e+00 
R6271t1052 n6272 n1053 R=3.057e+00 
R6271t2487 n6272 n2488 R=1.667e+01 
R6271t1698 n6272 n1699 R=5.005e+00 
R6272t3246 n6273 n3247 R=4.891e+00 
R6272t3526 n6273 n3527 R=4.988e+00 
R6272t5069 n6273 n5070 R=4.670e+00 
R6272t4153 n6273 n4154 R=6.760e+01 
R6273t2154 n6274 n2155 R=8.226e+00 
R6273t3536 n6274 n3537 R=2.734e+01 
R6274t1085 n6275 n1086 R=1.274e+01 
R6274t2079 n6275 n2080 R=1.386e+01 
R6274t700 n6275 n701 R=2.927e+00 
R6274t5002 n6275 n5003 R=2.380e+01 
R6274t3950 n6275 n3951 R=2.919e+00 
R6274t612 n6275 n613 R=9.109e+01 
R6275t2729 n6276 n2730 R=3.716e+01 
R6275t5945 n6276 n5946 R=5.199e+00 
R6275t1605 n6276 n1606 R=1.169e+01 
R6275t1894 n6276 n1895 R=3.790e+01 
R6276t383 n6277 n384 R=2.278e+01 
R6276t1474 n6277 n1475 R=3.798e+00 
R6277t3260 n6278 n3261 R=5.139e+01 
R6277t47 n6278 n48 R=2.538e+01 
R6277t6025 n6278 n6026 R=6.102e+00 
R6277t1673 n6278 n1674 R=5.620e+00 
R6278t4106 n6279 n4107 R=7.034e+00 
R6278t5191 n6279 n5192 R=7.782e+00 
R6278t3910 n6279 n3911 R=1.150e+01 
R6278t2273 n6279 n2274 R=7.423e+00 
R6278t5242 n6279 n5243 R=3.002e+02 
R6278t93 n6279 n94 R=1.381e+01 
R6278t3462 n6279 n3463 R=5.189e+00 
R6279t1482 n6280 n1483 R=2.504e+01 
R6279t400 n6280 n401 R=1.705e+01 
R6279t887 n6280 n888 R=6.088e+00 
R6279t3328 n6280 n3329 R=6.389e+00 
R6280t1229 n6281 n1230 R=7.539e+00 
R6280t5781 n6281 n5782 R=4.135e+00 
R6280t925 n6281 n926 R=4.625e+00 
R6281t291 n6282 n292 R=3.360e+00 
R6281t2569 n6282 n2570 R=4.368e+00 
R6281t4168 n6282 n4169 R=2.143e+02 
R6281t5866 n6282 n5867 R=3.321e+01 
R6282t2514 n6283 n2515 R=4.124e+01 
R6282t1277 n6283 n1278 R=4.799e+00 
R6282t5543 n6283 n5544 R=4.091e+00 
R6283t1750 n6284 n1751 R=6.309e+00 
R6283t5229 n6284 n5230 R=5.519e+00 
R6283t4811 n6284 n4812 R=1.496e+01 
R6283t5872 n6284 n5873 R=5.598e+00 
R6283t4194 n6284 n4195 R=1.010e+01 
R6283t3233 n6284 n3234 R=4.860e+01 
R6284t5195 n6285 n5196 R=5.849e+01 
R6284t1115 n6285 n1116 R=6.161e+00 
R6284t2996 n6285 n2997 R=3.590e+00 
R6284t46 n6285 n47 R=1.002e+01 
R6285t3772 n6286 n3773 R=4.079e+00 
R6285t4433 n6286 n4434 R=2.945e+01 
R6285t2342 n6286 n2343 R=4.197e+00 
R6285t3438 n6286 n3439 R=2.596e+01 
R6285t2731 n6286 n2732 R=2.745e+00 
R6286t1514 n6287 n1515 R=4.914e+02 
R6286t2581 n6287 n2582 R=3.432e+00 
R6286t243 n6287 n244 R=1.087e+01 
R6286t2902 n6287 n2903 R=9.832e+00 
R6286t4219 n6287 n4220 R=3.971e+00 
R6287t2704 n6288 n2705 R=3.030e+00 
R6287t915 n6288 n916 R=6.661e+00 
R6287t5447 n6288 n5448 R=2.816e+00 
R6287t4950 n6288 n4951 R=2.861e+01 
R6287t2885 n6288 n2886 R=1.185e+01 
R6288t2733 n6289 n2734 R=2.390e+00 
R6288t5136 n6289 n5137 R=2.084e+01 
R6288t38 n6289 n39 R=7.438e+00 
R6289t1726 n6290 n1727 R=1.129e+01 
R6289t4364 n6290 n4365 R=1.760e+01 
R6290t4207 n6291 n4208 R=3.970e+00 
R6290t4716 n6291 n4717 R=5.994e+00 
R6290t4230 n6291 n4231 R=1.028e+01 
R6291t5229 n6292 n5230 R=1.884e+02 
R6291t4605 n6292 n4606 R=2.050e+01 
R6291t2404 n6292 n2405 R=2.885e+01 
R6291t423 n6292 n424 R=1.300e+01 
R6291t4811 n6292 n4812 R=3.098e+00 
R6292t4070 n6293 n4071 R=5.862e+00 
R6292t4284 n6293 n4285 R=1.551e+01 
R6292t1001 n6293 n1002 R=3.340e+00 
R6292t3973 n6293 n3974 R=5.853e+01 
R6292t1477 n6293 n1478 R=6.754e+00 
R6293t1944 n6294 n1945 R=1.235e+01 
R6293t4454 n6294 n4455 R=3.709e+00 
R6293t2897 n6294 n2898 R=7.677e+00 
R6293t2894 n6294 n2895 R=4.198e+01 
R6294t331 n6295 n332 R=5.893e+00 
R6294t4363 n6295 n4364 R=1.688e+01 
R6294t1233 n6295 n1234 R=3.703e+00 
R6295t125 n6296 n126 R=4.690e+01 
R6295t4891 n6296 n4892 R=4.458e+00 
R6295t3876 n6296 n3877 R=1.082e+01 
R6295t2688 n6296 n2689 R=5.488e+00 
R6296t3761 n6297 n3762 R=1.895e+01 
R6296t3815 n6297 n3816 R=7.132e+00 
R6296t5342 n6297 n5343 R=5.290e+00 
R6296t436 n6297 n437 R=1.247e+01 
R6296t4808 n6297 n4809 R=1.177e+01 
R6297t950 n6298 n951 R=1.319e+02 
R6297t1831 n6298 n1832 R=1.088e+03 
R6297t5948 n6298 n5949 R=5.511e+01 
R6297t4634 n6298 n4635 R=2.794e+00 
R6297t4175 n6298 n4176 R=2.285e+01 
R6297t1417 n6298 n1418 R=2.016e+01 
R6298t2665 n6299 n2666 R=8.651e+00 
R6298t5279 n6299 n5280 R=3.828e+00 
R6298t4713 n6299 n4714 R=3.497e+00 
R6299t4610 n6300 n4611 R=4.824e+00 
R6299t4549 n6300 n4550 R=1.939e+00 
R6300t1216 n6301 n1217 R=1.839e+01 
R6300t4994 n6301 n4995 R=6.100e+00 
R6300t3903 n6301 n3904 R=3.467e+00 
R6300t955 n6301 n956 R=3.473e+02 
R6300t462 n6301 n463 R=8.024e+00 
R6302t1079 n6303 n1080 R=2.388e+01 
R6302t3031 n6303 n3032 R=6.188e+00 
R6302t5806 n6303 n5807 R=2.665e+01 
R6302t4528 n6303 n4529 R=1.143e+01 
R6303t737 n6304 n738 R=4.449e+00 
R6303t969 n6304 n970 R=2.356e+01 
R6303t3220 n6304 n3221 R=5.756e+00 
R6303t404 n6304 n405 R=2.294e+01 
R6303t4936 n6304 n4937 R=4.923e+01 
R6303t771 n6304 n772 R=6.597e+00 
R6304t3234 n6305 n3235 R=2.004e+00 
R6304t2575 n6305 n2576 R=1.185e+01 
R6304t4976 n6305 n4977 R=2.029e+01 
R6305t2415 n6306 n2416 R=4.889e+00 
R6306t2060 n6307 n2061 R=3.605e+00 
R6306t5971 n6307 n5972 R=9.166e+00 
R6306t4966 n6307 n4967 R=5.225e+00 
R6306t5228 n6307 n5229 R=7.058e+00 
R6307t5092 n6308 n5093 R=4.322e+00 
R6307t1034 n6308 n1035 R=3.319e+00 
R6307t5921 n6308 n5922 R=5.905e+00 
R6308t1059 n6309 n1060 R=3.927e+00 
R6308t4738 n6309 n4739 R=9.396e+00 
R6308t601 n6309 n602 R=6.011e+00 
R6308t496 n6309 n497 R=9.973e+00 
R6309t4974 n6310 n4975 R=5.838e+00 
R6310t5197 n6311 n5198 R=2.231e+00 
R6310t4635 n6311 n4636 R=5.924e+00 
R6311t5319 n6312 n5320 R=1.583e+02 
R6311t3719 n6312 n3720 R=3.868e+00 
R6311t3648 n6312 n3649 R=3.005e+00 
R6311t1886 n6312 n1887 R=2.056e+00 
R6311t4271 n6312 n4272 R=4.177e+01 
R6312t5367 n6313 n5368 R=5.979e+00 
R6312t5671 n6313 n5672 R=8.384e+00 
R6312t246 n6313 n247 R=1.039e+01 
R6312t3524 n6313 n3525 R=7.208e+00 
R6312t4814 n6313 n4815 R=7.246e+01 
R6312t5905 n6313 n5906 R=4.131e+00 
R6313t4945 n6314 n4946 R=2.058e+02 
R6313t258 n6314 n259 R=1.385e+01 
R6313t5336 n6314 n5337 R=4.287e+00 
R6313t655 n6314 n656 R=1.556e+01 
R6314t113 n6315 n114 R=4.227e+01 
R6314t5097 n6315 n5098 R=1.099e+01 
R6314t2621 n6315 n2622 R=4.684e+00 
R6314t5224 n6315 n5225 R=1.339e+01 
R6314t507 n6315 n508 R=5.732e+00 
R6314t3540 n6315 n3541 R=2.215e+01 
R6314t2108 n6315 n2109 R=6.864e+00 
R6315t4198 n6316 n4199 R=4.304e+01 
R6315t5504 n6316 n5505 R=5.033e+00 
R6315t214 n6316 n215 R=3.178e+00 
R6315t3460 n6316 n3461 R=4.363e+00 
R6316t1805 n6317 n1806 R=1.469e+01 
R6316t5843 n6317 n5844 R=4.062e+00 
R6317t235 n6318 n236 R=2.777e+01 
R6317t2104 n6318 n2105 R=2.388e+00 
R6317t4985 n6318 n4986 R=3.533e+01 
R6318t2965 n6319 n2966 R=7.596e+00 
R6318t4149 n6319 n4150 R=7.059e+00 
R6318t5826 n6319 n5827 R=2.584e+01 
R6318t2380 n6319 n2381 R=8.864e+01 
R6318t1945 n6319 n1946 R=4.340e+00 
R6318t4122 n6319 n4123 R=4.254e+01 
R6318t2158 n6319 n2159 R=1.408e+02 
R6319t2446 n6320 n1 R=6.390e+01 
R6319t1625 n6320 n1626 R=7.315e+00 
R6319t2614 n6320 n2615 R=1.271e+01 
R6319t1 n6320 n2 R=9.671e+00 
R6320t4027 n6321 n4028 R=2.893e+00 
R6320t4163 n6321 n4164 R=3.867e+00 
R6321t1116 n6322 n1117 R=2.275e+01 
R6321t4543 n6322 n4544 R=1.234e+01 
R6321t2565 n6322 n2566 R=5.153e+00 
R6321t4607 n6322 n4608 R=3.725e+01 
R6321t5844 n6322 n5845 R=3.922e+00 
R6321t524 n6322 n525 R=1.995e+01 
R6322t1088 n6323 n1089 R=4.152e+00 
R6322t2082 n6323 n2083 R=6.540e+00 
R6322t1409 n6323 n1410 R=7.276e+00 
R6323t430 n6324 n431 R=5.317e+01 
R6323t1546 n6324 n1547 R=4.426e+00 
R6323t147 n6324 n148 R=5.432e+00 
R6323t604 n6324 n605 R=3.511e+01 
R6324t4985 n6325 n4986 R=1.029e+01 
R6324t6078 n6325 n6079 R=4.358e+00 
R6324t3525 n6325 n3526 R=5.220e+00 
R6324t3163 n6325 n3164 R=1.362e+02 
R6325t521 n6326 n522 R=1.515e+01 
R6325t4594 n6326 n4595 R=8.169e+00 
R6325t6259 n6326 n6260 R=9.107e+00 
R6325t947 n6326 n948 R=2.861e+00 
R6326t3790 n6327 n3791 R=1.536e+01 
R6326t5789 n6327 n5790 R=5.008e+00 
R6326t1489 n6327 n1490 R=6.924e+00 
R6327t1731 n6328 n1732 R=6.765e+00 
R6327t5780 n6328 n5781 R=6.029e+00 
R6327t5907 n6328 n5908 R=1.540e+01 
R6327t5608 n6328 n5609 R=3.484e+01 
R6328t2512 n6329 n2513 R=4.308e+00 
R6329t701 n6330 n702 R=3.876e+01 
R6329t2739 n6330 n2740 R=3.691e+00 
R6329t1454 n6330 n1455 R=7.114e+00 
R6329t293 n6330 n294 R=5.035e+00 
R6330t579 n6331 n580 R=4.887e+00 
R6330t4831 n6331 n4832 R=3.734e+00 
R6331t424 n6332 n425 R=3.149e+01 
R6331t1752 n6332 n1753 R=2.671e+00 
R6331t2978 n6332 n2979 R=3.504e+00 
R6331t4735 n6332 n4736 R=1.407e+01 
R6332t1782 n6333 n1783 R=4.001e+00 
R6332t2635 n6333 n2636 R=3.579e+00 
R6332t3054 n6333 n3055 R=5.055e+00 
R6332t3405 n6333 n3406 R=1.800e+01 
R6333t2772 n6334 n2773 R=4.128e+00 
R6333t4243 n6334 n4244 R=7.768e+00 
R6334t1216 n6335 n1217 R=6.085e+00 
R6334t4275 n6335 n4276 R=6.811e+00 
R6334t5123 n6335 n5124 R=2.006e+01 
R6334t1357 n6335 n1358 R=4.925e+00 
R6334t5252 n6335 n5253 R=1.060e+01 
R6334t543 n6335 n544 R=2.881e+01 
R6334t3584 n6335 n3585 R=8.008e+00 
R6335t4309 n6336 n4310 R=4.482e+00 
R6335t4056 n6336 n4057 R=2.535e+00 
R6335t5054 n6336 n5055 R=5.222e+01 
R6335t25 n6336 n26 R=1.240e+01 
R6336t6126 n6337 n6127 R=6.128e+00 
R6337t206 n6338 n207 R=5.914e+00 
R6337t1022 n6338 n1023 R=3.214e+00 
R6337t5753 n6338 n5754 R=1.385e+02 
R6337t5733 n6338 n5734 R=9.577e+01 
R6337t842 n6338 n843 R=1.717e+01 
R6338t896 n6339 n897 R=3.172e+00 
R6338t2750 n6339 n2751 R=6.500e+01 
R6338t3865 n6339 n3866 R=3.518e+01 
R6338t6322 n6339 n6323 R=1.200e+01 
R6338t2082 n6339 n2083 R=2.645e+00 
R6339t2510 n6340 n2511 R=7.558e+00 
R6339t6279 n6340 n6280 R=4.071e+00 
R6339t1482 n6340 n1483 R=2.656e+01 
R6339t56 n6340 n57 R=2.058e+01 
R6340t156 n6341 n157 R=6.859e+00 
R6340t5487 n6341 n5488 R=9.460e+00 
R6341t2606 n6342 n2607 R=1.103e+01 
R6341t4247 n6342 n4248 R=2.801e+00 
R6341t2882 n6342 n2883 R=3.317e+00 
R6342t1670 n1 n1671 R=3.090e+01 
R6342t2506 n1 n2507 R=1.840e+01 
R6343t5035 n6344 n5036 R=2.349e+00 
R6343t5584 n6344 n5585 R=3.892e+00 
R6343t1356 n6344 n1357 R=9.030e+00 
R6344t4446 n6345 n4447 R=1.297e+00 
R6344t776 n6345 n777 R=1.600e+00 
R6344t2780 n6345 n2781 R=5.109e+02 
R6345t5396 n6346 n5397 R=4.979e+01 
R6345t210 n6346 n211 R=2.380e+00 
R6346t6320 n6347 n6321 R=8.001e+00 
R6346t4163 n6347 n4164 R=1.838e+01 
R6346t3589 n6347 n3590 R=3.861e+00 
R6346t1901 n6347 n1902 R=1.435e+01 
R6346t5180 n6347 n5181 R=4.315e+00 
R6347t3351 n6348 n3352 R=2.879e+00 
R6347t4488 n6348 n4489 R=2.095e+01 
R6347t1264 n6348 n1265 R=8.632e+00 
R6347t6085 n6348 n6086 R=1.874e+00 
R6348t6055 n6349 n6056 R=1.102e+01 
R6348t4612 n6349 n4613 R=1.640e+01 
R6348t3657 n6349 n3658 R=4.814e+00 
R6348t1887 n6349 n1888 R=9.716e+01 
R6348t1489 n6349 n1490 R=7.888e+00 
R6349t3568 n6350 n3569 R=7.792e+00 
R6349t5910 n6350 n5911 R=2.045e+00 
R6350t5979 n6351 n5980 R=9.101e+00 
R6350t3121 n6351 n3122 R=1.045e+01 
R6351t4849 n6352 n4850 R=3.423e+00 
R6351t5310 n6352 n5311 R=9.280e+00 
R6351t4056 n6352 n4057 R=1.201e+01 
R6351t6335 n6352 n6336 R=7.174e+00 
R6351t4309 n6352 n4310 R=1.995e+01 
R6351t2115 n6352 n2116 R=7.233e+01 
R6352t646 n6353 n647 R=1.130e+01 
R6352t1251 n6353 n1252 R=1.717e+01 
R6352t335 n6353 n336 R=1.892e+01 
R6353t4252 n6354 n4253 R=3.672e+00 
R6353t3778 n6354 n3779 R=9.876e+00 
R6354t3166 n6355 n3167 R=4.585e+00 
R6355t2277 n6356 n2278 R=1.104e+01 
R6355t403 n6356 n404 R=3.623e+00 
R6355t2112 n6356 n2113 R=1.977e+01 
R6356t1934 n6357 n1935 R=1.086e+01 
R6356t2753 n6357 n2754 R=6.218e+00 
R6357t5961 n6358 n5962 R=9.111e+00 
R6357t2396 n6358 n2397 R=5.211e+02 
R6357t1512 n6358 n1513 R=1.732e+02 
R6357t3261 n6358 n3262 R=3.941e+00 
R6358t2125 n6359 n2126 R=5.968e+00 
R6358t670 n6359 n671 R=5.061e+00 
R6358t2355 n6359 n2356 R=6.359e+00 
R6359t5439 n6360 n5440 R=3.618e+00 
R6359t1973 n6360 n1974 R=5.383e+01 
R6360t2312 n6361 n2313 R=6.478e+00 
R6360t3471 n6361 n3472 R=3.552e+00 
R6360t6131 n6361 n6132 R=2.472e+01 
R6360t2789 n6361 n2790 R=7.105e+00 
R6360t34 n6361 n35 R=6.248e+00 
R6361t1619 n6362 n1620 R=2.161e+00 
R6361t4109 n6362 n4110 R=4.282e+00 
R6361t4429 n6362 n4430 R=5.078e+00 
R6362t160 n6363 n161 R=6.539e+01 
R6362t4524 n6363 n4525 R=4.058e+01 
R6363t5207 n6364 n5208 R=5.204e+01 
R6363t554 n6364 n555 R=1.140e+01 
R6363t4495 n6364 n4496 R=7.537e+00 
R6364t470 n6365 n471 R=1.599e+01 
R6364t5316 n6365 n5317 R=5.048e+00 
R6364t1541 n6365 n1542 R=1.611e+01 
R6364t179 n6365 n180 R=9.812e+00 
R6364t5038 n6365 n5039 R=4.824e+00 
R6365t1447 n6366 n1448 R=7.168e+01 
R6365t795 n6366 n796 R=2.255e+00 
R6365t4122 n6366 n4123 R=1.295e+01 
R6365t1521 n6366 n1522 R=1.336e+01 
R6366t1722 n6367 n1723 R=3.297e+00 
R6366t2011 n6367 n2012 R=7.539e+00 
R6367t282 n6368 n283 R=5.941e+00 
R6367t4270 n6368 n4271 R=1.038e+01 
R6367t6246 n6368 n6247 R=1.908e+02 
R6367t5003 n6368 n5004 R=3.832e+00 
R6367t4580 n6368 n4581 R=1.093e+01 
R6367t4903 n6368 n4904 R=6.138e+00 
R6368t5824 n6369 n5825 R=8.450e+00 
R6368t2395 n6369 n1 R=3.416e+00 
R6368t5455 n6369 n5456 R=3.766e+00 
R6368t4425 n6369 n4426 R=1.208e+01 
R6369t427 n6370 n428 R=2.310e+00 
R6369t2072 n6370 n2073 R=2.836e+02 
R6370t2668 n6371 n2669 R=4.252e+01 
R6370t6363 n6371 n6364 R=1.388e+01 
R6370t5207 n6371 n5208 R=1.399e+02 
R6370t4025 n6371 n4026 R=4.511e+00 
R6370t4920 n6371 n4921 R=5.772e+00 
R6371t414 n6372 n415 R=6.979e+00 
R6371t4831 n6372 n4832 R=1.693e+01 
R6371t5122 n6372 n5123 R=3.756e+00 
R6371t6330 n6372 n6331 R=4.931e+00 
R6372t2497 n6373 n2498 R=3.658e+01 
R6372t2827 n6373 n2828 R=1.604e+00 
R6372t1087 n6373 n1088 R=6.145e+01 
R6372t5997 n6373 n5998 R=4.185e+00 
R6372t2838 n6373 n2839 R=3.081e+00 
R6373t458 n6374 n459 R=8.119e+00 
R6373t599 n6374 n600 R=7.235e+00 
R6373t1927 n6374 n1928 R=4.324e+01 
R6373t2005 n6374 n2006 R=4.119e+01 
R6373t3407 n6374 n3408 R=1.221e+01 
R6374t3977 n6375 n3978 R=4.791e+01 
R6374t5786 n6375 n5787 R=3.903e+01 
R6374t1159 n6375 n1160 R=6.172e+01 
R6374t4641 n6375 n4642 R=5.797e+01 
R6375t4177 n6376 n4178 R=2.862e+01 
R6375t6023 n6376 n6024 R=6.606e+00 
R6375t3849 n6376 n3850 R=2.816e+00 
R6375t5720 n6376 n5721 R=4.915e+02 
R6376t2497 n6377 n2498 R=4.580e+00 
R6376t6372 n6377 n6373 R=3.533e+01 
R6376t2838 n6377 n2839 R=9.616e+01 
R6376t1484 n6377 n1 R=1.012e+01 
R6376t3244 n6377 n3245 R=2.918e+02 
R6376t4577 n6377 n4578 R=1.833e+01 
R6376t627 n6377 n628 R=1.388e+01 
R6377t2676 n6378 n2677 R=1.662e+01 
R6377t2193 n6378 n2194 R=4.087e+00 
R6377t2806 n6378 n2807 R=2.157e+01 
R6378t5764 n6379 n5765 R=2.829e+01 
R6378t396 n6379 n397 R=4.259e+00 
R6378t3963 n6379 n3964 R=8.736e+00 
R6378t293 n6379 n294 R=1.114e+02 
R6379t1898 n6380 n1899 R=4.846e+00 
R6379t6181 n6380 n6182 R=7.621e+00 
R6379t1320 n6380 n1321 R=1.697e+01 
R6379t5656 n6380 n5657 R=1.128e+01 
R6379t2314 n6380 n2315 R=5.812e+01 
R6380t943 n6381 n944 R=8.866e+00 
R6380t1995 n6381 n1996 R=6.932e+00 
R6380t131 n6381 n132 R=1.139e+02 
R6381t3521 n6382 n3522 R=1.296e+01 
R6381t1426 n6382 n1427 R=7.572e+01 
R6381t6092 n6382 n6093 R=7.362e+01 
R6382t1720 n6383 n1721 R=1.375e+01 
R6382t4511 n6383 n4512 R=8.319e+00 
R6382t4985 n6383 n4986 R=5.455e+00 
R6382t6324 n6383 n6325 R=6.170e+00 
R6383t5173 n6384 n5174 R=1.508e+01 
R6383t5464 n6384 n5465 R=1.385e+01 
R6383t4538 n6384 n4539 R=2.649e+00 
R6383t4188 n6384 n4189 R=1.463e+01 
R6384t100 n6385 n101 R=7.202e+00 
R6384t4084 n6385 n4085 R=5.011e+00 
R6384t4262 n6385 n4263 R=8.765e+01 
R6384t5789 n6385 n5790 R=1.019e+01 
R6384t1430 n6385 n1431 R=2.463e+02 
R6385t4772 n6386 n4773 R=6.202e+00 
R6385t2018 n6386 n2019 R=4.436e+00 
R6385t2387 n6386 n2388 R=6.730e+00 
R6385t3435 n6386 n3436 R=1.988e+01 
R6386t3211 n6387 n3212 R=2.718e+00 
R6386t3148 n6387 n3149 R=2.867e+01 
R6387t785 n6388 n786 R=4.905e+00 
R6387t859 n6388 n860 R=7.832e+00 
R6387t2786 n6388 n2787 R=8.694e+00 
R6387t786 n6388 n787 R=6.926e+00 
R6387t5636 n6388 n5637 R=5.557e+01 
R6387t1202 n6388 n1203 R=7.993e+01 
R6387t541 n6388 n542 R=3.527e+01 
R6388t4393 n6389 n4394 R=3.854e+04 
R6388t4437 n6389 n4438 R=6.294e+00 
R6388t1135 n6389 n1136 R=5.979e+00 
R6388t414 n6389 n415 R=2.744e+01 
R6389t2019 n6390 n2020 R=3.551e+00 
R6389t5619 n6390 n5620 R=7.383e+00 
R6389t5289 n6390 n5290 R=6.125e+00 
R6389t1337 n6390 n1338 R=6.587e+00 
R6389t2514 n6390 n2515 R=5.081e+01 
R6390t2431 n6391 n2432 R=2.633e+01 
R6390t3126 n6391 n3127 R=4.490e+00 
R6390t5331 n6391 n5332 R=4.355e+00 
R6391t6280 n6392 n6281 R=2.589e+01 
R6391t1487 n6392 n1488 R=1.333e+01 
R6391t3901 n6392 n3902 R=7.067e+00 
R6391t5929 n6392 n5930 R=1.439e+01 
R6392t3105 n6393 n3106 R=1.772e+00 
R6392t845 n6393 n846 R=3.584e+00 
R6393t3350 n6394 n3351 R=6.576e+00 
R6393t3841 n6394 n3842 R=8.331e+00 
R6393t2599 n6394 n2600 R=3.863e+01 
R6393t3713 n6394 n3714 R=2.860e+00 
R6393t5612 n6394 n5613 R=2.342e+01 
R6393t4182 n6394 n4183 R=5.843e+00 
R6394t377 n6395 n378 R=1.423e+01 
R6394t2170 n6395 n2171 R=2.511e+00 
R6394t4033 n6395 n4034 R=3.907e+00 
R6394t155 n6395 n156 R=7.979e+00 
R6395t1073 n6396 n1074 R=6.054e+00 
R6395t5681 n6396 n5682 R=2.181e+00 
R6395t3250 n6396 n3251 R=3.440e+00 
R6396t1751 n6397 n1752 R=1.549e+01 
R6397t2821 n6398 n2822 R=1.433e+01 
R6397t1280 n6398 n1281 R=8.371e+00 
R6397t4299 n6398 n4300 R=3.652e+00 
R6398t2340 n6399 n2341 R=3.444e+00 
R6398t3218 n6399 n3219 R=8.407e+00 
R6398t3439 n6399 n3440 R=7.074e+01 
R6398t2374 n6399 n2375 R=5.695e+01 
R6398t5579 n6399 n5580 R=2.619e+00 
R6398t1479 n6399 n1480 R=2.484e+01 
R6399t1855 n6400 n1856 R=6.646e+00 
R6399t6198 n6400 n6199 R=2.148e+01 
R6400t5623 n6401 n5624 R=7.241e+00 
R6400t6088 n6401 n6089 R=1.169e+01 
R6400t2064 n6401 n2065 R=4.362e+00 
R6401t3399 n6402 n3400 R=2.445e+01 
R6402t3352 n6403 n3353 R=3.431e+01 
R6402t44 n6403 n45 R=2.630e+01 
R6403t781 n6404 n782 R=2.613e+00 
R6403t4341 n6404 n4342 R=2.208e+00 
R6403t5543 n6404 n5544 R=1.749e+01 
R6403t1277 n6404 n1278 R=1.968e+01 
R6404t5620 n6405 n5621 R=1.292e+01 
R6404t3976 n6405 n3977 R=9.329e+00 
R6404t512 n6405 n513 R=5.377e+00 
R6404t905 n6405 n906 R=1.676e+01 
R6404t5956 n6405 n5957 R=1.686e+01 
R6405t4830 n6406 n4831 R=1.274e+01 
R6405t3202 n6406 n3203 R=3.805e+00 
R6405t4301 n6406 n4302 R=6.876e+00 
R6405t1186 n6406 n1187 R=4.308e+01 
R6405t4478 n6406 n4479 R=9.743e+00 
R6405t3268 n6406 n3269 R=3.696e+00 
R6406t3923 n6407 n3924 R=2.978e+00 
R6406t874 n6407 n875 R=2.208e+01 
R6406t4014 n6407 n4015 R=1.049e+01 
R6407t5085 n6408 n5086 R=4.587e+00 
R6407t2670 n6408 n2671 R=3.851e+00 
R6407t4237 n6408 n4238 R=1.677e+01 
R6407t4746 n6408 n4747 R=8.122e+00 
R6407t1637 n6408 n1638 R=3.843e+01 
R6407t3737 n6408 n3738 R=9.646e+00 
R6408t745 n6409 n746 R=7.562e+00 
R6408t548 n6409 n549 R=1.111e+01 
R6408t5458 n6409 n5459 R=5.652e+00 
R6408t5742 n6409 n5743 R=5.436e+00 
R6408t5783 n6409 n5784 R=1.598e+01 
R6409t3188 n6410 n3189 R=1.372e+01 
R6409t5360 n6410 n5361 R=4.249e+00 
R6409t4479 n6410 n4480 R=9.271e+01 
R6410t3583 n6411 n3584 R=3.497e+01 
R6410t184 n6411 n185 R=3.528e+00 
R6410t4937 n6411 n4938 R=4.292e+01 
R6411t5880 n6412 n5881 R=1.304e+01 
R6412t4413 n6413 n4414 R=2.458e+00 
R6412t3725 n6413 n3726 R=1.272e+01 
R6412t658 n6413 n659 R=1.334e+01 
R6412t3424 n6413 n3425 R=1.991e+00 
R6413t331 n6414 n332 R=3.002e+00 
R6413t4363 n6414 n4364 R=5.208e+00 
R6414t1125 n6415 n1126 R=4.652e+00 
R6414t3053 n6415 n3054 R=1.318e+01 
R6414t5989 n6415 n5990 R=8.839e+00 
R6414t2316 n6415 n2317 R=3.183e+00 
R6415t3001 n6416 n3002 R=6.818e+01 
R6415t6004 n6416 n6005 R=9.226e+00 
R6415t2120 n6416 n2121 R=4.145e+01 
R6415t2364 n6416 n2365 R=1.233e+01 
R6416t5960 n6417 n5961 R=1.131e+01 
R6416t5885 n6417 n5886 R=1.775e+00 
R6416t3881 n6417 n3882 R=9.220e+01 
R6416t473 n6417 n474 R=1.821e+00 
R6417t1867 n6418 n1868 R=2.030e+01 
R6418t298 n6419 n299 R=1.369e+02 
R6418t4474 n6419 n4475 R=1.781e+00 
R6418t899 n6419 n900 R=1.415e+02 
R6418t2824 n6419 n2825 R=3.835e+00 
R6419t1844 n6420 n1845 R=3.845e+01 
R6419t4755 n6420 n4756 R=6.805e+00 
R6419t2867 n6420 n2868 R=3.420e+00 
R6419t3408 n6420 n3409 R=1.662e+01 
R6420t1386 n6421 n1387 R=4.993e+00 
R6420t730 n6421 n731 R=7.748e+00 
R6420t1311 n6421 n1312 R=6.957e+00 
R6421t1167 n6422 n1168 R=1.039e+01 
R6421t5573 n6422 n5574 R=6.066e+00 
R6421t1896 n6422 n1897 R=6.064e+00 
R6421t3996 n6422 n3997 R=1.104e+01 
R6422t4289 n6423 n4290 R=4.476e+00 
R6422t3226 n6423 n3227 R=6.146e+00 
R6422t1964 n6423 n1965 R=5.595e+01 
R6423t1295 n6424 n1296 R=8.694e+00 
R6423t1031 n6424 n1032 R=3.326e+00 
R6423t2459 n6424 n2460 R=9.296e+01 
R6423t6066 n6424 n6067 R=4.843e+00 
R6423t3157 n6424 n3158 R=3.973e+00 
R6424t912 n6425 n913 R=2.820e+00 
R6424t1576 n6425 n1577 R=5.634e+00 
R6424t3550 n6425 n3551 R=7.758e+01 
R6425t2721 n6426 n2722 R=2.300e+00 
R6425t3615 n6426 n3616 R=1.439e+01 
R6426t1285 n6427 n1286 R=8.860e+00 
R6426t2050 n6427 n2051 R=7.883e+00 
R6426t1554 n6427 n1555 R=3.977e+01 
R6426t4342 n6427 n4343 R=1.315e+01 
R6426t3446 n6427 n3447 R=1.778e+03 
R6427t1386 n6428 n1387 R=1.069e+01 
R6427t833 n6428 n834 R=7.669e+00 
R6427t724 n6428 n725 R=3.722e+00 
R6428t4584 n6429 n4585 R=5.024e+01 
R6428t4830 n6429 n4831 R=5.725e+00 
R6428t1780 n6429 n1781 R=3.188e+01 
R6428t4536 n6429 n4537 R=5.978e+00 
R6428t3494 n6429 n3495 R=3.792e+00 
R6428t1715 n6429 n1716 R=3.414e+01 
R6428t4647 n6429 n4648 R=2.606e+02 
R6428t3202 n6429 n3203 R=7.398e+00 
R6428t6405 n6429 n6406 R=4.258e+01 
R6429t3294 n6430 n3295 R=8.659e+00 
R6429t4146 n6430 n4147 R=1.373e+01 
R6429t1771 n6430 n1772 R=4.942e+01 
R6430t1367 n6431 n1368 R=4.994e+00 
R6430t3590 n6431 n3591 R=4.397e+00 
R6430t4235 n6431 n4236 R=2.830e+00 
R6431t228 n6432 n229 R=5.016e+00 
R6431t804 n6432 n805 R=5.617e+00 
R6431t3699 n6432 n3700 R=4.265e+00 
R6431t5254 n6432 n5255 R=7.307e+01 
R6432t882 n6433 n883 R=2.690e+00 
R6432t2034 n6433 n2035 R=9.322e+00 
R6432t5381 n6433 n5382 R=1.125e+01 
R6433t2197 n6434 n2198 R=7.480e+00 
R6433t5562 n6434 n5563 R=4.447e+00 
R6433t6122 n6434 n6123 R=8.789e+00 
R6433t6083 n6434 n6084 R=1.256e+01 
R6434t5116 n6435 n5117 R=5.265e+01 
R6434t4169 n6435 n4170 R=3.486e+00 
R6434t5659 n6435 n5660 R=9.936e+01 
R6435t421 n6436 n422 R=2.435e+00 
R6435t5688 n6436 n5689 R=1.472e+01 
R6435t3660 n6436 n3661 R=3.930e+00 
R6436t4673 n6437 n4674 R=1.114e+01 
R6436t5916 n6437 n5917 R=5.940e+00 
R6436t1660 n6437 n1661 R=9.559e+02 
R6436t1816 n6437 n1817 R=2.827e+00 
R6436t3741 n6437 n3742 R=3.628e+01 
R6436t950 n6437 n951 R=8.022e+00 
R6437t4873 n6438 n4874 R=2.812e+00 
R6437t4883 n6438 n4884 R=4.421e+02 
R6437t4215 n6438 n4216 R=5.764e+00 
R6438t5928 n6439 n5929 R=7.113e+00 
R6438t5406 n6439 n5407 R=5.347e+00 
R6438t1214 n6439 n1215 R=5.667e+00 
R6439t981 n6440 n982 R=1.805e+01 
R6439t6263 n6440 n6264 R=3.671e+00 
R6439t3784 n6440 n3785 R=2.613e+02 
R6439t3497 n6440 n3498 R=2.908e+00 
R6440t6352 n6441 n6353 R=7.951e+00 
R6440t335 n6441 n336 R=2.849e+00 
R6440t1172 n6441 n1173 R=1.591e+01 
R6441t1548 n6442 n1549 R=8.140e+00 
R6441t1677 n6442 n1678 R=5.556e+00 
R6441t4497 n6442 n4498 R=5.793e+00 
R6441t4076 n6442 n4077 R=1.478e+01 
R6441t317 n6442 n318 R=1.456e+01 
R6442t215 n6443 n216 R=7.267e+00 
R6442t4658 n6443 n4659 R=1.787e+01 
R6442t2175 n6443 n2176 R=5.561e+00 
R6442t4584 n6443 n4585 R=1.049e+01 
R6442t4450 n6443 n4451 R=4.668e+00 
R6442t2761 n6443 n2762 R=7.684e+00 
R6442t4254 n6443 n4255 R=2.644e+01 
R6443t3800 n6444 n3801 R=1.159e+01 
R6443t4039 n6444 n4040 R=1.640e+01 
R6444t768 n6445 n769 R=1.658e+01 
R6444t2099 n6445 n2100 R=7.883e+01 
R6444t4622 n6445 n4623 R=2.203e+00 
R6444t1901 n6445 n1902 R=1.086e+01 
R6445t3168 n6446 n1 R=4.938e+00 
R6445t6090 n6446 n6091 R=6.869e+01 
R6445t4778 n6446 n1 R=2.189e+00 
R6445t2850 n6446 n1 R=1.052e+01 
R6446t846 n6447 n847 R=5.533e+00 
R6446t6095 n6447 n6096 R=7.758e+00 
R6446t3035 n6447 n3036 R=3.520e+00 
R6446t2732 n6447 n2733 R=7.752e+00 
R6446t3501 n6447 n3502 R=6.275e+01 
R6447t4643 n6448 n4644 R=6.677e+00 
R6447t5815 n6448 n5816 R=1.196e+01 
R6448t900 n6449 n901 R=9.487e+01 
R6448t3969 n6449 n3970 R=4.239e+00 
R6448t5260 n6449 n5261 R=3.879e+00 
R6449t6194 n6450 n6195 R=1.154e+01 
R6449t1868 n6450 n1869 R=9.339e+00 
R6449t1341 n6450 n1342 R=3.596e+00 
R6449t5536 n6450 n5537 R=1.199e+03 
R6449t1382 n6450 n1383 R=6.708e+00 
R6450t195 n6451 n196 R=3.043e+00 
R6450t5851 n6451 n5852 R=8.667e+00 
R6450t3399 n6451 n3400 R=1.299e+01 
R6450t6401 n6451 n6402 R=3.417e+00 
R6451t3230 n6452 n3231 R=5.476e+00 
R6451t3406 n6452 n3407 R=2.761e+00 
R6451t1440 n6452 n1441 R=6.964e+00 
R6452t1864 n6453 n1865 R=8.870e+00 
R6452t149 n6453 n150 R=5.067e+00 
R6453t1651 n6454 n1652 R=2.042e+01 
R6453t3066 n6454 n3067 R=3.449e+00 
R6453t2712 n6454 n2713 R=4.348e+00 
R6453t3361 n6454 n3362 R=6.296e+00 
R6454t6175 n6455 n6176 R=1.412e+01 
R6454t30 n6455 n31 R=4.523e+00 
R6455t909 n6456 n910 R=7.520e+00 
R6455t5003 n6456 n5004 R=1.819e+01 
R6455t4203 n6456 n4204 R=5.500e+00 
R6455t2978 n6456 n2979 R=3.580e+00 
R6455t1127 n6456 n1128 R=1.978e+01 
R6456t6323 n6457 n6324 R=3.306e+00 
R6456t604 n6457 n605 R=3.864e+00 
R6456t3136 n6457 n3137 R=9.848e+00 
R6457t2530 n6458 n2531 R=5.064e+00 
R6458t5044 n6459 n5045 R=3.202e+01 
R6458t153 n6459 n154 R=2.064e+00 
R6459t5694 n6460 n5695 R=3.194e+01 
R6459t4295 n6460 n4296 R=5.712e+00 
R6460t4415 n6461 n4416 R=6.161e+00 
R6460t3189 n6461 n3190 R=2.229e+02 
R6460t1435 n6461 n1436 R=1.471e+01 
R6460t3026 n6461 n3027 R=6.904e+00 
R6460t3802 n6461 n3803 R=3.446e+01 
R6461t1987 n6462 n1988 R=7.600e+00 
R6461t5723 n6462 n5724 R=4.641e+00 
R6461t5485 n6462 n5486 R=7.390e+00 
R6461t4267 n6462 n4268 R=2.174e+01 
R6462t5593 n6463 n5594 R=2.856e+01 
R6462t5189 n6463 n5190 R=2.638e+00 
R6462t5419 n6463 n5420 R=6.143e+01 
R6462t2857 n6463 n2858 R=7.278e+00 
R6462t101 n6463 n102 R=1.181e+01 
R6462t5793 n6463 n5794 R=7.731e+00 
R6463t2786 n6464 n2787 R=2.004e+00 
R6463t859 n6464 n860 R=1.953e+01 
R6464t3932 n6465 n3933 R=7.963e+00 
R6464t6045 n6465 n6046 R=9.839e+00 
R6464t6001 n6465 n6002 R=7.658e+00 
R6464t5248 n6465 n5249 R=1.582e+02 
R6464t1237 n6465 n1238 R=4.409e+00 
R6464t1773 n6465 n1774 R=1.145e+01 
R6464t2697 n6465 n2698 R=1.107e+01 
R6464t2420 n6465 n2421 R=3.717e+01 
R6465t1997 n6466 n1998 R=3.065e+00 
R6465t4998 n6466 n4999 R=5.001e+01 
R6466t1446 n6467 n1447 R=1.378e+01 
R6466t1590 n6467 n1591 R=4.335e+00 
R6466t2572 n6467 n2573 R=3.124e+01 
R6466t2542 n6467 n2543 R=5.304e+00 
R6466t195 n6467 n196 R=9.451e+00 
R6466t2461 n6467 n2462 R=6.265e+00 
R6467t2955 n6468 n2956 R=3.960e+00 
R6467t5187 n6468 n5188 R=1.016e+01 
R6467t2094 n6468 n2095 R=2.297e+01 
R6467t1373 n6468 n1374 R=3.038e+00 
R6468t2281 n6469 n2282 R=2.516e+00 
R6468t4434 n6469 n4435 R=2.762e+01 
R6468t257 n6469 n258 R=1.232e+01 
R6468t761 n6469 n762 R=7.719e+00 
R6470t3542 n6471 n3543 R=2.147e+01 
R6470t5919 n6471 n5920 R=6.545e+00 
R6470t4835 n6471 n4836 R=5.635e+00 
R6471t5505 n6472 n5506 R=2.049e+00 
R6471t3198 n6472 n3199 R=6.293e+00 
R6471t87 n6472 n88 R=2.758e+00 
R6472t1968 n6473 n1969 R=2.523e+01 
R6472t2388 n6473 n2389 R=2.273e+01 
R6472t4521 n6473 n4522 R=5.310e+00 
R6472t3672 n6473 n3673 R=7.828e+00 
R6472t3837 n6473 n3838 R=2.171e+01 
R6473t864 n6474 n865 R=5.786e+00 
R6473t3430 n6474 n3431 R=8.469e+00 
R6474t3876 n6475 n3877 R=1.144e+01 
R6474t5351 n6475 n5352 R=8.914e+00 
R6474t6075 n6475 n6076 R=9.122e+00 
R6475t2817 n6476 n2818 R=3.103e+01 
R6475t5938 n6476 n5939 R=4.718e+00 
R6475t3680 n6476 n3681 R=1.090e+01 
R6476t6000 n6477 n6001 R=3.407e+00 
R6476t5933 n6477 n5934 R=3.894e+00 
R6477t2979 n6478 n2980 R=1.241e+01 
R6477t2026 n6478 n2027 R=4.667e+00 
R6477t5145 n6478 n5146 R=1.437e+01 
R6477t4679 n6478 n4680 R=3.662e+00 
R6477t815 n6478 n816 R=8.322e+01 
R6478t1881 n6479 n1882 R=4.006e+01 
R6478t3353 n6479 n3354 R=2.904e+00 
R6478t6242 n6479 n6243 R=7.604e+00 
R6478t4298 n6479 n4299 R=4.261e+00 
R6479t6148 n6480 n6149 R=2.114e+00 
R6479t4505 n6480 n4506 R=3.448e+01 
R6479t5190 n6480 n5191 R=3.116e+01 
R6479t5943 n6480 n5944 R=6.360e+00 
R6480t4040 n6481 n4041 R=1.487e+00 
R6480t5745 n6481 n5746 R=8.218e+00 
R6480t3601 n6481 n3602 R=1.952e+03 
R6480t1606 n6481 n1607 R=9.834e+00 
R6481t1122 n6482 n1123 R=7.630e+00 
R6481t5954 n6482 n5955 R=6.597e+00 
R6481t3086 n6482 n3087 R=2.509e+01 
R6481t5362 n6482 n5363 R=7.607e+00 
R6481t1204 n6482 n1205 R=4.831e+00 
R6482t6034 n6483 n6035 R=1.211e+01 
R6482t1954 n6483 n1955 R=3.367e+00 
R6482t3244 n6483 n3245 R=1.224e+01 
R6483t2686 n6484 n2687 R=5.559e+00 
R6483t3843 n6484 n3844 R=3.130e+01 
R6483t539 n6484 n540 R=1.586e+01 
R6483t2863 n6484 n2864 R=3.764e+00 
R6484t2903 n6485 n2904 R=2.263e+01 
R6484t6078 n6485 n6079 R=2.545e+01 
R6484t4985 n6485 n4986 R=6.260e+00 
R6484t6317 n6485 n6318 R=3.703e+00 
R6484t1249 n6485 n1250 R=9.942e+00 
R6484t1260 n6485 n1261 R=5.559e+00 
R6485t2099 n6486 n2100 R=3.551e+01 
R6485t5111 n6486 n5112 R=1.013e+02 
R6485t5216 n6486 n5217 R=3.209e+00 
R6485t4464 n6486 n4465 R=6.290e+00 
R6486t735 n6487 n736 R=7.102e+00 
R6486t4550 n6487 n4551 R=1.670e+01 
R6486t3627 n6487 n3628 R=2.765e+00 
R6487t1297 n6488 n1298 R=3.981e+00 
R6487t2462 n6488 n2463 R=9.754e+00 
R6487t5426 n6488 n5427 R=1.596e+01 
R6487t5888 n6488 n5889 R=1.268e+01 
R6487t6100 n6488 n6101 R=1.258e+01 
R6488t2032 n6489 n2033 R=1.199e+01 
R6488t2702 n6489 n2703 R=6.123e+00 
R6488t6452 n6489 n6453 R=2.973e+00 
R6488t1864 n6489 n1865 R=9.887e+02 
R6488t1458 n6489 n1459 R=5.043e+00 
R6489t711 n6490 n712 R=8.305e+00 
R6489t3034 n6490 n3035 R=1.081e+01 
R6489t350 n6490 n351 R=7.176e+00 
R6489t3343 n6490 n3344 R=6.649e+00 
R6489t6245 n6490 n6246 R=4.845e+01 
R6489t634 n6490 n635 R=6.146e+00 
R6490t3722 n6491 n3723 R=6.784e+00 
R6490t3186 n6491 n3187 R=4.406e+00 
R6490t2058 n6491 n2059 R=1.624e+02 
R6491t2960 n6492 n2961 R=2.477e+01 
R6491t4720 n6492 n4721 R=7.285e+00 
R6491t4539 n6492 n4540 R=4.003e+00 
R6491t3792 n6492 n3793 R=5.283e+00 
R6492t3792 n6493 n3793 R=6.749e+00 
R6492t414 n6493 n415 R=2.164e+00 
R6493t886 n6494 n887 R=1.300e+01 
R6493t3398 n6494 n3399 R=6.580e+00 
R6493t5002 n6494 n5003 R=1.576e+01 
R6493t6274 n6494 n6275 R=4.813e+00 
R6493t3950 n6494 n3951 R=8.211e+00 
R6493t612 n6494 n613 R=1.315e+01 
R6493t4710 n6494 n4711 R=3.714e+01 
R6494t973 n6495 n974 R=9.360e+00 
R6494t4948 n6495 n4949 R=4.306e+00 
R6494t324 n6495 n325 R=5.373e+00 
R6494t5886 n6495 n5887 R=2.095e+01 
R6494t3190 n6495 n3191 R=5.054e+00 
R6494t3417 n6495 n3418 R=2.900e+01 
R6494t2403 n6495 n2404 R=1.589e+02 
R6495t6132 n6496 n6133 R=1.662e+01 
R6496t1498 n6497 n1499 R=1.189e+01 
R6496t2774 n6497 n2775 R=6.104e+00 
R6496t2337 n6497 n2338 R=2.055e+01 
R6496t3726 n6497 n3727 R=1.644e+01 
R6496t2639 n6497 n2640 R=1.375e+01 
R6496t1794 n6497 n1795 R=3.599e+00 
R6497t763 n6498 n764 R=2.215e+00 
R6497t816 n6498 n817 R=1.566e+01 
R6497t6249 n6498 n6250 R=2.222e+01 
R6497t981 n6498 n982 R=1.345e+02 
R6497t586 n6498 n587 R=4.803e+00 
R6498t2455 n6499 n2456 R=1.386e+00 
R6498t3052 n6499 n3053 R=3.864e+01 
R6498t4418 n6499 n4419 R=3.195e+00 
R6499t2234 n6500 n2235 R=8.641e+00 
R6499t366 n6500 n367 R=2.776e+01 
R6499t869 n6500 n870 R=3.408e+00 
R6499t4192 n6500 n4193 R=9.201e+00 
R6499t2389 n6500 n2390 R=1.025e+02 
R6499t2300 n6500 n2301 R=2.808e+01 
R6499t5813 n6500 n5814 R=3.253e+00 
R6499t4660 n6500 n4661 R=2.862e+01 
R6500t3760 n6501 n3761 R=3.230e+00 
R6500t4238 n6501 n4239 R=2.587e+00 
R6500t2073 n6501 n2074 R=5.098e+00 
R6501t5114 n6502 n5115 R=9.846e+00 
R6502t4809 n6503 n4810 R=3.218e+00 
R6502t5808 n6503 n5809 R=8.982e+00 
R6502t3683 n6503 n3684 R=1.421e+01 
R6502t6058 n6503 n6059 R=1.161e+01 
R6502t3059 n6503 n3060 R=1.211e+01 
R6503t1334 n6504 n1335 R=2.570e+01 
R6503t3002 n6504 n3003 R=1.293e+01 
R6503t5380 n6504 n5381 R=1.767e+01 
R6503t3689 n6504 n3690 R=1.542e+01 
R6503t5027 n6504 n5028 R=2.105e+01 
R6503t3023 n6504 n3024 R=1.328e+01 
R6503t4852 n6504 n4853 R=1.203e+01 
R6503t5869 n6504 n5870 R=3.798e+01 
R6503t5673 n6504 n5674 R=5.407e+01 
R6503t36 n6504 n37 R=5.440e+00 
R6503t755 n6504 n756 R=2.331e+01 
R6504t4252 n6505 n4253 R=3.099e+01 
R6504t1504 n6505 n1505 R=2.768e+00 
R6504t647 n6505 n648 R=1.669e+01 
R6504t1872 n6505 n1873 R=1.180e+02 
R6505t555 n6506 n556 R=5.839e+00 
R6505t6086 n6506 n6087 R=1.797e+01 
R6505t5600 n6506 n5601 R=7.421e+00 
R6505t4369 n6506 n4370 R=2.345e+00 
R6505t3975 n6506 n3976 R=2.188e+01 
R6506t3211 n6507 n3212 R=1.188e+01 
R6506t6386 n6507 n6387 R=2.220e+01 
R6506t6159 n6507 n6160 R=7.404e+00 
R6506t1800 n6507 n1801 R=4.069e+00 
R6507t2243 n6508 n2244 R=1.181e+01 
R6507t4136 n6508 n4137 R=2.746e+00 
R6507t1892 n6508 n1893 R=1.011e+01 
R6507t3065 n6508 n3066 R=4.637e+00 
R6507t3730 n6508 n3731 R=1.225e+01 
R6508t3722 n6509 n3723 R=7.541e+00 
R6508t3186 n6509 n3187 R=3.194e+00 
R6508t2166 n6509 n2167 R=1.821e+01 
R6508t1820 n6509 n1821 R=3.882e+00 
R6509t730 n6510 n731 R=2.247e+01 
R6509t1386 n6510 n1387 R=9.282e+00 
R6509t6427 n6510 n6428 R=4.314e+00 
R6509t724 n6510 n725 R=1.408e+01 
R6509t2617 n6510 n2618 R=4.935e+01 
R6509t3915 n6510 n3916 R=3.913e+00 
R6509t2098 n6510 n2099 R=6.248e+00 
R6510t442 n6511 n443 R=8.525e+00 
R6510t2465 n6511 n2466 R=9.074e+00 
R6512t4437 n6513 n4438 R=1.047e+01 
R6512t4705 n6513 n4706 R=3.089e+00 
R6512t5439 n6513 n5440 R=5.984e+00 
R6512t1135 n6513 n1136 R=1.768e+01 
R6513t4752 n6514 n4753 R=1.554e+01 
R6513t4934 n6514 n4935 R=3.705e+00 
R6513t3532 n6514 n3533 R=4.698e+00 
R6513t1966 n6514 n1967 R=5.341e+00 
R6514t1178 n6515 n1179 R=2.973e+00 
R6514t1388 n6515 n1389 R=1.652e+01 
R6514t549 n6515 n550 R=1.313e+01 
R6514t4077 n6515 n4078 R=1.314e+01 
R6514t2424 n6515 n2425 R=3.341e+00 
R6515t5357 n6516 n5358 R=2.644e+01 
R6515t962 n6516 n963 R=9.441e+00 
R6515t1810 n6516 n1811 R=5.241e+00 
R6515t6061 n6516 n6062 R=1.182e+01 
R6516t3420 n6517 n3421 R=1.585e+01 
R6516t1197 n6517 n1198 R=2.884e+00 
R6517t5638 n6518 n5639 R=4.003e+00 
R6517t496 n6518 n497 R=8.862e+00 
R6517t6308 n6518 n6309 R=1.616e+01 
R6517t1059 n6518 n1060 R=5.508e+00 
R6518t1705 n6519 n1706 R=3.823e+00 
R6518t4446 n6519 n4447 R=8.490e+02 
R6518t2780 n6519 n2781 R=4.989e+00 
R6518t6344 n6519 n6345 R=1.278e+01 
R6519t1876 n6520 n1877 R=1.923e+00 
R6519t3008 n6520 n3009 R=1.003e+01 
R6519t1537 n6520 n1538 R=6.808e+00 
R6520t780 n6521 n781 R=2.956e+00 
R6521t830 n6522 n831 R=1.534e+01 
R6521t5226 n6522 n5227 R=1.712e+01 
R6521t516 n6522 n517 R=1.556e+01 
R6521t2153 n6522 n2154 R=2.301e+01 
R6522t5615 n6523 n5616 R=1.611e+01 
R6522t2931 n6523 n2932 R=5.629e+00 
R6522t2193 n6523 n2194 R=1.290e+01 
R6522t6222 n6523 n6223 R=1.464e+01 
R6523t4642 n6524 n4643 R=3.072e+01 
R6523t4870 n6524 n4871 R=4.294e+00 
R6523t365 n6524 n366 R=2.913e+01 
R6523t2422 n6524 n2423 R=8.106e+00 
R6523t3355 n6524 n3356 R=3.175e+01 
R6524t4199 n6525 n4200 R=1.695e+01 
R6524t4563 n6525 n4564 R=1.985e+01 
R6524t2077 n6525 n2078 R=5.251e+01 
R6524t136 n6525 n137 R=1.335e+01 
R6524t5235 n6525 n5236 R=3.702e+00 
R6524t5004 n6525 n5005 R=3.251e+00 
R6525t5058 n6526 n5059 R=6.508e+00 
R6525t4867 n6526 n4868 R=1.835e+01 
R6525t5846 n6526 n5847 R=3.247e+00 
R6525t914 n6526 n915 R=9.507e+01 
R6526t625 n6527 n626 R=4.777e+00 
R6526t5036 n6527 n5037 R=1.852e+01 
R6526t80 n6527 n81 R=2.173e+00 
R6526t4745 n6527 n4746 R=5.198e+02 
R6527t4601 n6528 n4602 R=3.663e+00 
R6527t3223 n6528 n1 R=6.150e+00 
R6527t6119 n6528 n1 R=5.572e+00 
R6527t2901 n6528 n2902 R=5.861e+01 
R6528t178 n6529 n179 R=7.094e+00 
R6528t4247 n6529 n4248 R=7.652e+00 
R6528t1320 n6529 n1321 R=2.312e+01 
R6528t5656 n6529 n5657 R=4.609e+00 
R6528t1188 n6529 n1189 R=6.183e+00 
R6529t5000 n6530 n5001 R=5.875e+00 
R6529t2947 n6530 n2948 R=6.632e+00 
R6529t5571 n6530 n5572 R=6.686e+00 
R6530t2481 n6531 n2482 R=3.245e+00 
R6530t2849 n6531 n2850 R=6.557e+00 
R6530t1663 n6531 n1664 R=2.734e+01 
R6531t1471 n6532 n1472 R=2.547e+00 
R6531t417 n6532 n418 R=3.809e+00 
R6531t5056 n6532 n5057 R=3.992e+01 
R6532t421 n6533 n422 R=7.375e+00 
R6532t6435 n6533 n6436 R=2.788e+01 
R6533t147 n6534 n148 R=6.151e+00 
R6533t435 n6534 n436 R=3.112e+00 
R6533t1546 n6534 n1547 R=1.621e+01 
R6533t5022 n6534 n5023 R=1.049e+01 
R6534t348 n6535 n349 R=9.306e+01 
R6534t3957 n6535 n3958 R=5.152e+00 
R6534t6011 n6535 n6012 R=9.678e+00 
R6534t1047 n6535 n1048 R=5.058e+00 
R6534t3102 n6535 n3103 R=3.121e+00 
R6535t464 n6536 n465 R=8.345e+00 
R6535t3906 n6536 n3907 R=4.738e+00 
R6535t2755 n6536 n2756 R=1.961e+01 
R6535t1359 n6536 n1360 R=4.815e+00 
R6535t6479 n6536 n6480 R=4.109e+01 
R6535t6148 n6536 n6149 R=3.961e+00 
R6536t167 n6537 n168 R=5.785e+02 
R6536t1629 n6537 n1630 R=1.352e+01 
R6536t1861 n6537 n1862 R=3.913e+00 
R6536t5155 n6537 n5156 R=3.798e+01 
R6536t2612 n6537 n2613 R=8.201e+00 
R6536t1365 n6537 n1366 R=9.030e+00 
R6537t318 n6538 n319 R=1.147e+01 
R6537t592 n6538 n593 R=3.466e+00 
R6537t2389 n6538 n2390 R=3.073e+00 
R6537t613 n6538 n614 R=7.498e+00 
R6537t55 n6538 n56 R=2.709e+01 
R6538t2129 n6539 n2130 R=4.026e+00 
R6538t5980 n6539 n5981 R=4.269e+01 
R6538t1571 n6539 n1572 R=1.220e+01 
R6538t3603 n6539 n3604 R=3.756e+00 
R6539t4354 n6540 n4355 R=4.734e+00 
R6539t3695 n6540 n3696 R=8.364e+00 
R6539t3070 n6540 n3071 R=3.706e+00 
R6540t372 n6541 n373 R=4.277e+00 
R6540t5171 n6541 n5172 R=4.312e+00 
R6540t5629 n6541 n5630 R=2.651e+00 
R6540t1194 n6541 n1195 R=4.032e+01 
R6540t4485 n6541 n4486 R=3.296e+01 
R6541t4608 n6542 n4609 R=3.309e+01 
R6541t5942 n6542 n5943 R=1.100e+03 
R6541t2179 n6542 n2180 R=1.824e+00 
R6541t1674 n6542 n1675 R=4.298e+01 
R6541t2913 n6542 n2914 R=1.739e+01 
R6541t5766 n6542 n5767 R=1.868e+00 
R6542t4945 n6543 n4946 R=5.973e+01 
R6542t6313 n6543 n6314 R=4.944e+00 
R6542t258 n6543 n259 R=3.147e+00 
R6542t5627 n6543 n5628 R=3.347e+00 
R6543t1712 n6544 n1713 R=1.159e+01 
R6543t5336 n6544 n5337 R=4.124e+01 
R6543t6313 n6544 n6314 R=7.233e+00 
R6543t3326 n6544 n3327 R=1.230e+02 
R6543t2565 n6544 n2566 R=1.003e+01 
R6543t6321 n6544 n6322 R=5.642e+00 
R6543t4607 n6544 n4608 R=5.916e+01 
R6543t6077 n6544 n6078 R=4.789e+00 
R6544t2206 n6545 n2207 R=5.403e+00 
R6544t1776 n6545 n1777 R=2.358e+01 
R6545t2551 n6546 n2552 R=2.645e+00 
R6546t3276 n6547 n3277 R=1.288e+01 
R6546t5680 n6547 n5681 R=6.096e+00 
R6547t1896 n6548 n1897 R=1.046e+01 
R6547t6421 n6548 n6422 R=2.585e+01 
R6547t5054 n6548 n5055 R=8.445e+00 
R6547t4056 n6548 n4057 R=3.037e+00 
R6547t5573 n6548 n5574 R=5.195e+00 
R6548t828 n6549 n829 R=1.792e+01 
R6548t5716 n6549 n5717 R=6.047e+00 
R6548t259 n6549 n260 R=5.981e+00 
R6548t1356 n6549 n1357 R=2.960e+00 
R6548t3167 n6549 n3168 R=5.185e+01 
R6549t3305 n6550 n3306 R=5.058e+00 
R6549t4588 n6550 n4589 R=7.713e+00 
R6549t5977 n6550 n5978 R=1.167e+01 
R6550t2741 n6551 n2742 R=5.695e+00 
R6550t3483 n6551 n3484 R=4.172e+00 
R6550t5641 n6551 n5642 R=4.725e+00 
R6550t5421 n6551 n5422 R=6.652e+00 
R6550t3082 n6551 n3083 R=1.340e+03 
R6550t2314 n6551 n2315 R=2.351e+01 
R6551t377 n6552 n378 R=2.821e+02 
R6551t270 n6552 n271 R=1.867e+01 
R6551t1089 n6552 n1090 R=5.213e+00 
R6551t6188 n6552 n6189 R=2.411e+01 
R6552t2848 n6553 n2849 R=1.344e+01 
R6552t2944 n6553 n2945 R=5.092e+00 
R6552t4817 n6553 n4818 R=8.518e+00 
R6552t5032 n6553 n5033 R=1.243e+01 
R6553t1405 n6554 n1406 R=6.548e+00 
R6553t3716 n6554 n3717 R=1.936e+00 
R6553t600 n6554 n601 R=1.549e+01 
R6554t4157 n6555 n4158 R=4.611e+00 
R6554t5048 n6555 n5049 R=6.292e+00 
R6554t4873 n6555 n4874 R=2.607e+01 
R6554t6437 n6555 n6438 R=1.951e+00 
R6554t4215 n6555 n4216 R=1.005e+02 
R6555t306 n6556 n307 R=4.162e+00 
R6555t1807 n6556 n1808 R=8.459e+00 
R6556t2935 n6557 n2936 R=3.307e+00 
R6556t5139 n6557 n5140 R=5.988e+01 
R6556t2293 n6557 n2294 R=7.425e+00 
R6557t4411 n6558 n4412 R=4.052e+00 
R6557t5981 n6558 n5982 R=5.213e+01 
R6558t1440 n6559 n1441 R=2.928e+01 
R6558t1475 n6559 n1476 R=8.397e+00 
R6558t3011 n6559 n3012 R=1.956e+00 
R6558t471 n6559 n472 R=9.747e+01 
R6558t4116 n6559 n4117 R=7.691e+00 
R6559t1891 n6560 n1892 R=4.797e+01 
R6559t5077 n6560 n5078 R=3.432e+00 
R6559t3270 n6560 n3271 R=4.007e+00 
R6560t3331 n6561 n3332 R=8.338e+00 
R6560t5344 n6561 n5345 R=1.204e+01 
R6561t2756 n6562 n2757 R=1.551e+02 
R6561t4796 n6562 n4797 R=1.356e+01 
R6561t5944 n6562 n5945 R=9.602e+00 
R6561t5124 n6562 n5125 R=4.331e+00 
R6561t3377 n6562 n3378 R=2.483e+00 
R6561t2149 n6562 n2150 R=1.526e+02 
R6562t1064 n6563 n1065 R=5.953e+01 
R6562t1432 n6563 n1433 R=4.440e+00 
R6562t2962 n6563 n2963 R=4.846e+00 
R6562t6227 n6563 n6228 R=1.400e+01 
R6562t1155 n6563 n1156 R=3.125e+01 
R6563t4054 n6564 n4055 R=8.955e+00 
R6563t5100 n6564 n5101 R=4.614e+00 
R6563t1715 n6564 n1716 R=1.170e+01 
R6563t4647 n6564 n4648 R=7.266e+01 
R6563t3352 n6564 n3353 R=4.495e+00 
R6564t110 n6565 n111 R=5.659e+00 
R6564t4416 n6565 n4417 R=8.250e+00 
R6564t1646 n6565 n1647 R=1.085e+01 
R6564t986 n6565 n987 R=7.242e+00 
R6564t4854 n6565 n4855 R=5.161e+00 
R6564t5078 n6565 n5079 R=1.109e+01 
R6565t2403 n6566 n2404 R=5.992e+00 
R6565t6166 n6566 n6167 R=4.591e+00 
R6566t4482 n6567 n4483 R=2.063e+01 
R6566t2099 n6567 n2100 R=2.213e+01 
R6566t1848 n6567 n1849 R=3.767e+00 
R6567t2529 n6568 n2530 R=4.963e+00 
R6567t5740 n6568 n5741 R=3.767e+00 
R6567t302 n6568 n303 R=4.810e+01 
R6568t5416 n6569 n5417 R=4.196e+00 
R6568t3633 n6569 n3634 R=3.270e+01 
R6568t2945 n6569 n2946 R=6.311e+00 
R6568t4646 n6569 n4647 R=1.005e+01 
R6569t1859 n6570 n1860 R=8.004e+00 
R6569t2588 n6570 n2589 R=4.211e+01 
R6569t5473 n6570 n5474 R=6.401e+00 
R6569t4239 n6570 n4240 R=1.523e+01 
R6569t3781 n6570 n3782 R=5.664e+00 
R6569t2884 n6570 n2885 R=3.111e+00 
R6570t317 n6571 n318 R=1.733e+01 
R6570t4373 n6571 n4374 R=2.456e+00 
R6570t5611 n6571 n5612 R=1.161e+01 
R6570t3720 n6571 n3721 R=2.198e+01 
R6571t3548 n6572 n3549 R=3.968e+00 
R6571t135 n6572 n136 R=4.186e+00 
R6572t1798 n6573 n1799 R=1.547e+01 
R6572t4071 n6573 n4072 R=4.027e+00 
R6572t4700 n6573 n4701 R=1.362e+01 
R6573t5440 n6574 n5441 R=4.827e+00 
R6573t3744 n6574 n3745 R=7.453e+00 
R6574t17 n6575 n18 R=5.052e+00 
R6574t822 n6575 n823 R=3.904e+00 
R6574t3204 n6575 n3205 R=3.634e+01 
R6574t649 n6575 n650 R=6.955e+00 
R6575t3179 n6576 n3180 R=4.718e+01 
R6576t814 n6577 n815 R=2.879e+01 
R6576t2411 n6577 n2412 R=8.771e+00 
R6576t3921 n6577 n3922 R=1.265e+01 
R6577t2070 n6578 n2071 R=1.930e+01 
R6577t4475 n6578 n4476 R=8.000e+00 
R6577t1468 n6578 n1469 R=1.439e+01 
R6578t113 n6579 n114 R=7.691e+00 
R6578t6314 n6579 n6315 R=2.184e+01 
R6578t2108 n6579 n2109 R=4.049e+00 
R6578t1742 n6579 n1743 R=1.520e+01 
R6578t4093 n6579 n4094 R=3.408e+00 
R6578t2116 n6579 n2117 R=5.132e+01 
R6579t1841 n6580 n1842 R=5.047e+00 
R6579t5502 n6580 n5503 R=5.332e+00 
R6579t2481 n6580 n2482 R=3.671e+00 
R6579t6530 n6580 n6531 R=1.033e+02 
R6580t3851 n6581 n3852 R=4.399e+00 
R6580t5320 n6581 n5321 R=3.490e+00 
R6580t3612 n6581 n3613 R=1.982e+01 
R6581t3075 n6582 n3076 R=3.839e+00 
R6581t3821 n6582 n3822 R=1.632e+01 
R6581t2872 n6582 n2873 R=4.476e+01 
R6581t1883 n6582 n1884 R=7.809e+00 
R6581t91 n6582 n92 R=2.580e+00 
R6582t5803 n6583 n5804 R=3.012e+00 
R6582t1663 n6583 n1664 R=4.354e+00 
R6582t2201 n6583 n2202 R=4.533e+01 
R6582t1899 n6583 n1900 R=7.787e+00 
R6583t517 n6584 n518 R=4.363e+00 
R6583t3981 n6584 n3982 R=5.964e+00 
R6584t6340 n6585 n6341 R=5.614e+00 
R6584t5487 n6585 n5488 R=1.816e+01 
R6584t5137 n6585 n5138 R=1.340e+01 
R6584t3311 n6585 n3312 R=3.134e+00 
R6585t2243 n6586 n2244 R=2.176e+00 
R6585t5484 n6586 n5485 R=3.374e+00 
R6585t3185 n6586 n3186 R=1.688e+01 
R6586t2294 n6587 n2295 R=2.710e+00 
R6586t2286 n6587 n2287 R=4.055e+00 
R6587t1121 n6588 n1122 R=2.075e+01 
R6587t5904 n6588 n5905 R=2.849e+00 
R6587t2333 n6588 n2334 R=1.252e+02 
R6587t2915 n6588 n2916 R=4.633e+00 
R6588t2688 n6589 n2689 R=3.010e+00 
R6588t2820 n6589 n2821 R=1.225e+01 
R6588t6075 n6589 n6076 R=4.893e+01 
R6588t4907 n6589 n4908 R=2.308e+00 
R6589t1870 n6590 n1871 R=2.673e+01 
R6589t4135 n6590 n4136 R=6.832e+00 
R6589t4747 n6590 n4748 R=2.541e+00 
R6590t5955 n6591 n5956 R=5.027e+00 
R6591t5408 n6592 n5409 R=4.077e+01 
R6591t5640 n6592 n5641 R=2.272e+00 
R6591t6248 n6592 n6249 R=1.768e+01 
R6591t1838 n6592 n1839 R=5.747e+00 
R6592t5947 n6593 n5948 R=9.915e+00 
R6592t6168 n6593 n6169 R=3.354e+00 
R6592t3522 n6593 n3523 R=1.335e+01 
R6593t3414 n6594 n3415 R=5.967e+00 
R6593t5428 n6594 n5429 R=2.774e+00 
R6593t5747 n6594 n5748 R=1.026e+01 
R6593t1230 n6594 n1231 R=4.153e+00 
R6594t1759 n6595 n1760 R=4.413e+00 
R6594t1172 n6595 n1173 R=1.328e+01 
R6594t6440 n6595 n6441 R=3.961e+00 
R6595t98 n6596 n99 R=4.813e+00 
R6595t4526 n6596 n4527 R=1.006e+01 
R6595t3090 n6596 n3091 R=1.679e+02 
R6595t2546 n6596 n2547 R=4.951e+01 
R6595t5110 n6596 n5111 R=4.186e+00 
R6595t108 n6596 n109 R=3.735e+01 
R6595t2331 n6596 n2332 R=9.006e+00 
R6596t3230 n6597 n3231 R=6.663e+00 
R6596t6451 n6597 n6452 R=1.776e+01 
R6596t1854 n6597 n1855 R=5.443e+00 
R6596t4056 n6597 n4057 R=4.070e+01 
R6596t6351 n6597 n6352 R=2.176e+01 
R6596t4849 n6597 n4850 R=4.140e+00 
R6596t3406 n6597 n3407 R=4.903e+02 
R6598t139 n6599 n140 R=1.128e+01 
R6598t972 n6599 n973 R=2.065e+00 
R6598t1592 n6599 n1593 R=5.348e+01 
R6598t2815 n6599 n2816 R=2.014e+01 
R6599t1391 n6600 n1392 R=4.855e+02 
R6599t1486 n6600 n1487 R=3.542e+00 
R6600t5805 n6601 n5806 R=3.775e+01 
R6600t2367 n6601 n2368 R=6.738e+00 
R6600t5533 n6601 n5534 R=1.041e+01 
R6600t676 n6601 n677 R=7.022e+00 
R6600t4150 n6601 n4151 R=7.605e+00 
R6601t4675 n6602 n4676 R=7.193e+01 
R6601t4361 n6602 n4362 R=6.222e+00 
R6601t4599 n6602 n4600 R=1.638e+01 
R6601t1672 n6602 n1673 R=6.111e+00 
R6602t74 n6603 n75 R=1.418e+01 
R6602t2692 n6603 n2693 R=5.416e+00 
R6602t841 n6603 n842 R=1.265e+01 
R6602t5403 n6603 n5404 R=3.203e+00 
R6603t4639 n6604 n4640 R=8.248e+01 
R6603t4942 n6604 n4943 R=1.322e+01 
R6603t1812 n6604 n1813 R=5.014e+00 
R6603t3634 n6604 n3635 R=2.386e+00 
R6604t4177 n6605 n4178 R=5.487e+00 
R6604t6375 n6605 n6376 R=2.932e+00 
R6605t872 n6606 n873 R=6.529e+00 
R6605t6476 n6606 n6477 R=6.083e+00 
R6605t5933 n6606 n5934 R=7.280e+01 
R6605t951 n6606 n952 R=9.496e+00 
R6606t1507 n6607 n1508 R=1.799e+01 
R6606t5650 n6607 n5651 R=8.113e+01 
R6606t2713 n6607 n2714 R=2.129e+01 
R6606t4320 n6607 n4321 R=7.470e+00 
R6606t1580 n6607 n1581 R=4.503e+00 
R6607t5542 n6608 n5543 R=6.106e+00 
R6607t4808 n6608 n4809 R=5.595e+01 
R6607t3709 n6608 n3710 R=6.932e+01 
R6607t4214 n6608 n4215 R=1.376e+00 
R6607t5635 n6608 n5636 R=1.406e+01 
R6607t4914 n6608 n4915 R=6.480e+01 
R6608t911 n6609 n912 R=6.260e+00 
R6608t6175 n6609 n6176 R=6.694e+00 
R6608t6454 n6609 n6455 R=8.305e+00 
R6608t6079 n6609 n6080 R=5.418e+00 
R6608t880 n6609 n881 R=1.917e+01 
R6609t4772 n6610 n4773 R=7.785e+00 
R6609t6385 n6610 n6386 R=1.027e+01 
R6609t2018 n6610 n2019 R=4.753e+01 
R6609t3478 n6610 n3479 R=3.249e+00 
R6610t2567 n6611 n2568 R=1.395e+01 
R6610t968 n6611 n969 R=1.932e+00 
R6611t28 n6612 n29 R=1.397e+01 
R6611t2042 n6612 n2043 R=7.524e+00 
R6611t5425 n6612 n5426 R=7.611e+00 
R6611t1230 n6612 n1231 R=1.700e+01 
R6612t5431 n6613 n5432 R=1.932e+01 
R6612t5040 n6613 n5041 R=3.158e+00 
R6612t1506 n6613 n1507 R=9.048e+00 
R6612t3587 n6613 n3588 R=2.188e+00 
R6612t6234 n6613 n6235 R=6.247e+01 
R6613t575 n6614 n576 R=1.933e+00 
R6613t6029 n6614 n6030 R=1.246e+01 
R6613t2276 n6614 n2277 R=2.526e+02 
R6613t1694 n6614 n1695 R=7.742e+00 
R6613t57 n6614 n58 R=9.336e+00 
R6613t393 n6614 n394 R=1.295e+01 
R6613t977 n6614 n978 R=3.462e+01 
R6614t6590 n6615 n6591 R=3.958e+01 
R6614t2832 n6615 n2833 R=4.608e+02 
R6614t5541 n6615 n5542 R=2.620e+00 
R6614t3507 n6615 n3508 R=4.369e+01 
R6615t5928 n6616 n5929 R=1.922e+01 
R6615t6438 n6616 n6439 R=1.006e+01 
R6615t3700 n6616 n3701 R=2.746e+00 
R6615t1801 n6616 n1802 R=7.654e+01 
R6615t5406 n6616 n5407 R=8.956e+00 
R6616t727 n6617 n728 R=4.163e+00 
R6616t2702 n6617 n2703 R=9.814e+01 
R6616t2032 n6617 n2033 R=6.502e+01 
R6616t4656 n6617 n4657 R=9.931e+00 
R6616t3800 n6617 n3801 R=8.199e+00 
R6616t2925 n6617 n2926 R=1.200e+01 
R6617t1276 n6618 n1277 R=1.836e+01 
R6617t4405 n6618 n4406 R=7.247e+00 
R6618t4503 n6619 n4504 R=3.239e+00 
R6618t5519 n6619 n5520 R=6.048e+00 
R6618t201 n6619 n202 R=1.253e+01 
R6618t578 n6619 n579 R=5.578e+00 
R6619t1483 n6620 n1484 R=4.737e+00 
R6619t6043 n6620 n6044 R=6.596e+00 
R6619t3166 n6620 n3167 R=1.205e+01 
R6619t6354 n6620 n6355 R=4.212e+01 
R6619t5233 n6620 n5234 R=1.252e+02 
R6620t620 n6621 n621 R=6.473e+01 
R6620t900 n6621 n901 R=4.886e+00 
R6620t939 n6621 n940 R=4.725e+01 
R6620t5425 n6621 n5426 R=3.126e+00 
R6620t6611 n6621 n6612 R=1.138e+01 
R6620t2042 n6621 n2043 R=7.495e+00 
R6621t3676 n6622 n3677 R=5.668e+00 
R6621t3228 n6622 n3229 R=4.064e+00 
R6621t3995 n6622 n3996 R=6.470e+00 
R6622t5947 n6623 n5948 R=2.361e+01 
R6622t6592 n6623 n6593 R=2.458e+00 
R6622t2038 n6623 n2039 R=2.914e+00 
R6623t3930 n6624 n3931 R=9.527e+00 
R6623t4876 n6624 n4877 R=1.082e+01 
R6623t3443 n6624 n3444 R=8.371e+00 
R6623t995 n6624 n996 R=3.481e+00 
R6623t2918 n6624 n2919 R=1.626e+01 
R6623t6147 n6624 n6148 R=1.232e+01 
R6624t2424 n6625 n2425 R=2.850e+00 
R6624t3112 n6625 n3113 R=5.336e+00 
R6624t2652 n6625 n2653 R=7.766e+00 
R6624t1368 n6625 n1369 R=4.208e+00 
R6625t1729 n6626 n1730 R=4.419e+01 
R6625t4181 n6626 n4182 R=2.403e+01 
R6625t1423 n6626 n1424 R=8.087e+00 
R6625t2238 n6626 n2239 R=5.827e+00 
R6626t5176 n6627 n5177 R=1.297e+01 
R6626t5318 n6627 n5319 R=1.337e+02 
R6626t5901 n6627 n5902 R=2.678e+00 
R6626t1162 n6627 n1163 R=1.599e+01 
R6626t242 n6627 n243 R=2.344e+00 
R6627t3309 n6628 n3310 R=5.094e+00 
R6627t140 n6628 n141 R=3.158e+01 
R6627t3740 n6628 n3741 R=4.570e+00 
R6627t765 n6628 n766 R=7.690e+00 
R6627t1808 n6628 n1809 R=9.445e+01 
R6628t208 n6629 n209 R=1.140e+01 
R6628t1460 n6629 n1461 R=5.746e+00 
R6628t5823 n6629 n5824 R=2.338e+01 
R6628t571 n6629 n572 R=2.298e+00 
R6628t4645 n6629 n4646 R=1.239e+01 
R6629t287 n6630 n288 R=5.299e+00 
R6629t3106 n6630 n3107 R=3.700e+00 
R6630t1532 n6631 n1533 R=4.045e+00 
R6630t4538 n6631 n4539 R=7.491e+00 
R6630t6383 n6631 n6384 R=5.616e+01 
R6630t4188 n6631 n4189 R=2.957e+00 
R6630t4484 n6631 n4485 R=2.971e+01 
R6630t2420 n6631 n2421 R=3.075e+01 
R6631t1511 n6632 n1512 R=6.272e+00 
R6631t4057 n6632 n4058 R=4.988e+00 
R6631t1456 n6632 n1457 R=2.146e+01 
R6631t1942 n6632 n1943 R=2.297e+01 
R6631t2348 n6632 n2349 R=8.940e+01 
R6632t117 n6633 n118 R=4.275e+00 
R6632t2346 n6633 n2347 R=1.255e+01 
R6632t5008 n6633 n5009 R=2.324e+02 
R6632t1461 n6633 n1462 R=3.292e+00 
R6632t2366 n6633 n2367 R=4.773e+00 
R6632t878 n6633 n879 R=1.763e+01 
R6633t2368 n6634 n2369 R=6.674e+00 
R6633t4751 n6634 n4752 R=3.270e+00 
R6633t5498 n6634 n5499 R=8.168e+00 
R6633t5592 n6634 n5593 R=5.797e+00 
R6634t5683 n6635 n5684 R=3.595e+00 
R6634t26 n6635 n27 R=4.256e+01 
R6634t819 n6635 n820 R=2.967e+00 
R6634t5908 n6635 n5909 R=6.425e+00 
R6635t944 n6636 n945 R=2.167e+00 
R6635t2707 n6636 n2708 R=1.051e+02 
R6635t131 n6636 n132 R=4.169e+00 
R6635t4412 n6636 n4413 R=6.411e+00 
R6635t3514 n6636 n3515 R=2.441e+02 
R6636t1838 n6637 n1839 R=2.666e+00 
R6636t6591 n6637 n6592 R=9.833e+01 
R6636t6248 n6637 n6249 R=3.639e+00 
R6636t1020 n6637 n1021 R=6.257e+00 
R6636t3743 n6637 n3744 R=2.089e+01 
R6636t2559 n6637 n2560 R=5.531e+01 
R6637t3302 n6638 n3303 R=3.774e+00 
R6637t6267 n6638 n6268 R=7.520e+00 
R6637t639 n6638 n640 R=2.107e+01 
R6637t5866 n6638 n5867 R=5.215e+00 
R6638t5423 n6639 n5424 R=1.874e+01 
R6638t5481 n6639 n5482 R=2.056e+01 
R6638t1369 n6639 n1370 R=7.006e+00 
R6638t5507 n6639 n5508 R=1.062e+02 
R6638t6301 n6639 n6302 R=2.868e+02 
R6639t6169 n6640 n6170 R=6.596e+00 
R6639t4153 n6640 n4154 R=3.624e+00 
R6639t2682 n6640 n2683 R=4.041e+00 
R6640t3868 n6641 n3869 R=3.923e+00 
R6640t4201 n6641 n4202 R=6.967e+00 
R6640t1770 n6641 n1771 R=7.011e+00 
R6641t3412 n6642 n3413 R=8.701e+00 
R6641t4885 n6642 n4886 R=1.537e+01 
R6641t3555 n6642 n3556 R=9.132e+00 
R6641t358 n6642 n359 R=4.259e+01 
R6641t671 n6642 n672 R=1.967e+01 
R6641t2487 n6642 n2488 R=6.894e+00 
R6641t6271 n6642 n6272 R=2.934e+00 
R6641t1052 n6642 n1053 R=1.173e+02 
R6641t1378 n6642 n1379 R=1.399e+02 
R6642t4614 n6643 n4615 R=7.836e+00 
R6642t1645 n6643 n1646 R=5.698e+00 
R6642t1812 n6643 n1813 R=3.869e+00 
R6642t3614 n6643 n3615 R=1.630e+02 
R6642t5506 n6643 n5507 R=2.948e+00 
R6642t2936 n6643 n2937 R=5.156e+01 
R6643t1418 n6644 n1419 R=1.316e+01 
R6643t4603 n6644 n4604 R=3.128e+00 
R6643t740 n6644 n741 R=1.993e+02 
R6644t5973 n6645 n5974 R=6.496e+00 
R6644t2399 n6645 n2400 R=1.619e+01 
R6644t4514 n6645 n4515 R=1.047e+01 
R6644t5350 n6645 n5351 R=1.263e+01 
R6644t4846 n6645 n4847 R=1.177e+01 
R6645t2689 n6646 n2690 R=3.077e+01 
R6645t5917 n6646 n5918 R=6.439e+00 
R6645t46 n6646 n47 R=2.056e+01 
R6645t4483 n6646 n4484 R=8.417e+00 
R6645t849 n6646 n850 R=3.168e+00 
R6647t3505 n6648 n3506 R=3.610e+00 
R6647t3776 n6648 n3777 R=5.050e+00 
R6648t1922 n6649 n1923 R=6.116e+00 
R6648t5817 n6649 n5818 R=1.143e+01 
R6648t4234 n6649 n4235 R=2.126e+01 
R6649t2538 n6650 n2539 R=6.117e+00 
R6649t5405 n6650 n5406 R=8.942e+00 
R6649t1195 n6650 n1196 R=2.347e+02 
R6649t1084 n6650 n1085 R=2.850e+01 
R6649t5483 n6650 n5484 R=5.606e+00 
R6649t2871 n6650 n2872 R=1.067e+01 
R6650t467 n6651 n468 R=5.815e+00 
R6650t213 n6651 n214 R=2.240e+01 
R6650t5968 n6651 n5969 R=1.006e+01 
R6650t2550 n6651 n2551 R=7.870e+00 
R6650t783 n6651 n784 R=1.492e+01 
R6650t244 n6651 n245 R=9.403e+01 
R6651t305 n6652 n306 R=1.170e+01 
R6651t5491 n6652 n5492 R=1.457e+01 
R6651t5469 n6652 n5470 R=1.442e+01 
R6651t4482 n6652 n4483 R=3.201e+01 
R6651t3531 n6652 n3532 R=1.492e+01 
R6652t2791 n6653 n2792 R=3.661e+00 
R6652t5335 n6653 n5336 R=6.090e+00 
R6652t3080 n6653 n3081 R=1.906e+00 
R6652t2762 n6653 n2763 R=5.978e+01 
R6653t5856 n6654 n5857 R=7.224e+00 
R6653t2028 n6654 n2029 R=1.929e+01 
R6653t6116 n6654 n6117 R=9.190e+00 
R6654t3900 n6655 n3901 R=1.935e+01 
R6654t4859 n6655 n4860 R=5.082e+00 
R6654t709 n6655 n710 R=4.015e+00 
R6654t977 n6655 n978 R=3.463e+00 
R6654t3397 n6655 n3398 R=1.374e+01 
R6655t991 n6656 n992 R=3.995e+00 
R6655t4730 n6656 n4731 R=4.094e+00 
R6655t6111 n6656 n6112 R=6.860e+00 
R6655t6000 n6656 n6001 R=1.051e+03 
R6656t1375 n6657 n1376 R=7.166e+00 
R6656t3928 n6657 n3929 R=2.924e+00 
R6656t5868 n6657 n5869 R=2.794e+00 
R6656t3656 n6657 n3657 R=1.871e+01 
R6657t1306 n6658 n1307 R=4.422e+00 
R6657t2663 n6658 n2664 R=1.395e+01 
R6657t337 n6658 n338 R=2.592e+00 
R6657t2326 n6658 n2327 R=3.423e+00 
R6658t919 n6659 n920 R=1.647e+00 
R6658t5936 n6659 n5937 R=3.872e+01 
R6658t1557 n6659 n1558 R=9.554e+00 
R6659t4908 n6660 n4909 R=6.093e+01 
R6659t3417 n6660 n3418 R=5.900e+00 
R6659t3190 n6660 n3191 R=6.588e+00 
R6659t2329 n6660 n2330 R=1.812e+01 
R6659t3673 n6660 n3674 R=4.285e+00 
R6660t1028 n6661 n1029 R=7.010e+00 
R6660t6192 n6661 n6193 R=6.369e+00 
R6660t5635 n6661 n5636 R=1.933e+01 
R6660t2443 n6661 n2444 R=1.023e+02 
R6660t1403 n6661 n1404 R=1.185e+02 
R6660t4227 n6661 n4228 R=1.185e+01 
R6660t1400 n6661 n1401 R=6.190e+00 
R6660t6180 n6661 n6181 R=6.020e+00 
R6661t1531 n6662 n1532 R=6.454e+00 
R6661t5493 n6662 n5494 R=3.188e+01 
R6661t5300 n6662 n5301 R=1.264e+01 
R6661t4406 n6662 n4407 R=8.317e+00 
R6661t2323 n6662 n2324 R=8.970e+00 
R6662t197 n6663 n198 R=2.799e+01 
R6662t4815 n6663 n4816 R=5.829e+00 
R6662t4555 n6663 n4556 R=1.295e+02 
R6662t6123 n6663 n6124 R=5.035e+00 
R6662t647 n6663 n648 R=6.400e+00 
R6663t2659 n6664 n2660 R=9.678e+00 
R6663t3653 n6664 n3654 R=6.110e+01 
R6663t5032 n6664 n5033 R=1.582e+00 
R6663t2188 n6664 n2189 R=1.072e+01 
R6663t1305 n6664 n1306 R=5.802e+00 
R6664t3357 n6665 n3358 R=7.997e+00 
R6664t4346 n6665 n4347 R=2.147e+01 
R6664t2279 n6665 n2280 R=8.899e+00 
R6664t4748 n6665 n4749 R=2.024e+01 
R6664t4024 n6665 n4025 R=3.317e+00 
R6665t1986 n6666 n1987 R=9.675e+00 
R6665t4697 n6666 n4698 R=1.201e+01 
R6665t3141 n6666 n3142 R=7.436e+00 
R6665t2925 n6666 n2926 R=3.556e+00 
R6666t78 n6667 n79 R=5.361e+00 
R6666t1097 n6667 n1098 R=5.580e+00 
R6666t1192 n6667 n1193 R=8.546e+00 
R6666t4585 n6667 n4586 R=7.399e+01 
R6666t5514 n6667 n5515 R=1.313e+01 
R6666t3393 n6667 n3394 R=2.137e+02 
R6666t4954 n6667 n4955 R=5.956e+00 
R6667t51 n6668 n52 R=3.787e+00 
R6667t367 n6668 n368 R=6.074e+00 
R6667t3409 n6668 n3410 R=1.955e+01 
R6668t1674 n6669 n1675 R=7.865e+00 
R6668t2913 n6669 n2914 R=1.176e+01 
R6668t5466 n6669 n5467 R=9.765e+00 
R6668t532 n6669 n533 R=5.446e+00 
R6668t5317 n6669 n5318 R=2.333e+01 
R6668t1569 n6669 n1570 R=2.205e+02 
R6668t3954 n6669 n3955 R=4.833e+00 
R6669t1970 n6670 n1971 R=1.126e+01 
R6669t58 n6670 n59 R=2.866e+00 
R6670t5172 n6671 n5173 R=8.110e+01 
R6670t3280 n6671 n3281 R=9.891e+00 
R6670t3121 n6671 n3122 R=1.647e+01 
R6671t1547 n6672 n1548 R=1.401e+01 
R6671t2764 n6672 n2765 R=3.614e+00 
R6672t6362 n6673 n6363 R=7.886e+00 
R6672t285 n6673 n286 R=1.013e+02 
R6672t4524 n6673 n4525 R=3.339e+00 
R6673t1450 n6674 n1451 R=3.736e+00 
R6673t5818 n6674 n5819 R=9.880e+00 
R6673t5699 n6674 n5700 R=4.189e+01 
R6673t1152 n6674 n1153 R=2.543e+01 
R6673t44 n6674 n45 R=3.596e+02 
R6674t1443 n6675 n1444 R=6.031e+00 
R6674t3956 n6675 n3957 R=4.750e+00 
R6674t2148 n6675 n2149 R=6.958e+00 
R6674t6122 n6675 n6123 R=2.820e+01 
R6674t2620 n6675 n2621 R=4.722e+01 
R6675t2810 n6676 n2811 R=2.343e+00 
R6675t417 n6676 n418 R=4.876e+00 
R6675t5056 n6676 n5057 R=6.156e+00 
R6676t2133 n6677 n2134 R=7.994e+00 
R6676t1865 n6677 n1866 R=5.094e+00 
R6677t666 n6678 n667 R=1.914e+01 
R6677t311 n6678 n312 R=2.212e+01 
R6677t5745 n6678 n5746 R=8.525e+00 
R6677t5284 n6678 n5285 R=3.454e+00 
R6678t3704 n6679 n3705 R=2.534e+02 
R6678t4652 n6679 n4653 R=4.339e+00 
R6678t1644 n6679 n1645 R=2.894e+00 
R6678t5390 n6679 n5391 R=2.301e+01 
R6678t5610 n6679 n5611 R=2.145e+00 
R6678t6172 n6679 n6173 R=5.597e+01 
R6679t365 n6680 n366 R=4.086e+00 
R6679t2441 n6680 n2442 R=3.038e+00 
R6679t6523 n6680 n6524 R=5.669e+00 
R6680t1404 n6681 n1405 R=1.021e+01 
R6680t2981 n6681 n2982 R=9.461e+00 
R6680t3639 n6681 n3640 R=7.608e+00 
R6681t1336 n6682 n1337 R=1.669e+00 
R6681t3444 n6682 n3445 R=6.492e+01 
R6681t2021 n6682 n2022 R=3.099e+00 
R6681t4840 n6682 n4841 R=7.127e+00 
R6681t5974 n6682 n5975 R=1.206e+01 
R6682t2876 n6683 n2877 R=6.667e+01 
R6682t5238 n6683 n5239 R=3.882e+00 
R6682t3611 n6683 n3612 R=6.429e+00 
R6683t202 n6684 n203 R=3.279e+00 
R6683t2647 n6684 n2648 R=8.222e+00 
R6683t3586 n6684 n3587 R=2.992e+00 
R6684t4731 n6685 n4732 R=8.229e+00 
R6684t52 n6685 n53 R=4.207e+00 
R6684t758 n6685 n759 R=1.009e+01 
R6685t225 n6686 n226 R=4.062e+00 
R6685t1261 n6686 n1262 R=8.439e+00 
R6685t5603 n6686 n5604 R=4.494e+00 
R6685t4249 n6686 n4250 R=7.093e+01 
R6686t408 n6687 n409 R=1.287e+01 
R6686t5412 n6687 n5413 R=2.428e+00 
R6686t5981 n6687 n5982 R=1.223e+01 
R6686t3195 n6687 n3196 R=3.262e+00 
R6687t6154 n6688 n6155 R=2.895e+00 
R6687t530 n6688 n531 R=1.444e+01 
R6687t1186 n6688 n1187 R=6.344e+00 
R6687t4301 n6688 n4302 R=5.744e+00 
R6688t1027 n6689 n1028 R=1.664e+00 
R6688t1756 n6689 n1757 R=8.035e+00 
R6688t2555 n6689 n2556 R=2.443e+01 
R6688t4615 n6689 n4616 R=3.719e+01 
R6689t3622 n6690 n3623 R=7.095e+01 
R6689t2363 n6690 n2364 R=3.386e+00 
R6689t5306 n6690 n5307 R=3.330e+00 
R6690t5852 n6691 n5853 R=2.325e+00 
R6691t3767 n6692 n3768 R=6.730e+00 
R6691t5442 n6692 n5443 R=4.731e+00 
R6691t5393 n6692 n5394 R=6.550e+00 
R6692t497 n6693 n498 R=3.639e+01 
R6692t5398 n6693 n5399 R=2.652e+00 
R6692t4640 n6693 n4641 R=4.212e+01 
R6693t579 n6694 n580 R=4.697e+01 
R6693t4624 n6694 n4625 R=5.951e+00 
R6693t5122 n6694 n5123 R=8.226e+00 
R6693t6371 n6694 n6372 R=1.414e+01 
R6693t6330 n6694 n6331 R=9.823e+00 
R6694t2687 n6695 n2688 R=2.562e+01 
R6694t1241 n6695 n1242 R=2.545e+01 
R6694t6273 n6695 n6274 R=4.990e+00 
R6695t2419 n6696 n2420 R=6.844e+00 
R6695t4440 n6696 n4441 R=4.309e+00 
R6695t1940 n6696 n1941 R=2.754e+00 
R6696t3804 n6697 n3805 R=2.047e+01 
R6696t3794 n6697 n3795 R=1.689e+01 
R6696t2839 n6697 n2840 R=2.587e+01 
R6697t3115 n6698 n3116 R=1.004e+01 
R6697t5946 n6698 n5947 R=3.438e+01 
R6697t3700 n6698 n3701 R=1.111e+01 
R6697t2027 n6698 n2028 R=2.176e+01 
R6697t3124 n6698 n3125 R=1.201e+01 
R6697t66 n6698 n67 R=6.098e+00 
R6698t1180 n6699 n1181 R=1.896e+01 
R6698t4618 n6699 n4619 R=5.303e+00 
R6698t2400 n6699 n2401 R=7.164e+00 
R6698t2991 n6699 n2992 R=6.671e+00 
R6698t3709 n6699 n3710 R=5.581e+00 
R6698t4808 n6699 n4809 R=1.354e+01 
R6699t4287 n6700 n4288 R=1.234e+02 
R6699t37 n6700 n38 R=1.796e+01 
R6700t1894 n6701 n1895 R=5.087e+00 
R6700t4541 n6701 n4542 R=3.674e+00 
R6700t6275 n6701 n6276 R=3.028e+00 
R6700t2729 n6701 n2730 R=7.155e+00 
R6701t985 n6702 n986 R=8.736e+01 
R6701t2007 n6702 n2008 R=1.526e+02 
R6701t733 n6702 n734 R=1.674e+01 
R6701t2016 n6702 n2017 R=2.697e+01 
R6702t23 n6703 n24 R=7.461e+00 
R6702t4749 n6703 n4750 R=6.588e+00 
R6702t1013 n6703 n1014 R=1.037e+01 
R6702t5226 n6703 n5227 R=1.536e+01 
R6702t6521 n6703 n6522 R=5.574e+00 
R6703t1048 n6704 n1049 R=3.142e+01 
R6703t6197 n6704 n6198 R=3.089e+00 
R6703t226 n6704 n227 R=1.564e+02 
R6703t168 n6704 n169 R=3.452e+00 
R6704t1959 n6705 n1960 R=4.017e+00 
R6704t4557 n6705 n4558 R=8.457e+00 
R6704t6097 n6705 n6098 R=5.300e+00 
R6705t6508 n6706 n6509 R=2.371e+01 
R6705t3722 n6706 n3723 R=5.600e+00 
R6705t924 n6706 n925 R=1.464e+02 
R6705t694 n6706 n695 R=1.069e+01 
R6706t3312 n6707 n3313 R=1.584e+01 
R6706t4414 n6707 n4415 R=4.178e+00 
R6707t4767 n6708 n4768 R=2.491e+00 
R6707t5146 n6708 n5147 R=4.126e+00 
R6707t2705 n6708 n2706 R=6.550e+00 
R6707t2567 n6708 n2568 R=3.103e+01 
R6708t1073 n6709 n1074 R=6.653e+00 
R6708t2404 n6709 n2405 R=6.247e+00 
R6708t419 n6709 n420 R=2.916e+01 
R6709t670 n6710 n671 R=9.441e+00 
R6709t5237 n6710 n5238 R=5.024e+00 
R6709t2723 n6710 n2724 R=9.512e+00 
R6709t2355 n6710 n2356 R=4.313e+00 
R6710t6344 n6711 n6345 R=1.463e+02 
R6710t6155 n6711 n6156 R=4.371e+00 
R6710t1897 n6711 n1898 R=3.107e+01 
R6710t4184 n6711 n4185 R=2.713e+02 
R6710t3191 n6711 n3192 R=3.521e+00 
R6710t2780 n6711 n2781 R=1.482e+01 
R6710t776 n6711 n777 R=1.111e+01 
R6711t5620 n6712 n5621 R=1.032e+01 
R6711t6404 n6712 n6405 R=8.868e+00 
R6711t5956 n6712 n5957 R=4.052e+00 
R6711t4288 n6712 n4289 R=2.303e+00 
R6712t369 n6713 n370 R=4.196e+00 
R6712t6127 n6713 n6128 R=4.585e+00 
R6712t1945 n6713 n1946 R=4.808e+00 
R6712t2380 n6713 n2381 R=9.312e+00 
R6712t4279 n6713 n4280 R=1.069e+01 
R6712t5280 n6713 n5281 R=2.124e+02 
R6713t2038 n6714 n2039 R=1.369e+01 
R6713t6622 n6714 n6623 R=4.188e+01 
R6713t6592 n6714 n6593 R=4.302e+02 
R6713t1408 n6714 n1409 R=1.402e+01 
R6714t5017 n6715 n5018 R=2.194e+00 
R6714t4193 n6715 n4194 R=1.808e+01 
R6714t4236 n6715 n4237 R=5.824e+00 
R6714t3684 n6715 n3685 R=4.440e+00 
R6715t1939 n6716 n1940 R=9.734e+00 
R6715t2873 n6716 n2874 R=1.546e+01 
R6715t2358 n6716 n2359 R=4.128e+00 
R6715t2764 n6716 n2765 R=9.188e+00 
R6715t6671 n6716 n6672 R=2.616e+01 
R6715t1547 n6716 n1548 R=1.439e+01 
R6715t3327 n6716 n3328 R=5.603e+00 
R6716t546 n6717 n547 R=7.245e+00 
R6716t3281 n6717 n3282 R=3.609e+00 
R6716t3144 n6717 n3145 R=4.202e+00 
R6717t25 n6718 n26 R=3.257e+01 
R6717t5191 n6718 n5192 R=4.095e+00 
R6718t3621 n6719 n3622 R=4.525e+01 
R6718t6643 n6719 n6644 R=9.002e+00 
R6718t1418 n6719 n1419 R=9.440e+00 
R6718t697 n6719 n698 R=3.683e+00 
R6719t4125 n6720 n4126 R=1.770e+01 
R6719t3862 n6720 n3863 R=2.278e+00 
R6719t2026 n6720 n2027 R=4.021e+01 
R6719t5920 n6720 n5921 R=2.473e+00 
R6720t6081 n6721 n6082 R=9.283e+00 
R6720t5143 n6721 n5144 R=1.798e+01 
R6720t963 n6721 n964 R=2.904e+00 
R6721t4072 n6722 n4073 R=1.003e+02 
R6721t4579 n6722 n4580 R=3.431e+00 
R6721t2641 n6722 n2642 R=2.705e+02 
R6721t1041 n6722 n1042 R=3.072e+00 
R6722t1678 n6723 n1679 R=7.528e+00 
R6722t4290 n6723 n4291 R=1.845e+01 
R6722t4487 n6723 n4488 R=3.095e+00 
R6722t3814 n6723 n3815 R=1.710e+01 
R6723t5281 n6724 n5282 R=3.210e+01 
R6723t143 n6724 n144 R=8.208e+00 
R6723t121 n6724 n122 R=3.522e+00 
R6723t1784 n6724 n1785 R=9.398e+00 
R6724t162 n6725 n163 R=3.018e+00 
R6724t1772 n6725 n1773 R=2.328e+01 
R6724t736 n6725 n737 R=4.640e+00 
R6725t2792 n6726 n2793 R=2.076e+00 
R6725t5352 n6726 n5353 R=1.729e+00 
R6725t1599 n6726 n1600 R=7.991e+00 
R6726t5626 n6727 n5627 R=2.206e+00 
R6726t2029 n6727 n2030 R=4.891e+00 
R6726t2798 n6727 n2799 R=1.272e+01 
R6726t774 n6727 n775 R=1.874e+01 
R6726t4889 n6727 n4890 R=1.616e+01 
R6727t5637 n6728 n5638 R=2.107e+00 
R6727t4477 n6728 n4478 R=2.451e+01 
R6727t189 n6728 n190 R=4.323e+00 
R6728t1252 n6729 n1253 R=5.578e+00 
R6728t5883 n6729 n5884 R=2.977e+00 
R6728t2139 n6729 n2140 R=1.196e+01 
R6728t1943 n6729 n1944 R=3.147e+01 
R6728t6112 n6729 n6113 R=4.834e+00 
R6729t3536 n6730 n3537 R=3.098e+00 
R6729t560 n6730 n561 R=9.792e+00 
R6729t4748 n6730 n4749 R=7.887e+00 
R6730t754 n6731 n755 R=3.138e+01 
R6730t1164 n6731 n1165 R=3.183e+01 
R6730t6253 n6731 n6254 R=3.421e+00 
R6730t412 n6731 n413 R=9.755e+01 
R6730t641 n6731 n642 R=3.397e+01 
R6731t5538 n6732 n5539 R=6.180e+00 
R6731t667 n6732 n668 R=6.945e+00 
R6731t5539 n6732 n5540 R=6.751e+00 
R6731t3142 n6732 n3143 R=1.463e+01 
R6732t494 n6733 n495 R=1.537e+01 
R6732t6187 n6733 n6188 R=2.722e+00 
R6732t2488 n6733 n2489 R=6.630e+00 
R6732t5133 n6733 n5134 R=8.236e+00 
R6733t1657 n6734 n1658 R=3.295e+00 
R6733t1676 n6734 n1677 R=1.430e+01 
R6733t1162 n6734 n1163 R=1.684e+01 
R6733t3194 n6734 n3195 R=1.763e+01 
R6733t4052 n6734 n4053 R=2.460e+01 
R6733t1123 n6734 n1124 R=1.939e+01 
R6734t1377 n6735 n1378 R=6.720e+00 
R6734t4358 n6735 n4359 R=1.260e+01 
R6734t2211 n6735 n2212 R=1.256e+01 
R6735t2693 n6736 n2694 R=1.261e+00 
R6735t948 n6736 n949 R=8.567e+00 
R6735t437 n6736 n438 R=2.464e+00 
R6736t770 n6737 n771 R=2.098e+01 
R6736t5027 n6737 n5028 R=3.927e+00 
R6736t1163 n6737 n1164 R=3.016e+00 
R6736t2335 n6737 n2336 R=6.188e+00 
R6737t583 n6738 n584 R=4.134e+00 
R6737t857 n6738 n858 R=3.344e+00 
R6737t3785 n6738 n3786 R=5.008e+00 
R6738t625 n6739 n626 R=1.898e+01 
R6738t6526 n6739 n6527 R=3.934e+00 
R6738t5036 n6739 n5037 R=7.935e+00 
R6739t3179 n6740 n3180 R=2.896e+01 
R6739t5677 n6740 n5678 R=2.917e+00 
R6739t2749 n6740 n2750 R=2.735e+00 
R6739t3497 n6740 n3498 R=3.300e+00 
R6740t6096 n6741 n6097 R=5.235e+00 
R6740t170 n6741 n171 R=1.010e+01 
R6740t2227 n6741 n2228 R=5.093e+00 
R6741t6362 n6742 n6363 R=1.606e+01 
R6741t6672 n6742 n6673 R=1.769e+00 
R6741t285 n6742 n286 R=8.574e+00 
R6742t5699 n6743 n5700 R=1.875e+01 
R6742t4114 n6743 n4115 R=3.693e+00 
R6742t1144 n6743 n1145 R=7.160e+00 
R6743t5332 n6744 n5333 R=1.146e+01 
R6743t6108 n6744 n6109 R=1.640e+00 
R6743t2369 n6744 n2370 R=3.001e+00 
R6743t5809 n6744 n5810 R=7.034e+00 
R6744t2252 n6745 n2253 R=1.907e+01 
R6744t6349 n6745 n6350 R=1.383e+01 
R6745t5508 n6746 n5509 R=8.491e+00 
R6745t518 n6746 n519 R=2.700e+00 
R6746t3439 n6747 n3440 R=2.166e+01 
R6746t4503 n6747 n4504 R=1.582e+01 
R6746t2374 n6747 n2375 R=1.039e+01 
R6746t3396 n6747 n3397 R=1.471e+01 
R6746t1775 n6747 n1776 R=5.159e+00 
R6747t2020 n6748 n2021 R=4.826e+00 
R6747t6170 n6748 n6171 R=3.916e+00 
R6748t2388 n6749 n2389 R=6.725e+00 
R6748t6149 n6749 n6150 R=5.515e+00 
R6748t6162 n6749 n6163 R=6.354e+01 
R6748t6526 n6749 n6527 R=1.403e+02 
R6748t625 n6749 n626 R=5.789e+00 
R6748t5156 n6749 n5157 R=9.818e+01 
R6748t818 n6749 n819 R=9.270e+01 
R6749t4098 n6750 n4099 R=6.419e+00 
R6749t5288 n6750 n5289 R=5.493e+00 
R6749t2631 n6750 n2632 R=1.188e+01 
R6749t2432 n6750 n2433 R=2.455e+01 
R6750t1624 n6751 n1625 R=7.910e+01 
R6750t1863 n6751 n1864 R=1.020e+01 
R6750t223 n6751 n224 R=2.978e+00 
R6750t3817 n6751 n3818 R=5.858e+01 
R6750t4292 n6751 n4293 R=6.745e+00 
R6750t5052 n6751 n5053 R=3.354e+01 
R6750t4319 n6751 n4320 R=3.094e+00 
R6751t2876 n6752 n2877 R=6.323e+01 
R6751t5238 n6752 n5239 R=4.280e+01 
R6751t4276 n6752 n4277 R=7.920e+00 
R6751t2629 n6752 n2630 R=3.770e+00 
R6752t1978 n6753 n1979 R=1.494e+01 
R6752t3028 n6753 n3029 R=2.893e+00 
R6752t2317 n6753 n2318 R=5.590e+00 
R6753t812 n6754 n813 R=5.888e+00 
R6753t5608 n6754 n5609 R=6.028e+00 
R6753t3279 n6754 n3280 R=3.234e+01 
R6753t928 n6754 n929 R=4.387e+00 
R6753t5973 n6754 n5974 R=1.349e+01 
R6754t6204 n6755 n6205 R=6.439e+00 
R6754t5219 n6755 n5220 R=4.366e+00 
R6754t2376 n6755 n2377 R=3.034e+01 
R6754t3574 n6755 n3575 R=5.156e+01 
R6754t3744 n6755 n3745 R=6.606e+00 
R6755t3166 n6756 n3167 R=4.328e+01 
R6755t3728 n6756 n3729 R=1.858e+00 
R6755t461 n6756 n462 R=1.455e+01 
R6755t6043 n6756 n6044 R=2.141e+00 
R6755t6619 n6756 n6620 R=9.241e+00 
R6756t5659 n6757 n5660 R=5.706e+00 
R6756t6434 n6757 n6435 R=6.353e+00 
R6756t2812 n6757 n2813 R=9.216e+00 
R6756t4197 n6757 n4198 R=6.205e+00 
R6756t4169 n6757 n4170 R=1.087e+01 
R6757t1324 n6758 n1325 R=1.919e+01 
R6757t2501 n6758 n2502 R=2.441e+00 
R6757t4400 n6758 n4401 R=6.498e+00 
R6757t6035 n6758 n6036 R=5.782e+00 
R6757t3339 n6758 n3340 R=2.736e+01 
R6757t5046 n6758 n5047 R=1.930e+01 
R6757t4469 n6758 n4470 R=1.674e+01 
R6758t1536 n6759 n1537 R=2.094e+01 
R6758t1549 n6759 n1550 R=7.644e+00 
R6758t3663 n6759 n3664 R=3.461e+01 
R6758t640 n6759 n641 R=2.852e+00 
R6758t2184 n6759 n2185 R=2.595e+01 
R6758t5622 n6759 n5623 R=5.511e+00 
R6759t2107 n6760 n2108 R=7.242e+00 
R6759t639 n6760 n640 R=1.489e+02 
R6759t291 n6760 n292 R=9.601e+00 
R6759t3645 n6760 n3646 R=2.298e+00 
R6760t640 n6761 n641 R=1.155e+01 
R6760t6758 n6761 n6759 R=5.076e+01 
R6760t2184 n6761 n2185 R=2.229e+00 
R6760t3603 n6761 n3604 R=5.124e+02 
R6760t5340 n6761 n5341 R=2.863e+00 
R6761t5090 n6762 n5091 R=6.005e+01 
R6761t3905 n6762 n3906 R=3.231e+00 
R6761t716 n6762 n717 R=5.349e+00 
R6762t3495 n6763 n3496 R=1.026e+01 
R6762t5467 n6763 n5468 R=4.214e+00 
R6762t1331 n6763 n1332 R=5.792e+00 
R6762t4023 n6763 n4024 R=2.593e+00 
R6763t224 n6764 n225 R=9.149e+00 
R6763t2511 n6764 n2512 R=2.136e+01 
R6763t3358 n6764 n3359 R=1.397e+01 
R6763t1402 n6764 n1403 R=5.910e+00 
R6764t560 n6765 n561 R=2.342e+01 
R6764t3536 n6765 n3537 R=3.431e+00 
R6764t2154 n6765 n2155 R=1.224e+01 
R6764t1620 n6765 n1621 R=3.449e+00 
R6765t1143 n6766 n1144 R=2.310e+00 
R6765t4317 n6766 n4318 R=6.211e+00 
R6765t4010 n6766 n4011 R=1.527e+01 
R6765t1023 n6766 n1024 R=2.580e+00 
R6766t4531 n6767 n4532 R=1.058e+01 
R6766t2225 n6767 n2226 R=8.366e+00 
R6766t5714 n6767 n5715 R=4.620e+00 
R6766t2205 n6767 n2206 R=1.060e+01 
R6767t4968 n6768 n4969 R=5.932e+01 
R6767t157 n6768 n158 R=2.339e+01 
R6767t451 n6768 n452 R=2.768e+02 
R6767t5601 n6768 n5602 R=7.278e+00 
R6767t6328 n6768 n6329 R=2.001e+02 
R6767t2512 n6768 n2513 R=1.453e+02 
R6768t6723 n6769 n6724 R=6.283e+01 
R6768t4414 n6769 n4415 R=4.723e+00 
R6768t4863 n6769 n4864 R=7.170e+01 
R6768t4005 n6769 n4006 R=1.020e+01 
R6768t2784 n6769 n2785 R=4.125e+00 
R6768t121 n6769 n122 R=1.588e+01 
R6769t2328 n6770 n2329 R=5.729e+01 
R6769t5803 n6770 n5804 R=1.283e+01 
R6769t2551 n6770 n2552 R=2.430e+02 
R6769t6530 n6770 n6531 R=7.829e+00 
R6769t1663 n6770 n1664 R=4.552e+00 
R6769t6582 n6770 n6583 R=9.127e+00 
R6770t1400 n6771 n1401 R=9.932e+00 
R6770t1583 n6771 n1584 R=9.636e+00 
R6770t3484 n6771 n3485 R=3.075e+00 
R6770t661 n6771 n662 R=2.922e+01 
R6770t798 n6771 n799 R=6.693e+00 
R6770t1829 n6771 n1830 R=1.120e+01 
R6771t2284 n6772 n2285 R=3.150e+02 
R6771t3436 n6772 n3437 R=1.799e+00 
R6771t5099 n6772 n5100 R=9.292e+01 
R6771t5732 n6772 n5733 R=2.542e+00 
R6771t3630 n6772 n3631 R=4.410e+00 
R6771t2203 n6772 n2204 R=9.286e+02 
R6771t340 n6772 n341 R=9.066e+00 
R6772t3830 n6773 n3831 R=1.506e+01 
R6772t4420 n6773 n4421 R=8.498e+01 
R6772t956 n6773 n957 R=2.114e+01 
R6772t3001 n6773 n3002 R=6.495e+00 
R6772t2662 n6773 n2663 R=5.899e+01 
R6772t304 n6773 n305 R=3.105e+00 
R6773t200 n6774 n201 R=4.320e+00 
R6773t875 n6774 n876 R=1.375e+01 
R6773t2353 n6774 n2354 R=6.166e+00 
R6773t3100 n6774 n3101 R=4.017e+01 
R6773t3637 n6774 n3638 R=3.401e+00 
R6774t228 n6775 n229 R=3.004e+01 
R6774t4344 n6775 n4345 R=8.884e+01 
R6774t6431 n6775 n6432 R=4.886e+00 
R6774t5254 n6775 n5255 R=4.471e+01 
R6774t5646 n6775 n5647 R=5.571e+00 
R6774t1915 n6775 n1916 R=3.916e+01 
R6775t2157 n6776 n2158 R=2.945e+00 
R6775t6080 n6776 n6081 R=6.483e+00 
R6775t3381 n6776 n3382 R=3.251e+00 
R6775t5986 n6776 n5987 R=6.744e+01 
R6775t938 n6776 n939 R=1.345e+01 
R6776t1290 n6777 n1291 R=1.639e+02 
R6776t3037 n6777 n3038 R=3.531e+00 
R6776t3245 n6777 n3246 R=7.781e+01 
R6776t1665 n6777 n1666 R=1.043e+01 
R6776t4419 n6777 n4420 R=1.036e+01 
R6776t192 n6777 n193 R=3.234e+00 
R6777t3067 n6778 n3068 R=1.357e+01 
R6777t1793 n6778 n1794 R=3.744e+00 
R6777t126 n6778 n127 R=5.256e+00 
R6777t3695 n6778 n3696 R=9.214e+00 
R6777t778 n6778 n779 R=1.005e+01 
R6778t3012 n6779 n3013 R=1.013e+01 
R6778t3750 n6779 n3751 R=1.249e+01 
R6778t5543 n6779 n5544 R=1.263e+01 
R6778t6282 n6779 n6283 R=2.768e+01 
R6778t3024 n6779 n3025 R=8.881e+00 
R6778t2648 n6779 n2649 R=7.708e+00 
R6779t1426 n6780 n1427 R=5.133e+00 
R6779t6381 n6780 n6382 R=1.564e+01 
R6779t866 n6780 n867 R=9.744e+00 
R6779t3105 n6780 n3106 R=3.203e+01 
R6779t845 n6780 n846 R=1.735e+01 
R6779t753 n6780 n754 R=5.352e+01 
R6779t1565 n6780 n1566 R=1.448e+01 
R6779t1361 n6780 n1362 R=5.008e+00 
R6780t2285 n6781 n2286 R=6.064e+01 
R6780t449 n6781 n450 R=6.358e+00 
R6780t5157 n6781 n5158 R=4.319e+00 
R6780t4911 n6781 n4912 R=9.137e+00 
R6781t5953 n6782 n5954 R=2.816e+00 
R6781t5859 n6782 n5860 R=4.052e+00 
R6781t4512 n6782 n4513 R=6.383e+00 
R6782t4061 n6783 n4062 R=4.397e+00 
R6782t1262 n6783 n1263 R=8.800e+02 
R6783t1343 n6784 n1344 R=2.179e+01 
R6783t3780 n6784 n3781 R=9.227e+00 
R6783t6693 n6784 n6694 R=8.301e+00 
R6783t5122 n6784 n5123 R=7.078e+00 
R6783t2937 n6784 n2938 R=4.708e+00 
R6784t1733 n6785 n1734 R=3.956e+00 
R6784t6221 n6785 n6222 R=3.380e+00 
R6784t4835 n6785 n4836 R=7.283e+00 
R6784t1054 n6785 n1055 R=4.712e+00 
R6785t2121 n6786 n2122 R=4.270e+00 
R6785t2522 n6786 n2523 R=6.632e+00 
R6785t5360 n6786 n5361 R=8.975e+00 
R6786t3893 n6787 n3894 R=5.688e+00 
R6786t4507 n6787 n4508 R=1.175e+01 
R6787t2481 n6788 n2482 R=7.667e+00 
R6787t4889 n6788 n4890 R=2.179e+00 
R6787t6726 n6788 n6727 R=3.845e+01 
R6788t244 n6789 n245 R=2.797e+01 
R6788t3857 n6789 n3858 R=4.753e+01 
R6788t4973 n6789 n4974 R=1.715e+01 
R6788t6279 n6789 n6280 R=1.443e+03 
R6789t2425 n6790 n2426 R=1.080e+01 
R6789t3999 n6790 n4000 R=1.189e+01 
R6789t2989 n6790 n2990 R=2.191e+01 
R6789t3790 n6790 n3791 R=5.842e+00 
R6789t2196 n6790 n2197 R=9.057e+00 
R6789t4769 n6790 n4770 R=1.691e+01 
R6790t1538 n6791 n1539 R=1.409e+01 
R6790t2421 n6791 n2422 R=9.100e+00 
R6790t5186 n6791 n5187 R=9.091e+00 
R6790t3247 n6791 n3248 R=1.034e+01 
R6790t668 n6791 n669 R=2.926e+00 
R6791t854 n6792 n855 R=1.335e+02 
R6791t2691 n6792 n2692 R=3.027e+00 
R6791t4245 n6792 n4246 R=8.213e+01 
R6791t751 n6792 n752 R=7.918e+01 
R6791t5023 n6792 n5024 R=3.449e+00 
R6791t519 n6792 n520 R=3.534e+01 
R6791t3318 n6792 n3319 R=6.743e+00 
R6791t2504 n6792 n2505 R=3.949e+01 
R6792t2530 n6793 n2531 R=1.661e+00 
R6792t233 n6793 n234 R=1.855e+01 
R6793t4375 n6794 n4376 R=9.336e+01 
R6793t5993 n6794 n5994 R=4.178e+00 
R6793t2594 n6794 n2595 R=1.240e+01 
R6793t2347 n6794 n2348 R=8.165e+00 
R6794t616 n6795 n617 R=5.687e+00 
R6794t5066 n6795 n5067 R=3.919e+00 
R6794t1219 n6795 n1220 R=2.901e+00 
R6795t5791 n6796 n5792 R=3.748e+00 
R6795t3914 n6796 n3915 R=1.179e+02 
R6795t5030 n6796 n5031 R=3.626e+00 
R6796t5191 n6797 n5192 R=2.078e+01 
R6796t6717 n6797 n6718 R=7.963e+00 
R6796t3462 n6797 n3463 R=2.139e+00 
R6796t6278 n6797 n6279 R=1.963e+01 
R6797t5289 n6798 n5290 R=6.097e+00 
R6797t4220 n6798 n4221 R=5.555e+00 
R6797t5619 n6798 n5620 R=2.515e+00 
R6797t6389 n6798 n6390 R=3.649e+02 
R6798t2998 n6799 n2999 R=1.839e+01 
R6799t5547 n6800 n5548 R=2.493e+00 
R6799t4095 n6800 n4096 R=1.493e+01 
R6799t5940 n6800 n5941 R=2.776e+00 
R6800t582 n6801 n583 R=4.695e+00 
R6800t1016 n6801 n1017 R=4.945e+00 
R6800t389 n6801 n390 R=2.664e+01 
R6801t160 n6802 n161 R=2.154e+01 
R6801t1236 n6802 n1237 R=1.182e+01 
R6801t5675 n6802 n5676 R=4.185e+00 
R6801t1611 n6802 n1612 R=5.234e+00 
R6801t5218 n6802 n5219 R=2.504e+00 
R6801t4524 n6802 n4525 R=4.808e+01 
R6802t1769 n6803 n1770 R=2.896e+01 
R6802t5076 n6803 n5077 R=1.526e+00 
R6802t3456 n6803 n3457 R=2.951e+01 
R6802t1872 n6803 n1873 R=1.780e+02 
R6802t3037 n6803 n3038 R=2.124e+01 
R6802t1290 n6803 n1291 R=4.140e+00 
R6802t1706 n6803 n1707 R=1.788e+01 
R6803t5254 n6804 n5255 R=1.089e+01 
R6803t375 n6804 n376 R=2.119e+00 
R6803t1055 n6804 n1056 R=2.554e+01 
R6803t2078 n6804 n2079 R=3.120e+01 
R6803t1915 n6804 n1916 R=8.052e+00 
R6804t459 n6805 n460 R=2.339e+01 
R6804t5489 n6805 n5490 R=5.137e+00 
R6804t2660 n6805 n2661 R=3.381e+00 
R6804t15 n6805 n16 R=2.957e+01 
R6804t5564 n6805 n5565 R=4.792e+01 
R6804t1975 n6805 n1976 R=2.961e+00 
R6805t3253 n6806 n3254 R=1.067e+01 
R6805t963 n6806 n964 R=5.702e+00 
R6805t4278 n6806 n4279 R=9.774e+00 
R6805t3441 n6806 n3442 R=4.251e+01 
R6805t4250 n6806 n4251 R=1.079e+01 
R6806t1815 n6807 n1816 R=6.800e+00 
R6806t3535 n6807 n3536 R=3.192e+01 
R6807t5724 n6808 n5725 R=4.766e+00 
R6807t3853 n6808 n3854 R=7.619e+00 
R6807t2319 n6808 n2320 R=1.783e+01 
R6808t2105 n6809 n2106 R=2.008e+01 
R6808t3803 n6809 n3804 R=5.326e+00 
R6808t3175 n6809 n3176 R=5.589e+01 
R6808t1537 n6809 n1538 R=4.819e+00 
R6808t6519 n6809 n6520 R=4.761e+01 
R6808t1876 n6809 n1877 R=1.641e+01 
R6808t1903 n6809 n1904 R=6.863e+00 
R6809t1615 n6810 n1616 R=3.757e+00 
R6809t5204 n6810 n5205 R=1.019e+01 
R6809t2172 n6810 n2173 R=3.733e+01 
R6809t3877 n6810 n3878 R=2.248e+00 
R6810t3733 n6811 n3734 R=1.206e+01 
R6810t1012 n6811 n1013 R=2.024e+00 
R6810t2716 n6811 n2717 R=3.688e+02 
R6810t3295 n6811 n3296 R=2.452e+01 
R6810t1860 n6811 n1861 R=3.817e+00 
R6811t3197 n6812 n3198 R=8.203e+00 
R6811t5714 n6812 n5715 R=6.340e+00 
R6811t2205 n6812 n2206 R=3.704e+00 
R6811t3094 n6812 n3095 R=3.529e+01 
R6811t2828 n6812 n2829 R=1.203e+01 
R6811t5245 n6812 n5246 R=7.028e+00 
R6812t3753 n6813 n3754 R=1.583e+03 
R6812t1748 n6813 n1749 R=4.294e+01 
R6812t1454 n6813 n1455 R=2.558e+01 
R6812t1067 n6813 n1068 R=6.350e+01 
R6813t2551 n6814 n2552 R=2.242e+01 
R6813t6545 n6814 n6546 R=7.945e+00 
R6813t163 n6814 n164 R=5.334e+00 
R6813t6128 n6814 n6129 R=1.567e+01 
R6813t2013 n6814 n2014 R=8.951e+00 
R6814t2995 n6815 n2996 R=3.237e+01 
R6814t5182 n6815 n5183 R=6.562e+00 
R6814t2597 n6815 n2598 R=4.769e+00 
R6814t5879 n6815 n5880 R=6.380e+00 
R6815t763 n6816 n764 R=3.620e+00 
R6815t1446 n6816 n1447 R=7.318e+00 
R6815t659 n6816 n660 R=2.302e+01 
R6815t3010 n6816 n3011 R=3.217e+00 
R6816t1121 n6817 n1122 R=9.607e+00 
R6816t6587 n6817 n6588 R=5.552e+00 
R6816t2915 n6817 n2916 R=2.427e+02 
R6816t5369 n6817 n5370 R=3.535e+00 
R6817t2594 n6818 n2595 R=4.257e+00 
R6817t5625 n6818 n5626 R=6.653e+00 
R6817t4375 n6818 n4376 R=3.172e+01 
R6817t3958 n6818 n3959 R=2.231e+00 
R6818t374 n6819 n375 R=2.685e+00 
R6818t6501 n6819 n6502 R=2.765e+00 
R6818t5114 n6819 n5115 R=1.401e+01 
R6819t4311 n6820 n4312 R=4.102e+00 
R6819t5102 n6820 n5103 R=8.338e+00 
R6819t780 n6820 n781 R=3.001e+01 
R6819t4810 n6820 n4811 R=2.174e+00 
R6819t1821 n6820 n1822 R=1.583e+01 
R6820t644 n6821 n645 R=2.948e+00 
R6820t1635 n6821 n1636 R=1.202e+01 
R6820t5845 n6821 n5846 R=5.874e+00 
R6820t2475 n6821 n2476 R=4.412e+00 
R6820t5682 n6821 n5683 R=1.049e+01 
R6821t3401 n6822 n3402 R=3.415e+00 
R6821t5976 n6822 n5977 R=9.344e+00 
R6821t4526 n6822 n4527 R=6.744e+00 
R6821t1999 n6822 n2000 R=1.502e+01 
R6821t5743 n6822 n5744 R=6.546e+00 
R6822t2020 n6823 n2021 R=3.993e+00 
R6822t6747 n6823 n6748 R=3.409e+00 
R6823t1846 n6824 n1847 R=6.463e+00 
R6823t3869 n6824 n3870 R=1.747e+01 
R6823t2568 n6824 n2569 R=1.309e+01 
R6823t1104 n6824 n1105 R=7.308e+00 
R6823t4930 n6824 n4931 R=1.094e+01 
R6824t298 n6825 n299 R=8.088e+00 
R6824t4383 n6825 n4384 R=2.126e+01 
R6824t5638 n6825 n5639 R=1.083e+01 
R6824t1059 n6825 n1060 R=3.545e+00 
R6824t4738 n6825 n4739 R=7.368e+00 
R6825t3258 n6826 n3259 R=8.775e+00 
R6825t5250 n6826 n5251 R=6.428e+00 
R6825t4152 n6826 n4153 R=9.160e+00 
R6825t2375 n6826 n2376 R=7.614e+00 
R6825t4165 n6826 n4166 R=4.176e+01 
R6826t1418 n6827 n1419 R=8.369e+00 
R6826t6643 n6827 n6644 R=5.485e+00 
R6826t740 n6827 n741 R=3.913e+00 
R6826t633 n6827 n634 R=4.337e+00 
R6827t10 n6828 n11 R=1.804e+01 
R6827t92 n6828 n93 R=2.766e+00 
R6827t4780 n6828 n4781 R=9.827e+00 
R6828t1371 n6829 n1372 R=3.800e+00 
R6828t4348 n6829 n4349 R=5.473e+00 
R6828t4267 n6829 n4268 R=6.830e+00 
R6828t2110 n6829 n2111 R=4.067e+01 
R6829t5107 n6830 n5108 R=4.306e+00 
R6829t6088 n6830 n6089 R=2.665e+01 
R6829t6544 n6830 n6545 R=1.046e+01 
R6830t1257 n6831 n1258 R=7.007e+00 
R6830t5109 n6831 n5110 R=1.312e+01 
R6830t5941 n6831 n5942 R=2.534e+00 
R6830t313 n6831 n314 R=7.700e+00 
R6830t3832 n6831 n3833 R=5.350e+00 
R6831t632 n6832 n633 R=4.021e+01 
R6831t2865 n6832 n2866 R=2.634e+00 
R6832t2862 n6833 n2863 R=2.656e+00 
R6832t3334 n6833 n3335 R=8.442e+00 
R6832t5598 n6833 n5599 R=1.510e+02 
R6832t5256 n6833 n5257 R=6.585e+00 
R6833t44 n6834 n45 R=8.931e+00 
R6833t4054 n6834 n4055 R=2.283e+00 
R6833t3352 n6834 n3353 R=9.047e+00 
R6833t6402 n6834 n6403 R=1.876e+00 
R6834t6731 n6835 n6732 R=2.680e+00 
R6834t3142 n6835 n3143 R=3.469e+01 
R6834t2204 n6835 n2205 R=6.402e+00 
R6834t1417 n6835 n1418 R=4.073e+00 
R6834t6297 n6835 n6298 R=1.923e+01 
R6835t5116 n6836 n5117 R=4.924e+00 
R6835t2618 n6836 n2619 R=5.142e+00 
R6835t5257 n6836 n5258 R=1.048e+01 
R6835t5888 n6836 n5889 R=1.061e+01 
R6836t5689 n6837 n5690 R=1.158e+01 
R6836t469 n6837 n470 R=1.127e+01 
R6836t3419 n6837 n3420 R=4.264e+00 
R6836t3788 n6837 n3789 R=1.851e+01 
R6836t535 n6837 n536 R=2.214e+01 
R6837t3559 n6838 n3560 R=3.496e+00 
R6837t5998 n6838 n5999 R=5.530e+00 
R6837t2893 n6838 n2894 R=5.992e+00 
R6837t2861 n6838 n2862 R=5.241e+00 
R6838t2181 n6839 n2182 R=2.279e+01 
R6838t2492 n6839 n2493 R=4.595e+00 
R6839t423 n6840 n424 R=8.405e+00 
R6839t1360 n6840 n1361 R=4.707e+00 
R6839t1441 n6840 n1442 R=1.089e+02 
R6839t1427 n6840 n1428 R=1.026e+01 
R6839t4556 n6840 n4557 R=1.575e+01 
R6839t1616 n6840 n1617 R=1.913e+01 
R6840t5381 n6841 n5382 R=8.067e+00 
R6840t5777 n6841 n5778 R=8.081e+00 
R6840t853 n6841 n854 R=1.964e+01 
R6840t2843 n6841 n2844 R=2.724e+01 
R6840t2034 n6841 n2035 R=4.443e+00 
R6841t3234 n6842 n3235 R=8.636e+00 
R6841t1232 n6842 n1233 R=6.710e+00 
R6841t4397 n6842 n4398 R=7.900e+01 
R6842t2015 n6843 n2016 R=3.368e+00 
R6842t3649 n6843 n3650 R=1.486e+01 
R6842t3432 n6843 n3433 R=3.578e+00 
R6842t5282 n6843 n5283 R=2.012e+01 
R6843t6386 n6844 n6387 R=4.533e+00 
R6843t6506 n6844 n6507 R=3.610e+00 
R6843t6159 n6844 n6160 R=3.079e+02 
R6843t3148 n6844 n3149 R=1.146e+01 
R6844t1951 n6845 n1952 R=1.271e+01 
R6844t5096 n6845 n5097 R=6.509e+00 
R6844t4229 n6845 n4230 R=2.585e+00 
R6845t2183 n6846 n2184 R=9.405e+00 
R6845t4999 n6846 n5000 R=4.385e+00 
R6845t1801 n6846 n1802 R=3.500e+01 
R6845t2768 n6846 n2769 R=7.089e+00 
R6845t302 n6846 n303 R=8.215e+00 
R6846t4718 n6847 n4719 R=7.171e+00 
R6846t5451 n6847 n5452 R=4.126e+00 
R6846t746 n6847 n747 R=6.605e+01 
R6846t5715 n6847 n5716 R=1.906e+00 
R6846t6145 n6847 n6146 R=1.716e+01 
R6846t1769 n6847 n1770 R=2.324e+01 
R6847t1229 n6848 n1230 R=3.136e+00 
R6847t6280 n6848 n6281 R=1.179e+01 
R6847t5781 n6848 n5782 R=4.416e+01 
R6847t1943 n6848 n1944 R=4.254e+00 
R6847t2244 n6848 n2245 R=8.375e+00 
R6847t1983 n6848 n1984 R=2.282e+01 
R6848t527 n6849 n528 R=1.087e+01 
R6848t4062 n6849 n4063 R=5.326e+00 
R6848t4196 n6849 n4197 R=3.872e+00 
R6849t446 n6850 n447 R=1.801e+01 
R6849t5071 n6850 n5072 R=3.805e+00 
R6849t5251 n6850 n5252 R=3.638e+00 
R6849t988 n6850 n989 R=2.249e+01 
R6850t3665 n6851 n3666 R=2.267e+00 
R6850t6085 n6851 n6086 R=4.098e+01 
R6850t1264 n6851 n1265 R=6.113e+00 
R6850t514 n6851 n515 R=3.792e+00 
R6851t152 n6852 n153 R=3.970e+00 
R6851t6065 n6852 n6066 R=4.509e+00 
R6851t6060 n6852 n6061 R=2.295e+01 
R6851t3151 n6852 n3152 R=1.007e+01 
R6852t1081 n6853 n1082 R=3.656e+00 
R6852t5079 n6853 n5080 R=2.528e+00 
R6852t1540 n6853 n1541 R=3.098e+01 
R6852t6216 n6853 n6217 R=8.614e+00 
R6852t3918 n6853 n3919 R=1.972e+01 
R6853t3257 n6854 n3258 R=5.489e+00 
R6853t1857 n6854 n1858 R=4.957e+00 
R6853t4045 n6854 n4046 R=8.478e+00 
R6853t3352 n6854 n3353 R=3.249e+01 
R6853t6402 n6854 n6403 R=2.094e+01 
R6854t728 n6855 n729 R=3.365e+00 
R6854t1563 n6855 n1564 R=3.988e+01 
R6854t2415 n6855 n2416 R=1.645e+01 
R6854t5348 n6855 n5349 R=2.614e+00 
R6855t2328 n6856 n2329 R=5.370e+00 
R6855t1149 n6856 n1150 R=5.087e+00 
R6855t3959 n6856 n3960 R=3.706e+01 
R6855t1328 n6856 n1329 R=6.999e+00 
R6856t2904 n6857 n2905 R=1.742e+01 
R6856t1323 n6857 n1324 R=4.115e+01 
R6856t5189 n6857 n5190 R=6.028e+00 
R6856t3935 n6857 n3936 R=9.934e+00 
R6857t277 n6858 n278 R=5.370e+00 
R6857t5259 n6858 n5260 R=7.840e+00 
R6857t6135 n6858 n6136 R=9.129e+00 
R6857t3561 n6858 n3562 R=7.146e+00 
R6857t1538 n6858 n1539 R=1.847e+02 
R6858t5650 n6859 n5651 R=8.282e+01 
R6858t3172 n6859 n3173 R=3.107e+01 
R6858t2470 n6859 n2471 R=1.180e+01 
R6858t5878 n6859 n5879 R=4.662e+01 
R6859t3532 n6860 n3533 R=2.321e+01 
R6859t1966 n6860 n1967 R=5.275e+00 
R6859t4845 n6860 n4846 R=2.056e+01 
R6859t4289 n6860 n4290 R=3.333e+00 
R6859t2718 n6860 n2719 R=3.929e+01 
R6860t705 n6861 n706 R=6.766e+00 
R6860t2229 n6861 n2230 R=1.408e+01 
R6860t2216 n6861 n2217 R=3.831e+00 
R6860t424 n6861 n425 R=8.168e+00 
R6860t4903 n6861 n4904 R=3.117e+02 
R6860t5520 n6861 n5521 R=6.407e+00 
R6860t1714 n6861 n1715 R=1.807e+01 
R6861t145 n6862 n146 R=1.505e+01 
R6861t1528 n6862 n1529 R=3.981e+00 
R6861t1771 n6862 n1772 R=4.701e+00 
R6861t6429 n6862 n6430 R=4.687e+00 
R6862t173 n6863 n174 R=2.740e+00 
R6862t2803 n6863 n2804 R=2.753e+01 
R6862t292 n6863 n293 R=1.831e+01 
R6862t904 n6863 n905 R=9.771e+00 
R6862t2715 n6863 n2716 R=6.903e+00 
R6863t6798 n6864 n6799 R=3.064e+00 
R6863t343 n6864 n344 R=1.181e+00 
R6864t1451 n6865 n1452 R=8.822e+02 
R6864t5 n6865 n6 R=4.500e+00 
R6865t5631 n6866 n5632 R=2.050e+02 
R6865t3982 n6866 n3983 R=2.314e+01 
R6865t3749 n6866 n3750 R=1.674e+01 
R6865t3138 n6866 n3139 R=8.684e+00 
R6865t1040 n6866 n1041 R=1.461e+02 
R6865t490 n6866 n491 R=2.503e+00 
R6866t2614 n6867 n2615 R=6.834e+00 
R6866t4340 n6867 n4341 R=5.353e+00 
R6866t1625 n6867 n1626 R=5.610e+00 
R6866t3039 n6867 n1 R=5.967e+01 
R6866t4202 n6867 n4203 R=3.411e+00 
R6867t3696 n6868 n3697 R=7.329e+01 
R6867t5461 n6868 n5462 R=1.551e+01 
R6867t2069 n6868 n2070 R=2.240e+00 
R6867t4013 n6868 n4014 R=4.868e+00 
R6867t6051 n6868 n6052 R=2.176e+01 
R6868t3019 n6869 n3020 R=1.482e+02 
R6868t1668 n6869 n1669 R=3.275e+00 
R6868t4710 n6869 n4711 R=1.346e+01 
R6868t4047 n6869 n4048 R=1.654e+01 
R6869t1695 n6870 n1696 R=4.680e+00 
R6869t5366 n6870 n5367 R=2.472e+01 
R6869t3134 n6870 n3135 R=3.852e+01 
R6869t5048 n6870 n5049 R=7.442e+00 
R6870t2741 n6871 n2742 R=2.898e+00 
R6870t3483 n6871 n3484 R=1.850e+01 
R6870t5641 n6871 n5642 R=9.724e+00 
R6870t6181 n6871 n6182 R=3.241e+00 
R6870t1898 n6871 n1899 R=9.022e+00 
R6871t4951 n6872 n4952 R=7.232e+00 
R6871t1998 n6872 n1999 R=5.068e+00 
R6871t4231 n6872 n4232 R=1.561e+01 
R6872t4051 n6873 n4052 R=1.492e+01 
R6872t5402 n6873 n5403 R=4.421e+00 
R6872t4104 n6873 n4105 R=4.849e+00 
R6872t5558 n6873 n5559 R=4.293e+01 
R6872t1281 n6873 n1282 R=1.395e+01 
R6873t2254 n6874 n2255 R=2.237e+01 
R6873t6447 n6874 n6448 R=5.194e+00 
R6873t5815 n6874 n5816 R=3.153e+01 
R6873t4002 n6874 n4003 R=4.622e+00 
R6874t1203 n6875 n1204 R=6.958e+00 
R6874t2246 n6875 n2247 R=7.855e+00 
R6874t1117 n6875 n1118 R=2.311e+01 
R6874t4087 n6875 n4088 R=2.414e+00 
R6874t5966 n6875 n5967 R=8.526e+00 
R6875t2301 n6876 n2302 R=2.089e+00 
R6875t2933 n6876 n2934 R=9.742e+00 
R6875t5740 n6876 n5741 R=7.881e+01 
R6875t1930 n6876 n1931 R=1.525e+01 
R6876t4939 n6877 n4940 R=1.262e+01 
R6876t6115 n6877 n6116 R=2.123e+00 
R6876t2014 n6877 n2015 R=2.603e+01 
R6876t1653 n6877 n1654 R=5.154e+00 
R6876t3991 n6877 n3992 R=8.369e+00 
R6877t1226 n6878 n1227 R=7.886e+00 
R6877t2050 n6878 n2051 R=5.388e+00 
R6877t1285 n6878 n1286 R=2.346e+00 
R6878t2292 n6879 n2293 R=7.290e+00 
R6878t4962 n6879 n4963 R=6.736e+01 
R6878t1041 n6879 n1042 R=1.236e+01 
R6878t3146 n6879 n3147 R=2.394e+00 
R6878t6250 n6879 n6251 R=1.190e+01 
R6879t1759 n6880 n1760 R=1.586e+01 
R6879t6594 n6880 n6595 R=4.629e+00 
R6879t4632 n6880 n4633 R=1.698e+01 
R6879t4832 n6880 n4833 R=4.389e+00 
R6879t948 n6880 n949 R=8.825e+00 
R6879t1963 n6880 n1964 R=7.915e+00 
R6879t6440 n6880 n6441 R=4.685e+01 
R6880t2322 n6881 n2323 R=3.439e+01 
R6880t5508 n6881 n5509 R=3.131e+00 
R6880t6745 n6881 n6746 R=2.892e+00 
R6881t317 n6882 n318 R=1.293e+01 
R6881t1644 n6882 n1645 R=2.695e+00 
R6881t5390 n6882 n5391 R=1.487e+01 
R6881t3720 n6882 n3721 R=9.619e+01 
R6881t6570 n6882 n6571 R=1.520e+00 
R6882t379 n6883 n380 R=3.225e+00 
R6882t5944 n6883 n5945 R=5.467e+00 
R6882t5124 n6883 n5125 R=3.087e+00 
R6882t1105 n6883 n1106 R=1.660e+01 
R6883t3463 n6884 n3464 R=3.818e+01 
R6883t1051 n6884 n1052 R=1.263e+01 
R6884t4324 n6885 n4325 R=3.544e+02 
R6884t5293 n6885 n5294 R=6.907e+00 
R6884t3266 n6885 n3267 R=9.125e+00 
R6885t209 n6886 n210 R=6.754e+00 
R6885t873 n6886 n874 R=7.284e+01 
R6885t6224 n6886 n6225 R=1.265e+01 
R6885t2432 n6886 n2433 R=7.369e+00 
R6886t2096 n6887 n2097 R=3.729e+00 
R6886t2533 n6887 n2534 R=3.583e+00 
R6887t3518 n6888 n3519 R=7.500e+00 
R6887t5747 n6888 n5748 R=3.776e+00 
R6887t6135 n6888 n6136 R=2.741e+01 
R6887t3561 n6888 n3562 R=5.062e+00 
R6887t2421 n6888 n2422 R=1.540e+01 
R6887t3032 n6888 n3033 R=2.247e+01 
R6887t5428 n6888 n5429 R=1.287e+01 
R6888t4519 n6889 n4520 R=1.083e+01 
R6888t6583 n6889 n6584 R=1.303e+01 
R6888t3981 n6889 n3982 R=5.661e+00 
R6888t5445 n6889 n5446 R=1.574e+01 
R6888t5007 n6889 n5008 R=4.122e+00 
R6889t2817 n6890 n2818 R=3.549e+00 
R6889t4790 n6890 n4791 R=3.464e+00 
R6889t4844 n6890 n4845 R=3.728e+01 
R6889t6475 n6890 n6476 R=7.002e+00 
R6890t1613 n6891 n1614 R=6.314e+00 
R6890t4241 n6891 n4242 R=7.871e+00 
R6890t1921 n6891 n1922 R=5.228e+00 
R6890t3403 n6891 n3404 R=3.805e+00 
R6890t3547 n6891 n3548 R=6.275e+01 
R6891t3257 n6892 n3258 R=1.837e+01 
R6891t1103 n6892 n1104 R=1.713e+01 
R6891t1242 n6892 n1243 R=5.298e+01 
R6891t5984 n6892 n5985 R=9.028e+00 
R6891t1857 n6892 n1858 R=1.035e+01 
R6891t6853 n6892 n6854 R=2.738e+01 
R6892t3822 n6893 n3823 R=3.231e+00 
R6892t5166 n6893 n5167 R=5.050e+00 
R6892t465 n6893 n466 R=2.699e+01 
R6893t2992 n6894 n2993 R=2.748e+00 
R6893t3863 n6894 n3864 R=9.403e+00 
R6893t5850 n6894 n5851 R=4.328e+00 
R6893t6267 n6894 n6268 R=5.435e+00 
R6894t882 n6895 n883 R=3.932e+00 
R6894t4120 n6895 n4121 R=4.629e+01 
R6894t382 n6895 n383 R=3.608e+02 
R6894t5522 n6895 n5523 R=3.721e+00 
R6894t5692 n6895 n5693 R=1.811e+01 
R6895t2790 n6896 n2791 R=7.937e+00 
R6895t5446 n6896 n5447 R=8.417e+00 
R6895t2636 n6896 n2637 R=9.866e+00 
R6895t2735 n6896 n2736 R=9.716e+00 
R6896t4354 n6897 n4355 R=3.421e+01 
R6896t4637 n6897 n4638 R=3.032e+00 
R6896t3701 n6897 n3702 R=3.303e+00 
R6897t1521 n6898 n1522 R=8.434e+00 
R6897t3014 n6898 n3015 R=3.230e+00 
R6897t827 n6898 n828 R=2.038e+00 
R6898t4834 n6899 n4835 R=9.723e+00 
R6898t685 n6899 n686 R=1.953e+01 
R6898t488 n6899 n489 R=7.810e+00 
R6899t4089 n6900 n4090 R=9.720e+00 
R6899t4864 n6900 n4865 R=2.827e+01 
R6899t2619 n6900 n2620 R=5.890e+00 
R6899t1681 n6900 n1682 R=5.187e+00 
R6900t2695 n6901 n2696 R=2.159e+00 
R6900t4097 n6901 n4098 R=5.761e+00 
R6900t760 n6901 n761 R=1.957e+00 
R6901t2018 n6902 n2019 R=7.517e+00 
R6901t706 n6902 n707 R=1.024e+01 
R6901t2387 n6902 n2388 R=4.909e+00 
R6902t6647 n6903 n6648 R=6.570e+00 
R6902t3505 n6903 n3506 R=1.860e+01 
R6903t2277 n6904 n2278 R=3.025e+01 
R6903t6355 n6904 n6356 R=2.988e+00 
R6903t5313 n6904 n5314 R=1.478e+01 
R6904t6221 n6905 n6222 R=2.008e+01 
R6904t5919 n6905 n5920 R=6.913e+01 
R6904t6470 n6905 n6471 R=7.523e+00 
R6904t4835 n6905 n4836 R=6.862e+00 
R6905t4288 n6906 n4289 R=3.931e+00 
R6905t6711 n6906 n6712 R=6.355e+01 
R6905t6067 n6906 n6068 R=1.485e+01 
R6905t1596 n6906 n1597 R=5.546e+00 
R6905t5956 n6906 n5957 R=2.356e+01 
R6906t2603 n6907 n2604 R=2.714e+01 
R6906t3068 n6907 n3069 R=1.832e+01 
R6906t3639 n6907 n3640 R=1.848e+01 
R6906t5262 n6907 n5263 R=2.261e+00 
R6906t3970 n6907 n3971 R=7.582e+01 
R6906t4663 n6907 n4664 R=6.412e+00 
R6906t1044 n6907 n1045 R=5.055e+00 
R6907t611 n6908 n612 R=1.949e+01 
R6907t4218 n6908 n4219 R=1.182e+01 
R6907t2460 n6908 n2461 R=3.208e+00 
R6907t4930 n6908 n4931 R=2.668e+01 
R6907t2971 n6908 n2972 R=2.446e+00 
R6907t1389 n6908 n1390 R=1.346e+01 
R6908t3468 n6909 n3469 R=4.720e+02 
R6909t1475 n6910 n1476 R=6.068e+00 
R6909t6558 n6910 n6559 R=6.306e+01 
R6909t3230 n6910 n3231 R=4.202e+00 
R6910t3937 n6911 n3938 R=4.945e+00 
R6911t1276 n6912 n1277 R=4.636e+00 
R6911t6617 n6912 n6618 R=5.095e+00 
R6911t1250 n6912 n1251 R=9.719e+00 
R6911t2716 n6912 n2717 R=5.905e+01 
R6912t2310 n6913 n2311 R=1.229e+01 
R6912t4930 n6913 n4931 R=5.308e+00 
R6912t2460 n6913 n2461 R=9.529e+01 
R6912t1474 n6913 n1475 R=2.725e+00 
R6912t725 n6913 n726 R=3.746e+01 
R6913t2475 n6914 n2476 R=6.732e+01 
R6913t4775 n6914 n4776 R=6.213e+00 
R6913t5666 n6914 n5667 R=6.535e+00 
R6913t2656 n6914 n2657 R=1.759e+00 
R6914t1883 n6915 n1884 R=1.377e+01 
R6914t2872 n6915 n2873 R=5.815e+00 
R6914t2568 n6915 n2569 R=1.709e+01 
R6914t3254 n6915 n3255 R=1.026e+01 
R6914t750 n6915 n751 R=4.746e+00 
R6915t4255 n6916 n4256 R=2.864e+00 
R6915t5279 n6916 n5280 R=4.248e+02 
R6915t6298 n6916 n6299 R=1.237e+01 
R6915t4713 n6916 n4714 R=1.800e+01 
R6915t1061 n6916 n1062 R=1.878e+01 
R6915t4719 n6916 n4720 R=5.130e+00 
R6916t686 n6917 n687 R=3.603e+01 
R6916t6133 n6917 n6134 R=1.938e+01 
R6916t4979 n6917 n4980 R=8.296e+00 
R6917t6864 n6918 n6865 R=6.658e+00 
R6917t2638 n6918 n2639 R=4.289e+00 
R6917t1592 n6918 n1593 R=2.300e+01 
R6917t681 n6918 n682 R=6.491e+00 
R6917t5 n6918 n6 R=9.873e+00 
R6918t3449 n6919 n3450 R=2.005e+01 
R6918t4534 n6919 n4535 R=5.787e+00 
R6918t1949 n6919 n1950 R=1.126e+01 
R6918t3712 n6919 n3713 R=1.268e+01 
R6918t5829 n6919 n5830 R=7.357e+00 
R6919t238 n6920 n239 R=3.587e+00 
R6919t1877 n6920 n1878 R=6.702e+01 
R6919t2804 n6920 n2805 R=9.968e+00 
R6919t5811 n6920 n5812 R=1.191e+01 
R6919t2452 n6920 n2453 R=6.990e+00 
R6920t1215 n6921 n1216 R=6.916e+00 
R6920t3571 n6921 n3572 R=9.030e+00 
R6920t5494 n6921 n5495 R=3.130e+01 
R6920t3289 n6921 n3290 R=2.776e+00 
R6920t5971 n6921 n5972 R=4.961e+01 
R6920t3074 n6921 n3075 R=5.037e+01 
R6920t1039 n6921 n1040 R=3.710e+00 
R6921t200 n6922 n201 R=4.106e+00 
R6921t875 n6922 n876 R=4.232e+01 
R6921t826 n6922 n827 R=1.164e+02 
R6921t4894 n6922 n4895 R=1.741e+00 
R6922t923 n6923 n924 R=3.170e+00 
R6922t5894 n6923 n5895 R=6.166e+00 
R6923t4287 n6924 n4288 R=3.487e+00 
R6923t6699 n6924 n6700 R=6.310e+01 
R6923t1325 n6924 n1326 R=9.403e+00 
R6923t2511 n6924 n2512 R=1.869e+01 
R6924t5914 n6925 n5915 R=6.598e+00 
R6924t3971 n6925 n3972 R=2.467e+01 
R6925t1358 n6926 n1359 R=3.800e+01 
R6925t5978 n6926 n5979 R=3.773e+00 
R6926t2825 n6927 n2826 R=3.135e+01 
R6926t5203 n6927 n5204 R=5.864e+00 
R6926t2531 n6927 n2532 R=1.148e+01 
R6926t130 n6927 n131 R=3.466e+00 
R6926t726 n6927 n727 R=6.345e+00 
R6927t474 n6928 n475 R=3.112e+01 
R6927t1964 n6928 n1965 R=3.283e+00 
R6927t6422 n6928 n6423 R=7.393e+00 
R6927t4289 n6928 n4290 R=2.405e+01 
R6927t4845 n6928 n4846 R=4.139e+00 
R6928t1292 n6929 n1293 R=1.477e+01 
R6928t4556 n6929 n4557 R=1.143e+01 
R6928t3099 n6929 n3100 R=6.766e+00 
R6928t4695 n6929 n4696 R=1.345e+01 
R6929t866 n6930 n867 R=1.166e+01 
R6929t1426 n6930 n1427 R=5.235e+00 
R6929t2191 n6930 n2192 R=2.068e+02 
R6930t974 n6931 n975 R=2.865e+00 
R6930t576 n6931 n577 R=3.485e+01 
R6930t5693 n6931 n5694 R=2.218e+01 
R6930t3449 n6931 n3450 R=3.756e+00 
R6930t5829 n6931 n5830 R=5.208e+00 
R6931t6822 n6932 n6823 R=1.563e+00 
R6931t6867 n6932 n6868 R=3.085e+01 
R6931t2069 n6932 n2070 R=2.835e+00 
R6931t4171 n6932 n4172 R=2.711e+01 
R6932t5010 n6933 n5011 R=8.688e+00 
R6932t5696 n6933 n5697 R=1.844e+00 
R6932t2430 n6933 n2431 R=2.350e+00 
R6933t2498 n6934 n2499 R=1.597e+01 
R6933t6077 n6934 n6078 R=9.159e+00 
R6933t4607 n6934 n4608 R=1.951e+00 
R6933t5574 n6934 n5575 R=1.533e+02 
R6933t3085 n6934 n3086 R=7.007e+00 
R6934t3405 n6935 n3406 R=5.541e+00 
R6934t5359 n6935 n5360 R=5.086e+00 
R6935t344 n6936 n345 R=9.231e+00 
R6935t4167 n6936 n4168 R=5.644e+00 
R6935t756 n6936 n757 R=4.614e+00 
R6935t3681 n6936 n3682 R=4.645e+01 
R6935t1110 n6936 n1111 R=3.788e+00 
R6936t2750 n6937 n2751 R=4.200e+00 
R6936t6338 n6937 n6339 R=2.142e+01 
R6936t2082 n6937 n2083 R=2.450e+01 
R6936t642 n6937 n643 R=9.825e+00 
R6936t1499 n6937 n1500 R=1.485e+01 
R6936t63 n6937 n64 R=9.891e+00 
R6936t5651 n6937 n5652 R=5.288e+02 
R6937t4653 n6938 n4654 R=1.427e+01 
R6937t241 n6938 n242 R=3.145e+02 
R6937t2397 n6938 n2398 R=5.872e+00 
R6937t681 n6938 n682 R=4.205e+00 
R6937t5198 n6938 n5199 R=4.114e+01 
R6938t5424 n6939 n5425 R=4.252e+01 
R6938t3387 n6939 n3388 R=4.907e+00 
R6938t4466 n6939 n4467 R=3.235e+01 
R6938t4871 n6939 n4872 R=1.293e+01 
R6938t5026 n6939 n5027 R=6.122e+00 
R6939t1811 n6940 n1812 R=3.540e+00 
R6939t3956 n6940 n3957 R=4.284e+00 
R6939t1443 n6940 n1444 R=2.630e+01 
R6939t1409 n6940 n1410 R=2.196e+00 
R6940t4 n6941 n5 R=7.154e+00 
R6940t970 n6941 n971 R=4.618e+00 
R6940t4285 n6941 n4286 R=1.063e+01 
R6940t1805 n6941 n1806 R=5.941e+00 
R6940t5923 n6941 n5924 R=3.267e+00 
R6941t5314 n6942 n5315 R=9.662e+00 
R6941t6162 n6942 n6163 R=2.115e+01 
R6941t3671 n6942 n3672 R=3.609e+00 
R6941t945 n6942 n946 R=1.866e+02 
R6941t2059 n6942 n2060 R=2.825e+00 
R6942t395 n6943 n396 R=3.275e+00 
R6942t4628 n6943 n4629 R=7.653e+00 
R6942t137 n6943 n138 R=2.105e+00 
R6942t4910 n6943 n4911 R=6.629e+01 
R6942t2379 n6943 n2380 R=1.504e+01 
R6943t2929 n6944 n2930 R=9.643e+00 
R6943t894 n6944 n895 R=1.416e+01 
R6943t3612 n6944 n3613 R=1.922e+01 
R6943t5320 n6944 n5321 R=3.331e+01 
R6943t65 n6944 n66 R=1.574e+01 
R6944t2463 n6945 n2464 R=4.618e+00 
R6944t4657 n6945 n4658 R=2.825e+01 
R6944t1273 n6945 n1 R=2.619e+01 
R6944t5209 n6945 n1 R=1.418e+01 
R6944t301 n6945 n302 R=6.691e+00 
R6945t4149 n6946 n4150 R=6.079e+00 
R6945t5372 n6946 n5373 R=3.359e+00 
R6945t4150 n6946 n4151 R=5.512e+00 
R6945t6600 n6946 n6601 R=1.609e+01 
R6945t676 n6946 n677 R=7.305e+00 
R6946t468 n6947 n469 R=1.190e+01 
R6946t507 n6947 n508 R=3.800e+00 
R6946t3540 n6947 n3541 R=1.889e+02 
R6946t433 n6947 n434 R=1.111e+01 
R6946t2628 n6947 n2629 R=3.249e+00 
R6946t3479 n6947 n3480 R=3.103e+01 
R6947t4300 n6948 n4301 R=6.189e+00 
R6948t5378 n6949 n5379 R=6.243e+00 
R6948t6037 n6949 n6038 R=8.474e+00 
R6948t3287 n6949 n3288 R=6.117e+00 
R6948t2651 n6949 n2652 R=1.200e+01 
R6949t400 n6950 n401 R=4.383e+00 
R6949t887 n6950 n888 R=3.258e+00 
R6949t1394 n6950 n1395 R=6.483e+00 
R6949t4973 n6950 n4974 R=5.040e+01 
R6950t1290 n6951 n1291 R=4.997e+00 
R6950t6776 n6951 n6777 R=2.686e+01 
R6950t192 n6951 n193 R=1.266e+01 
R6950t1706 n6951 n1707 R=6.955e+00 
R6951t28 n6952 n29 R=2.749e+00 
R6951t3562 n6952 n3563 R=3.719e+00 
R6951t118 n6952 n119 R=1.495e+01 
R6951t839 n6952 n840 R=2.235e+01 
R6951t266 n6952 n267 R=1.005e+02 
R6952t5863 n6953 n5864 R=4.334e+00 
R6952t4061 n6953 n4062 R=6.563e+00 
R6952t1262 n6953 n1263 R=4.381e+00 
R6953t6415 n6954 n6416 R=3.103e+00 
R6953t2120 n6954 n2121 R=7.353e+01 
R6953t5891 n6954 n5892 R=3.711e+00 
R6954t4519 n6955 n4520 R=5.819e+00 
R6954t6888 n6955 n6889 R=7.616e+00 
R6954t5007 n6955 n5008 R=2.531e+01 
R6954t3422 n6955 n3423 R=1.592e+01 
R6954t3415 n6955 n3416 R=7.928e+00 
R6955t1223 n6956 n1224 R=3.641e+01 
R6955t719 n6956 n720 R=7.319e+00 
R6955t2576 n6956 n2577 R=7.593e+00 
R6955t6049 n6956 n6050 R=4.262e+00 
R6955t1053 n6956 n1054 R=6.908e+00 
R6956t2390 n6957 n2391 R=9.942e+00 
R6956t2299 n6957 n2300 R=2.947e+00 
R6956t4901 n6957 n4902 R=1.793e+01 
R6956t3047 n6957 n3048 R=1.690e+01 
R6957t5655 n6958 n5656 R=8.664e+00 
R6957t3154 n6958 n3155 R=2.820e+00 
R6958t1287 n6959 n1288 R=6.830e+00 
R6958t4841 n6959 n4842 R=8.511e+00 
R6958t1355 n6959 n1356 R=1.764e+01 
R6958t2116 n6959 n2117 R=3.627e+00 
R6959t2107 n6960 n2108 R=4.024e+01 
R6959t2319 n6960 n2320 R=1.278e+01 
R6959t5604 n6960 n5605 R=4.810e+00 
R6959t6343 n6960 n6344 R=1.801e+01 
R6959t1356 n6960 n1357 R=2.103e+01 
R6959t3645 n6960 n3646 R=6.637e+00 
R6959t6759 n6960 n6760 R=1.231e+01 
R6960t1929 n6961 n1930 R=2.380e+01 
R6960t2191 n6961 n2192 R=6.934e+01 
R6960t1687 n6961 n1688 R=2.362e+00 
R6960t3641 n6961 n3642 R=3.031e+01 
R6960t3959 n6961 n3960 R=1.344e+01 
R6960t5363 n6961 n5364 R=3.474e+00 
R6960t1979 n6961 n1980 R=1.124e+01 
R6961t565 n6962 n566 R=1.803e+02 
R6961t3570 n6962 n3571 R=3.543e+00 
R6961t3139 n6962 n3140 R=4.833e+00 
R6962t2317 n6963 n2318 R=1.364e+02 
R6962t6794 n6963 n6795 R=8.937e+00 
R6962t616 n6963 n617 R=1.551e+01 
R6962t5797 n6963 n5798 R=4.036e+00 
R6963t1099 n6964 n1100 R=6.738e+00 
R6963t5509 n6964 n5510 R=5.237e+01 
R6963t29 n6964 n30 R=1.782e+01 
R6963t3443 n6964 n3444 R=6.338e+01 
R6963t3166 n6964 n3167 R=5.381e+00 
R6963t6354 n6964 n6355 R=1.949e+01 
R6964t4026 n6965 n4027 R=1.329e+01 
R6964t4062 n6965 n4063 R=1.395e+01 
R6964t5775 n6965 n5776 R=3.641e+00 
R6964t5864 n6965 n5865 R=1.960e+01 
R6965t4259 n6966 n4260 R=6.954e+00 
R6965t1614 n6966 n1615 R=5.429e+00 
R6965t2763 n6966 n2764 R=5.871e+00 
R6965t552 n6966 n553 R=7.689e+00 
R6967t2341 n6968 n2342 R=3.762e+00 
R6967t2883 n6968 n2884 R=5.204e+00 
R6967t4931 n6968 n4932 R=6.351e+00 
R6968t1015 n6969 n1016 R=1.216e+01 
R6968t4644 n6969 n4645 R=6.763e+00 
R6968t1761 n6969 n1762 R=1.790e+01 
R6968t3987 n6969 n3988 R=5.157e+00 
R6968t5084 n6969 n5085 R=5.656e+00 
R6969t171 n6970 n172 R=4.223e+00 
R6969t4509 n6970 n4510 R=9.081e+00 
R6969t5955 n6970 n5956 R=1.754e+01 
R6969t6590 n6970 n6591 R=3.376e+01 
R6969t2288 n6970 n2289 R=6.118e+01 
R6970t2321 n6971 n2322 R=1.703e+02 
R6970t4942 n6971 n4943 R=4.899e+00 
R6970t2805 n6971 n2806 R=2.389e+01 
R6970t3445 n6971 n3446 R=3.404e+01 
R6970t3178 n6971 n3179 R=2.369e+01 
R6970t5556 n6971 n5557 R=1.149e+01 
R6970t2444 n6971 n2445 R=3.960e+00 
R6971t2060 n6972 n2061 R=1.971e+01 
R6971t6306 n6972 n6307 R=7.030e+00 
R6971t997 n6972 n998 R=1.194e+02 
R6971t5228 n6972 n5229 R=3.340e+00 
R6972t517 n6973 n518 R=2.361e+02 
R6972t1497 n6973 n1498 R=1.874e+01 
R6972t261 n6973 n262 R=2.149e+00 
R6972t3734 n6973 n3735 R=1.407e+02 
R6972t4443 n6973 n4444 R=4.264e+00 
R6972t5432 n6973 n5433 R=5.878e+00 
R6972t3981 n6973 n3982 R=2.020e+01 
R6973t590 n6974 n591 R=5.237e+00 
R6973t6159 n6974 n6160 R=8.657e+01 
R6973t6506 n6974 n6507 R=2.486e+01 
R6973t1800 n6974 n1801 R=5.258e+00 
R6973t5071 n6974 n5072 R=5.893e+00 
R6973t4661 n6974 n4662 R=7.611e+00 
R6974t1177 n6975 n1178 R=2.836e+00 
R6974t4540 n6975 n4541 R=9.722e+01 
R6974t6022 n6975 n6023 R=2.403e+00 
R6974t4392 n6975 n4393 R=1.077e+01 
R6975t2278 n6976 n2279 R=7.577e+01 
R6975t5388 n6976 n5389 R=1.038e+02 
R6975t269 n6976 n270 R=3.572e+01 
R6975t3567 n6976 n3568 R=2.549e+01 
R6975t4380 n6976 n4381 R=1.010e+02 
R6975t229 n6976 n230 R=6.968e+00 
R6975t6093 n6976 n6094 R=7.592e+00 
R6976t2451 n6977 n2452 R=7.396e+00 
R6976t3306 n6977 n3307 R=4.452e+02 
R6976t154 n6977 n155 R=7.692e+00 
R6976t1679 n6977 n1680 R=9.993e+01 
R6976t1721 n6977 n1722 R=1.600e+01 
R6976t5072 n6977 n5073 R=4.493e+00 
R6977t3221 n6978 n3222 R=1.625e+01 
R6977t1128 n6978 n1129 R=2.483e+00 
R6977t1469 n6978 n1470 R=7.556e+01 
R6978t2626 n6979 n2627 R=7.595e+00 
R6978t6201 n6979 n6202 R=6.135e+00 
R6978t4532 n6979 n4533 R=7.816e+00 
R6978t2561 n6979 n2562 R=1.432e+01 
R6978t6705 n6979 n6706 R=9.252e+00 
R6978t694 n6979 n695 R=3.118e+01 
R6978t6179 n6979 n6180 R=6.045e+00 
R6979t6948 n6980 n6949 R=6.362e+00 
R6979t492 n6980 n493 R=8.064e+00 
R6979t314 n6980 n315 R=2.415e+01 
R6979t2986 n6980 n2987 R=9.966e+00 
R6980t3003 n6981 n3004 R=5.665e+00 
R6980t3315 n6981 n3316 R=2.294e+01 
R6980t5047 n6981 n5048 R=2.908e+00 
R6981t2248 n6982 n2249 R=2.755e+00 
R6981t6106 n6982 n6107 R=4.194e+00 
R6982t2823 n6983 n2824 R=6.147e+01 
R6982t2213 n6983 n2214 R=3.553e+00 
R6982t5384 n6983 n5385 R=5.166e+01 
R6982t5588 n6983 n5589 R=3.695e+00 
R6983t4099 n6984 n4100 R=5.428e+00 
R6983t5047 n6984 n5048 R=7.364e+00 
R6983t3315 n6984 n3316 R=5.341e+00 
R6984t4301 n6985 n4302 R=1.137e+01 
R6984t6687 n6985 n6688 R=7.437e+00 
R6984t6154 n6985 n6155 R=1.302e+01 
R6984t4045 n6985 n4046 R=1.493e+01 
R6985t6947 n6986 n6948 R=4.467e+01 
R6985t6221 n6986 n6222 R=4.035e+00 
R6985t6904 n6986 n6905 R=4.625e+00 
R6986t5936 n6987 n5937 R=6.631e+00 
R6986t6658 n6987 n6659 R=2.979e+00 
R6986t1557 n6987 n1558 R=4.706e+00 
R6986t937 n6987 n938 R=7.332e+00 
R6987t502 n6988 n503 R=2.294e+00 
R6987t4700 n6988 n4701 R=1.063e+01 
R6987t1423 n6988 n1424 R=3.112e+01 
R6987t6625 n6988 n6626 R=3.933e+00 
R6987t4181 n6988 n4182 R=3.332e+01 
R6988t3460 n6989 n3461 R=6.560e+00 
R6988t4824 n6989 n4825 R=2.321e+00 
R6988t2068 n6989 n2069 R=4.542e+01 
R6989t509 n6990 n510 R=3.018e+01 
R6989t2384 n6990 n2385 R=1.833e+01 
R6989t4304 n6990 n4305 R=2.415e+00 
R6989t775 n6990 n776 R=2.487e+00 
R6990t906 n6991 n907 R=9.455e+00 
R6990t5912 n6991 n5913 R=1.039e+01 
R6990t2225 n6991 n2226 R=5.924e+00 
R6990t5714 n6991 n5715 R=2.869e+01 
R6991t10 n6992 n11 R=4.303e+01 
R6991t5250 n6992 n5251 R=1.413e+02 
R6991t5065 n6992 n5066 R=2.118e+00 
R6991t4928 n6992 n4929 R=3.496e+02 
R6991t1057 n6992 n1058 R=7.496e+00 
R6992t2241 n6993 n2242 R=9.369e+00 
R6992t3677 n6993 n3678 R=7.699e+00 
R6992t1329 n6993 n1330 R=2.238e+01 
R6992t5050 n6993 n5051 R=9.583e+00 
R6992t1387 n6993 n1388 R=8.486e+00 
R6993t3892 n6994 n3893 R=4.860e+00 
R6993t43 n6994 n44 R=8.395e+00 
R6994t6229 n6995 n6230 R=2.933e+01 
R6994t6454 n6995 n6455 R=4.557e+00 
R6994t3227 n6995 n3228 R=3.003e+00 
R6995t1679 n6996 n1680 R=4.542e+00 
R6995t5805 n6996 n5806 R=4.083e+00 
R6995t1619 n6996 n1620 R=4.903e+01 
R6995t6031 n6996 n6032 R=6.932e+00 
R6995t3416 n6996 n3417 R=2.176e+01 
R6996t4146 n6997 n4147 R=9.951e+00 
R6996t143 n6997 n144 R=4.259e+00 
R6997t2669 n6998 n2670 R=1.029e+01 
R6997t5893 n6998 n5894 R=9.182e+00 
R6997t3746 n6998 n3747 R=2.674e+01 
R6997t5686 n6998 n5687 R=5.757e+00 
R6997t2842 n6998 n2843 R=1.880e+01 
R6997t5947 n6998 n5948 R=4.569e+00 
R6997t2698 n6998 n2699 R=1.888e+01 
R6998t3207 n6999 n3208 R=1.929e+01 
R6999t891 n7000 n892 R=3.356e+00 
R6999t3429 n7000 n3430 R=8.492e+00 
R6999t4842 n7000 n4843 R=1.295e+01 
R6999t5755 n7000 n5756 R=8.176e+00 
R6999t2435 n7000 n2436 R=1.760e+01 
R7000t253 n7001 n254 R=3.548e+01 
R7000t2559 n7001 n2560 R=4.518e+00 
R7000t3743 n7001 n3744 R=9.144e+01 
R7000t2134 n7001 n2135 R=4.884e+00 
R7000t2536 n7001 n2537 R=7.722e+00 
R7001t2848 n7002 n2849 R=4.982e+00 
R7001t6552 n7002 n6553 R=4.414e+00 
R7001t5032 n7002 n5033 R=1.243e+02 
R7001t1568 n7002 n1569 R=7.560e+00 
R7002t4567 n7003 n4568 R=1.596e+01 
R7002t4780 n7003 n4781 R=4.118e+00 
R7002t5578 n7003 n5579 R=1.115e+01 
R7002t4997 n7003 n4998 R=6.710e+00 
R7002t6977 n7003 n6978 R=1.294e+01 
R7003t3380 n7004 n3381 R=2.420e+00 
R7003t4071 n7004 n4072 R=2.013e+01 
R7004t4762 n7005 n4763 R=8.876e+00 
R7004t5485 n7005 n5486 R=2.423e+00 
R7004t2110 n7005 n2111 R=6.672e+00 
R7004t6828 n7005 n6829 R=8.232e+00 
R7004t4267 n7005 n4268 R=1.383e+02 
R7005t870 n7006 n871 R=3.132e+00 
R7005t3654 n7006 n3655 R=1.318e+01 
R7005t3327 n7006 n3328 R=7.408e+00 
R7006t1871 n7007 n1872 R=1.475e+01 
R7006t1309 n7007 n1310 R=6.238e+00 
R7006t2264 n7007 n2265 R=4.482e+00 
R7006t600 n7007 n601 R=1.761e+01 
R7006t6144 n7007 n6145 R=2.834e+00 
R7007t142 n7008 n143 R=2.545e+01 
R7007t3690 n7008 n3691 R=3.656e+00 
R7007t2822 n7008 n2823 R=1.262e+01 
R7008t5819 n7009 n5820 R=6.091e+00 
R7009t4731 n7010 n4732 R=6.623e+00 
R7009t4816 n7010 n4817 R=7.575e+00 
R7009t52 n7010 n53 R=1.972e+01 
R7009t6684 n7010 n6685 R=4.912e+00 
R7010t5550 n7011 n5551 R=3.007e+00 
R7010t3486 n7011 n3487 R=3.664e+01 
R7010t4261 n7011 n4262 R=8.673e+00 
R7010t3961 n7011 n3962 R=8.546e+00 
R7010t5904 n7011 n5905 R=7.835e+01 
R7010t6587 n7011 n6588 R=9.607e+00 
R7010t1121 n7011 n1122 R=4.888e+01 
R7011t364 n7012 n365 R=7.377e+00 
R7011t4549 n7012 n4550 R=9.031e+00 
R7011t6745 n7012 n6746 R=7.403e+00 
R7011t6880 n7012 n6881 R=1.017e+02 
R7012t3588 n7013 n3589 R=3.501e+00 
R7012t2367 n7013 n2368 R=2.917e+01 
R7012t5533 n7013 n5534 R=3.343e+00 
R7012t676 n7013 n677 R=1.522e+01 
R7012t2965 n7013 n2966 R=3.271e+01 
R7012t5826 n7013 n5827 R=2.123e+01 
R7013t2324 n7014 n2325 R=1.922e+02 
R7013t862 n7014 n863 R=4.602e+02 
R7013t3198 n7014 n3199 R=2.327e+01 
R7013t3125 n7014 n3126 R=2.562e+00 
R7014t1825 n7015 n1826 R=3.107e+00 
R7014t4318 n7015 n4319 R=3.075e+01 
R7014t362 n7015 n363 R=8.313e+00 
R7014t1680 n7015 n1681 R=5.348e+01 
R7014t4701 n7015 n4702 R=4.739e+00 
R7014t4770 n7015 n4771 R=3.980e+01 
R7015t854 n7016 n855 R=2.080e+01 
R7015t4179 n7016 n4180 R=4.722e+00 
R7015t2691 n7016 n2692 R=9.596e+00 
R7015t4245 n7016 n4246 R=8.268e+00 
R7015t4606 n7016 n4607 R=1.639e+01 
R7015t2543 n7016 n2544 R=7.851e+00 
R7016t6229 n7017 n6230 R=5.442e+00 
R7016t330 n7017 n331 R=1.386e+01 
R7016t4489 n7017 n4490 R=3.354e+00 
R7016t4114 n7017 n4115 R=7.780e+00 
R7017t1105 n7018 n1106 R=4.745e+00 
R7017t2556 n7018 n2557 R=1.485e+01 
R7017t6069 n7018 n6070 R=5.191e+00 
R7017t3470 n7018 n3471 R=4.313e+00 
R7018t93 n7019 n94 R=1.604e+01 
R7018t2147 n7019 n2148 R=2.249e+00 
R7018t3462 n7019 n3463 R=2.820e+01 
R7018t6796 n7019 n6797 R=3.745e+01 
R7018t6717 n7019 n6718 R=5.100e+00 
R7018t25 n7019 n26 R=4.787e+01 
R7019t39 n7020 n40 R=3.271e+00 
R7019t1748 n7020 n1749 R=4.882e+01 
R7019t1464 n7020 n1465 R=1.049e+01 
R7019t701 n7020 n702 R=9.662e+00 
R7019t6329 n7020 n6330 R=2.835e+00 
R7019t1454 n7020 n1455 R=1.729e+01 
R7020t4208 n7021 n4209 R=2.023e+01 
R7020t5937 n7021 n5938 R=4.175e+00 
R7020t4493 n7021 n4494 R=5.485e+00 
R7020t3472 n7021 n3473 R=8.622e+00 
R7020t3454 n7021 n3455 R=8.823e+00 
R7021t411 n7022 n412 R=8.079e+00 
R7021t862 n7022 n863 R=6.782e+02 
R7021t6236 n7022 n6237 R=3.117e+00 
R7021t6838 n7022 n6839 R=1.947e+01 
R7021t2181 n7022 n2182 R=3.128e+00 
R7022t2411 n7023 n2412 R=1.467e+01 
R7022t6576 n7023 n6577 R=2.421e+00 
R7022t814 n7023 n815 R=6.389e+00 
R7023t5144 n7024 n5145 R=3.161e+00 
R7023t5634 n7024 n5635 R=1.186e+01 
R7023t178 n7024 n179 R=4.240e+00 
R7023t4247 n7024 n4248 R=5.250e+02 
R7023t6341 n7024 n6342 R=7.571e+00 
R7024t4685 n7025 n4686 R=4.017e+00 
R7024t367 n7025 n368 R=2.711e+00 
R7025t4268 n7026 n4269 R=3.975e+00 
R7026t1390 n7027 n1391 R=7.114e+00 
R7026t2418 n7027 n2419 R=2.926e+00 
R7026t102 n7027 n103 R=8.511e+01 
R7026t2489 n7027 n2490 R=1.051e+02 
R7026t4722 n7027 n4723 R=3.012e+00 
R7027t4898 n7028 n4899 R=1.506e+01 
R7027t1818 n7028 n1819 R=5.217e+00 
R7028t403 n7029 n404 R=5.107e+00 
R7028t4663 n7029 n4664 R=6.419e+00 
R7028t3274 n7029 n3275 R=4.333e+01 
R7029t3956 n7030 n3957 R=5.220e+00 
R7029t4781 n7030 n4782 R=3.285e+01 
R7029t1719 n7030 n1720 R=6.244e+00 
R7029t2620 n7030 n2621 R=4.352e+00 
R7029t6674 n7030 n6675 R=2.077e+02 
R7030t285 n7031 n286 R=7.241e+01 
R7030t5218 n7031 n5219 R=4.317e+00 
R7030t5763 n7031 n5764 R=2.359e+00 
R7030t2132 n7031 n2133 R=4.088e+00 
R7031t5205 n7032 n5206 R=4.189e+01 
R7031t5227 n7032 n5228 R=3.870e+00 
R7031t5748 n7032 n5749 R=5.074e+00 
R7032t3395 n7033 n3396 R=2.207e+00 
R7032t4441 n7033 n4442 R=5.647e+00 
R7032t4106 n7033 n4107 R=1.332e+01 
R7032t851 n7033 n852 R=9.953e+00 
R7033t6084 n7034 n6085 R=5.772e+00 
R7033t4088 n7034 n4089 R=3.466e+00 
R7033t522 n7034 n523 R=1.471e+02 
R7033t2276 n7034 n2277 R=2.725e+01 
R7033t4081 n7034 n4082 R=8.197e+00 
R7033t5029 n7034 n5030 R=4.695e+00 
R7034t72 n7035 n73 R=3.978e+01 
R7034t4995 n7035 n4996 R=3.444e+00 
R7034t3179 n7035 n3180 R=2.023e+01 
R7034t6575 n7035 n6576 R=3.517e+00 
R7035t2823 n7036 n2824 R=3.662e+00 
R7035t3883 n7036 n3884 R=7.259e+00 
R7035t6982 n7036 n6983 R=5.540e+00 
R7036t1693 n7037 n1694 R=6.314e+00 
R7036t5185 n7037 n5186 R=4.138e+00 
R7036t2226 n7037 n2227 R=1.069e+01 
R7036t6406 n7037 n6407 R=7.395e+00 
R7037t2065 n7038 n2066 R=4.837e+00 
R7037t2224 n7038 n2225 R=5.414e+00 
R7037t5517 n7038 n5518 R=1.036e+02 
R7037t4563 n7038 n4564 R=4.684e+00 
R7037t4199 n7038 n4200 R=9.734e+00 
R7038t4033 n7039 n4034 R=5.766e+00 
R7038t6394 n7039 n6395 R=8.753e+00 
R7038t270 n7039 n271 R=1.056e+01 
R7038t377 n7039 n378 R=8.396e+00 
R7039t6429 n7040 n6430 R=3.315e+00 
R7039t4146 n7040 n4147 R=2.129e+02 
R7039t6996 n7040 n6997 R=1.118e+01 
R7039t143 n7040 n144 R=3.630e+00 
R7039t5870 n7040 n5871 R=9.114e+00 
R7040t128 n7041 n129 R=2.443e+00 
R7040t4324 n7041 n4325 R=6.982e+00 
R7041t3320 n7042 n3321 R=1.793e+01 
R7041t5082 n7042 n5083 R=3.311e+00 
R7041t6689 n7042 n6690 R=4.216e+00 
R7041t5306 n7042 n5307 R=2.039e+02 
R7041t2081 n7042 n2082 R=1.437e+01 
R7042t4339 n7043 n4340 R=5.918e+00 
R7042t424 n7043 n425 R=1.066e+02 
R7042t6860 n7043 n6861 R=2.593e+02 
R7042t2216 n7043 n2217 R=8.748e+00 
R7042t6328 n7043 n6329 R=4.027e+00 
R7042t2512 n7043 n2513 R=2.530e+01 
R7043t3795 n7044 n3796 R=8.453e+00 
R7043t3702 n7044 n3703 R=8.689e+02 
R7043t268 n7044 n269 R=3.835e+01 
R7043t3330 n7044 n3331 R=9.361e+00 
R7043t3143 n7044 n3144 R=8.169e+00 
R7043t2017 n7044 n2018 R=3.867e+01 
R7043t6049 n7044 n6050 R=1.990e+01 
R7044t2448 n7045 n2449 R=3.411e+00 
R7044t77 n7045 n78 R=1.785e+00 
R7044t1689 n7045 n1690 R=7.611e+00 
R7045t478 n7046 n479 R=4.493e+00 
R7045t1223 n7046 n1224 R=2.805e+00 
R7045t6955 n7046 n6956 R=9.296e+00 
R7045t1053 n7046 n1054 R=9.099e+00 
R7046t3054 n7047 n3055 R=3.000e+01 
R7046t3710 n7047 n3711 R=3.092e+00 
R7046t5835 n7047 n5836 R=3.649e+00 
R7047t1770 n7048 n1771 R=6.917e+00 
R7047t6640 n7048 n6641 R=1.250e+01 
R7047t3868 n7048 n3869 R=1.070e+01 
R7047t4313 n7048 n4314 R=2.402e+00 
R7048t4587 n7049 n4588 R=4.821e+00 
R7048t1310 n7049 n1311 R=6.159e+00 
R7048t4302 n7049 n4303 R=1.429e+01 
R7048t5278 n7049 n5279 R=9.418e+00 
R7048t3387 n7049 n3388 R=6.440e+00 
R7049t280 n7050 n281 R=2.286e+00 
R7049t2243 n7050 n2244 R=3.877e+02 
R7049t6585 n7050 n6586 R=7.311e+00 
R7049t5484 n7050 n5485 R=4.031e+00 
R7049t3367 n7050 n3368 R=3.642e+01 
R7049t2094 n7050 n2095 R=2.013e+01 
R7050t5870 n7051 n5871 R=1.200e+01 
R7051t6473 n7052 n6474 R=3.956e+00 
R7051t6426 n7052 n6427 R=2.998e+01 
R7051t1554 n7052 n1555 R=1.540e+00 
R7051t3430 n7052 n3431 R=1.175e+01 
R7052t3557 n7053 n3558 R=5.332e+01 
R7052t3606 n7053 n3607 R=4.138e+00 
R7052t3009 n7053 n3010 R=9.717e+00 
R7052t4416 n7053 n4417 R=1.866e+01 
R7052t110 n7053 n111 R=6.296e+00 
R7052t4860 n7053 n4861 R=8.588e+00 
R7053t3522 n7054 n3523 R=2.637e+02 
R7053t5298 n7054 n5299 R=1.868e+00 
R7053t6592 n7054 n6593 R=1.468e+01 
R7053t6713 n7054 n6714 R=2.094e+00 
R7053t5348 n7054 n5349 R=4.005e+01 
R7053t1563 n7054 n1564 R=1.356e+01 
R7054t1596 n7055 n1597 R=1.842e+01 
R7054t6905 n7055 n6906 R=9.536e+00 
R7054t419 n7055 n420 R=6.219e+01 
R7055t5576 n7056 n5577 R=4.552e+00 
R7055t6730 n7056 n6731 R=5.060e+00 
R7055t754 n7056 n755 R=1.129e+01 
R7055t3178 n7056 n3179 R=1.178e+01 
R7056t872 n7057 n873 R=4.973e+00 
R7056t6605 n7057 n6606 R=1.005e+01 
R7056t1350 n7057 n1351 R=3.834e+00 
R7056t951 n7057 n952 R=5.094e+00 
R7057t5151 n7058 n5152 R=4.220e+00 
R7057t5565 n7058 n5566 R=7.423e+00 
R7057t3338 n7058 n3339 R=9.978e+01 
R7057t2035 n7058 n2036 R=1.520e+01 
R7058t5475 n7059 n5476 R=2.150e+00 
R7058t662 n7059 n663 R=8.064e+00 
R7058t6059 n7059 n6060 R=4.384e+00 
R7058t3800 n7059 n3801 R=4.255e+01 
R7059t864 n7060 n865 R=6.535e+00 
R7059t481 n7060 n482 R=3.363e+01 
R7059t4912 n7060 n4913 R=1.012e+01 
R7059t4342 n7060 n4343 R=9.260e+00 
R7060t2646 n7061 n2647 R=4.859e+00 
R7060t4650 n7061 n4651 R=4.117e+00 
R7060t5645 n7061 n5646 R=2.568e+01 
R7060t497 n7061 n498 R=2.518e+01 
R7060t5398 n7061 n5399 R=4.805e+00 
R7060t4906 n7061 n4907 R=9.297e+01 
R7061t1538 n7062 n1539 R=2.058e+00 
R7061t6790 n7062 n6791 R=2.647e+01 
R7061t3561 n7062 n3562 R=1.089e+01 
R7061t2421 n7062 n2422 R=1.729e+00 
R7062t1360 n7063 n1361 R=8.881e+00 
R7062t5059 n7063 n5060 R=3.981e+00 
R7062t1616 n7063 n1617 R=4.278e+00 
R7062t5103 n7063 n5104 R=4.970e+00 
R7063t1368 n7064 n1369 R=2.861e+00 
R7063t3353 n7064 n3354 R=1.178e+01 
R7064t4819 n7065 n4820 R=2.696e+01 
R7064t6599 n7065 n6600 R=2.065e+01 
R7064t3136 n7065 n3137 R=6.346e+00 
R7064t3692 n7065 n3693 R=3.245e+00 
R7064t1981 n7065 n1982 R=1.862e+02 
R7065t2535 n7066 n2536 R=8.470e+00 
R7065t2557 n7066 n2558 R=9.230e+01 
R7065t6064 n7066 n6065 R=3.075e+00 
R7065t364 n7066 n365 R=1.272e+02 
R7066t3562 n7067 n3563 R=5.989e+00 
R7066t118 n7067 n119 R=3.543e+00 
R7067t435 n7068 n436 R=1.856e+01 
R7067t1557 n7068 n1558 R=2.297e+01 
R7067t6986 n7068 n6987 R=2.511e+01 
R7067t937 n7068 n938 R=6.896e+00 
R7067t604 n7068 n605 R=1.842e+01 
R7067t6323 n7068 n6324 R=1.135e+02 
R7067t147 n7068 n148 R=3.292e+00 
R7068t2162 n7069 n2163 R=5.864e+00 
R7068t5043 n7069 n5044 R=1.215e+00 
R7068t2088 n7069 n2089 R=4.106e+01 
R7068t3967 n7069 n3968 R=3.669e+00 
R7069t2710 n7070 n2711 R=3.797e+01 
R7069t5178 n7070 n5179 R=4.980e+02 
R7069t1822 n7070 n1823 R=1.940e+01 
R7069t2485 n7070 n2486 R=7.302e+01 
R7069t2773 n7070 n2774 R=5.016e+00 
R7069t1520 n7070 n1521 R=3.388e+01 
R7069t2184 n7070 n2185 R=9.309e+00 
R7069t6760 n7070 n6761 R=3.239e+01 
R7069t3603 n7070 n3604 R=4.700e+00 
R7069t654 n7070 n655 R=9.466e+00 
R7070t4573 n7071 n4574 R=4.259e+00 
R7070t4685 n7071 n4686 R=2.950e+01 
R7070t991 n7071 n992 R=5.989e+00 
R7070t6111 n7071 n6112 R=1.169e+01 
R7070t7024 n7071 n7025 R=6.156e+00 
R7071t1241 n7072 n1242 R=2.322e+01 
R7071t6694 n7072 n6695 R=1.355e+01 
R7071t5664 n7072 n5665 R=8.615e+00 
R7071t557 n7072 n558 R=1.462e+01 
R7072t6444 n7073 n6445 R=2.499e+01 
R7072t2373 n7073 n2374 R=8.322e+00 
R7072t5306 n7073 n5307 R=5.915e+00 
R7072t263 n7073 n264 R=1.794e+01 
R7072t1901 n7073 n1902 R=3.706e+00 
R7073t6279 n7074 n6280 R=9.631e+00 
R7073t6788 n7074 n6789 R=2.785e+00 
R7073t3328 n7074 n3329 R=2.438e+00 
R7073t4973 n7074 n4974 R=1.186e+01 
R7074t6234 n7075 n6235 R=1.212e+01 
R7075t5959 n7076 n5960 R=1.620e+01 
R7075t6546 n7076 n6547 R=1.173e+01 
R7075t5680 n7076 n5681 R=1.207e+01 
R7075t84 n7076 n85 R=1.005e+01 
R7076t2259 n7077 n2260 R=4.302e+00 
R7076t2810 n7077 n2811 R=1.561e+02 
R7076t6675 n7077 n6676 R=3.238e+01 
R7076t953 n7077 n954 R=1.883e+00 
R7077t5285 n7078 n5286 R=7.265e+02 
R7078t1531 n7079 n1532 R=9.119e+02 
R7078t1609 n7079 n1610 R=3.025e+00 
R7078t171 n7079 n172 R=8.584e+00 
R7078t2288 n7079 n2289 R=7.442e+00 
R7079t233 n7080 n234 R=5.953e+00 
R7079t2155 n7080 n2156 R=8.247e+00 
R7079t6792 n7080 n6793 R=4.632e+00 
R7079t4111 n7080 n4112 R=2.231e+01 
R7080t187 n7081 n188 R=3.083e+00 
R7080t5329 n7081 n5330 R=2.658e+02 
R7080t4924 n7081 n4925 R=1.681e+01 
R7080t4266 n7081 n4267 R=4.110e+00 
R7081t2876 n7082 n2877 R=4.310e+00 
R7081t6751 n7082 n6752 R=3.343e+00 
R7081t5238 n7082 n5239 R=1.768e+01 
R7081t6682 n7082 n6683 R=4.919e+00 
R7082t705 n7083 n706 R=4.389e+00 
R7082t1226 n7083 n1227 R=2.258e+01 
R7082t2229 n7083 n2230 R=1.146e+01 
R7082t1864 n7083 n1865 R=1.183e+01 
R7082t6452 n7083 n6453 R=5.197e+00 
R7082t149 n7083 n150 R=6.452e+00 
R7083t5945 n7084 n5946 R=1.223e+01 
R7083t875 n7084 n876 R=2.659e+00 
R7083t6773 n7084 n6774 R=1.240e+02 
R7083t2353 n7084 n2354 R=1.408e+01 
R7084t4540 n7085 n4541 R=2.790e+00 
R7084t6974 n7085 n6975 R=5.618e+00 
R7084t4548 n7085 n4549 R=8.083e+02 
R7084t5811 n7085 n5812 R=9.443e+01 
R7084t4984 n7085 n4985 R=3.954e+00 
R7084t1177 n7085 n1178 R=9.940e+00 
R7085t5661 n7086 n5662 R=1.890e+01 
R7085t2124 n7086 n2125 R=2.367e+00 
R7085t1487 n7086 n1488 R=7.309e+01 
R7085t5193 n7086 n5194 R=4.047e+00 
R7086t3071 n7087 n3072 R=1.115e+01 
R7086t5670 n7087 n5671 R=1.056e+01 
R7086t3581 n7087 n3582 R=1.758e+02 
R7086t4144 n7087 n4145 R=1.955e+01 
R7086t5525 n7087 n5526 R=2.898e+00 
R7086t4952 n7087 n4953 R=8.511e+00 
R7086t2644 n7087 n2645 R=4.401e+00 
R7087t249 n7088 n250 R=3.306e+00 
R7087t1751 n7088 n1752 R=8.436e+02 
R7087t6396 n7088 n6397 R=9.837e+00 
R7087t1298 n7088 n1299 R=6.523e+00 
R7088t569 n7089 n570 R=4.989e+00 
R7088t3585 n7089 n3586 R=8.047e+00 
R7088t3459 n7089 n3460 R=3.936e+00 
R7089t2051 n7090 n2052 R=1.005e+02 
R7089t4294 n7090 n4295 R=5.352e+00 
R7089t5370 n7090 n5371 R=1.221e+02 
R7089t2595 n7090 n2596 R=7.593e+00 
R7089t3890 n7090 n3891 R=9.697e+00 
R7090t2494 n7091 n2495 R=1.545e+01 
R7090t4893 n7091 n4894 R=9.572e+00 
R7090t4887 n7091 n4888 R=3.660e+00 
R7090t6069 n7091 n6070 R=3.354e+00 
R7091t2242 n7092 n2243 R=2.415e+01 
R7091t3774 n7092 n3775 R=5.890e+00 
R7091t3163 n7092 n3164 R=3.618e+02 
R7091t2347 n7092 n2348 R=9.214e+00 
R7092t3157 n7093 n3158 R=4.382e+00 
R7092t4347 n7093 n4348 R=8.122e+00 
R7093t6350 n7094 n6351 R=4.097e+00 
R7093t1423 n7094 n1424 R=1.543e+01 
R7093t3121 n7094 n3122 R=9.482e+01 
R7094t383 n7095 n384 R=7.545e+00 
R7094t4130 n7095 n4131 R=1.835e+02 
R7094t2460 n7095 n2461 R=2.459e+00 
R7094t1474 n7095 n1475 R=4.465e+01 
R7094t6276 n7095 n6277 R=2.970e+00 
R7095t3505 n7096 n3506 R=6.869e+00 
R7095t6902 n7096 n6903 R=1.155e+01 
R7096t2987 n7097 n2988 R=4.766e+00 
R7096t1255 n7097 n1256 R=4.579e+00 
R7097t1675 n7098 n1676 R=8.845e+00 
R7097t4945 n7098 n4946 R=1.089e+00 
R7097t4715 n7098 n4716 R=6.133e+00 
R7097t5627 n7098 n5628 R=1.335e+01 
R7097t6542 n7098 n6543 R=2.052e+01 
R7098t4358 n7099 n4359 R=9.108e+00 
R7098t2185 n7099 n2186 R=3.257e+01 
R7098t2187 n7099 n2188 R=4.287e+00 
R7098t2474 n7099 n2475 R=9.466e+00 
R7099t2049 n7100 n2050 R=1.130e+01 
R7099t6990 n7100 n6991 R=6.149e+00 
R7099t5714 n7100 n5715 R=5.393e+00 
R7099t3197 n7100 n3198 R=5.060e+01 
R7100t763 n7101 n764 R=3.087e+01 
R7100t1446 n7101 n1447 R=5.510e+01 
R7100t6497 n7101 n6498 R=5.042e+00 
R7100t586 n7101 n587 R=7.799e+00 
R7100t1590 n7101 n1591 R=2.042e+00 
R7100t6466 n7101 n6467 R=2.502e+01 
R7101t331 n7102 n332 R=1.490e+01 
R7101t657 n7102 n658 R=3.005e+00 
R7101t2076 n7102 n2077 R=1.434e+01 
R7101t6294 n7102 n6295 R=5.295e+00 
R7102t3530 n7103 n3531 R=2.490e+00 
R7102t3945 n7103 n3946 R=4.772e+01 
R7102t4630 n7103 n4631 R=3.655e+00 
R7103t6099 n7104 n6100 R=2.245e+01 
R7103t6904 n7104 n6905 R=3.468e+00 
R7103t5919 n7104 n5920 R=8.768e+00 
R7103t932 n7104 n933 R=6.541e+00 
R7104t178 n7105 n179 R=3.311e+01 
R7104t5132 n7105 n5133 R=6.407e+00 
R7104t1811 n7105 n1812 R=4.551e+00 
R7104t6939 n7105 n6940 R=6.170e+01 
R7104t1409 n7105 n1410 R=7.701e+02 
R7104t5641 n7105 n5642 R=1.670e+01 
R7104t6181 n7105 n6182 R=8.781e+00 
R7104t1320 n7105 n1321 R=5.597e+00 
R7105t848 n7106 n849 R=3.644e+00 
R7105t2287 n7106 n2288 R=6.092e+00 
R7105t3454 n7106 n3455 R=1.253e+01 
R7105t3472 n7106 n3473 R=2.928e+00 
R7106t2008 n7107 n2009 R=7.344e+00 
R7106t5994 n7107 n5995 R=6.325e+00 
R7106t5631 n7107 n5632 R=3.846e+00 
R7106t6865 n7107 n6866 R=8.339e+01 
R7106t3982 n7107 n3983 R=5.039e+00 
R7106t5744 n7107 n5745 R=1.196e+01 
R7107t1228 n7108 n1229 R=5.033e+00 
R7107t5391 n7108 n5392 R=3.283e+02 
R7107t2090 n7108 n2091 R=3.954e+00 
R7107t4747 n7108 n4748 R=6.218e+00 
R7108t1190 n7109 n1191 R=1.127e+01 
R7108t3420 n7109 n3421 R=7.372e+00 
R7108t5657 n7109 n5658 R=4.975e+00 
R7108t5862 n7109 n5863 R=1.889e+01 
R7108t906 n7109 n907 R=1.243e+01 
R7108t6990 n7109 n6991 R=2.017e+01 
R7109t51 n7110 n52 R=4.681e+01 
R7109t367 n7110 n368 R=5.044e+00 
R7109t2003 n7110 n2004 R=8.644e+00 
R7109t5935 n7110 n5936 R=4.137e+00 
R7109t2001 n7110 n2002 R=5.131e+01 
R7109t4825 n7110 n4826 R=2.122e+01 
R7110t1042 n7111 n1043 R=4.353e+00 
R7110t2537 n7111 n2538 R=5.458e+02 
R7110t6142 n7111 n6143 R=1.149e+01 
R7111t2417 n7112 n2418 R=6.948e+00 
R7111t5149 n7112 n5150 R=6.130e+00 
R7111t3983 n7112 n3984 R=5.701e+00 
R7112t1576 n7113 n1577 R=3.784e+00 
R7112t5802 n7113 n5803 R=7.603e+00 
R7112t5072 n7113 n5073 R=4.550e+00 
R7112t6032 n7113 n6033 R=1.221e+01 
R7112t2609 n7113 n2610 R=6.317e+00 
R7113t4639 n7114 n4640 R=5.029e+00 
R7113t6603 n7114 n6604 R=3.178e+00 
R7113t4515 n7114 n4516 R=1.335e+00 
R7113t1812 n7114 n1813 R=1.644e+01 
R7114t5087 n7115 n5088 R=4.924e+00 
R7114t2585 n7115 n2586 R=6.359e+00 
R7114t6114 n7115 n6115 R=4.589e+00 
R7115t5311 n7116 n5312 R=5.570e+00 
R7115t3195 n7116 n3196 R=1.952e+02 
R7115t3953 n7116 n3954 R=1.919e+01 
R7115t3652 n7116 n3653 R=6.982e+01 
R7116t5323 n7117 n5324 R=4.996e+01 
R7116t6210 n7117 n6211 R=8.718e+00 
R7116t4964 n7117 n4965 R=7.285e+00 
R7116t4323 n7117 n4324 R=4.292e+00 
R7117t1396 n7118 n1397 R=3.999e+00 
R7117t5580 n7118 n5581 R=6.940e+00 
R7117t796 n7118 n797 R=1.309e+01 
R7117t1642 n7118 n1643 R=2.922e+01 
R7117t328 n7118 n329 R=8.128e+00 
R7117t5760 n7118 n5761 R=5.773e+02 
R7118t322 n7119 n323 R=2.189e+00 
R7118t1691 n7119 n1692 R=3.214e+01 
R7118t2523 n7119 n2524 R=7.500e+00 
R7118t199 n7119 n200 R=5.237e+01 
R7118t373 n7119 n374 R=4.412e+00 
R7119t646 n7120 n647 R=8.297e+00 
R7119t6352 n7120 n6353 R=6.319e+00 
R7119t1251 n7120 n1252 R=3.200e+00 
R7119t3939 n7120 n3940 R=5.081e+00 
R7120t2540 n7121 n2541 R=3.315e+00 
R7120t5742 n7121 n5743 R=4.715e+00 
R7120t6408 n7121 n6409 R=1.558e+02 
R7120t6432 n7121 n6433 R=1.617e+01 
R7121t1182 n7122 n1183 R=3.075e+00 
R7121t4553 n7122 n4554 R=7.414e+00 
R7121t2073 n7122 n2074 R=1.271e+01 
R7121t1886 n7122 n1887 R=2.119e+00 
R7122t3450 n7123 n3451 R=3.487e+00 
R7122t4858 n7123 n4859 R=6.310e+00 
R7122t5047 n7123 n5048 R=6.676e+01 
R7122t6980 n7123 n6981 R=1.703e+01 
R7122t2516 n7123 n2517 R=1.648e+01 
R7123t5957 n7124 n5958 R=1.077e+01 
R7123t1333 n7124 n1334 R=2.673e+00 
R7124t1362 n7125 n1363 R=4.825e+00 
R7124t2794 n7125 n2795 R=1.315e+01 
R7124t5446 n7125 n5447 R=7.891e+00 
R7124t2636 n7125 n2637 R=8.418e+00 
R7124t1269 n7125 n1270 R=1.505e+01 
R7125t2340 n7126 n2341 R=7.330e+01 
R7125t5583 n7126 n5584 R=3.109e+00 
R7125t2904 n7126 n2905 R=2.438e+01 
R7125t341 n7126 n342 R=5.532e+00 
R7126t5978 n7127 n5979 R=1.517e+01 
R7126t6925 n7127 n6926 R=8.385e+00 
R7126t4822 n7127 n4823 R=2.891e+00 
R7127t2076 n7128 n2077 R=5.032e+01 
R7127t7101 n7128 n7102 R=6.972e+00 
R7127t3033 n7128 n3034 R=3.702e+00 
R7127t1233 n7128 n1234 R=1.607e+01 
R7127t6294 n7128 n6295 R=5.961e+00 
R7128t1679 n7129 n1680 R=4.006e+01 
R7128t1721 n7129 n1722 R=4.808e+00 
R7128t2942 n7129 n2943 R=5.205e+00 
R7128t5303 n7129 n5304 R=9.564e+00 
R7129t5237 n7130 n5238 R=1.072e+01 
R7129t6709 n7130 n6710 R=9.491e+00 
R7129t2723 n7130 n2724 R=7.654e+01 
R7129t1257 n7130 n1258 R=1.038e+01 
R7130t820 n7131 n821 R=1.092e+01 
R7130t1006 n7131 n1007 R=3.186e+00 
R7130t2791 n7131 n2792 R=4.229e+00 
R7130t6652 n7131 n6653 R=1.387e+01 
R7130t5335 n7131 n5336 R=2.871e+01 
R7131t6895 n7132 n6896 R=3.544e+01 
R7131t2790 n7132 n2791 R=4.636e+00 
R7131t2831 n7132 n2832 R=2.379e+01 
R7132t889 n7133 n890 R=4.364e+00 
R7132t975 n7133 n976 R=1.949e+01 
R7132t56 n7133 n57 R=1.395e+01 
R7132t3226 n7133 n3227 R=4.871e+00 
R7132t6422 n7133 n6423 R=6.404e+00 
R7133t1512 n7134 n1513 R=1.760e+00 
R7133t3733 n7134 n3734 R=7.152e+01 
R7133t3261 n7134 n3262 R=4.718e+01 
R7133t1860 n7134 n1861 R=3.721e+00 
R7133t6810 n7134 n6811 R=5.662e+00 
R7134t2852 n7135 n2853 R=3.679e+00 
R7134t419 n7135 n420 R=1.044e+01 
R7135t6299 n7136 n6300 R=5.552e+00 
R7135t4610 n7136 n4611 R=3.961e+00 
R7135t2076 n7136 n2077 R=1.337e+02 
R7135t797 n7136 n798 R=1.452e+01 
R7136t5880 n7137 n5881 R=6.076e+00 
R7136t3261 n7137 n3262 R=5.656e+00 
R7137t3422 n7138 n3423 R=6.999e+00 
R7137t6954 n7138 n6955 R=4.311e+00 
R7137t3415 n7138 n3416 R=7.662e+00 
R7138t3476 n7139 n3477 R=2.015e+00 
R7138t2734 n7139 n2735 R=5.315e+01 
R7138t323 n7139 n324 R=5.528e+00 
R7138t3342 n7139 n3343 R=9.724e+00 
R7139t1705 n7140 n1706 R=7.741e+00 
R7139t4476 n7140 n4477 R=5.133e+01 
R7139t2039 n7140 n2040 R=4.804e+00 
R7139t6518 n7140 n6519 R=1.982e+01 
R7140t2340 n7141 n2341 R=3.691e+00 
R7140t7125 n7141 n7126 R=3.942e+00 
R7140t1323 n7141 n1324 R=2.223e+01 
R7140t6856 n7141 n6857 R=3.397e+00 
R7140t2904 n7141 n2905 R=9.444e+00 
R7141t1246 n7142 n1247 R=1.086e+02 
R7141t3752 n7142 n3753 R=5.657e+01 
R7141t847 n7142 n848 R=2.890e+00 
R7141t4998 n7142 n4999 R=2.835e+00 
R7142t4406 n7143 n4407 R=2.176e+00 
R7142t6661 n7143 n6662 R=1.390e+01 
R7142t1289 n7143 n1290 R=4.072e+00 
R7142t2230 n7143 n2231 R=3.198e+01 
R7142t3775 n7143 n3776 R=1.495e+01 
R7143t3534 n7144 n3535 R=3.453e+00 
R7143t5110 n7144 n5111 R=6.669e+00 
R7143t5695 n7144 n5696 R=9.886e+00 
R7143t2360 n7144 n2361 R=7.160e+00 
R7143t6215 n7144 n6216 R=1.057e+01 
R7143t2546 n7144 n2547 R=2.140e+01 
R7144t921 n7145 n922 R=1.955e+01 
R7144t1173 n7145 n1174 R=7.153e+01 
R7144t2343 n7145 n2344 R=4.326e+00 
R7144t5934 n7145 n5935 R=1.117e+01 
R7144t1046 n7145 n1047 R=1.036e+01 
R7144t408 n7145 n409 R=2.028e+01 
R7144t3364 n7145 n3365 R=1.329e+01 
R7145t2770 n7146 n2771 R=6.794e+00 
R7145t1786 n7146 n1787 R=3.854e+00 
R7145t5838 n7146 n5839 R=1.005e+01 
R7145t1156 n7146 n1157 R=1.342e+01 
R7145t5329 n7146 n5330 R=2.600e+01 
R7145t5903 n7146 n5904 R=4.711e+00 
R7145t1387 n7146 n1388 R=1.511e+03 
R7146t4904 n7147 n4905 R=2.087e+01 
R7146t672 n7147 n673 R=1.751e+01 
R7146t3160 n7147 n3161 R=9.974e+00 
R7147t46 n7148 n47 R=1.732e+01 
R7147t6645 n7148 n6646 R=8.391e+00 
R7147t6284 n7148 n6285 R=1.866e+00 
R7147t5195 n7148 n5196 R=6.183e+03 
R7147t691 n7148 n692 R=1.604e+01 
R7147t5917 n7148 n5918 R=3.429e+00 
R7148t6838 n7149 n6839 R=1.033e+01 
R7148t2181 n7149 n2182 R=2.198e+00 
R7148t566 n7149 n567 R=3.495e+01 
R7148t520 n7149 n521 R=6.520e+00 
R7149t2165 n7150 n2166 R=1.981e+00 
R7149t5749 n7150 n5750 R=1.617e+01 
R7149t3761 n7150 n3762 R=9.039e+01 
R7149t3046 n7150 n3047 R=2.174e+00 
R7150t2405 n7151 n2406 R=1.867e+01 
R7150t3131 n7151 n3132 R=3.387e+01 
R7150t1302 n7151 n1303 R=8.341e+00 
R7150t2745 n7151 n2746 R=5.748e+00 
R7150t4779 n7151 n4780 R=4.815e+01 
R7150t6104 n7151 n6105 R=3.951e+00 
R7150t5990 n7151 n5991 R=1.080e+01 
R7151t855 n7152 n856 R=2.724e+01 
R7151t3214 n7152 n3215 R=2.934e+00 
R7151t1412 n7152 n1413 R=6.693e+00 
R7151t960 n7152 n961 R=6.021e+00 
R7152t4277 n7153 n4278 R=1.975e+01 
R7152t4754 n7153 n4755 R=2.485e+00 
R7152t5879 n7153 n5880 R=1.325e+01 
R7152t1063 n7153 n1064 R=1.257e+01 
R7153t1633 n7154 n1634 R=3.617e+00 
R7153t4371 n7154 n4372 R=3.192e+00 
R7153t6250 n7154 n6251 R=5.321e+00 
R7153t3146 n7154 n3147 R=3.098e+01 
R7154t2007 n7155 n2008 R=1.020e+01 
R7154t4410 n7155 n4411 R=4.143e+00 
R7154t3458 n7155 n3459 R=1.418e+01 
R7154t5527 n7155 n5528 R=1.352e+01 
R7155t2492 n7156 n2493 R=1.673e+01 
R7155t6838 n7156 n6839 R=6.418e+00 
R7155t7148 n7156 n7149 R=1.187e+01 
R7156t3624 n7157 n3625 R=2.323e+01 
R7156t4304 n7157 n4305 R=1.026e+02 
R7156t6989 n7157 n6990 R=1.020e+01 
R7156t775 n7157 n776 R=6.007e+00 
R7157t534 n7158 n535 R=1.273e+01 
R7157t4999 n7158 n5000 R=1.883e+01 
R7157t2183 n7158 n2184 R=3.092e+00 
R7157t1370 n7158 n1371 R=1.073e+01 
R7158t4242 n7159 n4243 R=2.791e+01 
R7158t1043 n7159 n1044 R=1.201e+01 
R7158t5528 n7159 n5529 R=1.542e+01 
R7158t4328 n7159 n4329 R=2.741e+00 
R7159t5200 n7160 n5201 R=9.296e+00 
R7159t4729 n7160 n4730 R=1.641e+01 
R7159t4040 n7160 n4041 R=9.169e+00 
R7159t5745 n7160 n5746 R=5.807e+01 
R7159t6677 n7160 n6678 R=1.030e+01 
R7159t311 n7160 n312 R=2.288e+00 
R7160t4286 n7161 n4287 R=9.042e+00 
R7160t3957 n7161 n3958 R=3.965e+00 
R7161t4442 n7162 n4443 R=3.660e+00 
R7161t5931 n7162 n5932 R=8.691e+00 
R7161t1444 n7162 n1445 R=7.887e+01 
R7161t653 n7162 n654 R=4.854e+01 
R7162t1410 n7163 n1411 R=7.510e+00 
R7162t6170 n7163 n6171 R=2.337e+00 
R7162t5302 n7163 n5303 R=3.754e+00 
R7162t2410 n7163 n2411 R=2.183e+01 
R7163t2960 n7164 n2961 R=1.237e+02 
R7163t161 n7164 n162 R=2.103e+00 
R7164t1178 n7165 n1179 R=4.812e+01 
R7164t4195 n7165 n4196 R=3.180e+01 
R7164t4271 n7165 n4272 R=2.941e+00 
R7164t6311 n7165 n6312 R=1.435e+02 
R7164t5319 n7165 n5320 R=4.542e+00 
R7164t438 n7165 n439 R=2.390e+00 
R7165t6610 n7166 n6611 R=1.043e+01 
R7165t968 n7166 n969 R=2.099e+01 
R7165t608 n7166 n609 R=5.835e+00 
R7165t5857 n7166 n5858 R=2.231e+01 
R7165t182 n7166 n183 R=7.096e+00 
R7166t5643 n7167 n5644 R=1.575e+01 
R7166t323 n7167 n324 R=3.833e+00 
R7166t5800 n7167 n5801 R=4.640e+00 
R7167t4776 n7168 n4777 R=7.528e+00 
R7167t1757 n7168 n1758 R=2.761e+00 
R7167t2043 n7168 n2044 R=1.427e+01 
R7167t3702 n7168 n3703 R=3.076e+02 
R7168t4975 n1 n4976 R=3.709e+01 
R7169t6433 n7170 n6434 R=2.452e+01 
R7169t3180 n7170 n3181 R=5.347e+01 
R7169t2520 n7170 n2521 R=5.970e+00 
R7169t6125 n7170 n6126 R=4.196e+00 
R7169t5562 n7170 n5563 R=6.660e+00 
R7170t1398 n7171 n1399 R=1.940e+01 
R7170t4516 n7171 n4517 R=9.728e+00 
R7170t4225 n7171 n4226 R=5.521e+00 
R7171t1480 n7172 n1481 R=2.252e+01 
R7171t2929 n7172 n2930 R=1.304e+01 
R7171t6943 n7172 n6944 R=4.371e+00 
R7172t4099 n7173 n4100 R=1.199e+01 
R7172t6983 n7173 n6984 R=7.899e+00 
R7172t307 n7173 n308 R=4.306e+00 
R7173t2960 n7174 n2961 R=1.217e+01 
R7173t7163 n7174 n7164 R=2.159e+00 
R7173t3792 n7174 n3793 R=5.477e+00 
R7173t6491 n7174 n6492 R=1.441e+01 
R7174t1502 n7175 n1503 R=3.551e+00 
R7174t2261 n7175 n2262 R=2.502e+01 
R7174t3940 n7175 n3941 R=2.187e+01 
R7174t2345 n7175 n2346 R=7.274e+00 
R7174t78 n7175 n79 R=1.525e+01 
R7174t4398 n7175 n4399 R=9.130e+00 
R7175t863 n7176 n864 R=3.763e+00 
R7175t3307 n7176 n3308 R=4.251e+02 
R7175t487 n7176 n488 R=3.819e+00 
R7175t1717 n7176 n1718 R=1.139e+01 
R7176t1275 n7177 n1276 R=6.898e+00 
R7176t5570 n7177 n1 R=2.720e+00 
R7176t3366 n7177 n3367 R=4.551e+00 
R7177t3797 n7178 n3798 R=9.830e+01 
R7177t4298 n7178 n4299 R=1.890e+00 
R7177t6478 n7178 n6479 R=2.060e+01 
R7178t581 n7179 n582 R=5.997e+02 
R7178t619 n7179 n620 R=1.411e+02 
R7178t2056 n7179 n2057 R=3.455e+00 
R7178t5763 n7179 n5764 R=1.425e+01 
R7178t7030 n7179 n7031 R=5.043e+01 
R7178t2132 n7179 n2133 R=1.305e+01 
R7178t1382 n7179 n1383 R=1.713e+01 
R7179t1191 n7180 n1192 R=1.193e+01 
R7179t3350 n7180 n3351 R=1.808e+01 
R7179t3996 n7180 n3997 R=7.663e+00 
R7179t5198 n7180 n5199 R=5.492e+01 
R7179t6937 n7180 n6938 R=8.217e+00 
R7179t681 n7180 n682 R=3.089e+01 
R7179t1640 n7180 n1641 R=3.486e+00 
R7180t2787 n7181 n2788 R=1.103e+01 
R7180t3138 n7181 n3139 R=1.106e+01 
R7180t6865 n7181 n6866 R=5.224e+00 
R7180t3749 n7181 n3750 R=5.462e+00 
R7181t4146 n7182 n4147 R=1.069e+01 
R7181t6996 n7182 n6997 R=1.956e+00 
R7181t143 n7182 n144 R=1.251e+01 
R7181t6723 n7182 n6724 R=1.802e+02 
R7182t4897 n7183 n4898 R=2.860e+01 
R7182t5257 n7183 n5258 R=6.271e+01 
R7182t5426 n7183 n5427 R=6.073e+00 
R7182t1781 n7183 n1782 R=3.273e+00 
R7183t3024 n7184 n3025 R=4.641e+01 
R7183t6778 n7184 n6779 R=1.491e+01 
R7183t6282 n7184 n6283 R=2.554e+00 
R7183t2514 n7184 n2515 R=1.176e+01 
R7184t669 n7185 n670 R=3.033e+00 
R7184t2105 n7185 n2106 R=2.180e+01 
R7184t1141 n7185 n1142 R=2.609e+00 
R7185t454 n7186 n455 R=2.535e+01 
R7185t658 n7186 n659 R=8.453e+00 
R7185t3424 n7186 n3425 R=3.660e+00 
R7185t4674 n7186 n4675 R=3.498e+01 
R7185t35 n7186 n36 R=1.190e+01 
R7185t445 n7186 n446 R=2.284e+01 
R7185t133 n7186 n134 R=6.987e+00 
R7186t20 n7187 n21 R=1.686e+01 
R7186t2737 n7187 n2738 R=7.142e+00 
R7186t1807 n7187 n1808 R=3.034e+01 
R7186t6555 n7187 n6556 R=3.525e+00 
R7186t306 n7187 n307 R=1.243e+01 
R7187t6305 n7188 n6306 R=3.563e+00 
R7187t2415 n7188 n2416 R=9.709e+00 
R7187t4195 n7188 n4196 R=1.061e+01 
R7187t4271 n7188 n4272 R=4.252e+00 
R7188t6928 n7189 n6929 R=1.215e+01 
R7188t4751 n7189 n4752 R=2.834e+00 
R7188t841 n7189 n842 R=1.706e+01 
R7188t2391 n7189 n2392 R=1.616e+01 
R7188t1978 n7189 n1979 R=3.708e+01 
R7188t3099 n7189 n3100 R=3.066e+00 
R7189t269 n7190 n270 R=2.910e+00 
R7189t6975 n7190 n6976 R=5.463e+00 
R7189t3119 n7190 n3120 R=2.849e+00 
R7190t1891 n7191 n1892 R=6.466e+00 
R7190t6559 n7191 n6560 R=2.752e+00 
R7190t3270 n7191 n3271 R=2.845e+02 
R7190t1624 n7191 n1625 R=8.508e+00 
R7190t5881 n7191 n5882 R=8.824e+00 
R7190t3583 n7191 n3584 R=9.579e+00 
R7191t4822 n7192 n4823 R=4.301e+00 
R7191t7126 n7192 n7127 R=2.307e+01 
R7191t5978 n7192 n5979 R=5.442e+00 
R7191t2837 n7192 n2838 R=1.489e+01 
R7191t3422 n7192 n3423 R=1.287e+02 
R7191t5239 n7192 n5240 R=4.973e+00 
R7191t2816 n7192 n2817 R=7.239e+00 
R7191t5950 n7192 n5951 R=1.758e+02 
R7192t4724 n7193 n4725 R=4.454e+00 
R7192t5995 n7193 n5996 R=2.769e+00 
R7193t4239 n7194 n4240 R=4.139e+02 
R7193t5828 n7194 n5829 R=2.248e+00 
R7193t835 n7194 n836 R=1.028e+01 
R7193t3045 n7194 n3046 R=2.865e+00 
R7194t312 n7195 n313 R=4.335e+00 
R7194t1578 n7195 n1579 R=1.256e+01 
R7194t244 n7195 n245 R=4.351e+00 
R7194t6650 n7195 n6651 R=1.122e+01 
R7194t467 n7195 n468 R=5.582e+00 
R7195t5332 n7196 n5333 R=6.868e+01 
R7195t5665 n7196 n5666 R=1.689e+00 
R7195t5847 n7196 n5848 R=1.815e+01 
R7195t1221 n7196 n1222 R=4.067e+01 
R7195t3496 n7196 n3497 R=1.228e+01 
R7195t6108 n7196 n6109 R=1.854e+01 
R7196t3723 n7197 n3724 R=1.069e+01 
R7196t4589 n7197 n4590 R=5.144e+00 
R7196t3962 n7197 n3963 R=8.433e+00 
R7197t2442 n7198 n2443 R=8.806e+01 
R7197t3697 n7198 n3698 R=4.014e+00 
R7197t5243 n7198 n1 R=7.889e+00 
R7197t2980 n7198 n2981 R=5.502e+01 
R7197t1500 n7198 n1501 R=3.828e+00 
R7198t1171 n7199 n1172 R=9.538e+00 
R7198t6082 n7199 n6083 R=1.768e+00 
R7198t884 n7199 n885 R=1.647e+01 
R7198t193 n7199 n194 R=3.542e+00 
R7198t5344 n7199 n5345 R=6.224e+01 
R7199t1325 n7200 n1326 R=1.857e+01 
R7199t6923 n7200 n6924 R=1.021e+01 
R7199t4287 n7200 n4288 R=6.584e+00 
R7199t2949 n7200 n2950 R=4.739e+00 
R7199t6247 n7200 n6248 R=1.184e+01 
R7199t5337 n7200 n5338 R=9.624e+00 
R7200t3188 n7201 n3189 R=1.373e+01 
R7200t6409 n7201 n6410 R=4.609e+00 
R7200t5360 n7201 n5361 R=9.762e+00 
R7200t6785 n7201 n6786 R=1.101e+01 
R7200t2121 n7201 n2122 R=9.245e+00 
R7201t604 n7202 n605 R=2.391e+00 
R7201t3547 n7202 n3548 R=5.072e+00 
R7202t188 n7203 n189 R=4.710e+00 
R7202t4906 n7203 n4907 R=7.627e+00 
R7202t6692 n7203 n6693 R=2.641e+01 
R7202t5398 n7203 n5399 R=3.450e+00 
R7202t7060 n7203 n7061 R=8.063e+00 
R7203t1161 n7204 n1162 R=2.959e+00 
R7203t1728 n7204 n1729 R=3.434e+00 
R7203t4982 n7204 n4983 R=3.973e+00 
R7204t4921 n7205 n4922 R=3.006e+00 
R7204t2154 n7205 n2155 R=4.433e+00 
R7204t3812 n7205 n3813 R=1.388e+01 
R7205t3101 n7206 n3102 R=7.140e+00 
R7205t1030 n7206 n1031 R=4.954e+00 
R7206t3221 n7207 n3222 R=5.705e+00 
R7206t6977 n7207 n6978 R=2.311e+01 
R7206t5500 n7207 n5501 R=7.696e+00 
R7206t4997 n7207 n4998 R=9.861e+00 
R7206t7002 n7207 n7003 R=7.984e+00 
R7207t4741 n7208 n4742 R=4.033e+00 
R7207t2899 n7208 n2900 R=7.940e+00 
R7207t5832 n7208 n5833 R=6.420e+01 
R7207t1433 n7208 n1434 R=3.362e+00 
R7208t982 n7209 n983 R=3.799e+01 
R7208t1568 n7209 n1569 R=1.983e+01 
R7208t7001 n7209 n7002 R=1.915e+01 
R7208t2848 n7209 n2849 R=1.027e+01 
R7208t1823 n7209 n1824 R=4.239e+00 
R7208t4353 n7209 n4354 R=1.159e+01 
R7209t5313 n7210 n5314 R=2.853e+01 
R7209t2352 n7210 n2353 R=3.989e+00 
R7209t5448 n7210 n5449 R=4.022e+00 
R7209t893 n7210 n894 R=8.734e+00 
R7210t391 n7211 n392 R=3.906e+00 
R7210t2355 n7211 n2356 R=3.440e+02 
R7210t6358 n7211 n6359 R=3.236e+00 
R7210t2125 n7211 n2126 R=2.031e+01 
R7210t3871 n7211 n3872 R=2.765e+01 
R7211t5812 n7212 n5813 R=6.869e+00 
R7211t7074 n7212 n7075 R=6.171e+01 
R7211t6234 n7212 n6235 R=3.727e+00 
R7211t6612 n7212 n6613 R=2.624e+01 
R7211t5431 n7212 n5432 R=2.872e+01 
R7211t1803 n7212 n1804 R=5.249e+00 
R7212t2336 n7213 n2337 R=8.375e+00 
R7212t3309 n7213 n3310 R=5.861e+00 
R7212t5185 n7213 n5186 R=3.524e+02 
R7212t2226 n7213 n2227 R=2.538e+01 
R7212t1808 n7213 n1809 R=2.435e+00 
R7212t6627 n7213 n6628 R=7.943e+00 
R7213t6229 n7214 n6230 R=1.488e+02 
R7213t7016 n7214 n7017 R=5.137e+00 
R7213t330 n7214 n331 R=1.533e+01 
R7213t3718 n7214 n3719 R=1.980e+01 
R7213t4572 n7214 n4573 R=8.090e+00 
R7213t30 n7214 n31 R=2.413e+01 
R7213t6454 n7214 n6455 R=3.156e+01 
R7213t6994 n7214 n6995 R=4.397e+00 
R7214t769 n7215 n770 R=1.858e+01 
R7214t2932 n7215 n2933 R=1.452e+02 
R7214t1764 n7215 n1765 R=4.544e+00 
R7215t5756 n7216 n5757 R=3.110e+00 
R7215t134 n7216 n135 R=1.302e+01 
R7215t7156 n7216 n7157 R=6.799e+00 
R7216t446 n7217 n447 R=3.952e+00 
R7216t6849 n7217 n6850 R=5.717e+00 
R7216t988 n7217 n989 R=1.020e+01 
R7216t472 n7217 n473 R=8.557e+00 
R7217t2684 n7218 n2685 R=2.219e+00 
R7217t3978 n7218 n3979 R=1.093e+01 
R7217t5373 n7218 n5374 R=2.042e+01 
R7217t5447 n7218 n5448 R=8.608e+01 
R7218t4117 n7219 n4118 R=2.355e+00 
R7218t4279 n7219 n4280 R=3.095e+01 
R7218t5280 n7219 n5281 R=2.447e+00 
R7218t1561 n7219 n1562 R=1.997e+01 
R7219t3403 n7220 n3404 R=4.456e+00 
R7219t4216 n7220 n4217 R=7.676e+00 
R7219t6890 n7220 n6891 R=1.954e+01 
R7219t3547 n7220 n3548 R=9.374e+00 
R7219t7201 n7220 n7202 R=2.292e+02 
R7220t3563 n7221 n3564 R=3.123e+01 
R7220t4878 n7221 n4879 R=1.153e+01 
R7220t5404 n7221 n5405 R=1.922e+01 
R7220t4253 n7221 n4254 R=2.857e+00 
R7220t3032 n7221 n3033 R=2.104e+01 
R7220t5186 n7221 n5187 R=2.678e+01 
R7220t4408 n7221 n4409 R=1.642e+01 
R7220t2742 n7221 n2743 R=1.939e+01 
R7220t1904 n7221 n1905 R=6.670e+00 
R7221t3402 n7222 n3403 R=2.191e+01 
R7221t6019 n7222 n6020 R=2.345e+01 
R7221t1133 n7222 n1134 R=5.914e+00 
R7221t3881 n7222 n3882 R=2.496e+03 
R7221t406 n7222 n407 R=3.359e+00 
R7222t1708 n7223 n1 R=5.340e+00 
R7222t3455 n7223 n3456 R=4.854e+00 
R7222t1827 n7223 n1828 R=8.468e+00 
R7222t4034 n7223 n4035 R=5.582e+00 
R7223t1339 n7224 n1340 R=3.016e+00 
R7223t3534 n7224 n3535 R=2.244e+01 
R7223t818 n7224 n819 R=1.436e+01 
R7223t5156 n7224 n5157 R=2.695e+00 
R7223t625 n7224 n626 R=2.883e+02 
R7223t27 n7224 n28 R=1.572e+01 
R7224t2843 n7225 n2844 R=2.057e+01 
R7224t5080 n7225 n5081 R=4.180e+00 
R7224t2435 n7225 n2436 R=2.804e+01 
R7224t891 n7225 n892 R=4.623e+01 
R7225t4877 n7226 n4878 R=1.628e+01 
R7225t207 n7226 n208 R=1.165e+01 
R7225t1481 n7226 n1482 R=3.031e+00 
R7225t1033 n7226 n1034 R=8.601e+00 
R7226t1155 n7227 n1156 R=1.539e+01 
R7226t1064 n7227 n1065 R=3.036e+00 
R7226t4537 n7227 n4538 R=1.044e+01 
R7226t4789 n7227 n4790 R=4.045e+01 
R7227t2240 n7228 n2241 R=3.794e+00 
R7227t5430 n7228 n5431 R=9.762e+00 
R7227t694 n7228 n695 R=4.084e+01 
R7227t525 n7228 n526 R=8.136e+00 
R7227t2685 n7228 n2686 R=6.177e+01 
R7228t542 n7229 n543 R=2.944e+00 
R7228t1081 n7229 n1082 R=1.564e+00 
R7228t3918 n7229 n3919 R=6.897e+00 
R7228t6852 n7229 n6853 R=1.057e+02 
R7229t1461 n7230 n1462 R=6.022e+00 
R7229t5008 n7230 n5009 R=1.589e+01 
R7229t713 n7230 n714 R=7.075e+00 
R7229t2202 n7230 n2203 R=4.873e+02 
R7229t651 n7230 n652 R=4.198e+00 
R7230t5743 n7231 n5744 R=4.372e+00 
R7230t5976 n7231 n5977 R=1.022e+01 
R7230t536 n7231 n537 R=3.837e+01 
R7230t3457 n7231 n3458 R=5.054e+01 
R7230t2951 n7231 n2952 R=8.702e+00 
R7230t58 n7231 n59 R=1.247e+01 
R7230t6669 n7231 n6670 R=9.400e+00 
R7231t322 n7232 n323 R=1.458e+01 
R7231t5486 n7232 n5487 R=4.330e+00 
R7231t7118 n7232 n7119 R=2.574e+01 
R7231t2523 n7232 n2524 R=5.417e+00 
R7231t4138 n7232 n4139 R=9.904e+01 
R7231t6177 n7232 n6178 R=1.125e+01 
R7232t2789 n7233 n2790 R=4.454e+00 
R7232t5678 n7233 n5679 R=8.434e+01 
R7232t4002 n7233 n4003 R=7.889e+00 
R7232t6873 n7233 n6874 R=5.036e+00 
R7232t2254 n7233 n2255 R=3.428e+00 
R7232t5682 n7233 n5683 R=4.505e+01 
R7233t7114 n7234 n7115 R=3.220e+01 
R7233t5087 n7234 n5088 R=2.750e+00 
R7233t965 n7234 n966 R=1.524e+02 
R7233t3962 n7234 n3963 R=8.245e+01 
R7233t7196 n7234 n7197 R=4.657e+00 
R7233t3723 n7234 n3724 R=8.261e+00 
R7234t2295 n7235 n2296 R=1.195e+01 
R7234t4574 n7235 n4575 R=4.866e+00 
R7234t2374 n7235 n2375 R=2.905e+01 
R7234t5579 n7235 n5580 R=3.841e+00 
R7234t1479 n7235 n1480 R=9.322e+00 
R7235t2971 n7236 n2972 R=2.522e+00 
R7235t4930 n7236 n4931 R=1.496e+01 
R7235t6823 n7236 n6824 R=7.592e+00 
R7235t1104 n7236 n1105 R=5.833e+00 
R7235t1389 n7236 n1390 R=1.661e+01 
R7236t5830 n7237 n5831 R=1.695e+01 
R7236t1103 n7237 n1104 R=5.094e+00 
R7236t6891 n7237 n6892 R=1.110e+01 
R7237t504 n7238 n505 R=2.478e+01 
R7237t2202 n7238 n2203 R=7.768e+00 
R7237t1926 n7238 n1927 R=2.900e+00 
R7237t1867 n7238 n1868 R=1.139e+01 
R7238t2765 n7239 n2766 R=9.349e+00 
R7238t1375 n7239 n1376 R=8.056e+02 
R7238t5939 n7239 n5940 R=6.153e+00 
R7239t4384 n7240 n4385 R=2.128e+01 
R7239t5642 n7240 n5643 R=4.353e+00 
R7239t6007 n7240 n6008 R=1.498e+01 
R7239t4786 n7240 n4787 R=5.195e+00 
R7239t4855 n7240 n4856 R=3.406e+02 
R7240t1726 n7241 n1727 R=2.946e+00 
R7240t6289 n7241 n6290 R=5.746e+00 
R7240t7080 n7241 n7081 R=3.650e+01 
R7240t187 n7241 n188 R=5.096e+00 
R7241t6352 n7242 n6353 R=1.920e+00 
R7241t6440 n7242 n6441 R=2.855e+01 
R7241t646 n7242 n647 R=2.619e+02 
R7241t6223 n7242 n6224 R=1.035e+01 
R7241t1963 n7242 n1964 R=1.682e+00 
R7241t6879 n7242 n6880 R=1.157e+02 
R7242t6766 n7243 n6767 R=2.295e+02 
R7242t2225 n7243 n2226 R=1.051e+01 
R7242t5912 n7243 n5913 R=1.029e+02 
R7242t569 n7243 n570 R=4.293e+01 
R7242t7088 n7243 n7089 R=6.009e+00 
R7242t3459 n7243 n3460 R=6.356e+01 
R7242t5873 n7243 n5874 R=6.943e+00 
R7242t2518 n7243 n2519 R=8.168e+00 
R7243t638 n7244 n639 R=1.051e+01 
R7243t1948 n7244 n1949 R=4.107e+01 
R7243t2134 n7244 n2135 R=1.611e+01 
R7243t7000 n7244 n7001 R=8.746e+00 
R7243t2536 n7244 n2537 R=5.493e+00 
R7243t2717 n7244 n2718 R=4.455e+01 
R7243t3458 n7244 n3459 R=2.914e+01 
R7243t7154 n7244 n7155 R=6.144e+00 
R7243t5356 n7244 n5357 R=8.225e+02 
R7244t1971 n7245 n1972 R=3.408e+00 
R7244t2856 n7245 n2857 R=1.341e+01 
R7244t5301 n7245 n5302 R=2.706e+00 
R7245t1536 n7246 n1537 R=1.809e+01 
R7245t4604 n7246 n4605 R=3.387e+01 
R7245t5842 n7246 n5843 R=3.555e+00 
R7245t802 n7246 n803 R=6.327e+00 
R7246t1045 n7247 n1046 R=1.186e+01 
R7246t3066 n7247 n3067 R=1.033e+02 
R7246t2799 n7247 n2800 R=1.802e+00 
R7247t1951 n7248 n1952 R=1.021e+01 
R7247t5354 n7248 n5355 R=1.261e+01 
R7247t218 n7248 n219 R=7.375e+00 
R7247t3229 n7248 n3230 R=3.240e+01 
R7248t4875 n7249 n4876 R=1.046e+01 
R7248t5663 n7249 n5664 R=8.173e+00 
R7248t4457 n7249 n4458 R=6.045e+00 
R7248t1704 n7249 n1705 R=7.055e+00 
R7248t5655 n7249 n5656 R=3.846e+00 
R7248t3821 n7249 n3822 R=2.894e+02 
R7248t3075 n7249 n3076 R=2.671e+01 
R7249t3261 n7250 n3262 R=3.775e+00 
R7249t7136 n7250 n7137 R=8.773e+01 
R7249t6357 n7250 n6358 R=6.712e+00 
R7250t3941 n7251 n3942 R=2.286e+01 
R7250t3173 n7251 n3174 R=1.735e+01 
R7250t4545 n7251 n4546 R=1.390e+01 
R7250t252 n7251 n253 R=8.250e+00 
R7250t1921 n7251 n1922 R=2.370e+01 
R7251t1691 n7252 n1692 R=3.197e+00 
R7251t6102 n7252 n6103 R=1.255e+01 
R7251t3029 n7252 n3030 R=6.660e+00 
R7251t373 n7252 n374 R=6.563e+00 
R7252t806 n7253 n807 R=5.877e+00 
R7252t4774 n7253 n4775 R=2.262e+01 
R7252t4449 n7253 n4450 R=4.231e+00 
R7252t4355 n7253 n4356 R=2.733e+00 
R7253t1566 n7254 n1567 R=4.523e+00 
R7253t3392 n7254 n3393 R=8.755e+00 
R7253t3605 n7254 n3606 R=2.959e+00 
R7253t5989 n7254 n5990 R=1.506e+01 
R7253t1686 n7254 n1687 R=7.368e+00 
R7254t2261 n7255 n2262 R=1.222e+01 
R7254t3940 n7255 n3941 R=3.154e+00 
R7254t3344 n7255 n3345 R=3.042e+00 
R7254t1875 n7255 n1876 R=7.647e+00 
R7255t441 n7256 n442 R=5.494e+00 
R7255t909 n7256 n910 R=8.701e+00 
R7255t6455 n7256 n6456 R=1.269e+01 
R7255t5003 n7256 n5004 R=1.480e+01 
R7255t4915 n7256 n4916 R=2.638e+00 
R7255t465 n7256 n466 R=8.553e+01 
R7255t868 n7256 n869 R=5.517e+00 
R7256t338 n7257 n339 R=1.036e+01 
R7256t1862 n7257 n1863 R=2.134e+01 
R7256t4756 n7257 n4757 R=3.265e+00 
R7256t3544 n7257 n3545 R=5.209e+00 
R7256t1263 n7257 n1264 R=4.906e+00 
R7257t2664 n7258 n2665 R=4.834e+00 
R7257t1763 n7258 n1764 R=2.179e+01 
R7257t2471 n7258 n2472 R=4.108e+01 
R7257t260 n7258 n261 R=1.358e+01 
R7257t3642 n7258 n3643 R=2.424e+01 
R7258t6186 n7259 n6187 R=9.731e+00 
R7258t6909 n7259 n6910 R=1.803e+01 
R7258t1475 n7259 n1476 R=4.162e+01 
R7258t73 n7259 n74 R=4.529e+00 
R7258t5814 n7259 n5815 R=9.924e+00 
R7258t2041 n7259 n2042 R=6.014e+01 
R7259t4162 n7260 n4163 R=1.550e+01 
R7259t3442 n7260 n3443 R=2.950e+00 
R7259t4801 n7260 n4802 R=1.641e+01 
R7259t678 n7260 n679 R=7.126e+00 
R7260t1422 n7261 n1423 R=4.713e+00 
R7260t6566 n7261 n6567 R=4.296e+00 
R7260t4482 n7261 n4483 R=3.392e+01 
R7260t6651 n7261 n6652 R=5.422e+00 
R7261t1057 n7262 n1058 R=3.061e+00 
R7261t5088 n7262 n5089 R=1.056e+01 
R7261t4928 n7262 n4929 R=1.644e+01 
R7261t3241 n7262 n3242 R=3.824e+00 
R7261t6183 n7262 n6184 R=1.358e+01 
R7262t3667 n7263 n3668 R=2.547e+01 
R7262t4553 n7263 n4554 R=1.047e+02 
R7262t4868 n7263 n4869 R=6.479e+00 
R7262t5348 n7263 n5349 R=4.701e+00 
R7262t7053 n7263 n7054 R=3.258e+02 
R7262t6713 n7263 n6714 R=5.336e+00 
R7262t1408 n7263 n1409 R=5.972e+00 
R7263t4492 n7264 n4493 R=3.782e+00 
R7263t5625 n7264 n5626 R=3.720e+00 
R7264t2310 n7265 n2311 R=1.885e+00 
R7264t6912 n7265 n6913 R=1.648e+01 
R7264t4372 n7265 n4373 R=1.485e+01 
R7264t3056 n7265 n3057 R=4.807e+00 
R7264t725 n7265 n726 R=9.234e+00 
R7265t2972 n7266 n2973 R=1.088e+01 
R7265t5678 n7266 n5679 R=2.235e+01 
R7265t2475 n7266 n2476 R=5.834e+00 
R7265t6913 n7266 n6914 R=7.962e+00 
R7265t2656 n7266 n2657 R=2.176e+01 
R7265t2873 n7266 n2874 R=1.791e+01 
R7265t127 n7266 n128 R=1.334e+01 
R7265t3466 n7266 n3467 R=5.099e+01 
R7265t3855 n7266 n3856 R=7.155e+00 
R7266t1095 n7267 n1096 R=8.320e+00 
R7266t5478 n7267 n5479 R=2.579e+00 
R7266t6130 n7267 n6131 R=2.206e+01 
R7266t6193 n7267 n6194 R=3.379e+00 
R7266t131 n7267 n132 R=7.508e+01 
R7266t4486 n7267 n4487 R=1.111e+01 
R7267t3234 n7268 n3235 R=6.178e+02 
R7267t2835 n7268 n2836 R=1.604e+01 
R7267t5875 n7268 n5876 R=5.007e+00 
R7267t5700 n7268 n5701 R=2.835e+00 
R7267t6841 n7268 n6842 R=4.353e+00 
R7268t1523 n7269 n1524 R=1.190e+01 
R7268t5610 n7269 n5611 R=4.167e+01 
R7268t1916 n7269 n1917 R=4.178e+00 
R7268t3523 n7269 n3524 R=1.346e+01 
R7269t19 n7270 n20 R=3.376e+01 
R7269t4847 n7270 n4848 R=1.735e+00 
R7269t2005 n7270 n2006 R=1.347e+01 
R7269t5444 n7270 n5445 R=5.831e+00 
R7270t4446 n7271 n4447 R=3.998e+01 
R7270t6344 n7271 n6345 R=2.623e+01 
R7270t6710 n7271 n6711 R=7.412e+00 
R7270t6155 n7271 n6156 R=6.149e+00 
R7270t3241 n7271 n3242 R=6.071e+00 
R7270t5217 n7271 n5218 R=3.968e+01 
R7270t2055 n7271 n2056 R=4.336e+00 
R7271t1073 n7272 n1074 R=2.869e+01 
R7271t7054 n7272 n7055 R=1.409e+01 
R7271t419 n7272 n420 R=4.100e+00 
R7271t6708 n7272 n6709 R=5.961e+00 
R7272t2165 n7273 n2166 R=4.958e+01 
R7272t5749 n7273 n5750 R=7.360e+00 
R7272t5630 n7273 n5631 R=4.165e+00 
R7272t4370 n7273 n4371 R=1.323e+01 
R7272t1833 n7273 n1834 R=6.196e+01 
R7272t782 n7273 n783 R=2.653e+00 
R7272t5542 n7273 n5543 R=4.618e+01 
R7273t281 n7274 n282 R=4.500e+00 
R7273t477 n7274 n478 R=6.198e+00 
R7273t351 n7274 n352 R=9.480e+01 
R7274t1334 n7275 n1335 R=4.169e+00 
R7274t2544 n7275 n2545 R=2.745e+01 
R7274t2894 n7275 n2895 R=3.758e+01 
R7274t5064 n7275 n5065 R=2.650e+00 
R7274t3870 n7275 n3871 R=2.628e+01 
R7274t36 n7275 n37 R=3.915e+01 
R7274t755 n7275 n756 R=4.864e+00 
R7275t1010 n7276 n1011 R=1.588e+00 
R7275t1949 n7276 n1950 R=3.751e+01 
R7276t1463 n7277 n1464 R=1.179e+01 
R7276t3409 n7277 n3410 R=2.356e+00 
R7276t5938 n7277 n5939 R=2.785e+00 
R7276t6475 n7277 n6476 R=1.776e+01 
R7276t3680 n7277 n3681 R=3.768e+01 
R7277t2886 n7278 n2887 R=2.532e+02 
R7277t3675 n7278 n3676 R=2.613e+00 
R7277t4986 n7278 n4987 R=3.394e+01 
R7278t2143 n7279 n2144 R=6.119e+01 
R7278t6580 n7279 n6581 R=6.242e+00 
R7278t3851 n7279 n3852 R=3.008e+01 
R7279t4082 n7280 n4083 R=1.418e+01 
R7279t5492 n7280 n5493 R=4.214e+00 
R7279t4774 n7280 n4775 R=2.887e+00 
R7279t433 n7280 n434 R=1.033e+01 
R7279t2628 n7280 n2629 R=1.664e+01 
R7280t5427 n7281 n5428 R=4.516e+00 
R7280t5945 n7281 n5946 R=3.843e+00 
R7280t6275 n7281 n6276 R=7.721e+00 
R7280t1605 n7281 n1606 R=1.693e+02 
R7281t180 n7282 n181 R=9.730e+00 
R7281t6336 n7282 n6337 R=2.854e+01 
R7281t6126 n7282 n6127 R=7.515e+00 
R7281t1457 n7282 n1458 R=3.362e+01 
R7281t4395 n7282 n4396 R=2.679e+01 
R7281t2883 n7282 n2884 R=1.126e+01 
R7281t6967 n7282 n6968 R=4.084e+00 
R7281t2341 n7282 n2342 R=2.105e+02 
R7282t3007 n7283 n3008 R=3.846e+00 
R7282t3686 n7283 n3687 R=6.201e+00 
R7282t3063 n7283 n3064 R=5.520e+02 
R7283t1121 n7284 n1122 R=4.214e+00 
R7283t6816 n7284 n6817 R=4.226e+00 
R7283t5369 n7284 n5370 R=1.858e+01 
R7283t2250 n7284 n2251 R=1.060e+02 
R7284t5151 n7285 n5152 R=4.769e+00 
R7284t5565 n7285 n5566 R=7.307e+00 
R7284t3338 n7285 n3339 R=7.095e+01 
R7284t1880 n7285 n1881 R=5.990e+01 
R7284t3919 n7285 n3920 R=1.753e+00 
R7284t3514 n7285 n3515 R=1.147e+03 
R7284t3464 n7285 n3465 R=1.233e+01 
R7285t2718 n7286 n2719 R=1.572e+01 
R7285t3765 n7286 n3766 R=1.991e+00 
R7285t6859 n7286 n6860 R=2.893e+01 
R7285t3532 n7286 n3533 R=1.227e+00 
R7285t556 n7286 n557 R=2.477e+01 
R7286t6800 n7287 n6801 R=2.575e+01 
R7286t2010 n7287 n2011 R=1.055e+01 
R7286t5448 n7287 n5449 R=1.178e+01 
R7286t7209 n7287 n7210 R=5.887e+01 
R7286t2352 n7287 n2353 R=3.127e+01 
R7286t563 n7287 n564 R=4.542e+00 
R7287t1639 n7288 n1640 R=5.968e+00 
R7287t483 n7288 n1 R=6.008e+00 
R7287t4969 n7288 n4970 R=5.472e+00 
R7288t6591 n7289 n6592 R=8.569e+00 
R7288t2559 n7289 n2560 R=2.353e+01 
R7288t7000 n7289 n7001 R=3.879e+01 
R7288t253 n7289 n254 R=5.051e+00 
R7288t2410 n7289 n2411 R=1.145e+02 
R7289t915 n7290 n916 R=1.009e+01 
R7289t5307 n7290 n5308 R=8.807e+00 
R7289t5447 n7290 n5448 R=4.661e+00 
R7289t2684 n7290 n2685 R=1.188e+01 
R7289t917 n7290 n918 R=5.648e+00 
R7290t996 n7291 n997 R=6.350e+00 
R7290t4935 n7291 n4936 R=1.517e+01 
R7290t1312 n7291 n1313 R=1.365e+01 
R7291t1038 n7292 n1039 R=4.123e+00 
R7291t1876 n7292 n1877 R=6.479e+00 
R7291t4155 n7292 n4156 R=3.243e+01 
R7291t2545 n7292 n2546 R=6.123e+00 
R7291t2685 n7292 n2686 R=2.059e+01 
R7291t1903 n7292 n1904 R=4.543e+00 
R7292t5900 n7293 n5901 R=2.132e+01 
R7292t6504 n7293 n6505 R=1.811e+01 
R7292t1872 n7293 n1873 R=3.393e+00 
R7292t3245 n7293 n3246 R=7.844e+00 
R7293t5369 n7294 n5370 R=3.581e+02 
R7293t1364 n7294 n1365 R=1.979e+01 
R7293t1517 n7294 n1518 R=7.946e+00 
R7293t4612 n7294 n4613 R=1.327e+01 
R7293t3657 n7294 n3658 R=6.497e+01 
R7294t909 n7295 n910 R=4.750e+00 
R7294t6455 n7295 n6456 R=2.052e+01 
R7294t1127 n7295 n1128 R=3.017e+00 
R7294t1766 n7295 n1767 R=3.617e+00 
R7294t5752 n7295 n5753 R=1.749e+01 
R7295t4418 n7296 n4419 R=1.017e+01 
R7295t6498 n7296 n6499 R=4.572e+00 
R7295t2772 n7296 n2773 R=1.815e+01 
R7295t6333 n7296 n6334 R=1.868e+01 
R7295t3052 n7296 n3053 R=2.213e+01 
R7296t3909 n7297 n3910 R=9.024e+00 
R7296t5265 n7297 n5266 R=3.893e+00 
R7296t2369 n7297 n2370 R=2.767e+01 
R7296t5809 n7297 n5810 R=5.194e+00 
R7297t5966 n7298 n5967 R=1.035e+01 
R7297t6874 n7298 n6875 R=3.844e+01 
R7297t4230 n7298 n4231 R=3.311e+01 
R7297t1319 n7298 n1320 R=1.332e+01 
R7297t5501 n7298 n5502 R=3.170e+00 
R7297t4087 n7298 n4088 R=2.828e+01 
R7298t728 n7299 n729 R=1.291e+01 
R7298t3578 n7299 n3579 R=3.029e+01 
R7298t1961 n7299 n1962 R=3.322e+00 
R7299t207 n7300 n208 R=1.878e+01 
R7299t1598 n7300 n1599 R=3.385e+00 
R7299t2427 n7300 n2428 R=2.691e+02 
R7299t9 n7300 n10 R=9.661e+00 
R7299t1991 n7300 n1992 R=3.521e+01 
R7300t6244 n7301 n6245 R=3.531e+00 
R7300t381 n7301 n382 R=6.522e+00 
R7300t4968 n7301 n4969 R=6.522e+00 
R7300t3310 n7301 n3311 R=9.839e+00 
R7301t2795 n7302 n2796 R=1.027e+01 
R7301t4251 n7302 n4252 R=3.589e+00 
R7301t5902 n7302 n5903 R=2.815e+00 
R7301t2221 n7302 n2222 R=2.312e+01 
R7301t5068 n7302 n5069 R=2.437e+02 
R7301t5975 n7302 n5976 R=1.392e+01 
R7302t4452 n1 n4453 R=8.375e+01 
R7302t5997 n1 n5998 R=4.381e+00 
R7302t2838 n1 n2839 R=6.945e+00 
R7303t3969 n7304 n3970 R=5.977e+00 
R7303t6448 n7304 n6449 R=2.584e+01 
R7303t5260 n7304 n5261 R=8.816e+00 
R7303t933 n7304 n934 R=1.929e+01 
R7303t1442 n7304 n1443 R=5.538e+00 
R7303t2272 n7304 n2273 R=5.894e+00 
R7303t3599 n7304 n3600 R=1.349e+01 
R7304t5082 n7305 n5083 R=8.325e+00 
R7304t1967 n7305 n1968 R=3.887e+00 
R7304t2081 n7305 n2082 R=4.642e+00 
R7305t3699 n7306 n3700 R=1.831e+01 
R7305t4773 n7306 n4774 R=9.958e+00 
R7305t550 n7306 n551 R=2.603e+00 
R7306t6182 n7307 n6183 R=1.300e+01 
R7306t1594 n7307 n1595 R=2.305e+01 
R7307t4586 n7308 n4587 R=2.122e+01 
R7307t2708 n7308 n2709 R=1.289e+01 
R7307t4913 n7308 n4914 R=8.715e+00 
R7307t5916 n7308 n5917 R=8.280e+01 
R7307t5437 n7308 n5438 R=3.578e+00 
R7308t4347 n7309 n4348 R=2.228e+02 
R7308t777 n7309 n778 R=2.356e+00 
R7309t6783 n7310 n6784 R=3.419e+01 
R7309t7161 n7310 n7162 R=4.949e+00 
R7309t5122 n7310 n5123 R=6.004e+00 
R7310t5458 n7311 n5459 R=6.481e+00 
R7310t6408 n7311 n6409 R=1.441e+02 
R7310t7120 n7311 n7121 R=2.521e+00 
R7310t6432 n7311 n6433 R=4.703e+00 
R7310t2034 n7311 n2035 R=7.219e+00 
R7310t2843 n7311 n2844 R=2.669e+01 
R7311t3524 n7312 n3525 R=1.187e+01 
R7311t4814 n7312 n4815 R=4.915e+00 
R7311t7134 n7312 n7135 R=8.927e+00 
R7311t2852 n7312 n2853 R=6.353e+01 
R7311t3383 n7312 n3384 R=9.075e+00 
R7312t6910 n7313 n6911 R=4.026e+00 
R7312t3937 n7313 n3938 R=1.083e+01 
R7312t913 n7313 n914 R=3.106e+00 
R7313t234 n7314 n235 R=7.032e+00 
R7313t1153 n7314 n1154 R=3.959e+00 
R7313t1603 n7314 n1604 R=4.405e+00 
R7313t1758 n7314 n1759 R=3.224e+00 
R7314t985 n7315 n986 R=2.573e+01 
R7314t6701 n7315 n6702 R=5.264e+00 
R7314t4621 n7315 n4622 R=1.198e+01 
R7314t3998 n7315 n3999 R=3.920e+00 
R7314t4410 n7315 n4411 R=1.140e+01 
R7315t4325 n7316 n4326 R=2.230e+01 
R7315t4877 n7316 n4878 R=4.767e+01 
R7315t3004 n7316 n3005 R=4.727e+00 
R7315t1977 n7316 n1978 R=9.832e+00 
R7315t1033 n7316 n1034 R=8.669e+00 
R7316t1852 n7317 n1853 R=3.766e+01 
R7316t5768 n7317 n5769 R=1.034e+01 
R7316t5044 n7317 n5045 R=3.151e+00 
R7316t18 n7317 n19 R=3.205e+00 
R7317t3004 n7318 n3005 R=4.261e+01 
R7317t7315 n7318 n7316 R=5.086e+00 
R7317t1977 n7318 n1978 R=3.020e+01 
R7317t481 n7318 n482 R=4.370e+00 
R7317t493 n7318 n494 R=1.771e+01 
R7318t4366 n7319 n4367 R=4.306e+02 
R7318t831 n7319 n832 R=1.230e+01 
R7318t4235 n7319 n4236 R=4.119e+02 
R7318t773 n7319 n774 R=5.676e+00 
R7318t3985 n7319 n3986 R=1.380e+01 
R7319t1419 n7320 n1420 R=1.212e+01 
R7319t3689 n7320 n3690 R=1.282e+01 
R7319t770 n7320 n771 R=4.074e+00 
R7319t2306 n7320 n2307 R=8.668e+00 
R7319t4034 n7320 n4035 R=4.246e+00 
R7320t7277 n7321 n7278 R=3.340e+00 
R7320t4986 n7321 n4987 R=2.865e+03 
R7320t903 n7321 n904 R=2.059e+00 
R7320t4611 n7321 n4612 R=3.009e+01 
R7321t439 n7322 n440 R=3.021e+00 
R7321t2009 n7322 n2010 R=7.698e+00 
R7321t810 n7322 n811 R=2.329e+01 
R7322t3296 n7323 n3297 R=6.698e+00 
R7322t5718 n7323 n5719 R=3.678e+00 
R7322t1869 n7323 n1870 R=3.025e+00 
R7322t4602 n7323 n4603 R=7.081e+00 
R7323t7246 n7324 n7247 R=5.511e+00 
R7323t3485 n7324 n3486 R=4.465e+00 
R7324t1100 n7325 n1101 R=3.861e+00 
R7324t6230 n7325 n6231 R=5.186e+00 
R7324t2846 n7325 n2847 R=4.043e+01 
R7324t872 n7325 n873 R=1.829e+01 
R7324t6605 n7325 n6606 R=1.809e+03 
R7324t914 n7325 n915 R=5.082e+01 
R7325t189 n7326 n190 R=3.978e+00 
R7325t2674 n7326 n2675 R=7.028e+00 
R7325t5196 n7326 n5197 R=2.327e+01 
R7325t1187 n7326 n1188 R=3.592e+00 
R7326t6673 n7327 n6674 R=3.809e+00 
R7326t602 n7327 n603 R=4.447e+00 
R7326t1017 n7327 n1018 R=1.122e+01 
R7326t1152 n7327 n1153 R=3.828e+01 
R7327t2968 n7328 n2969 R=4.332e+01 
R7327t5130 n7328 n5131 R=5.605e+00 
R7327t532 n7328 n533 R=1.663e+01 
R7328t327 n7329 n328 R=2.600e+02 
R7328t1273 n7329 n1 R=2.709e+00 
R7328t6944 n7329 n6945 R=9.289e+00 
R7328t4657 n7329 n4658 R=4.204e+00 
R7329t1434 n7330 n1435 R=1.793e+01 
R7329t4316 n7330 n4317 R=5.198e+01 
R7329t1113 n7330 n1114 R=1.752e+01 
R7329t3149 n7330 n3150 R=7.339e+00 
R7329t4391 n7330 n4392 R=7.556e+01 
R7330t97 n7331 n98 R=9.915e+00 
R7330t381 n7331 n382 R=1.857e+02 
R7330t5790 n7331 n5791 R=3.410e+00 
R7330t2266 n7331 n2267 R=2.521e+01 
R7331t6980 n7332 n6981 R=5.990e+00 
R7331t5321 n7332 n5322 R=1.451e+01 
R7331t1235 n7332 n1236 R=7.306e+00 
R7331t2778 n7332 n2779 R=2.867e+01 
R7331t1224 n7332 n1225 R=2.657e+01 
R7332t6355 n7333 n6356 R=2.886e+01 
R7332t6903 n7333 n6904 R=6.193e+00 
R7332t5313 n7333 n5314 R=5.079e+00 
R7332t3751 n7333 n3752 R=5.306e+01 
R7332t7028 n7333 n7029 R=6.771e+01 
R7332t403 n7333 n404 R=3.244e+01 
R7333t180 n7334 n181 R=1.555e+01 
R7333t1564 n7334 n1565 R=8.013e+00 
R7333t6336 n7334 n6337 R=8.472e+00 
R7333t7281 n7334 n7282 R=5.611e+00 
R7334t1824 n7335 n1825 R=3.678e+00 
R7334t5326 n7335 n5327 R=2.813e+00 
R7334t3367 n7335 n3368 R=5.904e+00 
R7335t3429 n7336 n3430 R=2.858e+00 
R7335t5196 n7336 n5197 R=1.421e+02 
R7335t2882 n7336 n2883 R=8.244e+00 
R7335t1623 n7336 n1624 R=2.379e+00 
R7336t2662 n7337 n2663 R=5.146e+01 
R7336t3001 n7337 n3002 R=3.839e+00 
R7336t6415 n7337 n6416 R=1.550e+01 
R7336t6953 n7337 n6954 R=2.588e+01 
R7337t4605 n7338 n4606 R=2.780e+01 
R7337t3250 n7338 n3251 R=9.728e+00 
R7337t2404 n7338 n2405 R=5.545e+00 
R7337t6291 n7338 n6292 R=4.646e+00 
R7338t1657 n7339 n1658 R=9.925e+00 
R7338t6733 n7339 n6734 R=1.387e+01 
R7338t1123 n7339 n1124 R=7.061e+00 
R7338t5781 n7339 n5782 R=7.873e+00 
R7338t6847 n7339 n6848 R=4.075e+01 
R7338t1943 n7339 n1944 R=1.129e+01 
R7338t2139 n7339 n2140 R=1.204e+01 
R7339t4017 n7340 n4018 R=2.729e+00 
R7339t6009 n7340 n6010 R=4.801e+01 
R7339t4726 n7340 n4727 R=1.265e+01 
R7339t6042 n7340 n6043 R=4.603e+00 
R7339t1406 n7340 n1407 R=1.178e+01 
R7340t7278 n7341 n7279 R=2.571e+00 
R7340t7311 n7341 n7312 R=6.449e+00 
R7340t4814 n7341 n4815 R=8.349e+00 
R7340t3612 n7341 n3613 R=1.551e+01 
R7340t6580 n7341 n6581 R=3.297e+01 
R7341t4086 n7342 n4087 R=2.868e+00 
R7341t1021 n7342 n1022 R=9.544e+00 
R7342t1114 n7343 n1115 R=5.568e+00 
R7342t3591 n7343 n3592 R=1.069e+01 
R7342t5546 n7343 n5547 R=3.479e+00 
R7343t2298 n7344 n2299 R=2.840e+00 
R7343t2926 n7344 n2927 R=5.140e+00 
R7343t5401 n7344 n5402 R=7.795e+01 
R7344t2970 n7345 n2971 R=5.323e+00 
R7344t837 n7345 n838 R=1.970e+01 
R7344t3635 n7345 n3636 R=3.737e+00 
R7345t4126 n7346 n4127 R=2.532e+00 
R7345t1605 n7346 n1606 R=2.904e+01 
R7345t1894 n7346 n1895 R=3.757e+00 
R7345t5731 n7346 n5732 R=1.688e+01 
R7345t1431 n7346 n1432 R=3.866e+01 
R7346t675 n7347 n676 R=3.910e+00 
R7346t1340 n7347 n1341 R=5.314e+00 
R7346t1164 n7347 n1165 R=3.944e+00 
R7346t6253 n7347 n6254 R=8.854e+01 
R7346t840 n7347 n841 R=5.549e+00 
R7346t714 n7347 n715 R=4.378e+02 
R7347t2013 n7348 n2014 R=6.606e+00 
R7347t2307 n7348 n2308 R=7.688e+00 
R7347t2849 n7348 n2850 R=3.859e+00 
R7347t1385 n7348 n1386 R=2.433e+01 
R7348t4248 n7349 n4249 R=6.866e+00 
R7348t5972 n7349 n5973 R=4.039e+00 
R7348t1166 n7349 n1167 R=1.374e+01 
R7349t4453 n7350 n4454 R=1.729e+01 
R7349t5574 n7350 n5575 R=9.584e+01 
R7349t2163 n7350 n2164 R=1.181e+01 
R7349t32 n7350 n33 R=3.427e+01 
R7349t4916 n7350 n4917 R=3.401e+00 
R7350t3015 n7351 n3016 R=5.412e+00 
R7350t3243 n7351 n3244 R=1.030e+01 
R7350t422 n7351 n423 R=5.741e+01 
R7350t5753 n7351 n5754 R=9.866e+00 
R7351t1835 n7352 n1836 R=1.599e+01 
R7351t3329 n7352 n3330 R=1.134e+01 
R7351t1087 n7352 n1088 R=1.598e+01 
R7351t2850 n7352 n1 R=2.189e+01 
R7351t6445 n7352 n6446 R=4.117e+01 
R7351t2407 n7352 n2408 R=3.220e+01 
R7352t3357 n7353 n3358 R=4.219e+01 
R7352t6664 n7353 n6665 R=4.950e+01 
R7352t4024 n7353 n4025 R=4.969e+00 
R7352t5664 n7353 n5665 R=4.276e+00 
R7352t574 n7353 n575 R=2.135e+01 
R7353t1853 n7354 n1854 R=9.421e+00 
R7353t5502 n7354 n5503 R=1.506e+01 
R7353t774 n7354 n775 R=4.978e+00 
R7353t2798 n7354 n2799 R=1.113e+02 
R7353t1282 n7354 n1283 R=6.003e+00 
R7353t793 n7354 n794 R=1.011e+01 
R7353t3602 n7354 n3603 R=1.110e+01 
R7354t1922 n7355 n1923 R=5.359e+00 
R7354t3912 n7355 n3913 R=5.135e+00 
R7354t1813 n7355 n1814 R=2.087e+00 
R7355t3335 n7356 n3336 R=8.432e+00 
R7355t3574 n7356 n3575 R=6.862e+00 
R7355t1684 n7356 n1685 R=1.243e+01 
R7355t5061 n7356 n5062 R=4.047e+00 
R7355t265 n7356 n266 R=7.521e+00 
R7356t1254 n7357 n1255 R=3.767e+01 
R7356t5307 n7357 n5308 R=6.023e+00 
R7356t1024 n7357 n1025 R=8.188e+00 
R7356t3440 n7357 n3441 R=1.252e+01 
R7356t789 n7357 n790 R=3.415e+00 
R7356t917 n7357 n918 R=6.513e+01 
R7357t6556 n7358 n6557 R=5.450e+00 
R7357t1581 n7358 n1582 R=7.095e+00 
R7358t4504 n1 n4505 R=2.626e+01 
R7358t4626 n1 n4627 R=1.413e+01 
R7358t4771 n1 n4772 R=9.620e+00 
R7358t4862 n1 n4863 R=8.261e+00 
R7358t4969 n1 n4970 R=7.940e+01 
R7358t7287 n1 n7288 R=5.687e+00 
R7359t1491 n7360 n1492 R=6.052e+00 
R7359t4623 n7360 n4624 R=6.759e+00 
R7359t1345 n7360 n1346 R=7.564e+01 
R7359t5662 n7360 n5663 R=9.545e+00 
R7359t2648 n7360 n2649 R=5.993e+00 
R7360t593 n7361 n594 R=9.393e+00 
R7360t4209 n7361 n4210 R=7.738e+01 
R7360t5099 n7361 n5100 R=2.848e+00 
R7360t329 n7361 n330 R=8.204e+00 
R7360t5504 n7361 n5505 R=7.003e+00 
R7360t2720 n7361 n2721 R=2.614e+01 
R7361t3917 n7362 n3918 R=5.348e+00 
R7361t5393 n7362 n5394 R=2.042e+00 
R7361t5435 n7362 n5436 R=7.074e+01 
R7361t4795 n7362 n4796 R=2.887e+00 
R7362t2325 n7363 n2326 R=9.807e+00 
R7362t4800 n7363 n4801 R=4.439e+00 
R7362t5906 n7363 n5907 R=5.390e+00 
R7362t3180 n7363 n3181 R=8.148e+01 
R7362t3887 n7363 n3888 R=5.232e+00 
R7363t1956 n7364 n1957 R=3.068e+00 
R7363t3556 n7364 n3557 R=1.052e+01 
R7363t6680 n7364 n6681 R=3.883e+01 
R7363t1404 n7364 n1405 R=4.374e+00 
R7363t6171 n7364 n6172 R=1.200e+01 
R7364t2222 n7365 n2223 R=2.446e+00 
R7364t2864 n7365 n2865 R=4.913e+01 
R7364t1341 n7365 n1342 R=2.149e+00 
R7364t1868 n7365 n1869 R=1.845e+01 
R7364t366 n7365 n367 R=2.357e+01 
R7364t869 n7365 n870 R=6.918e+00 
R7365t1849 n7366 n1850 R=2.901e+00 
R7365t4912 n7366 n4913 R=5.102e+01 
R7365t1481 n7366 n1482 R=2.980e+00 
R7365t2151 n7366 n2152 R=6.439e+00 
R7366t5720 n7367 n5721 R=3.099e+00 
R7366t5869 n7367 n5870 R=4.085e+01 
R7366t1068 n7367 n1069 R=3.511e+00 
R7366t5513 n7367 n5514 R=9.357e+00 
R7366t3870 n7367 n3871 R=6.453e+00 
R7366t5673 n7367 n5674 R=4.825e+01 
R7367t2941 n7368 n2942 R=6.631e+00 
R7367t3917 n7368 n3918 R=1.197e+01 
R7367t4597 n7368 n4598 R=2.504e+01 
R7367t5951 n7368 n5952 R=1.456e+01 
R7367t5613 n7368 n5614 R=1.070e+01 
R7367t4480 n7368 n4481 R=6.906e+00 
R7368t6783 n7369 n6784 R=1.772e+01 
R7368t7309 n7369 n7310 R=4.131e+00 
R7368t2937 n7369 n2938 R=7.187e+00 
R7368t5931 n7369 n5932 R=3.294e+00 
R7368t7161 n7369 n7162 R=1.425e+01 
R7369t924 n7370 n925 R=9.820e+00 
R7369t6705 n7370 n6706 R=4.247e+00 
R7369t2496 n7370 n2497 R=3.725e+00 
R7369t2561 n7370 n2562 R=7.170e+00 
R7369t6978 n7370 n6979 R=1.007e+01 
R7370t3886 n7371 n3887 R=3.640e+01 
R7370t4174 n7371 n4175 R=3.616e+01 
R7370t4274 n7371 n4275 R=2.937e+00 
R7370t2266 n7371 n2267 R=1.052e+01 
R7370t97 n7371 n98 R=1.464e+01 
R7371t45 n7372 n46 R=9.359e+00 
R7371t2888 n7372 n2889 R=3.411e+00 
R7371t767 n7372 n768 R=1.514e+01 
R7371t4630 n7372 n4631 R=8.331e+00 
R7372t2319 n7373 n2320 R=3.739e+01 
R7372t5604 n7373 n5605 R=3.070e+00 
R7373t4024 n7374 n4025 R=6.449e+00 
R7373t4748 n7374 n4749 R=5.812e+00 
R7373t6729 n7374 n6730 R=6.304e+00 
R7373t5664 n7374 n5665 R=1.912e+01 
R7374t5214 n7375 n5215 R=9.344e+00 
R7374t4390 n7375 n4391 R=5.413e+01 
R7375t2327 n7376 n2328 R=3.075e+01 
R7375t5113 n7376 n5114 R=5.874e+00 
R7376t5268 n7377 n5269 R=2.113e+01 
R7376t4780 n7377 n4781 R=6.190e+00 
R7376t6827 n7377 n6828 R=2.825e+01 
R7376t92 n7377 n93 R=6.138e+00 
R7377t1531 n7378 n1532 R=4.376e+01 
R7377t2715 n7378 n2716 R=1.221e+01 
R7377t151 n7378 n152 R=3.724e+00 
R7377t6164 n7378 n6165 R=8.740e+00 
R7378t2330 n7379 n2331 R=3.948e+00 
R7378t5166 n7379 n5167 R=3.511e+01 
R7378t3217 n7379 n3218 R=3.218e+00 
R7378t6892 n7379 n6893 R=8.993e+00 
R7379t2370 n7380 n2371 R=1.921e+01 
R7379t540 n7380 n541 R=4.289e+00 
R7379t3832 n7380 n3833 R=2.851e+01 
R7379t313 n7380 n314 R=3.871e+00 
R7379t1832 n7380 n1833 R=3.023e+02 
R7380t5676 n7381 n5677 R=1.517e+01 
R7380t1622 n7381 n1623 R=1.076e+01 
R7381t1634 n7382 n1635 R=3.260e+01 
R7381t865 n7382 n866 R=2.319e+00 
R7381t5981 n7382 n5982 R=7.656e+00 
R7381t6557 n7382 n6558 R=1.657e+00 
R7382t4707 n7383 n4708 R=7.579e+00 
R7382t6161 n7383 n6162 R=1.037e+01 
R7383t7323 n7384 n7324 R=1.192e+01 
R7383t2295 n7384 n2296 R=1.928e+01 
R7383t4574 n7384 n4575 R=1.055e+01 
R7383t43 n7384 n44 R=1.008e+01 
R7384t3977 n7385 n3978 R=2.127e+00 
R7384t6374 n7385 n6375 R=7.546e+00 
R7384t4641 n7385 n4642 R=4.094e+01 
R7384t4501 n7385 n4502 R=6.339e+00 
R7384t538 n7385 n539 R=1.514e+01 
R7385t1385 n7386 n1386 R=1.853e+01 
R7385t1866 n7386 n1867 R=3.897e+00 
R7385t4281 n7386 n4282 R=2.257e+01 
R7385t6264 n7386 n6265 R=6.488e+00 
R7386t6309 n7387 n6310 R=4.890e+01 
R7386t4689 n7387 n4690 R=1.345e+02 
R7386t3122 n7387 n3123 R=3.958e+00 
R7386t3035 n7387 n3036 R=3.168e+01 
R7386t6446 n7387 n6447 R=6.575e+01 
R7386t6095 n7387 n6096 R=6.468e+00 
R7387t716 n7388 n717 R=3.695e+00 
R7387t994 n7388 n995 R=2.186e+01 
R7387t2138 n7388 n2139 R=4.450e+00 
R7387t3905 n7388 n3906 R=2.527e+01 
R7388t6490 n7389 n6491 R=6.314e+00 
R7388t3722 n7389 n3723 R=2.455e+01 
R7388t3617 n7389 n3618 R=2.607e+00 
R7389t3204 n7390 n3205 R=5.598e+01 
R7389t4936 n7390 n4937 R=2.692e+00 
R7389t6303 n7390 n6304 R=7.860e+00 
R7389t771 n7390 n772 R=1.996e+01 
R7389t3735 n7390 n3736 R=2.790e+00 
R7389t2067 n7390 n2068 R=9.490e+00 
R7390t2735 n7391 n2736 R=4.021e+00 
R7390t2719 n7391 n2720 R=2.537e+01 
R7390t4750 n7391 n4751 R=2.298e+01 
R7390t2089 n7391 n2090 R=2.247e+00 
R7390t4518 n7391 n4519 R=7.503e+01 
R7391t6744 n7392 n6745 R=3.046e+00 
R7391t3273 n7392 n3274 R=1.743e+00 
R7391t4799 n7392 n4800 R=6.136e+01 
R7391t5910 n7392 n5911 R=8.264e+00 
R7391t6349 n7392 n6350 R=8.000e+01 
R7392t1006 n7393 n1007 R=1.847e+01 
R7392t1985 n7393 n1986 R=7.297e+00 
R7392t139 n7393 n140 R=1.423e+01 
R7392t5414 n7393 n5415 R=5.313e+01 
R7392t1747 n7393 n1748 R=5.872e+00 
R7392t5335 n7393 n5336 R=5.106e+00 
R7392t7130 n7393 n7131 R=2.440e+01 
R7393t3804 n7394 n3805 R=1.700e+02 
R7393t2933 n7394 n2934 R=3.223e+00 
R7393t6696 n7394 n6697 R=1.878e+00 
R7394t2076 n7395 n2077 R=4.547e+01 
R7394t2491 n7395 n2492 R=3.612e+00 
R7394t7135 n7395 n7136 R=1.195e+01 
R7394t797 n7395 n798 R=1.318e+00 
R7394t1762 n7395 n1763 R=1.821e+02 
R7394t2667 n7395 n2668 R=3.677e+01 
R7394t181 n7395 n182 R=6.128e+00 
R7395t99 n7396 n100 R=6.763e+00 
R7395t2084 n7396 n2085 R=1.159e+01 
R7396t3551 n7397 n3552 R=5.821e+00 
R7396t5967 n7397 n5968 R=1.457e+03 
R7396t1234 n7397 n1235 R=9.944e+00 
R7396t4734 n7397 n4735 R=1.013e+01 
R7396t4234 n7397 n4235 R=1.385e+01 
R7396t6648 n7397 n6649 R=5.189e+00 
R7396t1922 n7397 n1923 R=1.216e+02 
R7396t7354 n7397 n7355 R=1.059e+01 
R7396t1813 n7397 n1814 R=7.134e+01 
R7397t7025 n7398 n7026 R=7.829e+00 
R7397t4268 n7398 n4269 R=8.175e+00 
R7397t5395 n7398 n5396 R=1.807e+00 
R7397t943 n7398 n944 R=9.981e+00 
R7397t6380 n7398 n6381 R=1.566e+01 
R7398t4014 n7399 n4015 R=4.690e+00 
R7398t5112 n7399 n5113 R=7.439e+00 
R7398t4977 n7399 n4978 R=1.204e+01 
R7398t874 n7399 n875 R=2.991e+00 
R7399t6133 n7400 n6134 R=1.276e+01 
R7399t1055 n7400 n1056 R=2.848e+01 
R7399t3360 n7400 n3361 R=1.322e+01 
R7399t4979 n7400 n4980 R=9.033e+00 
R7399t6916 n7400 n6917 R=3.917e+00 
R7400t5449 n7401 n5450 R=1.304e+01 
R7400t2896 n7401 n2897 R=5.470e+00 
R7400t3571 n7401 n3572 R=5.075e+00 
R7400t5794 n7401 n5795 R=1.565e+01 
R7401t3301 n7402 n3302 R=4.064e+00 
R7401t5451 n7402 n5452 R=7.407e+00 
R7401t660 n7402 n661 R=7.798e+00 
R7401t3454 n7402 n3455 R=7.868e+02 
R7401t2287 n7402 n2288 R=2.410e+00 
R7402t1994 n7403 n1995 R=1.452e+01 
R7402t4884 n7403 n4885 R=8.947e+00 
R7402t1471 n7403 n1472 R=3.698e+01 
R7402t1770 n7403 n1771 R=4.251e+00 
R7402t6640 n7403 n6641 R=7.593e+00 
R7403t2228 n7404 n2229 R=1.473e+01 
R7403t7152 n7404 n7153 R=3.771e+00 
R7403t5879 n7404 n5880 R=5.106e+00 
R7404t2919 n7405 n2920 R=1.135e+01 
R7404t5019 n7405 n5020 R=2.530e+01 
R7404t5459 n7405 n5460 R=3.906e+00 
R7404t931 n7405 n932 R=3.886e+01 
R7404t4315 n7405 n4316 R=1.647e+01 
R7404t561 n7405 n562 R=3.304e+00 
R7405t6341 n7406 n6342 R=2.775e+01 
R7405t7023 n7406 n7024 R=7.661e+00 
R7405t5144 n7406 n5145 R=2.291e+01 
R7405t1604 n7406 n1605 R=5.537e+00 
R7405t1680 n7406 n1681 R=5.324e+01 
R7406t93 n7407 n94 R=4.406e+00 
R7406t5242 n7407 n5243 R=3.162e+00 
R7406t3500 n7407 n3501 R=1.324e+01 
R7406t222 n7407 n223 R=5.502e+01 
R7407t2 n7408 n3 R=5.618e+01 
R7407t5954 n7408 n5955 R=4.673e+01 
R7407t6481 n7408 n6482 R=9.841e+00 
R7407t3086 n7408 n3087 R=5.711e+00 
R7408t4818 n7409 n4819 R=3.475e+01 
R7408t2616 n7409 n2617 R=1.539e+01 
R7408t2000 n7409 n2001 R=1.306e+01 
R7409t1951 n7410 n1952 R=5.472e+00 
R7409t6844 n7410 n6845 R=3.784e+00 
R7409t7247 n7410 n7248 R=4.259e+00 
R7409t5354 n7410 n5355 R=4.791e+00 
R7409t4229 n7410 n4230 R=3.730e+01 
R7410t3173 n7411 n3174 R=4.685e+01 
R7410t3941 n7411 n3942 R=9.120e+00 
R7411t2109 n7412 n2110 R=9.471e+00 
R7411t2162 n7412 n2163 R=6.100e+00 
R7411t5067 n7412 n5068 R=3.543e+01 
R7411t2160 n7412 n2161 R=1.781e+01 
R7411t3967 n7412 n3968 R=7.295e+00 
R7412t1380 n7413 n1381 R=1.867e+01 
R7412t2833 n7413 n2834 R=8.661e+00 
R7412t6568 n7413 n6569 R=2.652e+01 
R7412t5416 n7413 n5417 R=7.780e+00 
R7412t3882 n7413 n3883 R=4.296e+00 
R7413t6289 n7414 n6290 R=8.512e+00 
R7413t6884 n7414 n6885 R=3.276e+00 
R7413t3266 n7414 n3267 R=2.767e+01 
R7414t19 n7415 n20 R=2.457e+01 
R7414t2199 n7415 n2200 R=5.694e+00 
R7414t1036 n7415 n1037 R=1.815e+01 
R7414t2313 n7415 n2314 R=1.037e+01 
R7415t5106 n7416 n5107 R=3.191e+00 
R7415t5470 n7416 n5471 R=9.323e+00 
R7415t5410 n7416 n5411 R=2.898e+01 
R7415t4723 n7416 n4724 R=6.363e+00 
R7415t232 n7416 n233 R=2.095e+02 
R7415t6199 n7416 n6200 R=1.192e+01 
R7415t2713 n7416 n2714 R=1.054e+01 
R7416t301 n7417 n302 R=9.026e+00 
R7416t6944 n7417 n6945 R=1.974e+01 
R7416t5209 n7417 n1 R=2.947e+00 
R7416t2900 n7417 n1 R=6.776e+00 
R7417t3088 n7418 n3089 R=3.712e+00 
R7417t3164 n7418 n3165 R=4.094e+01 
R7417t4057 n7418 n4058 R=1.663e+01 
R7417t1456 n7418 n1457 R=1.295e+01 
R7417t6152 n7418 n6153 R=4.509e+00 
R7417t1709 n7418 n1710 R=1.578e+01 
R7417t85 n7418 n86 R=9.475e+00 
R7418t6486 n7419 n6487 R=2.808e+00 
R7418t3974 n7419 n3975 R=3.570e+00 
R7418t5051 n7419 n5052 R=6.606e+02 
R7418t1094 n7419 n1095 R=5.064e+00 
R7418t4550 n7419 n4551 R=2.396e+01 
R7419t3559 n7420 n3560 R=2.575e+01 
R7419t5998 n7420 n5999 R=7.767e+00 
R7419t1893 n7420 n1894 R=4.786e+01 
R7419t1209 n7420 n1210 R=2.375e+01 
R7419t4206 n7420 n4207 R=4.263e+00 
R7420t1984 n7421 n1985 R=5.281e+02 
R7420t2352 n7421 n2353 R=4.814e+00 
R7421t61 n7422 n62 R=9.324e+00 
R7421t91 n7422 n92 R=2.142e+01 
R7421t5960 n7422 n5961 R=5.970e+00 
R7421t6416 n7422 n6417 R=3.241e+01 
R7421t473 n7422 n474 R=1.195e+01 
R7422t3145 n7423 n3146 R=1.217e+01 
R7422t5415 n7423 n5416 R=7.875e+00 
R7422t3128 n7423 n3129 R=8.734e+00 
R7422t1051 n7423 n1052 R=3.221e+00 
R7422t501 n7423 n502 R=1.789e+01 
R7422t5801 n7423 n5802 R=3.031e+01 
R7423t2030 n7424 n2031 R=3.607e+00 
R7423t2299 n7424 n2300 R=1.195e+01 
R7423t6956 n7424 n6957 R=2.400e+01 
R7423t4980 n7424 n4981 R=2.191e+00 
R7424t944 n7425 n945 R=1.087e+02 
R7424t2707 n7425 n2708 R=2.480e+01 
R7424t506 n7425 n507 R=3.237e+00 
R7424t1880 n7425 n1881 R=1.998e+02 
R7424t3919 n7425 n3920 R=1.623e+00 
R7424t3514 n7425 n3515 R=5.151e+00 
R7425t1289 n7426 n1290 R=7.402e+00 
R7425t1681 n7426 n1682 R=9.914e+00 
R7425t7142 n7426 n7143 R=6.930e+00 
R7425t6661 n7426 n6662 R=2.864e+01 
R7425t2323 n7426 n2324 R=1.301e+01 
R7425t4702 n7426 n4703 R=4.207e+00 
R7426t3069 n7427 n3070 R=7.882e+00 
R7426t5202 n7427 n5203 R=4.826e+00 
R7426t3724 n7427 n3725 R=4.582e+00 
R7426t3799 n7427 n3800 R=2.448e+00 
R7427t2825 n7428 n2826 R=4.466e+00 
R7427t5992 n7428 n5993 R=3.902e+00 
R7427t4001 n7428 n4002 R=4.118e+00 
R7428t4 n7429 n5 R=5.483e+00 
R7428t148 n7429 n149 R=3.770e+00 
R7428t970 n7429 n971 R=8.189e+01 
R7428t2237 n7429 n2238 R=1.678e+02 
R7428t3219 n7429 n3220 R=2.780e+00 
R7428t54 n7429 n55 R=1.228e+01 
R7429t5794 n7430 n5795 R=7.100e+01 
R7429t5494 n7430 n5495 R=5.124e+00 
R7429t3289 n7430 n3290 R=2.693e+02 
R7429t4966 n7430 n4967 R=5.965e+00 
R7429t5228 n7430 n5229 R=2.209e+01 
R7429t997 n7430 n998 R=1.580e+01 
R7429t6184 n7430 n6185 R=6.570e+00 
R7429t3426 n7430 n3427 R=3.194e+01 
R7430t1120 n7431 n1121 R=4.694e+00 
R7430t6829 n7431 n6830 R=1.187e+02 
R7430t6544 n7431 n6545 R=4.058e+00 
R7430t1776 n7431 n1777 R=3.766e+00 
R7431t6463 n7432 n6464 R=1.383e+00 
R7431t5548 n7432 n5549 R=5.697e+00 
R7431t859 n7432 n860 R=2.063e+01 
R7432t3050 n7433 n3051 R=6.150e+00 
R7432t3272 n7433 n3273 R=4.876e+00 
R7432t2135 n7433 n2136 R=2.426e+00 
R7432t1009 n7433 n1010 R=1.298e+01 
R7433t3202 n7434 n3203 R=4.290e+00 
R7433t4045 n7434 n4046 R=3.793e+01 
R7433t4647 n7434 n4648 R=3.078e+00 
R7434t440 n7435 n441 R=2.965e+01 
R7434t961 n7435 n962 R=1.664e+00 
R7434t3985 n7435 n3986 R=1.211e+02 
R7434t773 n7435 n774 R=1.025e+02 
R7434t53 n7435 n54 R=1.970e+01 
R7434t2548 n7435 n2549 R=2.756e+00 
R7435t982 n7436 n983 R=6.216e+00 
R7435t3953 n7436 n3954 R=1.075e+01 
R7436t3428 n7437 n3429 R=5.107e+00 
R7436t748 n7437 n749 R=1.707e+01 
R7436t5385 n7437 n5386 R=1.680e+01 
R7436t3550 n7437 n3551 R=4.300e+00 
R7436t912 n7437 n913 R=3.806e+00 
R7437t5615 n7438 n5616 R=1.656e+01 
R7437t6522 n7438 n6523 R=7.999e+00 
R7437t6222 n7438 n6223 R=3.598e+00 
R7437t1873 n7438 n1874 R=8.976e+00 
R7437t2936 n7438 n2937 R=5.662e+00 
R7438t6396 n7439 n6397 R=3.803e+00 
R7438t2171 n7439 n2172 R=8.166e+00 
R7438t1751 n7439 n1752 R=2.875e+00 
R7439t2718 n7440 n2719 R=1.227e+01 
R7439t556 n7440 n557 R=5.142e+00 
R7439t3539 n7440 n3540 R=1.855e+00 
R7439t677 n7440 n678 R=3.016e+01 
R7440t3278 n7441 n3279 R=3.622e+00 
R7440t7103 n7441 n7104 R=4.440e+01 
R7440t6904 n7441 n6905 R=5.447e+01 
R7440t6985 n7441 n6986 R=2.770e+00 
R7441t3751 n7442 n3752 R=6.339e+00 
R7441t7420 n7442 n7421 R=1.413e+02 
R7441t5313 n7442 n5314 R=2.330e+01 
R7442t3889 n7443 n3890 R=4.703e+00 
R7442t4599 n7443 n4600 R=6.826e+00 
R7442t4361 n7443 n4362 R=1.029e+01 
R7443t443 n7444 n444 R=1.308e+03 
R7443t3978 n7444 n3979 R=3.646e+02 
R7443t4581 n7444 n4582 R=2.031e+00 
R7443t2329 n7444 n2330 R=2.060e+01 
R7443t3626 n7444 n3627 R=2.380e+00 
R7444t5808 n7445 n5809 R=2.740e+00 
R7444t1185 n7445 n1186 R=2.091e+01 
R7444t493 n7445 n494 R=9.349e+00 
R7444t7317 n7445 n7318 R=5.270e+00 
R7444t481 n7445 n482 R=1.073e+01 
R7445t87 n7446 n88 R=1.527e+02 
R7445t6459 n7446 n6460 R=1.147e+01 
R7445t4295 n7446 n4296 R=3.435e+00 
R7445t156 n7446 n157 R=2.956e+01 
R7445t5526 n7446 n5527 R=4.738e+00 
R7445t4007 n7446 n4008 R=2.737e+01 
R7446t4160 n7447 n4161 R=1.042e+02 
R7446t5780 n7447 n5781 R=5.735e+00 
R7446t6327 n7447 n6328 R=8.273e+00 
R7446t5907 n7447 n5908 R=5.968e+00 
R7446t498 n7447 n499 R=3.953e+00 
R7446t4044 n7447 n4045 R=8.289e+00 
R7447t2490 n7448 n2491 R=5.306e+00 
R7447t2250 n7448 n2251 R=1.044e+01 
R7447t6157 n7448 n6158 R=4.567e+00 
R7447t447 n7448 n448 R=1.073e+01 
R7447t5468 n7448 n5469 R=2.930e+01 
R7448t1345 n7449 n1346 R=6.063e+00 
R7448t5918 n7449 n5919 R=7.536e+00 
R7448t5654 n7449 n5655 R=1.494e+01 
R7448t1474 n7449 n1475 R=5.020e+01 
R7448t6912 n7449 n6913 R=6.130e+00 
R7448t725 n7449 n726 R=4.969e+00 
R7449t3302 n7450 n3303 R=1.034e+01 
R7449t6267 n7450 n6268 R=3.603e+00 
R7449t6637 n7450 n6638 R=7.493e+00 
R7450t904 n7451 n905 R=6.513e+00 
R7450t5273 n7451 n5274 R=5.414e+00 
R7450t2323 n7451 n2324 R=1.195e+01 
R7450t6164 n7451 n6165 R=4.157e+00 
R7451t4389 n7452 n4390 R=5.001e+00 
R7451t4392 n7452 n4393 R=4.993e+01 
R7451t6974 n7452 n6975 R=3.350e+01 
R7451t1177 n7452 n1178 R=3.195e+00 
R7451t3337 n7452 n3338 R=3.865e+01 
R7451t6087 n7452 n6088 R=1.405e+03 
R7451t463 n7452 n464 R=8.845e+00 
R7451t1429 n7452 n1430 R=6.235e+00 
R7452t2188 n7453 n2189 R=3.520e+00 
R7452t3652 n7453 n3653 R=9.204e+00 
R7452t1305 n7453 n1306 R=7.265e+00 
R7453t4055 n7454 n4056 R=3.595e+00 
R7453t5779 n7454 n5780 R=5.957e+00 
R7453t6249 n7454 n6250 R=1.308e+01 
R7453t981 n7454 n982 R=3.977e+01 
R7453t6263 n7454 n6264 R=1.561e+01 
R7453t1529 n7454 n1530 R=7.483e+00 
R7453t2381 n7454 n2382 R=1.444e+01 
R7454t4785 n7455 n4786 R=5.856e+00 
R7454t1947 n7455 n1948 R=3.051e+00 
R7455t7408 n7456 n7409 R=9.408e+00 
R7455t4818 n7456 n4819 R=2.143e+00 
R7455t3084 n7456 n3085 R=1.624e+01 
R7455t2381 n7456 n2382 R=2.454e+00 
R7455t1529 n7456 n1530 R=2.629e+01 
R7455t959 n7456 n960 R=4.411e+02 
R7456t212 n7457 n213 R=1.951e+00 
R7456t3052 n7457 n3053 R=1.135e+01 
R7456t4060 n7457 n4061 R=3.623e+01 
R7456t3259 n7457 n3260 R=2.147e+00 
R7457t200 n7458 n201 R=8.501e+00 
R7457t6921 n7458 n6922 R=4.071e+00 
R7457t6773 n7458 n6774 R=1.175e+02 
R7457t3637 n7458 n3638 R=1.167e+01 
R7457t2895 n7458 n2896 R=2.533e+00 
R7457t3946 n7458 n3947 R=2.847e+01 
R7457t826 n7458 n827 R=1.790e+01 
R7458t1620 n7459 n1621 R=1.276e+01 
R7459t87 n7460 n88 R=3.413e+01 
R7459t7445 n7460 n7446 R=7.481e+00 
R7459t6471 n7460 n6472 R=7.403e+00 
R7459t5505 n7460 n5506 R=3.634e+00 
R7459t6459 n7460 n6460 R=3.731e+00 
R7460t2402 n7461 n2403 R=2.827e+00 
R7460t2667 n7461 n2668 R=1.233e+02 
R7461t1285 n7462 n1286 R=8.738e+00 
R7461t6877 n7462 n6878 R=1.899e+01 
R7461t5628 n7462 n5629 R=9.570e+00 
R7461t3044 n7462 n3045 R=6.105e+00 
R7461t710 n7462 n711 R=9.904e+00 
R7462t5464 n7463 n5465 R=2.558e+02 
R7462t4113 n7463 n4114 R=4.661e+00 
R7462t219 n7463 n220 R=1.716e+01 
R7462t3000 n7463 n3001 R=1.251e+02 
R7462t1142 n7463 n1143 R=4.318e+00 
R7462t3314 n7463 n3315 R=1.368e+01 
R7463t3204 n7464 n3205 R=8.037e+00 
R7463t5658 n7464 n5659 R=7.350e+00 
R7463t1582 n7464 n1583 R=1.614e+03 
R7463t3934 n7464 n3935 R=5.138e+00 
R7464t3514 n7465 n3515 R=4.009e+00 
R7464t7284 n7465 n7285 R=2.241e+01 
R7464t3464 n7465 n3465 R=3.679e+00 
R7464t1783 n7465 n1784 R=6.020e+00 
R7464t3942 n7465 n3943 R=1.551e+01 
R7464t4412 n7465 n4413 R=1.511e+01 
R7465t546 n7466 n547 R=3.471e+01 
R7465t4561 n7466 n4562 R=4.211e+00 
R7465t6716 n7466 n6717 R=1.099e+01 
R7465t3144 n7466 n3145 R=3.398e+00 
R7465t5056 n7466 n5057 R=3.101e+01 
R7465t6675 n7466 n6676 R=1.065e+01 
R7465t7076 n7466 n7077 R=8.503e+01 
R7465t953 n7466 n954 R=2.221e+01 
R7465t1225 n7466 n1226 R=2.242e+01 
R7466t1123 n7467 n1124 R=2.470e+00 
R7466t7338 n7467 n7339 R=1.362e+01 
R7466t5781 n7467 n5782 R=3.675e+00 
R7466t925 n7467 n926 R=4.355e+00 
R7467t1621 n7468 n1622 R=3.953e+00 
R7467t2726 n7468 n2727 R=2.136e+02 
R7467t5353 n7468 n5354 R=1.012e+01 
R7467t3846 n7468 n3847 R=1.027e+01 
R7467t852 n7468 n853 R=9.621e+00 
R7468t3415 n7469 n3416 R=3.966e+00 
R7468t1081 n7469 n1082 R=5.275e+00 
R7468t1313 n7469 n1314 R=5.815e+00 
R7469t2113 n7470 n2114 R=8.157e+00 
R7469t3057 n7470 n3058 R=2.392e+02 
R7469t3679 n7470 n3680 R=3.421e+00 
R7469t2238 n7470 n2239 R=2.694e+00 
R7470t3876 n7471 n3877 R=8.122e+00 
R7470t6295 n7471 n6296 R=3.899e+00 
R7470t2688 n7471 n2689 R=8.928e+00 
R7470t6075 n7471 n6076 R=1.474e+01 
R7470t6474 n7471 n6475 R=4.104e+00 
R7471t1117 n7472 n1118 R=2.555e+00 
R7471t5427 n7472 n5428 R=5.607e+00 
R7472t1130 n7473 n1131 R=2.478e+00 
R7472t4682 n7473 n4683 R=2.590e+01 
R7472t1492 n7473 n1493 R=5.976e+00 
R7472t5361 n7473 n5362 R=2.520e+00 
R7473t7027 n7474 n7028 R=1.069e+01 
R7473t1818 n7474 n1819 R=5.286e+01 
R7473t3170 n7474 n3171 R=8.635e+00 
R7473t1508 n7474 n1509 R=4.441e+00 
R7473t2153 n7474 n2154 R=1.967e+01 
R7473t830 n7474 n831 R=7.398e+01 
R7474t3511 n7475 n3512 R=7.514e+00 
R7474t4904 n7475 n4905 R=5.043e+00 
R7474t3804 n7475 n3805 R=3.917e+00 
R7474t7393 n7475 n7394 R=3.031e+01 
R7474t2933 n7475 n2934 R=5.371e+00 
R7475t1390 n7476 n1391 R=1.254e+01 
R7475t1941 n7476 n1942 R=6.252e+00 
R7475t3070 n7476 n3071 R=1.004e+02 
R7475t6539 n7476 n6540 R=6.412e+00 
R7475t5554 n7476 n5555 R=2.861e+01 
R7476t2025 n7477 n2026 R=7.092e+00 
R7476t5195 n7477 n5196 R=5.442e+00 
R7476t1150 n7477 n1151 R=3.098e+01 
R7476t3835 n7477 n3836 R=3.941e+00 
R7476t723 n7477 n724 R=4.073e+00 
R7477t1041 n7478 n1042 R=3.103e+01 
R7477t6878 n7478 n6879 R=1.560e+01 
R7477t5366 n7478 n5367 R=4.896e+00 
R7477t2738 n7478 n2739 R=6.282e+00 
R7478t622 n7479 n623 R=1.566e+01 
R7478t3469 n7479 n3470 R=4.162e+00 
R7479t3305 n7480 n3306 R=9.633e+00 
R7479t5006 n7480 n5007 R=6.623e+00 
R7479t2070 n7480 n2071 R=6.043e+00 
R7479t4588 n7480 n4589 R=3.047e+00 
R7479t6549 n7480 n6550 R=2.511e+01 
R7480t379 n7481 n380 R=1.103e+01 
R7480t5944 n7481 n5945 R=8.914e+00 
R7480t5532 n7481 n5533 R=7.067e+00 
R7480t2999 n7481 n3000 R=4.185e+00 
R7481t478 n7482 n479 R=1.041e+02 
R7481t3386 n7482 n3387 R=7.252e+00 
R7481t4232 n7482 n4233 R=4.027e+00 
R7482t5168 n7483 n5169 R=6.675e+00 
R7482t128 n7483 n129 R=1.610e+01 
R7482t7040 n7483 n7041 R=1.339e+01 
R7482t4324 n7483 n4325 R=8.190e+00 
R7483t6467 n7484 n6468 R=3.544e+00 
R7483t4076 n7484 n4077 R=5.767e+01 
R7483t5611 n7484 n5612 R=1.510e+01 
R7483t5187 n7484 n5188 R=5.836e+00 
R7484t4333 n7485 n4334 R=2.411e+00 
R7484t5575 n7485 n5576 R=9.798e+01 
R7484t533 n7485 n534 R=1.194e+01 
R7485t1783 n7486 n1784 R=6.003e+00 
R7485t3048 n7486 n3049 R=7.407e+00 
R7485t4909 n7486 n4910 R=7.551e+00 
R7485t3096 n7486 n3097 R=4.892e+00 
R7485t6120 n7486 n6121 R=8.658e+01 
R7485t3464 n7486 n3465 R=1.202e+01 
R7485t7464 n7486 n7465 R=3.611e+01 
R7486t3176 n7487 n3177 R=3.497e+00 
R7486t2504 n7487 n2505 R=4.126e+00 
R7487t6127 n7488 n6128 R=2.060e+01 
R7487t1945 n7488 n1946 R=7.466e+00 
R7487t6318 n7488 n6319 R=4.086e+00 
R7487t4122 n7488 n4123 R=2.157e+00 
R7488t4325 n7489 n4326 R=4.656e+00 
R7488t5154 n7489 n5155 R=1.008e+01 
R7488t1991 n7489 n1992 R=1.297e+01 
R7488t7299 n7489 n7300 R=7.200e+00 
R7489t5986 n7490 n5987 R=1.994e+03 
R7489t7447 n7490 n7448 R=6.135e+01 
R7489t2250 n7490 n2251 R=2.958e+00 
R7490t1650 n7491 n1651 R=2.710e+00 
R7490t3580 n7491 n3581 R=1.839e+01 
R7490t6002 n7491 n6003 R=1.471e+01 
R7491t1152 n7492 n1153 R=8.874e+00 
R7491t7326 n7492 n7327 R=3.040e+01 
R7491t1017 n7492 n1018 R=2.920e+00 
R7491t5830 n7492 n5831 R=3.833e+01 
R7491t7236 n7492 n7237 R=2.002e+01 
R7491t1103 n7492 n1104 R=4.973e+00 
R7492t4904 n7493 n4905 R=3.666e+00 
R7492t7146 n7493 n7147 R=1.106e+01 
R7492t5820 n7493 n5821 R=7.597e+00 
R7493t3253 n7494 n3254 R=1.002e+01 
R7493t2257 n7494 n2258 R=4.280e+00 
R7493t4533 n7494 n4534 R=3.678e+01 
R7493t6805 n7494 n6806 R=4.211e+00 
R7494t877 n7495 n878 R=1.926e+01 
R7494t1519 n7495 n1520 R=3.761e+00 
R7494t894 n7495 n895 R=4.855e+00 
R7494t6943 n7495 n6944 R=7.344e+00 
R7494t7171 n7495 n7172 R=9.673e+00 
R7495t1534 n7496 n1535 R=1.651e+02 
R7495t3299 n7496 n3300 R=1.031e+01 
R7495t2819 n7496 n2820 R=9.836e+00 
R7495t3316 n7496 n3317 R=6.294e+00 
R7496t4506 n7497 n4507 R=3.443e+00 
R7496t3263 n7497 n3264 R=8.566e+01 
R7496t3108 n7497 n3109 R=6.251e+01 
R7496t1308 n7497 n1309 R=2.094e+00 
R7497t2586 n7498 n2587 R=2.249e+01 
R7497t3262 n7498 n3263 R=3.827e+01 
R7497t288 n7498 n289 R=2.762e+00 
R7497t5053 n7498 n5054 R=3.287e+00 
R7497t14 n7498 n15 R=8.100e+00 
R7498t1276 n7499 n1277 R=3.229e+02 
R7498t2601 n7499 n2602 R=1.658e+01 
R7498t6411 n7499 n6412 R=1.118e+02 
R7498t616 n7499 n617 R=8.094e+00 
R7498t4405 n7499 n4406 R=2.770e+00 
R7499t2739 n7500 n2740 R=1.220e+01 
R7499t6378 n7500 n6379 R=6.573e+00 
R7499t5764 n7500 n5765 R=2.046e+00 
R7500t23 n7501 n24 R=9.146e+00 
R7500t6702 n7501 n6703 R=2.197e+01 
R7500t6521 n7501 n6522 R=6.061e+00 
R7500t3491 n7501 n3492 R=8.255e+00 
R7500t6105 n7501 n6106 R=1.376e+01 
R7502t1896 n7503 n1897 R=1.728e+01 
R7502t5198 n7503 n5199 R=2.046e+01 
R7502t2349 n7503 n2350 R=5.435e+00 
R7502t2147 n7503 n2148 R=8.415e+00 
R7502t25 n7503 n26 R=1.506e+01 
R7502t5054 n7503 n5055 R=7.406e+00 
R7503t4731 n7504 n4732 R=1.735e+01 
R7503t3865 n7504 n3866 R=7.194e+01 
R7503t896 n7504 n897 R=6.835e+00 
R7503t2750 n7504 n2751 R=8.392e+01 
R7503t5651 n7504 n5652 R=2.514e+01 
R7504t1371 n7505 n1372 R=7.885e+00 
R7504t5827 n7505 n5828 R=3.744e+00 
R7504t2110 n7505 n2111 R=2.272e+00 
R7504t6828 n7505 n6829 R=2.945e+01 
R7505t4333 n7506 n4334 R=6.215e+00 
R7505t4451 n7506 n4452 R=2.566e+01 
R7505t7484 n7506 n7485 R=3.963e+02 
R7505t533 n7506 n534 R=4.115e+00 
R7505t6156 n7506 n6157 R=7.688e+00 
R7505t3349 n7506 n3350 R=3.885e+00 
R7506t4904 n7507 n4905 R=1.415e+01 
R7506t7146 n7507 n7147 R=5.303e+00 
R7506t3160 n7507 n3161 R=4.910e+00 
R7506t1157 n7507 n1158 R=1.096e+01 
R7506t3804 n7507 n3805 R=9.953e+01 
R7506t3511 n7507 n3512 R=4.753e+00 
R7507t3306 n7508 n3307 R=3.231e+02 
R7507t2100 n7508 n2101 R=6.712e+00 
R7507t3025 n7508 n3026 R=3.328e+00 
R7507t2209 n7508 n2210 R=8.834e+00 
R7508t3061 n7509 n3062 R=6.619e+00 
R7508t4867 n7509 n4868 R=4.604e+00 
R7508t3139 n7509 n3140 R=4.540e+00 
R7509t2809 n7510 n2810 R=3.355e+00 
R7509t5818 n7510 n5819 R=7.687e+00 
R7509t4078 n7510 n4079 R=1.220e+01 
R7509t3811 n7510 n3812 R=8.279e+00 
R7509t1450 n7510 n1451 R=3.755e+00 
R7510t1176 n7511 n1177 R=8.257e+00 
R7510t2176 n7511 n2177 R=1.322e+01 
R7510t2177 n7511 n2178 R=2.472e+02 
R7510t2690 n7511 n2691 R=2.529e+01 
R7510t2995 n7511 n2996 R=7.665e+01 
R7510t2597 n7511 n2598 R=3.665e+00 
R7510t6814 n7511 n6815 R=3.425e+01 
R7510t3955 n7511 n3956 R=2.246e+01 
R7510t1111 n7511 n1112 R=1.241e+01 
R7511t1782 n7512 n1783 R=6.065e+00 
R7511t2635 n7512 n2636 R=8.859e+01 
R7511t5639 n7512 n5640 R=1.202e+01 
R7512t5031 n7513 n5032 R=2.082e+01 
R7512t4387 n7513 n4388 R=5.200e+00 
R7512t2880 n7513 n2881 R=8.462e+00 
R7513t1896 n7514 n1897 R=6.715e+00 
R7513t6421 n7514 n6422 R=6.333e+00 
R7513t7502 n7514 n7503 R=7.876e+00 
R7513t5198 n7514 n5199 R=1.017e+01 
R7513t3996 n7514 n3997 R=3.935e+00 
R7514t6231 n1 n6232 R=3.754e+00 
R7514t5708 n1 n5709 R=6.847e+00 
R7515t3456 n7516 n3457 R=3.486e+00 
R7515t6145 n7516 n6146 R=1.440e+02 
R7515t6353 n7516 n6354 R=1.180e+01 
R7515t3778 n7516 n3779 R=4.394e+00 
R7515t5715 n7516 n5716 R=5.801e+00 
R7515t6846 n7516 n6847 R=7.899e+01 
R7516t7376 n7517 n7377 R=3.474e+00 
R7516t6217 n7517 n6218 R=1.250e+00 
R7516t92 n7517 n93 R=2.021e+01 
R7517t4605 n7518 n4606 R=3.252e+00 
R7517t3712 n7518 n3713 R=4.084e+00 
R7517t6918 n7518 n6919 R=9.426e+00 
R7517t5829 n7518 n5830 R=7.023e+00 
R7518t2226 n7519 n2227 R=4.735e+00 
R7518t1808 n7519 n1809 R=1.876e+01 
R7519t4937 n7520 n4938 R=4.232e+00 
R7519t5244 n7520 n5245 R=9.196e+00 
R7519t5881 n7520 n5882 R=3.177e+01 
R7520t2319 n7521 n2320 R=1.611e+01 
R7520t6807 n7521 n6808 R=2.947e+01 
R7520t7372 n7521 n7373 R=2.860e+00 
R7521t5254 n7522 n5255 R=2.815e+00 
R7521t7305 n7522 n7306 R=3.389e+00 
R7521t3699 n7522 n3700 R=8.888e+00 
R7522t4397 n7523 n4398 R=1.812e+01 
R7522t5582 n7523 n5583 R=2.255e+00 
R7522t6841 n7523 n6842 R=1.742e+00 
R7522t3234 n7523 n3235 R=4.570e+01 
R7522t3651 n7523 n3652 R=1.330e+01 
R7523t1587 n7524 n1588 R=2.606e+00 
R7523t3054 n7524 n3055 R=2.526e+01 
R7523t6185 n7524 n6186 R=3.918e+00 
R7523t5702 n7524 n5703 R=5.158e+00 
R7524t2529 n7525 n2530 R=3.656e+01 
R7524t5820 n7525 n5821 R=6.426e+00 
R7524t7492 n7525 n7493 R=7.005e+00 
R7524t6875 n7525 n6876 R=7.092e+01 
R7524t5740 n7525 n5741 R=2.901e+00 
R7524t6567 n7525 n6568 R=2.560e+01 
R7525t34 n7526 n35 R=3.117e+00 
R7525t2972 n7526 n2973 R=5.034e+00 
R7525t4829 n7526 n4830 R=2.095e+02 
R7525t5726 n7526 n5727 R=4.366e+00 
R7525t3855 n7526 n3856 R=5.716e+00 
R7526t826 n7527 n827 R=5.427e+00 
R7526t6137 n7527 n6138 R=8.504e+00 
R7526t2729 n7527 n2730 R=1.638e+02 
R7526t4541 n7527 n4542 R=4.290e+00 
R7526t357 n7527 n358 R=3.926e+00 
R7526t3300 n7527 n3301 R=1.493e+01 
R7527t408 n7528 n409 R=2.115e+00 
R7527t6686 n7528 n6687 R=5.125e+01 
R7527t7144 n7528 n7145 R=6.210e+01 
R7527t3953 n7528 n3954 R=7.661e+00 
R7527t3195 n7528 n3196 R=1.163e+02 
R7528t3723 n7529 n3724 R=1.583e+01 
R7528t7233 n7529 n7234 R=8.645e+00 
R7528t7114 n7529 n7115 R=1.016e+01 
R7528t6114 n7529 n6115 R=4.345e+00 
R7528t2038 n7529 n2039 R=4.466e+01 
R7529t3331 n7530 n3332 R=1.528e+01 
R7529t6082 n7530 n6083 R=1.508e+00 
R7529t6560 n7530 n6561 R=2.540e+00 
R7529t5344 n7530 n5345 R=8.550e+00 
R7530t4629 n7531 n4630 R=2.875e+00 
R7530t6006 n7531 n6007 R=1.317e+01 
R7530t1364 n7531 n1365 R=6.143e+00 
R7531t4066 n7532 n4067 R=8.465e+00 
R7531t682 n7532 n683 R=2.809e+01 
R7531t4290 n7532 n4291 R=6.115e+01 
R7531t1710 n7532 n1711 R=3.903e+00 
R7532t5325 n7533 n5326 R=3.130e+01 
R7532t3106 n7533 n3107 R=2.424e+01 
R7532t6629 n7533 n6630 R=4.293e+01 
R7532t287 n7533 n288 R=2.091e+01 
R7532t3911 n7533 n3912 R=2.401e+00 
R7532t2547 n7533 n2548 R=3.922e+01 
R7532t3620 n7533 n3621 R=4.208e+00 
R7533t4607 n7534 n4608 R=3.997e+01 
R7533t5844 n7534 n5845 R=5.386e+00 
R7533t5574 n7534 n5575 R=4.387e+00 
R7533t524 n7534 n525 R=1.256e+01 
R7534t6019 n7535 n6020 R=8.559e+00 
R7534t7221 n7535 n7222 R=4.754e+00 
R7534t3283 n7535 n3284 R=2.657e+00 
R7534t2846 n7535 n2847 R=1.665e+01 
R7534t5660 n7535 n5661 R=6.779e+00 
R7535t5926 n7536 n5927 R=2.155e+01 
R7535t3584 n7536 n3585 R=1.734e+01 
R7535t543 n7536 n544 R=2.474e+00 
R7535t1735 n7536 n1736 R=1.194e+01 
R7536t4259 n7537 n4260 R=5.473e+00 
R7536t6965 n7537 n6966 R=2.357e+01 
R7536t4707 n7537 n4708 R=1.094e+01 
R7536t7382 n7537 n7383 R=6.422e+00 
R7536t6161 n7537 n6162 R=2.952e+01 
R7536t552 n7537 n553 R=3.418e+00 
R7537t4511 n7538 n4512 R=7.207e+00 
R7537t5691 n7538 n5692 R=7.713e+00 
R7537t4675 n7538 n4676 R=7.381e+00 
R7537t3525 n7538 n3526 R=1.086e+01 
R7537t6324 n7538 n6325 R=2.289e+01 
R7537t6382 n7538 n6383 R=4.597e+00 
R7538t8 n7539 n9 R=2.927e+00 
R7538t5346 n7539 n5347 R=1.318e+01 
R7538t6871 n7539 n6872 R=1.745e+01 
R7538t4951 n7539 n4952 R=1.946e+04 
R7539t6782 n7540 n6783 R=6.447e+00 
R7540t1436 n7541 n1437 R=1.987e+00 
R7540t5969 n7541 n5970 R=7.466e+00 
R7541t1423 n7542 n1424 R=5.446e+00 
R7541t5364 n7542 n5365 R=2.087e+02 
R7541t7093 n7542 n7094 R=3.389e+00 
R7541t3121 n7542 n3122 R=6.442e+02 
R7541t3280 n7542 n3281 R=7.135e+00 
R7541t5172 n7542 n5173 R=4.176e+00 
R7541t2093 n7542 n2094 R=2.166e+01 
R7542t3169 n7543 n3170 R=1.137e+01 
R7542t7471 n7543 n7472 R=6.333e+01 
R7542t5427 n7543 n5428 R=1.279e+01 
R7542t7280 n7543 n7281 R=4.064e+00 
R7543t7216 n7544 n7217 R=3.106e+01 
R7543t446 n7544 n447 R=4.394e+00 
R7543t4299 n7544 n4300 R=2.475e+01 
R7543t2061 n7544 n2062 R=6.783e+00 
R7543t1034 n7544 n1035 R=6.498e+00 
R7543t5921 n7544 n5922 R=1.076e+03 
R7544t3195 n7545 n3196 R=4.252e+00 
R7544t6686 n7545 n6687 R=5.875e+00 
R7544t7115 n7545 n7116 R=3.274e+00 
R7544t5311 n7545 n5312 R=1.807e+01 
R7544t865 n7545 n866 R=2.183e+01 
R7544t5981 n7545 n5982 R=4.193e+01 
R7545t4656 n7546 n4657 R=4.770e+00 
R7545t6616 n7546 n6617 R=5.330e+00 
R7545t5249 n7546 n5250 R=6.282e+00 
R7545t3800 n7546 n3801 R=4.229e+00 
R7546t3830 n7547 n3831 R=2.683e+00 
R7546t6772 n7547 n6773 R=2.566e+02 
R7546t1217 n7547 n1218 R=3.173e+00 
R7546t3801 n7547 n3802 R=7.377e+00 
R7546t464 n7547 n465 R=9.893e+00 
R7547t594 n7548 n595 R=1.234e+01 
R7547t2150 n7548 n2151 R=5.215e+01 
R7547t4028 n7548 n4029 R=3.693e+00 
R7547t1198 n7548 n1199 R=5.115e+00 
R7548t4456 n7549 n4457 R=2.429e+01 
R7548t898 n7549 n899 R=2.584e+00 
R7548t4310 n7549 n4311 R=1.562e+01 
R7549t291 n7550 n292 R=1.622e+01 
R7549t6281 n7550 n6282 R=1.174e+01 
R7549t5866 n7550 n5867 R=5.926e+00 
R7549t639 n7550 n640 R=2.796e+00 
R7549t6759 n7550 n6760 R=5.891e+00 
R7550t6798 n7551 n6799 R=2.081e+01 
R7550t6863 n7551 n6864 R=1.290e+02 
R7550t2998 n7551 n2999 R=4.158e+01 
R7550t4938 n7551 n4939 R=4.946e+00 
R7550t5564 n7551 n5565 R=5.171e+00 
R7550t2231 n7551 n2232 R=6.029e+00 
R7550t343 n7551 n344 R=7.053e+00 
R7551t94 n7552 n95 R=7.870e+00 
R7551t5609 n7552 n5610 R=3.446e+00 
R7551t3310 n7552 n3311 R=5.816e+01 
R7551t2512 n7552 n2513 R=6.465e+00 
R7551t1752 n7552 n1753 R=6.925e+00 
R7551t6331 n7552 n6332 R=2.013e+01 
R7551t2978 n7552 n2979 R=3.907e+01 
R7552t6074 n7553 n6075 R=4.245e+01 
R7552t4567 n7553 n4568 R=3.061e+00 
R7552t7002 n7553 n7003 R=2.813e+01 
R7552t6977 n7553 n6978 R=2.974e+00 
R7552t1469 n7553 n1470 R=5.340e+00 
R7553t2027 n7554 n2028 R=3.355e+00 
R7553t3700 n7554 n3701 R=4.072e+00 
R7553t6697 n7554 n6698 R=3.225e+00 
R7554t7328 n7555 n7329 R=5.580e+00 
R7554t2080 n7555 n2081 R=1.726e+01 
R7554t4657 n7555 n4658 R=4.045e+00 
R7555t5282 n7556 n5283 R=4.949e+00 
R7555t6842 n7556 n6843 R=1.001e+01 
R7555t1082 n7556 n1083 R=5.921e+00 
R7555t3303 n7556 n3304 R=2.183e+01 
R7555t3432 n7556 n3433 R=5.876e+00 
R7556t4687 n7557 n4688 R=4.949e+00 
R7556t5770 n7557 n5771 R=1.047e+01 
R7556t150 n7557 n151 R=7.454e+00 
R7557t2896 n7558 n2897 R=4.811e+01 
R7557t1272 n7558 n1273 R=4.167e+00 
R7557t3655 n7558 n3656 R=5.897e+01 
R7557t2754 n7558 n2755 R=1.889e+01 
R7557t524 n7558 n525 R=1.393e+02 
R7558t1927 n7559 n1928 R=2.718e+00 
R7558t2392 n7559 n2393 R=5.822e+00 
R7558t2005 n7559 n2006 R=9.817e+00 
R7558t6373 n7559 n6374 R=3.873e+00 
R7559t272 n7560 n273 R=3.308e+00 
R7559t378 n7560 n379 R=1.003e+01 
R7559t1303 n7560 n1304 R=3.212e+00 
R7559t1950 n7560 n1951 R=3.028e+01 
R7560t3572 n7561 n3573 R=6.462e+00 
R7560t5359 n7561 n5360 R=1.621e+01 
R7560t6185 n7561 n6186 R=2.682e+01 
R7560t1571 n7561 n1572 R=4.828e+00 
R7561t9 n7562 n10 R=3.327e+00 
R7561t1826 n7562 n1827 R=3.381e+00 
R7562t3878 n7563 n3879 R=2.915e+00 
R7563t879 n7564 n880 R=3.976e+00 
R7563t1128 n7564 n1129 R=2.403e+00 
R7563t5201 n7564 n5202 R=1.575e+01 
R7563t4075 n7564 n4076 R=4.634e+00 
R7564t2505 n7565 n2506 R=1.285e+01 
R7564t3007 n7565 n3008 R=4.706e+00 
R7564t4165 n7565 n4166 R=1.862e+01 
R7564t335 n7565 n336 R=2.188e+01 
R7564t1251 n7565 n1252 R=5.429e+00 
R7564t3686 n7565 n3687 R=4.115e+01 
R7565t3215 n7566 n3216 R=2.123e+01 
R7565t2560 n7566 n2561 R=4.209e+01 
R7565t2703 n7566 n2704 R=1.218e+01 
R7565t4258 n7566 n4259 R=2.109e+01 
R7565t5624 n7566 n5625 R=1.082e+01 
R7565t1789 n7566 n1790 R=2.863e+00 
R7566t495 n7567 n496 R=7.786e+00 
R7566t3537 n7567 n3538 R=4.092e+01 
R7566t5377 n7567 n5378 R=3.083e+00 
R7566t214 n7567 n215 R=1.351e+01 
R7566t1556 n7567 n1557 R=2.075e+01 
R7567t5252 n7568 n5253 R=1.275e+00 
R7567t6334 n7568 n6335 R=2.237e+01 
R7567t543 n7568 n544 R=1.471e+01 
R7567t4159 n7568 n4160 R=3.782e+00 
R7567t390 n7568 n391 R=2.564e+01 
R7567t2521 n7568 n2522 R=1.078e+01 
R7568t411 n7569 n412 R=2.587e+03 
R7568t862 n7569 n863 R=7.068e+00 
R7568t7013 n7569 n7014 R=2.708e+00 
R7568t3198 n7569 n3199 R=8.156e+00 
R7569t1660 n7570 n1661 R=6.338e+01 
R7570t1203 n7571 n1204 R=9.538e+00 
R7570t2246 n7571 n2247 R=1.580e+01 
R7570t3311 n7571 n3312 R=6.870e+00 
R7570t6584 n7571 n6585 R=6.911e+02 
R7570t5137 n7571 n5138 R=5.170e+00 
R7571t4905 n7572 n4906 R=2.980e+00 
R7571t7003 n7572 n7004 R=1.363e+00 
R7572t3207 n7573 n3208 R=1.649e+01 
R7572t4576 n7573 n4577 R=2.348e+01 
R7572t1588 n7573 n1589 R=5.729e+00 
R7572t4078 n7573 n4079 R=9.868e+00 
R7572t4023 n7573 n4024 R=1.185e+01 
R7572t5952 n7573 n5953 R=5.311e+00 
R7572t5015 n7573 n5016 R=7.919e+01 
R7573t2526 n7574 n2527 R=2.195e+01 
R7573t4627 n7574 n4628 R=1.413e+01 
R7573t6081 n7574 n6082 R=3.706e+00 
R7574t1912 n7575 n1913 R=7.424e+00 
R7574t4032 n7575 n4033 R=2.967e+00 
R7574t5572 n7575 n5573 R=4.952e+01 
R7574t1389 n7575 n1390 R=2.370e+00 
R7574t1104 n7575 n1105 R=1.103e+01 
R7575t809 n7576 n810 R=2.624e+00 
R7575t5500 n7576 n5501 R=3.473e+01 
R7575t4184 n7576 n4185 R=5.992e+00 
R7576t828 n7577 n829 R=3.975e+00 
R7576t6548 n7577 n6549 R=1.751e+01 
R7576t1232 n7577 n1233 R=4.940e+01 
R7576t5950 n7577 n5951 R=1.108e+01 
R7576t3167 n7577 n3168 R=2.603e+00 
R7577t2694 n7578 n2695 R=4.833e+00 
R7577t3304 n7578 n3305 R=1.179e+01 
R7577t849 n7578 n850 R=2.282e+01 
R7577t6645 n7578 n6646 R=2.759e+01 
R7577t2689 n7578 n2690 R=7.828e+00 
R7577t1843 n7578 n1844 R=5.052e+00 
R7577t4714 n7578 n4715 R=1.201e+02 
R7577t3706 n7578 n3707 R=1.027e+01 
R7578t1382 n7579 n1383 R=3.320e+00 
R7578t7178 n7579 n7179 R=1.152e+01 
R7579t1835 n7580 n1836 R=8.836e+00 
R7579t4575 n7580 n4576 R=3.313e+01 
R7579t2185 n7580 n2186 R=4.388e+00 
R7579t7098 n7580 n7099 R=2.196e+01 
R7579t2140 n7580 n2141 R=6.585e+00 
R7579t2407 n7580 n2408 R=1.051e+01 
R7580t1361 n7581 n1362 R=4.509e+00 
R7580t1565 n7581 n1566 R=1.422e+01 
R7580t3334 n7581 n3335 R=2.363e+01 
R7580t4902 n7581 n4903 R=1.898e+01 
R7580t7074 n7581 n7075 R=5.329e+00 
R7581t6895 n7582 n6896 R=7.975e+00 
R7581t7131 n7582 n7132 R=3.069e+00 
R7581t4518 n7582 n4519 R=3.763e+02 
R7581t7390 n7582 n7391 R=3.120e+00 
R7581t2735 n7582 n2736 R=1.173e+01 
R7582t1462 n7583 n1463 R=5.066e+00 
R7582t3985 n7583 n3986 R=7.706e+01 
R7582t732 n7583 n733 R=2.476e+00 
R7582t2118 n7583 n2119 R=5.623e+02 
R7583t4519 n7584 n4520 R=4.350e+00 
R7583t6888 n7584 n6889 R=1.896e+02 
R7583t6583 n7584 n6584 R=4.916e+00 
R7583t517 n7584 n518 R=5.500e+01 
R7583t3607 n7584 n3608 R=3.492e+01 
R7583t3715 n7584 n3716 R=4.158e+01 
R7583t1407 n7584 n1408 R=4.479e+00 
R7584t780 n7585 n781 R=9.539e+00 
R7584t6857 n7585 n6858 R=6.831e+00 
R7584t6135 n7585 n6136 R=2.160e+01 
R7584t320 n7585 n321 R=2.167e+01 
R7584t144 n7585 n145 R=8.203e+00 
R7584t4810 n7585 n4811 R=1.498e+01 
R7585t1693 n7586 n1694 R=1.250e+01 
R7585t3810 n7586 n3811 R=4.654e+00 
R7585t5621 n7586 n5622 R=5.802e+00 
R7586t6072 n7587 n6073 R=2.275e+00 
R7586t1266 n7587 n1267 R=4.643e+00 
R7587t1942 n7588 n1943 R=1.018e+01 
R7587t6631 n7588 n6632 R=3.363e+00 
R7587t387 n7588 n388 R=3.963e+00 
R7587t2348 n7588 n2349 R=4.297e+00 
R7588t3530 n7589 n3531 R=1.389e+01 
R7588t3594 n7589 n3595 R=2.159e+00 
R7588t7102 n7589 n7103 R=7.386e+00 
R7588t544 n7589 n545 R=7.571e+00 
R7589t1275 n7590 n1276 R=2.244e+01 
R7589t3366 n7590 n3367 R=4.756e+00 
R7589t1827 n7590 n1828 R=4.405e+00 
R7589t39 n7590 n40 R=2.102e+00 
R7590t4884 n7591 n4885 R=4.759e+00 
R7590t7402 n7591 n7403 R=5.631e+00 
R7590t1471 n7591 n1472 R=6.728e+00 
R7590t1175 n7591 n1176 R=4.507e+00 
R7591t4333 n7592 n4334 R=2.956e+01 
R7591t4826 n7592 n4827 R=5.293e+00 
R7591t7484 n7592 n7485 R=2.267e+00 
R7591t5575 n7592 n5576 R=4.115e+00 
R7592t742 n7593 n743 R=1.621e+00 
R7592t1587 n7593 n1588 R=2.041e+01 
R7592t3054 n7593 n3055 R=2.297e+01 
R7592t7046 n7593 n7047 R=2.590e+00 
R7592t5835 n7593 n5836 R=8.658e+00 
R7592t4241 n7593 n4242 R=1.607e+01 
R7592t3692 n7593 n3693 R=1.260e+03 
R7592t1981 n7593 n1982 R=8.329e+00 
R7593t6326 n7594 n6327 R=6.534e+00 
R7593t3790 n7594 n3791 R=4.585e+00 
R7593t6789 n7594 n6790 R=3.818e+01 
R7593t2989 n7594 n2990 R=7.140e+01 
R7593t1701 n7594 n1702 R=5.177e+00 
R7593t5571 n7594 n5572 R=4.136e+01 
R7593t6529 n7594 n6530 R=8.060e+00 
R7594t2782 n7595 n2783 R=4.745e+00 
R7594t5362 n7595 n5363 R=8.361e+01 
R7594t3086 n7595 n3087 R=5.481e+00 
R7594t4784 n7595 n4785 R=6.835e+00 
R7595t301 n7596 n302 R=6.634e+01 
R7595t2463 n7596 n2464 R=6.701e+02 
R7595t6901 n7596 n6902 R=5.150e+02 
R7595t5275 n7596 n5276 R=3.303e+00 
R7595t5512 n7596 n5513 R=2.966e+00 
R7596t4291 n7597 n4292 R=1.252e+02 
R7596t6206 n7597 n6207 R=5.341e+00 
R7596t5219 n7597 n5220 R=3.338e+01 
R7596t6204 n7597 n6205 R=7.140e+01 
R7596t6792 n7597 n6793 R=7.190e+00 
R7596t7079 n7597 n7080 R=4.083e+00 
R7596t4111 n7597 n4112 R=7.588e+01 
R7596t2440 n7597 n2441 R=6.550e+00 
R7597t1160 n7598 n1161 R=7.276e+00 
R7597t2891 n7598 n2892 R=5.818e+00 
R7597t3777 n7598 n3778 R=8.211e+00 
R7597t332 n7598 n333 R=1.014e+03 
R7598t1578 n7599 n1579 R=2.584e+03 
R7598t2484 n7599 n2485 R=2.544e+00 
R7598t7194 n7599 n7195 R=4.263e+01 
R7598t244 n7599 n245 R=3.808e+00 
R7598t6788 n7599 n6789 R=2.420e+01 
R7599t4342 n7600 n4343 R=1.255e+01 
R7599t4912 n7600 n4913 R=6.852e+00 
R7599t2973 n7600 n2974 R=4.439e+00 
R7599t1690 n7600 n1691 R=1.630e+01 
R7599t150 n7600 n151 R=7.188e+00 
R7599t3446 n7600 n3447 R=1.820e+01 
R7600t1761 n7601 n1762 R=9.823e+00 
R7600t4644 n7601 n4645 R=2.851e+00 
R7600t2662 n7601 n2663 R=9.643e+00 
R7600t7336 n7601 n7337 R=5.509e+00 
R7601t687 n7602 n688 R=2.325e+01 
R7601t5547 n7602 n5548 R=6.424e+00 
R7601t6799 n7602 n6800 R=2.005e+01 
R7601t5940 n7602 n5941 R=1.611e+01 
R7601t4949 n7602 n4950 R=4.374e+00 
R7601t3864 n7602 n3865 R=2.050e+00 
R7602t39 n7603 n40 R=2.537e+02 
R7602t1748 n7603 n1749 R=2.620e+00 
R7602t7589 n7603 n7590 R=2.006e+01 
R7602t1827 n7603 n1828 R=7.415e+00 
R7602t5152 n7603 n5153 R=2.543e+00 
R7603t2043 n7604 n2044 R=2.647e+00 
R7603t4009 n7604 n4010 R=1.091e+01 
R7603t3702 n7604 n3703 R=6.751e+00 
R7603t7167 n7604 n7168 R=7.714e+01 
R7604t4434 n7605 n4435 R=5.302e+00 
R7604t6468 n7605 n6469 R=6.033e+00 
R7604t761 n7605 n762 R=5.993e+00 
R7604t2947 n7605 n2948 R=2.787e+01 
R7604t5571 n7605 n5572 R=6.708e+00 
R7604t2989 n7605 n2990 R=3.477e+01 
R7605t498 n7606 n499 R=2.627e+00 
R7605t2655 n7606 n2656 R=1.403e+01 
R7605t4044 n7606 n4045 R=4.331e+01 
R7605t3986 n7606 n3987 R=1.315e+01 
R7605t349 n7606 n350 R=4.046e+00 
R7606t7342 n7607 n7343 R=1.938e+01 
R7606t3947 n7607 n3948 R=6.088e+00 
R7606t5865 n7607 n5866 R=6.858e+00 
R7606t5546 n7607 n5547 R=1.375e+01 
R7607t1741 n7608 n1742 R=2.223e+01 
R7607t2364 n7608 n2365 R=1.317e+01 
R7607t5751 n7608 n5752 R=9.662e+00 
R7607t5480 n7608 n5481 R=3.979e+00 
R7607t3018 n7608 n3019 R=5.131e+00 
R7608t377 n7609 n378 R=8.544e+01 
R7608t2170 n7609 n2171 R=2.262e+00 
R7608t4272 n7609 n4273 R=1.048e+01 
R7608t836 n7609 n837 R=3.859e+00 
R7608t890 n7609 n891 R=1.313e+01 
R7608t155 n7609 n156 R=1.479e+01 
R7609t6618 n7610 n6619 R=1.349e+01 
R7609t967 n7610 n968 R=3.713e+01 
R7609t2168 n7610 n2169 R=7.641e+00 
R7609t201 n7610 n202 R=3.659e+00 
R7610t2970 n7611 n2971 R=9.126e+01 
R7610t5317 n7611 n5318 R=2.689e+00 
R7610t532 n7611 n533 R=2.417e+01 
R7610t7327 n7611 n7328 R=4.996e+00 
R7610t5130 n7611 n5131 R=4.392e+00 
R7611t6556 n7612 n6557 R=1.238e+01 
R7611t7357 n7612 n7358 R=7.572e+00 
R7611t1581 n7612 n1582 R=4.407e+00 
R7611t5599 n7612 n5600 R=1.873e+01 
R7611t6112 n7612 n6113 R=1.146e+01 
R7611t2244 n7612 n2245 R=6.306e+00 
R7611t2293 n7612 n2294 R=9.165e+00 
R7612t6141 n7613 n6142 R=3.436e+00 
R7612t7486 n7613 n7487 R=3.188e+00 
R7612t3176 n7613 n3177 R=1.040e+02 
R7613t935 n7614 n936 R=1.209e+01 
R7613t1636 n7614 n1637 R=5.112e+00 
R7613t2878 n7614 n2879 R=5.367e+00 
R7613t4619 n7614 n4620 R=2.413e+01 
R7614t843 n7615 n844 R=7.445e+00 
R7614t2651 n7615 n2652 R=2.227e+01 
R7614t209 n7615 n210 R=1.039e+01 
R7614t6749 n7615 n6750 R=4.162e+00 
R7614t4098 n7615 n4099 R=1.345e+01 
R7614t425 n7615 n426 R=1.765e+02 
R7615t664 n7616 n665 R=1.034e+01 
R7615t5323 n7616 n5324 R=2.652e+01 
R7615t2311 n7616 n2312 R=2.020e+01 
R7615t4762 n7616 n4763 R=1.104e+01 
R7615t7004 n7616 n7005 R=1.693e+01 
R7615t2110 n7616 n2111 R=3.244e+00 
R7615t2117 n7616 n2118 R=4.453e+00 
R7616t2619 n7617 n2620 R=6.925e+00 
R7616t6899 n7617 n6900 R=6.924e+00 
R7616t4992 n7617 n4993 R=3.799e+01 
R7616t4089 n7617 n4090 R=6.666e+00 
R7617t1266 n7618 n1267 R=1.414e+01 
R7617t5772 n7618 n5773 R=1.224e+01 
R7617t5766 n7618 n5767 R=4.050e+01 
R7617t6541 n7618 n6542 R=6.948e+01 
R7617t4608 n7618 n4609 R=3.293e+00 
R7617t4817 n7618 n4818 R=1.459e+01 
R7617t2944 n7618 n2945 R=2.417e+01 
R7618t436 n7619 n437 R=6.426e+00 
R7618t762 n7619 n763 R=2.687e+01 
R7618t3538 n7619 n3539 R=7.714e+00 
R7618t636 n7619 n637 R=4.645e+00 
R7618t5290 n7619 n5291 R=8.715e+00 
R7619t7408 n7620 n7409 R=2.825e+00 
R7619t1600 n7620 n1601 R=3.190e+00 
R7619t4818 n7620 n4819 R=8.012e+00 
R7620t6379 n7621 n6380 R=5.663e+01 
R7620t881 n7621 n882 R=1.796e+01 
R7620t3029 n7621 n3030 R=1.114e+01 
R7621t248 n7622 n249 R=2.256e+01 
R7621t3182 n7622 n3183 R=9.282e+00 
R7621t984 n7622 n985 R=4.080e+00 
R7621t7573 n7622 n7574 R=5.019e+00 
R7621t2526 n7622 n2527 R=4.595e+01 
R7621t2736 n7622 n2737 R=3.032e+01 
R7622t408 n7623 n409 R=3.287e+00 
R7622t5471 n7623 n5472 R=1.873e+00 
R7622t1046 n7623 n1047 R=4.182e+00 
R7623t1872 n7624 n1873 R=5.246e+00 
R7623t3456 n7624 n3457 R=1.580e+01 
R7623t6504 n7624 n6505 R=3.557e+00 
R7623t4252 n7624 n4253 R=4.894e+01 
R7623t6353 n7624 n6354 R=6.682e+00 
R7623t7515 n7624 n7516 R=1.275e+01 
R7624t4740 n7625 n4741 R=1.869e+01 
R7624t235 n7625 n236 R=1.402e+02 
R7624t6317 n7625 n6318 R=5.282e+00 
R7624t6484 n7625 n6485 R=4.454e+01 
R7625t103 n7626 n104 R=9.110e+00 
R7625t5865 n7626 n5866 R=3.140e+00 
R7625t7606 n7626 n7607 R=2.358e+01 
R7625t3947 n7626 n3948 R=1.249e+01 
R7626t3591 n7627 n3592 R=9.567e+00 
R7626t4943 n7627 n4944 R=4.189e+00 
R7626t1535 n7627 n1536 R=9.996e+01 
R7626t1738 n7627 n1739 R=4.991e+00 
R7626t1108 n7627 n1109 R=8.883e+00 
R7627t4496 n7628 n4497 R=4.185e+00 
R7627t3794 n7628 n3795 R=5.391e+00 
R7627t6260 n7628 n6261 R=9.893e+01 
R7627t5011 n7628 n5012 R=5.159e+00 
R7628t274 n7629 n275 R=1.669e+01 
R7628t3644 n7629 n3645 R=2.917e+01 
R7628t4654 n7629 n4655 R=1.894e+00 
R7628t2641 n7629 n2642 R=4.076e+01 
R7628t5150 n7629 n5151 R=2.715e+00 
R7628t3152 n7629 n3153 R=3.744e+01 
R7629t4492 n7630 n4493 R=1.026e+02 
R7629t2594 n7630 n2595 R=9.961e+00 
R7629t6793 n7630 n6794 R=2.816e+00 
R7629t2347 n7630 n2348 R=1.413e+01 
R7629t2242 n7630 n2243 R=2.669e+00 
R7630t1160 n7631 n1161 R=6.857e+01 
R7630t4874 n7631 n4875 R=1.461e+01 
R7630t6975 n7631 n6976 R=1.086e+01 
R7630t7189 n7631 n7190 R=1.069e+01 
R7630t3119 n7631 n3120 R=1.216e+02 
R7630t3647 n7631 n3648 R=4.266e+00 
R7630t332 n7631 n333 R=4.529e+01 
R7631t3934 n7632 n3935 R=1.978e+00 
R7631t7463 n7632 n7464 R=5.078e+01 
R7631t2953 n7632 n2954 R=7.588e+00 
R7632t997 n7633 n998 R=1.104e+01 
R7632t5036 n7633 n5037 R=4.831e+00 
R7632t80 n7633 n81 R=7.087e+00 
R7632t2294 n7633 n2295 R=2.167e+02 
R7632t6184 n7633 n6185 R=5.271e+00 
R7632t7429 n7633 n7430 R=8.448e+00 
R7633t1806 n7634 n1807 R=4.815e+00 
R7633t3885 n7634 n3886 R=9.110e+00 
R7633t1247 n7634 n1248 R=7.558e+00 
R7633t5627 n7634 n5628 R=3.024e+01 
R7633t3875 n7634 n3876 R=4.649e+00 
R7633t2874 n7634 n2875 R=1.175e+01 
R7634t1148 n7635 n1149 R=1.276e+01 
R7634t579 n7635 n580 R=7.473e+00 
R7634t5842 n7635 n5843 R=1.712e+01 
R7634t7245 n7635 n7246 R=1.667e+01 
R7634t2111 n7635 n2112 R=6.668e+00 
R7635t4277 n7636 n4278 R=7.212e+00 
R7635t4754 n7636 n4755 R=1.393e+02 
R7635t1063 n7636 n1064 R=4.963e+00 
R7635t6232 n7636 n6233 R=3.862e+01 
R7636t1530 n7637 n1531 R=5.869e+00 
R7636t137 n7637 n138 R=1.941e+00 
R7636t6109 n7637 n6110 R=1.320e+01 
R7636t1069 n7637 n1070 R=4.340e+00 
R7637t1860 n7638 n1861 R=1.274e+01 
R7637t7133 n7638 n7134 R=1.775e+01 
R7637t1585 n7638 n1586 R=3.965e+00 
R7637t3295 n7638 n3296 R=1.178e+01 
R7637t5880 n7638 n5881 R=1.360e+01 
R7637t7136 n7638 n7137 R=3.796e+00 
R7637t3261 n7638 n3262 R=2.556e+01 
R7638t2466 n7639 n2467 R=7.626e+00 
R7638t3362 n7639 n3363 R=1.188e+01 
R7638t3774 n7639 n3775 R=2.133e+01 
R7638t3451 n7639 n3452 R=3.629e+00 
R7639t1136 n7640 n1137 R=1.635e+02 
R7639t3611 n7640 n3612 R=2.229e+01 
R7639t6682 n7640 n6683 R=8.376e+00 
R7639t4224 n7640 n4225 R=1.921e+00 
R7640t4911 n7641 n4912 R=5.129e+00 
R7640t3604 n7641 n3605 R=4.976e+00 
R7640t2033 n7641 n2034 R=4.984e+02 
R7640t196 n7641 n197 R=7.967e+00 
R7641t2601 n7642 n2602 R=3.219e+00 
R7641t7498 n7642 n7499 R=1.438e+01 
R7641t5880 n7642 n5881 R=8.275e+00 
R7641t6411 n7642 n6412 R=2.279e+00 
R7642t4789 n7643 n4790 R=9.208e+01 
R7642t2232 n7643 n2233 R=2.416e+01 
R7643t2384 n7644 n2385 R=2.525e+01 
R7643t2783 n7644 n2784 R=3.772e+00 
R7643t5515 n7644 n5516 R=8.954e+00 
R7643t4304 n7644 n4305 R=5.116e+00 
R7643t6989 n7644 n6990 R=5.088e+01 
R7644t5097 n7645 n5098 R=1.345e+01 
R7644t5518 n7645 n5519 R=4.884e+00 
R7644t5224 n7645 n5225 R=6.793e+00 
R7644t2621 n7645 n2622 R=9.749e+00 
R7645t3198 n7646 n3199 R=7.866e+00 
R7645t6471 n7646 n6472 R=7.243e+01 
R7645t5505 n7646 n5506 R=3.648e+01 
R7645t4684 n7646 n4685 R=2.715e+00 
R7645t4380 n7646 n4381 R=9.219e+01 
R7645t3567 n7646 n3568 R=1.606e+01 
R7645t296 n7646 n297 R=1.679e+01 
R7645t3125 n7646 n3126 R=7.485e+00 
R7645t7013 n7646 n7014 R=1.203e+02 
R7646t1282 n7647 n1283 R=1.760e+00 
R7646t5722 n7647 n5723 R=3.110e+01 
R7646t2798 n7647 n2799 R=3.525e+00 
R7646t6136 n7647 n6137 R=6.198e+00 
R7647t434 n7648 n435 R=7.824e+00 
R7647t1448 n7648 n1449 R=1.240e+01 
R7647t1442 n7648 n1443 R=4.371e+00 
R7647t4204 n7648 n4205 R=2.456e+01 
R7648t5059 n7649 n5060 R=7.977e+00 
R7648t5728 n7649 n5729 R=4.613e+00 
R7648t2811 n7649 n2812 R=1.022e+01 
R7648t1513 n7649 n1514 R=2.524e+00 
R7648t4128 n7649 n4129 R=7.829e+01 
R7649t1292 n7650 n1293 R=6.013e+00 
R7649t6928 n7650 n6929 R=5.561e+00 
R7649t7188 n7650 n7189 R=2.867e+01 
R7649t4751 n7650 n4752 R=9.007e+00 
R7650t5116 n7651 n5117 R=1.002e+01 
R7650t6434 n7651 n6435 R=7.246e+00 
R7650t5888 n7651 n5889 R=1.031e+01 
R7650t6100 n7651 n6101 R=6.343e+00 
R7650t5659 n7651 n5660 R=7.285e+00 
R7651t1362 n7652 n1363 R=1.571e+01 
R7651t3319 n7652 n3320 R=2.656e+00 
R7651t5446 n7652 n5447 R=1.100e+01 
R7651t2790 n7652 n2791 R=5.959e+00 
R7651t2831 n7652 n2832 R=1.003e+01 
R7651t2382 n7652 n2383 R=5.225e+01 
R7651t2794 n7652 n2795 R=8.472e+00 
R7652t347 n7653 n348 R=3.643e+00 
R7652t6064 n7653 n6065 R=3.235e+01 
R7652t3489 n7653 n3490 R=1.891e+01 
R7652t4549 n7653 n4550 R=2.417e+01 
R7652t7065 n7653 n7066 R=7.815e+00 
R7653t5736 n7654 n5737 R=6.599e+00 
R7653t3320 n7654 n3321 R=3.146e+02 
R7653t1755 n7654 n1756 R=1.943e+02 
R7653t4542 n7654 n4543 R=3.885e+00 
R7653t4394 n7654 n4395 R=1.519e+01 
R7654t1798 n7655 n1799 R=2.206e+00 
R7654t6132 n7655 n6133 R=7.180e+00 
R7654t799 n7655 n800 R=1.592e+00 
R7654t4071 n7655 n4072 R=1.961e+01 
R7655t1645 n7656 n1646 R=1.056e+01 
R7655t678 n7656 n679 R=2.503e+00 
R7655t7259 n7656 n7260 R=1.116e+01 
R7656t2356 n1 n2357 R=6.668e+01 
R7656t1728 n1 n1729 R=9.920e+00 
R7656t4982 n1 n4983 R=4.633e+00 
R7657t1692 n7658 n1693 R=5.172e+00 
R7657t5767 n7658 n5768 R=5.229e+00 
R7658t3110 n7659 n3111 R=3.205e+00 
R7658t2534 n7659 n2535 R=1.330e+01 
R7658t3212 n7659 n3213 R=4.261e+00 
R7658t3714 n7659 n3715 R=9.955e+00 
R7659t4806 n7660 n4807 R=3.522e+00 
R7659t6225 n7660 n6226 R=5.546e+00 
R7659t985 n7660 n986 R=8.330e+00 
R7659t1732 n7660 n1733 R=2.440e+01 
R7659t5603 n7660 n5604 R=4.754e+00 
R7660t3386 n7661 n3387 R=9.120e+00 
R7660t7481 n7661 n7482 R=5.317e+00 
R7660t3883 n7661 n3884 R=9.746e+00 
R7660t4185 n7661 n4186 R=2.632e+01 
R7660t4191 n7661 n4192 R=9.259e+00 
R7660t4105 n7661 n4106 R=7.705e+00 
R7660t204 n7661 n205 R=1.214e+01 
R7661t3305 n7662 n3306 R=2.097e+01 
R7661t3426 n7662 n3427 R=4.375e+01 
R7661t2294 n7662 n2295 R=2.206e+01 
R7661t6586 n7662 n6587 R=4.927e+00 
R7661t2286 n7662 n2287 R=1.578e+01 
R7661t3038 n7662 n3039 R=6.082e+00 
R7661t530 n7662 n531 R=3.337e+00 
R7663t2649 n7664 n2650 R=1.156e+01 
R7663t876 n7664 n877 R=3.466e+00 
R7663t5795 n7664 n5796 R=7.850e+00 
R7663t3277 n7664 n3278 R=6.011e+01 
R7664t5440 n7665 n5441 R=6.004e+00 
R7664t6573 n7665 n6574 R=9.167e+00 
R7664t3744 n7665 n3745 R=1.713e+01 
R7664t6754 n7665 n6755 R=1.290e+01 
R7664t6204 n7665 n6205 R=4.827e+00 
R7664t111 n7665 n112 R=8.096e+00 
R7665t5824 n1 n5825 R=2.748e+00 
R7665t6368 n1 n6369 R=9.812e+01 
R7665t4758 n1 n4759 R=4.674e+01 
R7665t3437 n1 n3438 R=2.441e+01 
R7666t859 n7667 n860 R=1.111e+01 
R7666t7431 n7667 n7432 R=4.290e+00 
R7666t5548 n7667 n5549 R=8.970e+00 
R7666t888 n7667 n889 R=3.994e+00 
R7666t4215 n7667 n4216 R=7.765e+01 
R7666t3321 n7667 n3322 R=7.290e+00 
R7667t711 n7668 n712 R=5.488e+00 
R7667t3784 n7668 n3785 R=5.864e+00 
R7667t1314 n7668 n1315 R=3.401e+01 
R7667t959 n7668 n960 R=4.188e+00 
R7668t2200 n7669 n2201 R=2.464e+00 
R7668t2903 n7669 n2904 R=1.570e+01 
R7668t2347 n7669 n2348 R=1.985e+01 
R7668t6793 n7669 n6794 R=7.435e+00 
R7668t5993 n7669 n5994 R=5.083e+00 
R7668t1260 n7669 n1261 R=1.100e+02 
R7669t543 n7670 n544 R=1.936e+00 
R7669t3805 n7670 n3806 R=3.016e+00 
R7669t7567 n7670 n7568 R=2.857e+01 
R7669t4159 n7670 n4160 R=2.739e+00 
R7670t6173 n7671 n6174 R=4.292e+00 
R7670t6629 n7671 n6630 R=2.966e+00 
R7670t3702 n7671 n3703 R=1.256e+01 
R7671t3091 n1 n3092 R=3.786e+00 
R7671t6231 n1 n6232 R=2.795e+00 
R7672t2185 n7673 n2186 R=6.466e+00 
R7672t2187 n7673 n2188 R=3.063e+01 
R7672t4575 n7673 n4576 R=5.802e+00 
R7672t6153 n7673 n6154 R=6.182e+00 
R7672t6258 n7673 n6259 R=1.347e+01 
R7673t2466 n7674 n2467 R=7.496e+01 
R7673t7638 n7674 n7639 R=1.659e+01 
R7673t4360 n7674 n4361 R=6.732e+00 
R7673t2190 n7674 n2191 R=3.891e+00 
R7674t5794 n7675 n5795 R=2.152e+00 
R7674t5977 n7675 n5978 R=2.819e+00 
R7675t3801 n7676 n3802 R=2.607e+01 
R7675t6148 n7676 n6149 R=8.345e+01 
R7675t6479 n7676 n6480 R=6.719e+00 
R7675t4505 n7676 n4506 R=3.077e+00 
R7676t1328 n7677 n1329 R=3.588e+01 
R7676t163 n7677 n164 R=5.651e+00 
R7676t2916 n7677 n2917 R=3.794e+00 
R7676t735 n7677 n736 R=4.232e+01 
R7677t1048 n7678 n1049 R=6.882e+00 
R7677t3778 n7678 n3779 R=3.224e+00 
R7677t5715 n7678 n5716 R=1.032e+01 
R7677t746 n7678 n747 R=8.960e+00 
R7678t4782 n7679 n4783 R=3.075e+00 
R7678t4740 n7679 n4741 R=1.529e+01 
R7679t3021 n7680 n3022 R=6.007e+00 
R7679t3284 n7680 n3285 R=4.560e+00 
R7679t3365 n7680 n3366 R=1.163e+02 
R7679t2745 n7680 n2746 R=5.010e+00 
R7680t3661 n7681 n3662 R=2.444e+00 
R7680t3717 n7681 n3718 R=5.054e+00 
R7680t4314 n7681 n4315 R=1.185e+02 
R7680t279 n7681 n280 R=2.802e+00 
R7680t370 n7681 n371 R=1.113e+02 
R7681t1038 n7682 n1039 R=3.698e+02 
R7681t5173 n7682 n5174 R=4.747e+00 
R7681t2855 n7682 n2856 R=9.201e+00 
R7681t4538 n7682 n4539 R=3.346e+01 
R7681t6383 n7682 n6384 R=3.965e+00 
R7682t4897 n7683 n4898 R=2.643e+00 
R7682t7182 n7683 n7183 R=2.476e+01 
R7682t5292 n7683 n5293 R=1.509e+01 
R7683t2451 n7684 n2452 R=2.173e+00 
R7683t6976 n7684 n6977 R=4.830e+01 
R7683t5072 n7684 n5073 R=1.411e+01 
R7683t1576 n7684 n1577 R=6.639e+00 
R7683t6424 n7684 n6425 R=8.862e+01 
R7684t1959 n7685 n1960 R=2.816e+00 
R7684t3425 n7685 n3426 R=7.687e+00 
R7684t1001 n7685 n1002 R=7.917e+01 
R7685t1861 n7686 n1862 R=2.341e+01 
R7685t5155 n7686 n5156 R=4.156e+00 
R7685t2644 n7686 n2645 R=1.444e+01 
R7685t4952 n7686 n4953 R=1.396e+01 
R7685t5736 n7686 n5737 R=2.123e+00 
R7686t919 n7687 n920 R=4.733e+00 
R7686t3055 n7687 n3056 R=8.355e+00 
R7686t3098 n7687 n3099 R=3.392e+00 
R7686t537 n7687 n538 R=1.641e+01 
R7686t861 n7687 n862 R=5.088e+00 
R7686t1557 n7687 n1558 R=1.285e+02 
R7687t2962 n7688 n2963 R=1.645e+01 
R7687t6562 n7688 n6563 R=7.441e+00 
R7688t4877 n7689 n4878 R=1.006e+01 
R7688t7225 n7689 n7226 R=4.895e+00 
R7688t207 n7689 n208 R=6.356e+00 
R7688t1598 n7689 n1599 R=2.916e+00 
R7688t1991 n7689 n1992 R=3.310e+01 
R7689t4726 n7690 n4727 R=5.422e+00 
R7689t2862 n7690 n2863 R=2.112e+01 
R7690t3649 n7691 n3650 R=9.615e+00 
R7690t4952 n7691 n4953 R=5.799e+00 
R7691t435 n7692 n436 R=9.984e+00 
R7691t6533 n7692 n6534 R=3.964e+00 
R7691t5022 n7692 n5023 R=1.963e+02 
R7691t3431 n7692 n3432 R=1.076e+01 
R7691t2587 n7692 n2588 R=2.597e+00 
R7691t1634 n7692 n1635 R=1.629e+02 
R7691t861 n7692 n862 R=1.272e+01 
R7692t4461 n7693 n4462 R=1.661e+01 
R7692t4895 n7693 n4896 R=3.113e+01 
R7692t292 n7693 n293 R=4.535e+00 
R7692t904 n7693 n905 R=4.988e+00 
R7692t116 n7693 n117 R=2.963e+00 
R7693t4234 n7694 n4235 R=8.464e+01 
R7693t6648 n7694 n6649 R=3.472e+00 
R7693t5817 n7694 n5818 R=5.339e+00 
R7694t2706 n7695 n2707 R=1.392e+01 
R7694t3653 n7695 n3654 R=4.924e+00 
R7694t1569 n7695 n1570 R=7.730e+00 
R7694t1305 n7695 n1306 R=2.852e+00 
R7694t6663 n7695 n6664 R=1.410e+02 
R7695t684 n7696 n685 R=6.990e+00 
R7695t6530 n7696 n6531 R=7.820e+01 
R7695t6579 n7696 n6580 R=6.135e+00 
R7696t1370 n7697 n1371 R=1.382e+01 
R7696t5896 n7697 n5897 R=1.276e+01 
R7696t1035 n7697 n1036 R=5.688e+00 
R7697t3094 n7698 n3095 R=6.469e+00 
R7697t4352 n7698 n4353 R=2.875e+00 
R7697t6811 n7698 n6812 R=1.416e+02 
R7697t2205 n7698 n2206 R=2.939e+00 
R7698t3061 n7699 n3062 R=1.124e+01 
R7698t914 n7699 n915 R=7.788e+00 
R7698t5846 n7699 n5847 R=8.713e+00 
R7698t4867 n7699 n4868 R=4.750e+00 
R7699t1661 n7700 n1662 R=3.656e+00 
R7699t4264 n7700 n4265 R=2.400e+01 
R7699t3848 n7700 n3849 R=3.338e+01 
R7699t3112 n7700 n3113 R=6.669e+00 
R7699t4077 n7700 n4078 R=1.265e+01 
R7699t549 n7700 n550 R=4.774e+00 
R7700t4887 n7701 n4888 R=5.747e+00 
R7700t7090 n7701 n7091 R=2.306e+01 
R7700t2897 n7701 n2898 R=6.865e+00 
R7700t1744 n7701 n1745 R=6.089e+00 
R7700t79 n7701 n80 R=5.146e+00 
R7700t4893 n7701 n4894 R=1.444e+01 
R7701t2463 n7702 n2464 R=5.504e+00 
R7701t2080 n7702 n2081 R=6.609e+01 
R7701t7554 n7702 n7555 R=2.373e+01 
R7701t4657 n7702 n4658 R=3.421e+00 
R7701t6944 n7702 n6945 R=2.960e+02 
R7702t372 n7703 n373 R=3.673e+00 
R7702t5171 n7703 n5172 R=8.016e+02 
R7702t838 n7703 n839 R=1.428e+01 
R7702t3423 n7703 n3424 R=1.102e+02 
R7702t592 n7703 n593 R=5.810e+00 
R7702t318 n7703 n319 R=4.063e+00 
R7703t2867 n7704 n2868 R=8.616e+00 
R7703t6419 n7704 n6420 R=8.992e+00 
R7703t3500 n7704 n3501 R=2.623e+00 
R7703t222 n7704 n223 R=2.004e+01 
R7703t3408 n7704 n3409 R=3.205e+00 
R7704t3141 n7705 n3142 R=3.369e+00 
R7704t6665 n7705 n6666 R=2.484e+01 
R7704t3861 n7705 n3862 R=7.149e+00 
R7704t1574 n7705 n1575 R=2.449e+01 
R7704t4409 n7705 n4410 R=7.998e+00 
R7704t2925 n7705 n2926 R=1.665e+01 
R7705t3193 n7706 n3194 R=3.190e+02 
R7705t5821 n7706 n5822 R=1.973e+00 
R7705t2099 n7706 n2100 R=2.763e+01 
R7705t6566 n7706 n6567 R=2.437e+00 
R7705t7260 n7706 n7261 R=2.750e+01 
R7705t1422 n7706 n1423 R=1.427e+01 
R7706t3253 n7707 n3254 R=4.997e+00 
R7706t7493 n7707 n7494 R=1.044e+01 
R7706t2257 n7707 n2258 R=1.423e+01 
R7706t4386 n7707 n4387 R=2.744e+01 
R7706t5545 n7707 n5546 R=6.347e+00 
R7707t4465 n7708 n4466 R=9.380e+01 
R7707t4997 n7708 n4998 R=3.717e+00 
R7707t7206 n7708 n7207 R=6.316e+00 
R7707t5500 n7708 n5501 R=5.922e+00 
R7707t3546 n7708 n3547 R=4.184e+00 
R7708t4153 n7709 n4154 R=7.153e+00 
R7708t3958 n7709 n3959 R=1.434e+01 
R7708t132 n7709 n133 R=2.689e+01 
R7708t5069 n7709 n5070 R=7.231e+01 
R7708t6272 n7709 n6273 R=4.223e+00 
R7709t5063 n7710 n5064 R=1.535e+01 
R7709t1399 n7710 n1400 R=8.126e+00 
R7709t3089 n7710 n3090 R=9.543e+00 
R7709t6241 n7710 n6242 R=5.244e+00 
R7710t1633 n7711 n1634 R=1.769e+01 
R7710t6250 n7711 n6251 R=5.865e+00 
R7710t3989 n7711 n3990 R=2.399e+01 
R7710t4807 n7711 n1 R=6.005e+01 
R7710t3223 n7711 n1 R=9.164e+00 
R7710t6527 n7711 n6528 R=4.474e+00 
R7710t4601 n7711 n4602 R=3.170e+02 
R7711t4731 n7712 n4732 R=6.137e+02 
R7711t7009 n7712 n7010 R=6.203e+00 
R7711t4816 n7712 n4817 R=6.803e+00 
R7711t823 n7712 n824 R=8.429e+00 
R7711t3865 n7712 n3866 R=7.551e+00 
R7711t7503 n7712 n7504 R=3.126e+00 
R7712t1912 n7713 n1913 R=2.114e+01 
R7712t4032 n7713 n4033 R=3.413e+00 
R7712t5572 n7713 n5573 R=6.892e+01 
R7712t4012 n7713 n4013 R=6.481e+00 
R7712t5463 n7713 n5464 R=5.561e+00 
R7712t4900 n7713 n4901 R=4.808e+01 
R7712t2539 n7713 n2540 R=9.618e+00 
R7713t3751 n7714 n3752 R=3.418e+01 
R7713t949 n7714 n950 R=3.602e+00 
R7713t4676 n7714 n4677 R=5.095e+01 
R7713t2562 n7714 n2563 R=2.028e+00 
R7714t7380 n7715 n7381 R=3.531e+00 
R7714t1622 n7715 n1623 R=7.673e+00 
R7714t1607 n7715 n1608 R=3.172e+00 
R7714t3780 n7715 n3781 R=1.358e+01 
R7715t5149 n7716 n5150 R=1.595e+01 
R7715t2894 n7716 n2895 R=5.098e+00 
R7715t2544 n7716 n2545 R=3.529e+00 
R7716t1910 n7717 n1911 R=1.993e+01 
R7716t4156 n7717 n4157 R=1.564e+01 
R7716t1647 n7717 n1648 R=9.014e+00 
R7716t3051 n7717 n3052 R=1.538e+01 
R7716t2639 n7717 n2640 R=8.231e+00 
R7717t4604 n7718 n4605 R=6.965e+00 
R7717t4645 n7718 n4646 R=1.326e+01 
R7718t5585 n7719 n5586 R=1.900e+01 
R7718t3265 n7719 n3266 R=7.686e+00 
R7718t2917 n7719 n2918 R=2.300e+00 
R7719t1871 n7720 n1872 R=1.966e+01 
R7719t6144 n7720 n6145 R=5.822e+00 
R7719t600 n7720 n601 R=1.253e+01 
R7719t6553 n7720 n6554 R=4.935e+00 
R7719t1405 n7720 n1406 R=1.529e+01 
R7720t3067 n7721 n3068 R=2.372e+00 
R7720t427 n7721 n428 R=3.707e+00 
R7721t969 n7722 n970 R=5.477e+00 
R7721t5296 n7722 n5297 R=1.888e+01 
R7721t7578 n7722 n7579 R=3.018e+01 
R7721t2447 n7722 n2448 R=4.371e+00 
R7722t4195 n7723 n4196 R=9.268e+00 
R7722t7187 n7723 n7188 R=4.464e+01 
R7722t1227 n7723 n1228 R=3.941e+01 
R7722t4363 n7723 n4364 R=8.615e+00 
R7722t1233 n7723 n1234 R=4.017e+00 
R7722t3578 n7723 n3579 R=2.193e+01 
R7722t1961 n7723 n1962 R=3.304e+01 
R7722t2415 n7723 n2416 R=4.012e+00 
R7723t1085 n7724 n1086 R=6.670e+00 
R7723t700 n7724 n701 R=2.257e+01 
R7723t5002 n7724 n5003 R=1.634e+01 
R7723t2555 n7724 n2556 R=3.893e+00 
R7723t6688 n7724 n6689 R=9.363e+00 
R7723t5413 n7724 n5414 R=2.981e+01 
R7724t367 n7725 n368 R=2.470e+01 
R7724t4685 n7725 n4686 R=6.744e+00 
R7724t1551 n7725 n1552 R=2.215e+00 
R7724t2450 n7725 n2451 R=8.779e+00 
R7724t824 n7725 n825 R=4.930e+00 
R7725t5966 n7726 n5967 R=6.027e+00 
R7725t4716 n7726 n4717 R=5.046e+00 
R7725t1908 n7726 n1909 R=1.025e+01 
R7725t415 n7726 n416 R=4.273e+00 
R7726t2379 n7727 n2380 R=1.752e+01 
R7726t5277 n7727 n5278 R=1.118e+01 
R7726t1189 n7727 n1190 R=3.189e+00 
R7726t2448 n7727 n2449 R=3.665e+01 
R7726t7044 n7727 n7045 R=2.452e+01 
R7726t1689 n7727 n1690 R=1.949e+00 
R7727t2277 n7728 n2278 R=4.523e+00 
R7727t893 n7728 n894 R=3.712e+00 
R7728t3384 n7729 n3385 R=3.385e+00 
R7728t4453 n7729 n4454 R=5.690e+00 
R7729t6717 n7730 n6718 R=5.352e+00 
R7729t6796 n7730 n6797 R=2.695e+00 
R7729t7018 n7730 n7019 R=3.178e+00 
R7730t426 n7731 n427 R=9.677e+00 
R7730t4286 n7731 n4287 R=2.345e+00 
R7730t6011 n7731 n6012 R=4.366e+00 
R7730t3957 n7731 n3958 R=2.488e+02 
R7730t7160 n7731 n7161 R=1.171e+01 
R7731t299 n7732 n300 R=1.764e+01 
R7731t1193 n7732 n1194 R=3.100e+02 
R7731t5018 n7732 n5019 R=3.921e+00 
R7731t3388 n7732 n3389 R=9.851e+00 
R7731t221 n7732 n222 R=1.403e+01 
R7731t942 n7732 n943 R=2.751e+01 
R7732t908 n7733 n909 R=9.476e+00 
R7732t4725 n7733 n4726 R=4.248e+00 
R7732t838 n7733 n839 R=3.608e+01 
R7732t5769 n7733 n5770 R=4.530e+00 
R7733t1081 n7734 n1082 R=4.476e+01 
R7733t7468 n7734 n7469 R=4.352e+01 
R7733t1313 n7734 n1314 R=1.515e+01 
R7733t158 n7734 n159 R=3.271e+00 
R7733t4090 n7734 n4091 R=3.155e+01 
R7733t5079 n7734 n5080 R=2.934e+00 
R7733t6852 n7734 n6853 R=2.138e+01 
R7734t1722 n7735 n1723 R=6.077e+01 
R7734t6366 n7735 n6367 R=6.344e+00 
R7734t1671 n7735 n1672 R=1.508e+01 
R7734t2990 n7735 n2991 R=4.108e+00 
R7734t3134 n7735 n3135 R=4.654e+01 
R7735t7547 n7736 n7548 R=2.394e+01 
R7735t594 n7736 n595 R=6.473e+00 
R7735t2030 n7736 n2031 R=1.521e+01 
R7735t7423 n7736 n7424 R=4.665e+01 
R7735t4980 n7736 n4981 R=1.265e+01 
R7735t677 n7736 n678 R=1.849e+02 
R7735t213 n7736 n214 R=8.874e+00 
R7735t6650 n7736 n6651 R=5.656e+01 
R7736t2334 n7737 n2335 R=2.036e+01 
R7736t5314 n7737 n5315 R=8.813e+00 
R7736t3671 n7737 n3672 R=1.051e+01 
R7736t3427 n7737 n3428 R=8.702e+00 
R7736t1857 n7737 n1858 R=3.391e+00 
R7736t6891 n7737 n6892 R=2.468e+01 
R7736t5984 n7737 n5985 R=1.820e+02 
R7736t1814 n7737 n1815 R=1.355e+01 
R7736t1713 n7737 n1714 R=5.001e+02 
R7736t3829 n7737 n3830 R=9.328e+00 
R7737t813 n7738 n814 R=8.495e+00 
R7737t3812 n7738 n3813 R=1.326e+01 
R7737t7204 n7738 n7205 R=8.834e+00 
R7737t2154 n7738 n2155 R=1.254e+01 
R7737t6273 n7738 n6274 R=7.210e+00 
R7738t1455 n7739 n1456 R=2.028e+00 
R7738t6269 n7739 n6270 R=2.961e+01 
R7738t4156 n7739 n4157 R=6.105e+00 
R7738t1647 n7739 n1648 R=3.114e+00 
R7739t2787 n7740 n2788 R=1.436e+01 
R7739t2994 n7740 n2995 R=3.164e+00 
R7739t5382 n7740 n5383 R=1.338e+01 
R7739t825 n7740 n826 R=9.882e+00 
R7740t7478 n7741 n7479 R=4.650e+00 
R7740t7406 n7741 n7407 R=6.933e+00 
R7740t93 n7741 n94 R=1.447e+01 
R7741t6210 n7742 n6211 R=3.430e+00 
R7741t3807 n7742 n3808 R=1.060e+01 
R7741t3813 n7742 n3814 R=6.938e+00 
R7741t1997 n7742 n1998 R=8.689e+00 
R7741t6465 n7742 n6466 R=5.588e+00 
R7742t6680 n7743 n6681 R=1.074e+01 
R7742t5262 n7743 n5263 R=5.956e+01 
R7742t2409 n7743 n2410 R=4.614e+00 
R7742t1956 n7743 n1957 R=1.378e+01 
R7742t7363 n7743 n7364 R=1.173e+01 
R7743t1377 n7744 n1378 R=4.017e+00 
R7743t6734 n7744 n6735 R=7.794e+00 
R7743t2211 n7744 n2212 R=4.433e+01 
R7743t2670 n7744 n2671 R=4.504e+00 
R7743t6407 n7744 n6408 R=1.475e+01 
R7743t5085 n7744 n5086 R=1.939e+01 
R7743t4992 n7744 n4993 R=1.842e+01 
R7743t4367 n7744 n4368 R=3.384e+01 
R7744t2291 n7745 n2292 R=3.704e+00 
R7744t2532 n7745 n2533 R=2.193e+01 
R7744t476 n7745 n477 R=1.120e+01 
R7744t4856 n7745 n4857 R=1.931e+01 
R7744t2145 n7745 n2146 R=6.525e+00 
R7744t709 n7745 n710 R=5.992e+00 
R7744t977 n7745 n978 R=3.148e+01 
R7745t2875 n7746 n2876 R=3.509e+01 
R7745t629 n7746 n630 R=4.619e+00 
R7745t1019 n7746 n1020 R=2.976e+01 
R7745t6575 n7746 n6576 R=2.010e+01 
R7746t4364 n7747 n4365 R=7.889e+00 
R7746t1107 n7747 n1108 R=1.534e+01 
R7746t1527 n7747 n1528 R=1.212e+01 
R7746t6167 n7747 n6168 R=2.526e+02 
R7747t5741 n7748 n5742 R=5.409e+01 
R7747t3468 n7748 n3469 R=1.610e+01 
R7747t1911 n7748 n1912 R=4.095e+01 
R7747t3137 n7748 n3138 R=7.667e+00 
R7748t1651 n7749 n1652 R=2.806e+00 
R7748t6453 n7749 n6454 R=2.300e+01 
R7748t440 n7749 n441 R=2.021e+01 
R7748t7434 n7749 n7435 R=4.132e+00 
R7748t2548 n7749 n2549 R=3.780e+00 
R7748t3361 n7749 n3362 R=1.497e+01 
R7749t1480 n7750 n1481 R=7.104e+01 
R7749t7171 n7750 n7172 R=3.611e+00 
R7749t7494 n7750 n7495 R=2.702e+01 
R7749t1519 n7750 n1520 R=7.190e+00 
R7749t631 n7750 n632 R=7.588e+00 
R7749t5892 n7750 n5893 R=4.596e+00 
R7750t432 n7751 n433 R=3.082e+00 
R7750t4566 n7751 n4567 R=1.327e+01 
R7750t1807 n7751 n1808 R=1.723e+01 
R7750t2737 n7751 n2738 R=8.907e+00 
R7750t4390 n7751 n4391 R=2.354e+00 
R7751t10 n7752 n11 R=1.301e+01 
R7751t6827 n7752 n6828 R=2.674e+00 
R7751t4780 n7752 n4781 R=3.282e+01 
R7751t7002 n7752 n7003 R=9.637e+01 
R7751t5578 n7752 n5579 R=3.176e+00 
R7751t4570 n7752 n4571 R=5.414e+00 
R7752t3138 n7753 n3139 R=1.974e+01 
R7752t2435 n7753 n2436 R=4.445e+00 
R7752t7224 n7753 n7225 R=7.498e+00 
R7752t3369 n7753 n3370 R=8.531e+00 
R7753t1788 n7754 n1789 R=4.129e+02 
R7753t6340 n7754 n6341 R=2.829e+01 
R7753t156 n7754 n157 R=1.600e+00 
R7753t4295 n7754 n4296 R=1.890e+01 
R7754t3725 n7755 n3726 R=1.100e+01 
R7754t658 n7755 n659 R=1.290e+01 
R7754t3896 n7755 n3897 R=8.794e+00 
R7754t5206 n7755 n5207 R=5.711e+00 
R7754t926 n7755 n927 R=5.602e+00 
R7755t2832 n7756 n2833 R=4.185e+00 
R7755t5541 n7756 n5542 R=8.885e+01 
R7755t2775 n7756 n2776 R=3.992e+01 
R7755t1488 n7756 n1489 R=5.154e+01 
R7755t4641 n7756 n4642 R=1.666e+00 
R7755t7384 n7756 n7385 R=1.270e+01 
R7755t4501 n7756 n4502 R=6.216e+00 
R7756t2070 n7757 n2071 R=4.128e+00 
R7756t5006 n7757 n5007 R=1.157e+01 
R7756t2643 n7757 n2644 R=5.201e+00 
R7756t5358 n7757 n5359 R=1.080e+01 
R7757t6761 n7758 n6762 R=1.589e+01 
R7757t7050 n7758 n7051 R=2.968e+01 
R7757t1528 n7758 n1529 R=7.566e+00 
R7757t145 n7758 n146 R=6.312e+00 
R7757t716 n7758 n717 R=1.799e+01 
R7758t331 n7759 n332 R=9.166e+00 
R7758t4610 n7759 n4611 R=5.034e+00 
R7758t657 n7759 n658 R=5.074e+00 
R7758t7101 n7759 n7102 R=1.497e+01 
R7759t5323 n7760 n5324 R=2.603e+01 
R7759t7116 n7760 n7117 R=5.757e+01 
R7759t4323 n7760 n4324 R=1.362e+01 
R7759t905 n7760 n906 R=3.706e+00 
R7759t6404 n7760 n6405 R=8.197e+00 
R7759t512 n7760 n513 R=1.818e+01 
R7759t2311 n7760 n2312 R=1.100e+01 
R7759t664 n7760 n665 R=1.462e+01 
R7760t74 n7761 n75 R=4.253e+01 
R7760t1584 n7761 n1585 R=2.488e+02 
R7760t4694 n7761 n4695 R=9.987e+00 
R7760t3772 n7761 n3773 R=2.101e+01 
R7760t2731 n7761 n2732 R=6.952e+00 
R7760t1586 n7761 n1587 R=1.966e+00 
R7761t621 n7762 n622 R=2.389e+00 
R7761t4463 n7762 n4464 R=1.462e+01 
R7761t3731 n7762 n3732 R=1.535e+01 
R7761t3797 n7762 n3798 R=4.768e+01 
R7761t7177 n7762 n7178 R=7.132e+00 
R7762t2618 n7763 n2619 R=3.625e+00 
R7762t6228 n7763 n6229 R=1.509e+01 
R7762t5257 n7763 n5258 R=1.153e+01 
R7762t7182 n7763 n7183 R=1.142e+01 
R7762t7682 n7763 n7683 R=4.210e+00 
R7762t5292 n7763 n5293 R=8.225e+00 
R7763t1036 n7764 n1037 R=6.255e+00 
R7763t7414 n7764 n7415 R=7.993e+00 
R7763t455 n7764 n456 R=8.495e+00 
R7763t1834 n7764 n1835 R=1.102e+01 
R7763t4908 n7764 n4909 R=2.842e+00 
R7763t3440 n7764 n3441 R=2.732e+01 
R7764t7083 n7765 n7084 R=2.051e+01 
R7764t5945 n7765 n5946 R=5.818e+01 
R7764t5427 n7765 n5428 R=2.577e+00 
R7764t7570 n7765 n7571 R=1.333e+01 
R7764t3311 n7765 n3312 R=3.651e+00 
R7764t1788 n7765 n1789 R=7.498e+01 
R7765t7129 n7766 n7130 R=4.026e+00 
R7765t2723 n7766 n2724 R=2.501e+00 
R7767t5717 n7768 n5718 R=4.732e+00 
R7767t35 n7768 n36 R=3.014e+00 
R7767t445 n7768 n446 R=2.261e+00 
R7768t6957 n7769 n6958 R=1.311e+01 
R7768t6782 n7769 n6783 R=4.527e+00 
R7768t4061 n7769 n4062 R=6.658e+00 
R7768t4401 n7769 n4402 R=1.984e+01 
R7768t3154 n7769 n3155 R=8.725e+00 
R7769t6701 n7770 n6702 R=6.574e+00 
R7769t7314 n7770 n7315 R=4.363e+00 
R7769t4410 n7770 n4411 R=8.584e+00 
R7769t2007 n7770 n2008 R=3.433e+00 
R7770t6670 n7771 n6671 R=4.334e+00 
R7770t5971 n7771 n5972 R=5.391e+00 
R7770t6920 n7771 n6921 R=2.759e+02 
R7770t3074 n7771 n3075 R=1.438e+00 
R7770t2678 n7771 n2679 R=6.519e+01 
R7771t1881 n7772 n1882 R=3.549e+00 
R7771t3353 n7772 n3354 R=6.232e+00 
R7771t1368 n7772 n1369 R=3.600e+00 
R7771t6624 n7772 n6625 R=4.467e+01 
R7772t896 n7773 n897 R=3.340e+00 
R7772t2750 n7773 n2751 R=2.080e+00 
R7772t7503 n7773 n7504 R=4.714e+00 
R7773t1539 n7774 n1540 R=9.290e+00 
R7773t5475 n7774 n5476 R=7.512e+00 
R7773t662 n7774 n663 R=5.089e+00 
R7773t2785 n7774 n2786 R=3.252e+00 
R7774t3302 n7775 n3303 R=4.455e+00 
R7774t4249 n7775 n4250 R=1.644e+01 
R7774t5926 n7775 n5927 R=5.756e+00 
R7774t3584 n7775 n3585 R=1.471e+01 
R7774t354 n7775 n355 R=9.666e+00 
R7774t5866 n7775 n5867 R=1.476e+01 
R7774t6637 n7775 n6638 R=2.543e+01 
R7775t8 n7776 n9 R=2.958e+01 
R7775t5324 n7776 n5325 R=9.528e+00 
R7775t4848 n7776 n4849 R=8.834e+00 
R7775t4951 n7776 n4952 R=5.508e+00 
R7775t7538 n7776 n7539 R=8.419e+00 
R7776t1797 n7777 n1798 R=4.296e+02 
R7776t3891 n7777 n3892 R=2.154e+01 
R7776t4529 n7777 n4530 R=8.625e+00 
R7776t6868 n7777 n6869 R=9.496e+00 
R7776t2633 n7777 n2634 R=1.100e+01 
R7776t631 n7777 n632 R=1.041e+01 
R7777t2550 n7778 n2551 R=6.592e+00 
R7777t5968 n7778 n5969 R=7.899e+02 
R7777t2510 n7778 n2511 R=2.494e+01 
R7777t975 n7778 n976 R=1.169e+01 
R7777t889 n7778 n890 R=7.324e+00 
R7777t7439 n7778 n7440 R=8.263e+00 
R7777t677 n7778 n678 R=1.147e+01 
R7778t3992 n7779 n3993 R=1.445e+01 
R7778t1733 n7779 n1734 R=1.252e+01 
R7778t1054 n7779 n1055 R=9.704e+00 
R7778t3147 n7779 n3148 R=9.085e+00 
R7779t911 n7780 n912 R=7.266e+00 
R7779t6175 n7780 n6176 R=9.878e+00 
R7779t1796 n7780 n1797 R=6.442e+01 
R7779t6014 n7780 n6015 R=4.919e+00 
R7779t2385 n7780 n2386 R=2.277e+01 
R7779t880 n7780 n881 R=1.601e+01 
R7780t3707 n7781 n3708 R=2.257e+01 
R7780t4700 n7781 n4701 R=2.932e+00 
R7780t6987 n7781 n6988 R=8.236e+00 
R7780t1423 n7781 n1424 R=1.478e+01 
R7780t5596 n7781 n5597 R=3.600e+00 
R7781t4695 n7782 n4696 R=5.926e+00 
R7781t2317 n7782 n2318 R=1.742e+01 
R7781t6752 n7782 n6753 R=6.126e+00 
R7781t1978 n7782 n1979 R=5.564e+01 
R7782t6924 n7783 n6925 R=9.488e+00 
R7782t5014 n7783 n5015 R=3.549e+01 
R7782t1486 n7783 n1487 R=1.064e+01 
R7782t3248 n7783 n3249 R=4.001e+00 
R7782t5914 n7783 n5915 R=1.135e+01 
R7783t3773 n7784 n3774 R=5.916e+00 
R7783t1973 n7784 n1974 R=9.906e+00 
R7783t6359 n7784 n6360 R=3.237e+00 
R7784t598 n7785 n599 R=4.586e+01 
R7784t2640 n7785 n2641 R=6.712e+00 
R7784t4743 n7785 n4744 R=2.020e+01 
R7784t635 n7785 n636 R=1.336e+01 
R7785t360 n7786 n361 R=6.062e+00 
R7785t185 n7786 n186 R=1.141e+01 
R7785t4999 n7786 n5000 R=2.451e+01 
R7785t6845 n7786 n6846 R=1.018e+01 
R7785t302 n7786 n303 R=5.374e+00 
R7785t6567 n7786 n6568 R=9.936e+00 
R7786t6412 n7787 n6413 R=5.400e+01 
R7786t9 n7787 n10 R=5.048e+01 
R7786t7561 n7787 n7562 R=7.259e+00 
R7786t1826 n7787 n1827 R=1.906e+01 
R7786t4674 n7787 n4675 R=5.775e+00 
R7786t3424 n7787 n3425 R=4.125e+01 
R7787t355 n7788 n356 R=2.868e+00 
R7787t4423 n7788 n4424 R=1.547e+01 
R7787t4767 n7788 n4768 R=4.264e+00 
R7787t6707 n7788 n6708 R=1.533e+01 
R7787t5146 n7788 n5147 R=1.527e+01 
R7787t4265 n7788 n4266 R=7.696e+00 
R7787t4377 n7788 n4378 R=4.104e+01 
R7788t1862 n7789 n1863 R=1.552e+01 
R7788t3285 n7789 n3286 R=1.171e+01 
R7788t6251 n7789 n6252 R=5.052e+00 
R7788t3491 n7789 n3492 R=2.663e+00 
R7788t7500 n7789 n7501 R=1.755e+01 
R7788t1263 n7789 n1264 R=6.109e+00 
R7789t513 n7790 n514 R=5.156e+00 
R7789t6631 n7790 n6632 R=1.461e+01 
R7789t2348 n7790 n2349 R=3.522e+00 
R7790t1216 n7791 n1217 R=5.462e+00 
R7790t6300 n7791 n6301 R=3.990e+00 
R7790t4275 n7791 n4276 R=1.203e+01 
R7790t462 n7791 n463 R=6.614e+00 
R7791t7414 n7792 n7415 R=2.845e+00 
R7791t7763 n7792 n7764 R=5.625e+01 
R7791t2313 n7792 n2314 R=7.904e+01 
R7791t3140 n7792 n3141 R=4.839e+00 
R7791t455 n7792 n456 R=3.533e+00 
R7792t1065 n7793 n1066 R=1.432e+01 
R7792t4902 n7793 n4903 R=2.741e+01 
R7792t2862 n7793 n2863 R=5.397e+00 
R7792t7689 n7793 n7690 R=7.319e+00 
R7792t405 n7793 n406 R=1.763e+01 
R7793t1403 n7794 n1404 R=3.526e+01 
R7793t4227 n7794 n4228 R=2.172e+01 
R7793t5225 n7794 n5226 R=2.284e+00 
R7794t88 n7795 n89 R=3.858e+00 
R7794t3897 n7795 n3898 R=2.939e+00 
R7794t5897 n7795 n5898 R=1.847e+00 
R7795t7059 n7796 n7060 R=3.128e+00 
R7795t481 n7796 n482 R=5.544e+00 
R7795t7444 n7796 n7445 R=2.165e+01 
R7795t5808 n7796 n5809 R=3.672e+01 
R7796t4605 n7797 n4606 R=9.879e+01 
R7796t7517 n7797 n7518 R=1.029e+01 
R7796t3712 n7797 n3713 R=3.145e+00 
R7796t1949 n7797 n1950 R=5.213e+01 
R7796t7275 n7797 n7276 R=2.615e+00 
R7796t7337 n7797 n7338 R=8.513e+00 
R7797t1367 n7798 n1368 R=5.395e+00 
R7797t6430 n7798 n6431 R=8.879e+00 
R7797t5841 n7798 n5842 R=1.452e+01 
R7797t831 n7798 n832 R=5.767e+00 
R7797t7318 n7798 n7319 R=5.144e+00 
R7797t4235 n7798 n4236 R=1.208e+01 
R7798t5344 n7799 n5345 R=1.232e+01 
R7798t1937 n7799 n1938 R=1.582e+01 
R7798t2035 n7799 n2036 R=8.791e+00 
R7798t7057 n7799 n7058 R=3.057e+01 
R7798t3338 n7799 n3339 R=6.547e+00 
R7799t2876 n7800 n2877 R=3.367e+00 
R7799t3697 n7800 n3698 R=3.388e+00 
R7799t7197 n7800 n7198 R=3.765e+01 
R7800t3392 n7801 n3393 R=8.636e+00 
R7800t4513 n7801 n4514 R=9.154e+00 
R7800t24 n7801 n25 R=6.612e+01 
R7800t4190 n7801 n4191 R=5.079e+00 
R7800t1566 n7801 n1567 R=1.605e+01 
R7801t6761 n7802 n6762 R=2.488e+00 
R7801t7757 n7802 n7758 R=1.384e+01 
R7801t4761 n7802 n4762 R=5.142e+02 
R7801t5090 n7802 n5091 R=6.307e+00 
R7802t3396 n7803 n3397 R=7.603e+00 
R7802t3892 n7803 n3893 R=2.531e+01 
R7802t6746 n7803 n6747 R=2.762e+00 
R7802t6993 n7803 n6994 R=2.912e+00 
R7803t3516 n7804 n3517 R=6.256e+00 
R7803t4520 n7804 n4521 R=3.686e+00 
R7803t4006 n7804 n4007 R=2.809e+01 
R7803t4699 n7804 n4700 R=1.874e+00 
R7804t889 n7805 n890 R=6.039e+00 
R7804t7132 n7805 n7133 R=3.949e+01 
R7804t6422 n7805 n6423 R=1.579e+01 
R7804t4289 n7805 n4290 R=8.682e+00 
R7804t2718 n7805 n2719 R=3.660e+00 
R7804t7439 n7805 n7440 R=5.589e+01 
R7804t7777 n7805 n7778 R=6.937e+00 
R7805t3694 n7806 n3695 R=1.168e+01 
R7805t4688 n7806 n4689 R=5.844e+01 
R7805t5681 n7806 n5682 R=4.411e+01 
R7805t6395 n7806 n6396 R=7.129e+00 
R7805t3250 n7806 n3251 R=1.291e+01 
R7805t7337 n7806 n7338 R=5.982e+00 
R7805t7796 n7806 n7797 R=1.489e+01 
R7805t7275 n7806 n7276 R=1.442e+01 
R7805t1010 n7806 n1011 R=1.313e+01 
R7807t3720 n7808 n3721 R=4.903e+00 
R7807t5390 n7808 n5391 R=9.320e+00 
R7807t646 n7808 n647 R=6.038e+00 
R7807t7008 n7808 n7009 R=4.254e+00 
R7807t5819 n7808 n5820 R=2.346e+02 
R7808t10 n7809 n11 R=6.852e+00 
R7808t489 n7809 n490 R=3.682e+00 
R7808t6827 n7809 n6828 R=1.828e+02 
R7808t92 n7809 n93 R=3.940e+00 
R7808t3984 n7809 n3985 R=8.473e+00 
R7809t17 n7810 n18 R=7.202e+00 
R7809t3545 n7810 n3546 R=9.789e+00 
R7809t3583 n7810 n3584 R=4.932e+00 
R7809t6410 n7810 n6411 R=5.094e+00 
R7809t184 n7810 n185 R=2.252e+01 
R7809t884 n7810 n885 R=8.391e+00 
R7810t1292 n7811 n1293 R=1.206e+01 
R7810t5103 n7811 n5104 R=7.941e+00 
R7810t4128 n7811 n4129 R=2.686e+00 
R7810t5498 n7811 n5499 R=1.060e+02 
R7810t6633 n7811 n6634 R=6.221e+01 
R7810t4751 n7811 n4752 R=1.019e+01 
R7810t7649 n7811 n7650 R=3.581e+00 
R7811t334 n7812 n335 R=1.324e+02 
R7811t365 n7812 n366 R=5.280e+01 
R7811t3169 n7812 n3170 R=5.229e+00 
R7811t7542 n7812 n7543 R=4.478e+00 
R7811t7280 n7812 n7281 R=1.742e+01 
R7811t1605 n7812 n1606 R=2.628e+00 
R7812t7500 n7813 n7501 R=5.877e+00 
R7812t7788 n7813 n7789 R=1.214e+02 
R7812t1263 n7813 n1264 R=7.037e+00 
R7812t3544 n7813 n3545 R=6.293e+00 
R7813t5039 n7814 n5040 R=3.994e+00 
R7813t6150 n7814 n6151 R=8.537e+00 
R7813t4491 n7814 n4492 R=7.678e+00 
R7813t2857 n7814 n2858 R=8.079e+00 
R7814t1159 n7815 n1160 R=3.181e+00 
R7814t6374 n7815 n6375 R=1.793e+01 
R7814t1488 n7815 n1489 R=8.505e+00 
R7814t4641 n7815 n4642 R=1.470e+00 
R7815t825 n7816 n826 R=1.440e+01 
R7815t5777 n7816 n5778 R=5.842e+00 
R7816t3077 n7817 n3078 R=1.836e+01 
R7816t5554 n7817 n5555 R=3.071e+00 
R7816t7475 n7817 n7476 R=7.873e+00 
R7816t6539 n7817 n6540 R=5.244e+00 
R7816t4354 n7817 n4355 R=1.453e+01 
R7817t7459 n7818 n7460 R=2.113e+02 
R7817t4684 n7818 n4685 R=5.590e+00 
R7817t7645 n7818 n7646 R=1.506e+01 
R7817t5505 n7818 n5506 R=5.066e+00 
R7818t6235 n7819 n6236 R=2.590e+01 
R7818t6910 n7819 n6911 R=5.735e+00 
R7818t6501 n7819 n6502 R=1.515e+01 
R7818t5343 n7819 n5344 R=6.366e+00 
R7819t5277 n7820 n5278 R=5.542e+00 
R7819t5832 n7820 n5833 R=2.986e+01 
R7819t2379 n7820 n2380 R=1.893e+01 
R7819t395 n7820 n396 R=1.373e+01 
R7819t1011 n7820 n1012 R=9.863e+00 
R7819t5581 n7820 n5582 R=1.301e+01 
R7819t3101 n7820 n3102 R=5.209e+02 
R7819t7205 n7820 n7206 R=3.318e+00 
R7820t4949 n7821 n4950 R=6.894e+00 
R7820t5940 n7821 n5941 R=5.966e+00 
R7820t4095 n7821 n4096 R=1.867e+01 
R7820t2676 n7821 n2677 R=8.476e+00 
R7820t2223 n7821 n2224 R=4.901e+00 
R7821t211 n7822 n212 R=3.710e+00 
R7821t2818 n7822 n2819 R=3.094e+01 
R7821t1509 n7822 n1510 R=5.151e+00 
R7821t4785 n7822 n4786 R=6.130e+00 
R7822t862 n7823 n863 R=4.288e+00 
R7822t4882 n7823 n4883 R=4.749e+00 
R7822t7013 n7823 n7014 R=5.346e+00 
R7822t2324 n7823 n2325 R=5.718e+00 
R7823t1838 n7824 n1839 R=4.406e+00 
R7823t6591 n7824 n6592 R=3.678e+01 
R7823t7288 n7824 n7289 R=2.664e+00 
R7823t2559 n7824 n2560 R=2.691e+00 
R7824t3932 n7825 n3933 R=1.085e+01 
R7824t6001 n7825 n6002 R=3.351e+00 
R7824t3079 n7825 n3080 R=6.712e+00 
R7824t1025 n7825 n1026 R=4.944e+00 
R7825t3455 n1 n3456 R=9.543e+00 
R7826t5709 n7827 n5710 R=9.474e+00 
R7826t6298 n7827 n6299 R=1.086e+01 
R7826t4713 n7827 n4714 R=5.465e+00 
R7826t2023 n7827 n2024 R=3.009e+01 
R7827t122 n7828 n123 R=4.236e+01 
R7827t2839 n7828 n2840 R=1.851e+01 
R7827t6696 n7828 n6697 R=3.437e+00 
R7827t3794 n7828 n3795 R=2.545e+00 
R7828t3021 n7829 n3022 R=3.803e+00 
R7828t7679 n7829 n7680 R=1.328e+02 
R7828t2745 n7829 n2746 R=8.901e+00 
R7828t1302 n7829 n1303 R=2.973e+00 
R7828t2836 n7829 n2837 R=5.279e+00 
R7829t372 n7830 n373 R=1.706e+01 
R7829t838 n7830 n839 R=2.909e+00 
R7829t7732 n7830 n7733 R=6.385e+00 
R7829t4485 n7830 n4486 R=1.405e+01 
R7830t5281 n7831 n5282 R=2.435e+00 
R7830t6723 n7831 n6724 R=1.052e+01 
R7830t143 n7831 n144 R=8.476e+00 
R7830t5870 n7831 n5871 R=4.734e+00 
R7830t7427 n7831 n7428 R=5.663e+01 
R7830t5992 n7831 n5993 R=1.856e+01 
R7831t4587 n7832 n4588 R=3.664e+00 
R7831t7048 n7832 n7049 R=2.365e+01 
R7831t2515 n7832 n2516 R=7.157e+00 
R7831t4506 n7832 n4507 R=1.109e+01 
R7831t4466 n7832 n4467 R=8.749e+01 
R7831t6938 n7832 n6939 R=4.117e+00 
R7831t3387 n7832 n3388 R=4.377e+01 
R7832t5115 n7833 n5116 R=3.818e+00 
R7832t1689 n7833 n1690 R=1.123e+01 
R7832t77 n7833 n78 R=7.713e+01 
R7833t1413 n7834 n1414 R=5.446e+00 
R7833t2660 n7834 n2661 R=4.423e+00 
R7834t1798 n7835 n1799 R=3.666e+00 
R7834t3575 n7835 n3576 R=2.262e+00 
R7834t4700 n7835 n4701 R=1.401e+02 
R7834t6572 n7835 n6573 R=4.631e+00 
R7835t1381 n7836 n1382 R=1.519e+01 
R7835t4974 n7836 n4975 R=4.548e+00 
R7835t4992 n7836 n4993 R=2.905e+00 
R7835t7616 n7836 n7617 R=4.162e+01 
R7835t6309 n7836 n6310 R=1.056e+01 
R7836t74 n7837 n75 R=1.246e+01 
R7836t4694 n7837 n4695 R=7.905e+00 
R7836t4433 n7837 n4434 R=1.390e+01 
R7836t6226 n7837 n6227 R=2.838e+00 
R7836t2692 n7837 n2693 R=1.005e+01 
R7836t6602 n7837 n6603 R=6.858e+00 
R7837t1826 n7838 n1827 R=2.976e+00 
R7837t2437 n7838 n2438 R=4.902e+01 
R7837t4742 n7838 n4743 R=1.302e+01 
R7837t5351 n7838 n5352 R=5.274e+00 
R7838t3928 n7839 n3929 R=1.882e+00 
R7838t5524 n7839 n5525 R=1.076e+01 
R7838t1375 n7839 n1376 R=1.317e+01 
R7839t2050 n7840 n2051 R=1.998e+01 
R7839t6426 n7840 n6427 R=1.431e+01 
R7839t1554 n7840 n1555 R=2.337e+01 
R7839t5211 n7840 n5212 R=3.377e+00 
R7839t3988 n7840 n3989 R=2.112e+01 
R7839t2032 n7840 n2033 R=1.397e+01 
R7839t6488 n7840 n6489 R=1.171e+01 
R7839t6452 n7840 n6453 R=1.285e+01 
R7839t149 n7840 n150 R=1.751e+01 
R7840t1726 n7841 n1727 R=2.768e+00 
R7840t4364 n7841 n4365 R=1.079e+01 
R7840t7746 n7841 n7747 R=4.757e+00 
R7840t2590 n7841 n2591 R=1.323e+01 
R7840t187 n7841 n188 R=1.978e+01 
R7840t7240 n7841 n7241 R=7.025e+01 
R7841t6194 n7842 n6195 R=3.076e+01 
R7841t1868 n7842 n1869 R=6.797e+00 
R7841t808 n7842 n809 R=7.318e+00 
R7842t55 n7843 n56 R=8.452e+00 
R7842t2453 n7843 n2454 R=5.591e+00 
R7842t6195 n7843 n6196 R=4.201e+00 
R7842t3573 n7843 n3574 R=6.124e+02 
R7843t4531 n7844 n4532 R=4.329e+00 
R7843t5704 n7844 n5705 R=3.449e+01 
R7843t2518 n7844 n2519 R=1.192e+01 
R7844t3 n7845 n4 R=4.724e+00 
R7844t3552 n7845 n3553 R=4.322e+01 
R7844t1383 n7845 n1384 R=2.906e+00 
R7845t6336 n7846 n6337 R=5.153e+00 
R7845t7333 n7846 n7334 R=6.033e+00 
R7845t1620 n7846 n1621 R=5.942e+00 
R7845t6764 n7846 n6765 R=1.390e+01 
R7846t4897 n7847 n4898 R=8.572e+01 
R7846t7682 n7847 n7683 R=5.261e+00 
R7846t5292 n7847 n5293 R=1.760e+01 
R7846t2904 n7847 n2905 R=6.705e+00 
R7847t7478 n7848 n7479 R=6.665e+01 
R7847t7740 n7848 n7741 R=1.540e+01 
R7847t7406 n7848 n7407 R=7.804e+00 
R7847t222 n7848 n223 R=3.052e+00 
R7847t3469 n7848 n3470 R=5.472e+00 
R7848t6017 n7849 n6018 R=1.103e+02 
R7848t6200 n7849 n6201 R=8.816e+00 
R7848t3774 n7849 n3775 R=6.844e+01 
R7848t7638 n7849 n7639 R=5.239e+00 
R7848t7673 n7849 n7674 R=4.528e+00 
R7848t7562 n7849 n7563 R=7.077e+00 
R7848t3878 n7849 n3879 R=5.914e+00 
R7849t1743 n7850 n1744 R=4.260e+00 
R7849t1335 n7850 n1336 R=4.326e+01 
R7849t4399 n7850 n4400 R=6.018e+00 
R7849t1293 n7850 n1294 R=8.553e+00 
R7850t3987 n7851 n3988 R=1.390e+00 
R7850t2608 n7851 n2609 R=2.613e+00 
R7850t1761 n7851 n1762 R=4.237e+01 
R7851t648 n7852 n649 R=3.909e+00 
R7851t5586 n7852 n5587 R=1.294e+01 
R7851t913 n7852 n914 R=4.092e+02 
R7851t3937 n7852 n3938 R=7.836e+01 
R7851t2797 n7852 n2798 R=7.856e+00 
R7851t5606 n7852 n5607 R=3.836e+00 
R7851t787 n7852 n788 R=9.618e+00 
R7852t5618 n7853 n5619 R=1.668e+02 
R7852t1656 n7853 n1657 R=2.202e+01 
R7852t4325 n7853 n4326 R=7.741e+02 
R7852t7488 n7853 n7489 R=5.758e+01 
R7852t2743 n7853 n2744 R=3.114e+01 
R7852t5129 n7853 n5130 R=2.210e+00 
R7853t4094 n7854 n4095 R=5.707e+00 
R7853t5915 n7854 n5916 R=1.803e+01 
R7853t2719 n7854 n2720 R=4.790e+00 
R7853t3932 n7854 n3933 R=4.219e+00 
R7853t7824 n7854 n7825 R=9.760e+00 
R7853t1025 n7854 n1026 R=2.140e+01 
R7854t374 n7855 n375 R=3.185e+00 
R7854t6818 n7855 n6819 R=8.669e+01 
R7854t2490 n7855 n2491 R=6.558e+00 
R7854t7447 n7855 n7448 R=5.998e+01 
R7854t5468 n7855 n5469 R=8.009e+00 
R7855t7216 n7856 n7217 R=6.750e+00 
R7855t472 n7856 n473 R=6.105e+00 
R7855t2280 n7856 n2281 R=1.433e+01 
R7855t6255 n7856 n6256 R=4.677e+00 
R7856t2112 n7857 n2113 R=7.517e+00 
R7856t6115 n7857 n6116 R=2.750e+00 
R7856t712 n7857 n713 R=3.092e+00 
R7856t3991 n7857 n3992 R=1.002e+01 
R7857t2908 n7858 n2909 R=6.468e+00 
R7857t4727 n7858 n4728 R=1.725e+01 
R7857t4784 n7858 n4785 R=2.309e+00 
R7857t2782 n7858 n2783 R=2.405e+02 
R7857t4439 n7858 n4440 R=1.267e+01 
R7857t1197 n7858 n1198 R=6.524e+01 
R7857t6516 n7858 n6517 R=8.609e+00 
R7858t423 n7859 n424 R=1.806e+01 
R7858t6839 n7859 n6840 R=3.333e+00 
R7858t1441 n7859 n1442 R=6.186e+00 
R7858t4194 n7859 n4195 R=1.957e+01 
R7858t5872 n7859 n5873 R=2.310e+00 
R7859t6169 n7860 n6170 R=1.955e+01 
R7859t6639 n7860 n6640 R=7.645e+00 
R7859t4153 n7860 n4154 R=1.068e+01 
R7859t7708 n7860 n7709 R=5.949e+00 
R7859t2361 n7860 n2362 R=5.253e+00 
R7860t2084 n7861 n2085 R=5.251e+00 
R7860t7395 n7861 n7396 R=2.483e+00 
R7860t3229 n7861 n3230 R=4.326e+00 
R7861t5966 n7862 n5967 R=8.395e+01 
R7861t7297 n7862 n7298 R=2.258e+00 
R7861t4230 n7862 n4231 R=9.190e+00 
R7861t6290 n7862 n6291 R=3.403e+00 
R7861t4716 n7862 n4717 R=5.771e+00 
R7861t7725 n7862 n7726 R=5.770e+01 
R7862t3196 n7863 n3197 R=5.958e+00 
R7862t112 n7863 n113 R=1.515e+01 
R7862t3324 n7863 n3325 R=4.907e+00 
R7862t5389 n7863 n5390 R=7.069e+00 
R7863t2818 n7864 n2819 R=9.867e+00 
R7863t7821 n7864 n7822 R=3.177e+00 
R7863t1947 n7864 n1948 R=2.445e+01 
R7863t7454 n7864 n7455 R=1.259e+01 
R7863t4785 n7864 n4786 R=5.783e+00 
R7864t916 n7865 n917 R=5.354e+00 
R7864t1283 n7865 n1284 R=4.624e+01 
R7864t2552 n7865 n2553 R=6.823e+00 
R7864t971 n7865 n972 R=2.773e+00 
R7864t2592 n7865 n2593 R=3.050e+00 
R7865t745 n7866 n746 R=1.764e+02 
R7865t6916 n7866 n6917 R=4.898e+01 
R7865t4979 n7866 n4980 R=1.050e+01 
R7865t5783 n7866 n5784 R=2.369e+00 
R7865t6408 n7866 n6409 R=1.924e+01 
R7866t2677 n7867 n2678 R=7.498e+00 
R7866t1856 n7867 n1857 R=4.033e+01 
R7866t6269 n7867 n6270 R=3.653e+00 
R7867t2758 n7868 n2759 R=3.441e+01 
R7867t1196 n7868 n1197 R=1.931e+01 
R7867t2771 n7868 n2772 R=7.486e+00 
R7867t4853 n7868 n4854 R=4.117e+00 
R7867t2304 n7868 n2305 R=1.482e+01 
R7868t1098 n7869 n1099 R=1.055e+02 
R7868t5867 n7869 n5868 R=6.718e+00 
R7868t5553 n7869 n5554 R=2.481e+01 
R7868t2355 n7869 n2356 R=1.955e+01 
R7868t391 n7869 n392 R=4.465e+00 
R7869t3817 n7870 n3818 R=5.821e+00 
R7869t6750 n7870 n6751 R=2.325e+02 
R7869t2277 n7870 n2278 R=2.149e+01 
R7869t7727 n7870 n7728 R=1.321e+01 
R7869t893 n7870 n894 R=1.120e+01 
R7869t5448 n7870 n5449 R=2.534e+01 
R7869t2097 n7870 n2098 R=8.124e+00 
R7869t223 n7870 n224 R=3.435e+00 
R7870t4553 n7871 n4554 R=6.569e+00 
R7870t7262 n7871 n7263 R=1.072e+01 
R7870t1408 n7871 n1409 R=1.597e+01 
R7870t3723 n7871 n3724 R=2.629e+02 
R7870t3668 n7871 n3669 R=3.105e+00 
R7871t6475 n7872 n6476 R=1.365e+02 
R7871t6889 n7872 n6890 R=1.301e+01 
R7871t4026 n7872 n4027 R=4.745e+01 
R7871t4686 n7872 n4687 R=3.949e+01 
R7871t4844 n7872 n4845 R=2.935e+00 
R7872t5207 n7873 n5208 R=3.465e+00 
R7872t6363 n7873 n6364 R=5.688e+00 
R7872t182 n7873 n183 R=2.004e+01 
R7872t554 n7873 n555 R=4.664e+00 
R7873t7624 n7874 n7625 R=1.976e+01 
R7873t6484 n7874 n6485 R=3.525e+01 
R7873t1249 n7874 n1250 R=2.238e+00 
R7873t440 n7874 n441 R=7.867e+00 
R7874t1696 n7875 n1697 R=1.471e+01 
R7874t3102 n7875 n3103 R=6.324e+00 
R7874t1047 n7875 n1048 R=1.112e+02 
R7875t2132 n7876 n2133 R=3.194e+01 
R7875t7178 n7876 n7179 R=5.946e+00 
R7875t5296 n7876 n5297 R=4.990e+00 
R7875t7721 n7876 n7722 R=4.302e+00 
R7875t7578 n7876 n7579 R=5.451e+00 
R7876t1427 n7877 n1428 R=3.497e+00 
R7876t4556 n7877 n4557 R=5.680e+00 
R7876t4695 n7877 n4696 R=4.156e+00 
R7876t6928 n7877 n6929 R=6.362e+00 
R7877t4586 n7878 n4587 R=7.460e+00 
R7877t1935 n7878 n1936 R=1.049e+01 
R7877t1381 n7878 n1382 R=4.009e+00 
R7877t3737 n7878 n3738 R=1.252e+01 
R7877t1637 n7878 n1638 R=7.328e+01 
R7877t1774 n7878 n1775 R=5.615e+00 
R7878t5680 n7879 n5681 R=3.834e+01 
R7878t6240 n7879 n6241 R=5.233e+00 
R7878t3081 n7879 n3082 R=2.964e+00 
R7878t4756 n7879 n4757 R=8.406e+00 
R7879t3507 n7880 n3508 R=5.566e+01 
R7879t6614 n7880 n6615 R=2.629e+01 
R7879t1533 n7880 n1534 R=3.253e+00 
R7879t237 n7880 n238 R=3.586e+01 
R7880t1761 n7881 n1762 R=1.112e+02 
R7880t7600 n7881 n7601 R=6.975e+01 
R7880t6953 n7881 n6954 R=3.557e+00 
R7880t7336 n7881 n7337 R=2.930e+00 
R7881t4761 n7882 n4762 R=1.128e+01 
R7881t7801 n7882 n7802 R=2.606e+00 
R7881t7757 n7882 n7758 R=1.201e+01 
R7881t7050 n7882 n7051 R=1.409e+01 
R7881t4001 n7882 n4002 R=3.072e+01 
R7881t3453 n7882 n3454 R=4.716e+00 
R7882t5585 n7883 n5586 R=3.541e+00 
R7882t7718 n7883 n7719 R=3.180e+01 
R7882t2922 n7883 n2923 R=1.028e+01 
R7883t2048 n7884 n2049 R=1.426e+01 
R7883t2579 n7884 n2580 R=2.701e+01 
R7883t2268 n7884 n2269 R=3.895e+00 
R7883t3961 n7884 n3962 R=7.831e+00 
R7884t378 n7885 n379 R=1.931e+01 
R7884t4896 n7885 n4897 R=1.405e+01 
R7884t1424 n7885 n1425 R=8.316e+00 
R7884t5668 n7885 n5669 R=5.966e+00 
R7884t1299 n7885 n1300 R=5.261e+00 
R7885t4546 n7886 n4547 R=1.395e+00 
R7885t3217 n7886 n3218 R=2.725e+00 
R7886t3105 n7887 n3106 R=8.482e+00 
R7886t6392 n7887 n6393 R=3.984e+00 
R7886t3959 n7887 n3960 R=1.078e+02 
R7886t6855 n7887 n6856 R=7.353e+00 
R7886t1149 n7887 n1150 R=5.609e+00 
R7886t845 n7887 n846 R=1.609e+01 
R7887t244 n7888 n245 R=5.685e+00 
R7887t1060 n7888 n1061 R=4.839e+00 
R7887t2510 n7888 n2511 R=3.198e+01 
R7887t6339 n7888 n6340 R=4.972e+00 
R7887t6279 n7888 n6280 R=1.288e+01 
R7887t6788 n7888 n6789 R=7.518e+00 
R7888t497 n7889 n498 R=1.428e+01 
R7888t6692 n7889 n6693 R=2.357e+00 
R7888t3916 n7889 n3917 R=4.168e+01 
R7888t1847 n7889 n1848 R=2.787e+00 
R7888t4640 n7889 n4641 R=6.032e+00 
R7889t3548 n7890 n3549 R=1.378e+01 
R7889t4190 n7890 n4191 R=3.553e+01 
R7889t115 n7890 n116 R=8.255e+00 
R7889t5019 n7890 n5020 R=3.382e+00 
R7889t5459 n7890 n5460 R=1.715e+01 
R7890t1448 n7891 n1449 R=1.331e+01 
R7890t6456 n7891 n6457 R=8.537e+00 
R7890t3136 n7891 n3137 R=4.783e+00 
R7891t992 n7892 n993 R=3.280e+01 
R7891t1018 n7892 n1019 R=4.160e+00 
R7891t5387 n7892 n5388 R=3.475e+00 
R7891t5476 n7892 n5477 R=4.009e+00 
R7892t5885 n7893 n5886 R=2.638e+01 
R7892t5960 n7893 n5961 R=9.971e+00 
R7892t1315 n7893 n1316 R=8.840e+00 
R7892t4396 n7893 n4397 R=3.240e+00 
R7893t7227 n7894 n7228 R=1.264e+01 
R7893t2657 n7894 n2658 R=3.711e+00 
R7893t6201 n7894 n6202 R=3.711e+00 
R7893t6179 n7894 n6180 R=2.333e+01 
R7893t525 n7894 n526 R=1.038e+01 
R7894t2281 n7895 n2282 R=3.773e+01 
R7894t4434 n7895 n4435 R=6.841e+00 
R7894t4382 n7895 n4383 R=4.495e+00 
R7894t5632 n7895 n5633 R=6.028e+00 
R7894t500 n7895 n501 R=1.369e+01 
R7894t5521 n7895 n5522 R=7.808e+01 
R7894t5559 n7895 n5560 R=1.860e+01 
R7895t5168 n7896 n5169 R=3.085e+00 
R7895t4324 n7896 n4325 R=1.642e+01 
R7895t6884 n7896 n6885 R=5.293e+00 
R7896t4316 n7897 n4317 R=1.498e+01 
R7896t7329 n7897 n7330 R=3.780e+00 
R7896t4391 n7897 n4392 R=6.397e+00 
R7896t2962 n7897 n2963 R=2.357e+01 
R7896t7687 n7897 n7688 R=5.744e+00 
R7897t3061 n7898 n3062 R=1.064e+01 
R7897t6140 n7898 n6141 R=5.808e+00 
R7897t3766 n7898 n3767 R=7.950e+00 
R7897t5127 n7898 n5128 R=3.820e+00 
R7897t358 n7898 n359 R=5.001e+01 
R7897t764 n7898 n765 R=2.000e+01 
R7898t6122 n7899 n6123 R=1.188e+01 
R7898t6674 n7899 n6675 R=1.291e+01 
R7898t3577 n7899 n3578 R=4.324e+00 
R7898t6083 n7899 n6084 R=7.991e+00 
R7899t4411 n7900 n4412 R=6.518e+01 
R7899t1543 n7900 n1544 R=4.902e+00 
R7899t4760 n7900 n4761 R=3.631e+00 
R7900t978 n7901 n979 R=1.823e+02 
R7900t4037 n7901 n4038 R=7.211e+00 
R7900t3826 n7901 n3827 R=4.262e+00 
R7900t5661 n7901 n5662 R=7.463e+00 
R7900t7085 n7901 n7086 R=5.184e+00 
R7900t2124 n7901 n2125 R=1.751e+01 
R7900t5796 n7901 n5797 R=8.519e+01 
R7901t968 n7902 n969 R=7.740e+00 
R7901t632 n7902 n633 R=3.778e+00 
R7901t4788 n7902 n4789 R=1.598e+02 
R7901t444 n7902 n445 R=2.091e+00 
R7902t2503 n7903 n2504 R=1.465e+03 
R7902t3249 n7903 n3250 R=2.419e+00 
R7902t1061 n7903 n1062 R=9.460e+00 
R7902t4713 n7903 n4714 R=2.165e+00 
R7902t2023 n7903 n2024 R=1.059e+01 
R7903t2382 n7904 n2383 R=2.596e+02 
R7903t5982 n7904 n5983 R=3.991e+00 
R7903t2267 n7904 n2268 R=7.061e+00 
R7903t3493 n7904 n3494 R=9.520e+00 
R7903t3786 n7904 n3787 R=4.492e+00 
R7903t2831 n7904 n2832 R=1.257e+01 
R7904t5639 n7905 n5640 R=5.144e+00 
R7904t5877 n7905 n5878 R=2.674e+01 
R7904t1571 n7905 n1572 R=3.773e+02 
R7904t6538 n7905 n6539 R=3.209e+00 
R7904t5980 n7905 n5981 R=1.429e+01 
R7905t3385 n7906 n3386 R=1.061e+02 
R7905t5332 n7906 n5333 R=3.897e+00 
R7906t3463 n7907 n3464 R=3.101e+00 
R7906t6883 n7907 n6884 R=1.850e+00 
R7906t1051 n7907 n1052 R=1.914e+01 
R7906t5591 n7907 n5592 R=9.783e+00 
R7907t605 n7908 n606 R=2.580e+01 
R7907t3286 n7908 n3287 R=5.743e+00 
R7907t1095 n7908 n1096 R=1.112e+01 
R7907t5148 n7908 n5149 R=8.992e+00 
R7907t2453 n7908 n2454 R=6.080e+01 
R7908t997 n7909 n998 R=2.948e+01 
R7908t6971 n7909 n6972 R=2.361e+00 
R7908t7827 n7909 n7828 R=1.021e+01 
R7908t122 n7909 n123 R=1.584e+01 
R7908t2060 n7909 n2061 R=2.701e+01 
R7909t1762 n7910 n1763 R=2.469e+01 
R7909t7631 n7910 n7632 R=1.579e+01 
R7909t2953 n7910 n2954 R=4.049e+00 
R7909t2667 n7910 n2668 R=4.028e+00 
R7910t3357 n7911 n3358 R=5.954e+00 
R7910t7352 n7911 n7353 R=3.620e+00 
R7910t313 n7911 n314 R=4.977e+01 
R7910t5941 n7911 n5942 R=4.984e+00 
R7910t574 n7911 n575 R=7.033e+00 
R7911t1564 n7912 n1565 R=1.040e+01 
R7911t4027 n7912 n4028 R=1.629e+01 
R7911t7333 n7912 n7334 R=5.580e+00 
R7911t7845 n7912 n7846 R=4.604e+01 
R7911t1620 n7912 n1621 R=1.367e+01 
R7911t7458 n7912 n7459 R=2.609e+00 
R7912t6307 n7913 n6308 R=8.038e+01 
R7912t5921 n7913 n5922 R=6.356e+00 
R7912t1082 n7913 n1083 R=6.058e+00 
R7912t4600 n7913 n4601 R=1.121e+01 
R7913t4290 n7914 n4291 R=1.151e+01 
R7913t5640 n7914 n5641 R=3.878e+00 
R7913t6722 n7914 n6723 R=8.064e+00 
R7914t44 n7915 n45 R=1.363e+01 
R7914t4054 n7915 n4055 R=6.711e+00 
R7914t7141 n7915 n7142 R=1.628e+02 
R7915t6214 n7916 n6215 R=1.744e+01 
R7915t6915 n7916 n6916 R=1.887e+01 
R7915t4719 n7916 n4720 R=6.262e+00 
R7916t4211 n7917 n4212 R=2.701e+00 
R7916t5836 n7917 n5837 R=5.814e+01 
R7916t4513 n7917 n4514 R=1.845e+00 
R7917t6740 n7918 n6741 R=5.250e+00 
R7917t4724 n7918 n4725 R=6.795e+00 
R7917t2468 n7918 n2469 R=3.901e+01 
R7917t2227 n7918 n2228 R=1.548e+01 
R7918t411 n7919 n412 R=4.868e+00 
R7918t7568 n7919 n7569 R=3.230e+00 
R7918t87 n7919 n88 R=1.735e+01 
R7918t3198 n7919 n3199 R=5.041e+00 
R7919t3629 n7920 n3630 R=6.104e+00 
R7919t6374 n7920 n6375 R=4.053e+00 
R7919t1159 n7920 n1160 R=3.692e+00 
R7920t1786 n7921 n1787 R=5.324e+00 
R7920t3101 n7921 n3102 R=3.608e+00 
R7920t5581 n7921 n5582 R=1.339e+01 
R7920t5138 n7921 n5139 R=6.189e+00 
R7921t6694 n7922 n6695 R=1.937e+01 
R7921t7071 n7922 n7072 R=5.537e+00 
R7921t5664 n7922 n5665 R=6.786e+00 
R7921t7373 n7922 n7374 R=4.823e+00 
R7922t5646 n7923 n5647 R=3.572e+00 
R7922t5254 n7923 n5255 R=6.376e+00 
R7922t6803 n7923 n6804 R=3.396e+00 
R7922t1915 n7923 n1916 R=6.587e+00 
R7923t3205 n7924 n3206 R=2.196e+01 
R7923t3316 n7924 n3317 R=2.498e+01 
R7923t5084 n7924 n5085 R=1.248e+01 
R7923t3987 n7924 n3988 R=4.303e+01 
R7923t7850 n7924 n7851 R=9.243e+00 
R7923t2608 n7924 n2609 R=5.156e+01 
R7923t5167 n7924 n5168 R=6.043e+00 
R7923t1168 n7924 n1169 R=1.262e+01 
R7923t5568 n7924 n5569 R=2.587e+01 
R7923t5482 n7924 n5483 R=4.469e+00 
R7924t6673 n7925 n6674 R=2.659e+02 
R7924t7326 n7925 n7327 R=5.435e+00 
R7924t602 n7925 n603 R=6.316e+00 
R7924t3664 n7925 n3665 R=5.273e+01 
R7924t4967 n7925 n4968 R=6.115e+00 
R7924t5699 n7925 n5700 R=2.855e+00 
R7925t2359 n7926 n2360 R=7.388e+00 
R7925t5170 n7926 n5171 R=2.658e+00 
R7925t5589 n7926 n5590 R=2.606e+01 
R7926t533 n7927 n534 R=3.596e+00 
R7926t7484 n7927 n7485 R=2.840e+01 
R7926t3501 n7927 n3502 R=4.200e+00 
R7926t2732 n7927 n2733 R=7.254e+00 
R7926t5575 n7927 n5576 R=7.055e+00 
R7927t2214 n7928 n2215 R=5.606e+01 
R7927t2614 n7928 n2615 R=3.366e+01 
R7927t3171 n7928 n3172 R=4.525e+00 
R7927t5599 n7928 n5600 R=4.460e+00 
R7927t7611 n7928 n7612 R=2.274e+03 
R7927t1581 n7928 n1582 R=1.994e+00 
R7928t7196 n7929 n7197 R=1.858e+01 
R7928t3962 n7929 n3963 R=1.621e+01 
R7928t4620 n7929 n4621 R=3.740e+00 
R7928t2829 n7929 n2830 R=2.730e+01 
R7929t1403 n7930 n1404 R=2.133e+01 
R7929t5225 n7930 n5226 R=3.841e+00 
R7929t7793 n7930 n7794 R=8.207e+00 
R7929t2751 n7930 n2752 R=4.155e+00 
R7930t1074 n7931 n1075 R=5.232e+00 
R7930t3488 n7931 n3489 R=3.804e+00 
R7930t5797 n7931 n5798 R=3.487e+00 
R7930t576 n7931 n577 R=1.212e+01 
R7930t747 n7931 n748 R=2.820e+01 
R7931t5847 n7932 n5848 R=5.283e+00 
R7931t6142 n7932 n6143 R=5.511e+00 
R7931t1653 n7932 n1654 R=1.033e+01 
R7931t618 n7932 n619 R=3.036e+01 
R7932t311 n7933 n312 R=2.642e+00 
R7932t2180 n7933 n2181 R=2.819e+01 
R7932t5996 n7933 n5997 R=5.781e+00 
R7932t666 n7933 n667 R=3.633e+00 
R7933t2073 n7934 n2074 R=3.309e+00 
R7933t3084 n7934 n3085 R=5.144e+01 
R7933t6500 n7934 n6501 R=1.211e+02 
R7933t4238 n7934 n4239 R=1.712e+01 
R7933t1600 n7934 n1601 R=1.123e+01 
R7933t4818 n7934 n4819 R=1.712e+00 
R7934t285 n7935 n286 R=3.831e+01 
R7934t7030 n7935 n7031 R=7.778e+00 
R7934t1992 n7935 n1993 R=8.890e+00 
R7934t4471 n7935 n4472 R=4.571e+01 
R7934t1749 n7935 n1750 R=3.374e+00 
R7934t5763 n7935 n5764 R=1.556e+01 
R7935t3941 n7936 n3942 R=4.687e+00 
R7935t4216 n7936 n4217 R=4.399e+00 
R7935t3403 n7936 n3404 R=2.040e+01 
R7935t1921 n7936 n1922 R=6.691e+00 
R7935t7250 n7936 n7251 R=6.126e+00 
R7936t4553 n7937 n4554 R=2.345e+00 
R7936t7121 n7937 n7122 R=1.017e+02 
R7936t2073 n7937 n2074 R=1.868e+01 
R7936t3668 n7937 n3669 R=7.366e+00 
R7936t7870 n7937 n7871 R=7.621e+00 
R7937t2513 n7938 n2514 R=6.849e+01 
R7937t3719 n7938 n3720 R=4.401e+01 
R7937t3648 n7938 n3649 R=3.314e+01 
R7937t3760 n7938 n3761 R=5.213e+00 
R7937t4238 n7938 n4239 R=5.539e+01 
R7937t4917 n7938 n4918 R=6.155e+00 
R7937t69 n7938 n70 R=1.499e+01 
R7937t1597 n7938 n1598 R=3.358e+00 
R7937t2541 n7938 n2542 R=1.381e+01 
R7938t6319 n1 n6320 R=3.265e+00 
R7939t1385 n7940 n1386 R=5.705e+01 
R7939t1866 n7940 n1867 R=9.131e+00 
R7939t2849 n7940 n2850 R=3.525e+00 
R7939t6264 n7940 n6265 R=7.760e+00 
R7940t1539 n7941 n1540 R=9.663e+00 
R7940t5294 n7941 n5295 R=1.248e+01 
R7940t1810 n7941 n1811 R=4.695e+00 
R7940t6515 n7941 n6516 R=1.393e+01 
R7940t962 n7941 n963 R=1.442e+01 
R7940t1957 n7941 n1958 R=3.285e+00 
R7941t1804 n7942 n1805 R=3.621e+00 
R7941t5376 n7942 n5377 R=3.191e+00 
R7942t6934 n7943 n6935 R=2.249e+01 
R7942t3405 n7943 n3406 R=3.105e+01 
R7942t1782 n7943 n1783 R=1.797e+01 
R7942t7511 n7943 n7512 R=2.578e+00 
R7942t5639 n7943 n5640 R=2.387e+01 
R7942t3572 n7943 n3573 R=3.408e+00 
R7943t6518 n7944 n6519 R=5.590e+00 
R7943t7139 n7944 n7140 R=3.467e+00 
R7944t2425 n7945 n2426 R=1.079e+00 
R7944t3999 n7945 n4000 R=3.062e+00 
R7944t6789 n7945 n6790 R=6.627e+01 
R7945t4432 n7946 n4433 R=7.143e+00 
R7945t6171 n7946 n6172 R=6.052e+00 
R7945t5954 n7946 n5955 R=7.272e+00 
R7945t7407 n7946 n7408 R=6.072e+00 
R7945t2 n7946 n3 R=6.025e+00 
R7946t933 n7947 n934 R=2.305e+00 
R7946t4204 n7947 n4205 R=4.600e+03 
R7946t217 n7947 n218 R=2.023e+01 
R7946t6098 n7947 n6099 R=1.672e+00 
R7946t620 n7947 n621 R=4.534e+01 
R7946t5260 n7947 n5261 R=3.164e+01 
R7947t1363 n7948 n1364 R=1.122e+01 
R7947t3248 n7948 n3249 R=1.049e+01 
R7947t7782 n7948 n7783 R=1.253e+01 
R7947t1486 n7948 n1487 R=2.335e+01 
R7947t6599 n7948 n6600 R=5.812e+00 
R7948t1021 n7949 n1022 R=9.004e+00 
R7948t2345 n7949 n2346 R=5.080e+00 
R7948t7341 n7949 n7342 R=3.373e+00 
R7948t5128 n7949 n5129 R=7.827e+00 
R7949t2333 n7950 n2334 R=5.810e+00 
R7949t6587 n7950 n6588 R=3.551e+01 
R7949t3893 n7950 n3894 R=1.584e+01 
R7949t6786 n7950 n6787 R=5.225e+00 
R7949t5904 n7950 n5905 R=1.472e+01 
R7950t6492 n7951 n6493 R=5.189e+00 
R7950t3792 n7951 n3793 R=2.017e+01 
R7951t5031 n7952 n5032 R=5.476e+00 
R7951t7512 n7952 n7513 R=3.835e+00 
R7951t1411 n7952 n1412 R=3.743e+01 
R7951t7684 n7952 n7685 R=2.689e+00 
R7951t4387 n7952 n4388 R=8.849e+00 
R7952t4531 n7953 n4532 R=4.384e+00 
R7952t6766 n7953 n6767 R=3.316e+00 
R7952t7242 n7953 n7243 R=3.958e+00 
R7952t2518 n7953 n2519 R=2.714e+01 
R7953t4665 n7954 n4666 R=7.470e+00 
R7953t5935 n7954 n5936 R=9.009e+01 
R7953t2003 n7954 n2004 R=3.305e+00 
R7953t4143 n7954 n4144 R=2.445e+00 
R7953t996 n7954 n997 R=3.370e+01 
R7954t169 n7955 n170 R=2.842e+00 
R7954t1470 n7955 n1471 R=9.162e+00 
R7954t4858 n7955 n4859 R=1.251e+01 
R7954t2516 n7955 n2517 R=5.183e+00 
R7955t1870 n7956 n1871 R=2.908e+00 
R7955t6589 n7956 n6590 R=1.907e+01 
R7955t3693 n7956 n3694 R=5.021e+00 
R7955t2627 n7956 n2628 R=1.902e+02 
R7955t2090 n7956 n2091 R=4.743e+00 
R7955t7107 n7956 n7108 R=1.961e+01 
R7955t4747 n7956 n4748 R=4.091e+01 
R7956t91 n7957 n92 R=5.121e+00 
R7956t7421 n7957 n7422 R=4.413e+00 
R7956t3402 n7957 n3403 R=1.292e+01 
R7956t406 n7957 n407 R=4.058e+00 
R7956t473 n7957 n474 R=6.648e+00 
R7957t1073 n7958 n1074 R=2.340e+00 
R7957t5681 n7958 n5682 R=1.680e+02 
R7957t5839 n7958 n5840 R=3.196e+00 
R7957t661 n7958 n662 R=7.455e+00 
R7958t5349 n7959 n5350 R=1.057e+02 
R7958t4274 n7959 n4275 R=5.453e+00 
R7958t6288 n7959 n6289 R=1.657e+01 
R7958t38 n7959 n39 R=4.956e+00 
R7959t743 n7960 n744 R=5.646e+00 
R7959t6677 n7960 n6678 R=2.783e+01 
R7959t5284 n7960 n5285 R=4.578e+00 
R7959t385 n7960 n386 R=1.912e+01 
R7959t2615 n7960 n2616 R=2.301e+00 
R7960t1002 n7961 n1003 R=1.324e+01 
R7960t3322 n7961 n3323 R=3.712e+01 
R7960t3858 n7961 n3859 R=1.604e+01 
R7960t5911 n7961 n5912 R=6.198e+00 
R7960t1077 n7961 n1078 R=3.787e+00 
R7960t3899 n7961 n3900 R=2.086e+01 
R7961t2481 n7962 n2482 R=2.943e+01 
R7961t6530 n7962 n6531 R=1.643e+01 
R7961t1663 n7962 n1664 R=1.249e+01 
R7961t2201 n7962 n2202 R=2.860e+00 
R7961t5626 n7962 n5627 R=7.454e+01 
R7961t6726 n7962 n6727 R=1.020e+03 
R7961t6787 n7962 n6788 R=1.842e+00 
R7962t1498 n7963 n1499 R=5.488e+00 
R7962t6496 n7963 n6497 R=1.873e+01 
R7962t535 n7963 n536 R=7.781e+00 
R7962t6836 n7963 n6837 R=6.977e+00 
R7963t686 n7964 n687 R=5.485e+01 
R7963t6916 n7964 n6917 R=2.863e+00 
R7963t7865 n7964 n7866 R=3.553e+00 
R7963t745 n7964 n746 R=2.008e+00 
R7964t4335 n7965 n4336 R=9.065e+00 
R7964t5524 n7965 n5525 R=7.784e+00 
R7964t7838 n7965 n7839 R=1.694e+01 
R7964t1375 n7965 n1376 R=5.616e+00 
R7965t3710 n7966 n3711 R=2.783e+00 
R7965t4241 n7966 n4242 R=2.997e+01 
R7965t6890 n7966 n6891 R=1.726e+01 
R7965t1921 n7966 n1922 R=2.510e+01 
R7965t729 n7966 n730 R=1.679e+01 
R7965t4559 n7966 n4560 R=4.143e+00 
R7965t2635 n7966 n2636 R=1.348e+02 
R7965t6332 n7966 n6333 R=2.206e+01 
R7965t3054 n7966 n3055 R=1.876e+01 
R7966t3725 n7967 n3726 R=4.828e+01 
R7966t4413 n7967 n4414 R=2.016e+01 
R7966t2800 n7967 n2801 R=5.588e+00 
R7966t2427 n7967 n2428 R=3.123e+00 
R7967t5112 n7968 n5113 R=4.320e+02 
R7967t4014 n7968 n4015 R=2.917e+00 
R7967t1802 n7968 n1803 R=2.365e+01 
R7967t203 n7968 n204 R=3.181e+01 
R7968t647 n7969 n648 R=3.448e+00 
R7968t6504 n7969 n6505 R=2.177e+01 
R7968t6123 n7969 n6124 R=3.840e+01 
R7968t4417 n7969 n4418 R=6.076e+00 
R7968t7292 n7969 n7293 R=6.876e+00 
R7969t4227 n7970 n4228 R=5.383e+00 
R7969t7793 n7970 n7794 R=2.622e+00 
R7969t1583 n7970 n1584 R=2.822e+00 
R7969t5746 n7970 n5747 R=5.163e+01 
R7969t2751 n7970 n2752 R=1.008e+02 
R7969t7929 n7970 n7930 R=1.584e+01 
R7970t2274 n7971 n2275 R=5.945e+00 
R7970t499 n7971 n500 R=3.538e+01 
R7970t5893 n7971 n5894 R=8.902e+00 
R7970t3746 n7971 n3747 R=8.368e+00 
R7971t1674 n7972 n1675 R=4.106e+00 
R7971t2659 n7972 n2660 R=3.736e+01 
R7971t6668 n7972 n6669 R=9.081e+00 
R7971t3954 n7972 n3955 R=3.104e+00 
R7972t186 n7973 n187 R=6.118e+00 
R7972t321 n7973 n322 R=1.028e+01 
R7972t319 n7973 n320 R=5.702e+00 
R7972t5148 n7973 n5149 R=2.605e+01 
R7972t1095 n7973 n1096 R=6.743e+01 
R7972t5478 n7973 n5479 R=3.042e+00 
R7972t4407 n7973 n4408 R=3.706e+01 
R7973t5118 n7974 n5119 R=6.666e+00 
R7973t2666 n7974 n2667 R=1.344e+01 
R7973t1902 n7974 n1903 R=4.234e+01 
R7973t617 n7974 n618 R=5.552e+00 
R7973t6400 n7974 n6401 R=2.556e+01 
R7973t2064 n7974 n2065 R=5.482e+01 
R7974t7501 n7975 n7502 R=1.957e+00 
R7974t5280 n7975 n5281 R=3.072e+02 
R7974t1561 n7975 n1562 R=6.848e+00 
R7974t1785 n7975 n1786 R=1.385e+01 
R7975t2152 n7976 n2153 R=8.305e+00 
R7975t7298 n7976 n7299 R=4.590e+00 
R7975t3578 n7976 n3579 R=2.931e+00 
R7975t5544 n7976 n5545 R=5.897e+00 
R7976t1454 n7977 n1455 R=3.064e+00 
R7976t3963 n7977 n3964 R=2.332e+01 
R7976t6812 n7977 n6813 R=4.428e+00 
R7976t1067 n7977 n1068 R=2.780e+00 
R7977t1148 n7978 n1149 R=1.265e+01 
R7977t4393 n7978 n4394 R=6.833e+00 
R7977t4437 n7978 n4438 R=1.101e+01 
R7977t4705 n7978 n4706 R=3.919e+00 
R7978t4990 n7979 n4991 R=3.478e+00 
R7978t3676 n7979 n3677 R=3.167e+00 
R7979t509 n7980 n510 R=5.737e+00 
R7979t2675 n7980 n2676 R=5.897e+00 
R7979t5470 n7980 n5471 R=7.222e+00 
R7979t3465 n7980 n3466 R=3.968e+00 
R7980t3598 n7981 n3599 R=1.533e+00 
R7980t3704 n7981 n3705 R=3.730e+01 
R7980t6057 n7981 n6058 R=7.604e+00 
R7980t1211 n7981 n1212 R=2.426e+00 
R7981t2068 n7982 n2069 R=2.780e+00 
R7982t3853 n7983 n3854 R=1.455e+01 
R7982t4352 n7983 n4353 R=6.033e+00 
R7982t6807 n7983 n6808 R=2.378e+01 
R7982t7520 n7983 n7521 R=4.517e+00 
R7982t2696 n7983 n2697 R=6.767e+00 
R7982t7697 n7983 n7698 R=4.212e+01 
R7983t1391 n7984 n1392 R=5.533e+01 
R7984t1676 n7985 n1677 R=2.744e+00 
R7984t5176 n7985 n5177 R=5.944e+01 
R7984t6733 n7985 n6734 R=7.385e+00 
R7984t1162 n7985 n1163 R=3.896e+00 
R7984t5901 n7985 n5902 R=9.594e+00 
R7985t650 n7986 n651 R=1.227e+01 
R7985t721 n7986 n722 R=4.742e+00 
R7985t203 n7986 n204 R=1.109e+01 
R7986t5985 n7987 n5986 R=8.453e+00 
R7986t6264 n7987 n6265 R=2.300e+00 
R7986t4281 n7987 n4282 R=4.697e+00 
R7986t553 n7987 n554 R=1.404e+01 
R7987t1675 n7988 n1676 R=5.254e+01 
R7987t5358 n7988 n5359 R=5.241e+00 
R7987t7756 n7988 n7757 R=1.659e+02 
R7988t1696 n7989 n1697 R=8.079e+00 
R7988t2795 n7989 n2796 R=4.025e+00 
R7988t3102 n7989 n3103 R=4.114e+00 
R7988t7874 n7989 n7875 R=4.004e+00 
R7989t1141 n7990 n1142 R=1.863e+00 
R7989t694 n7990 n695 R=2.636e+02 
R7989t5430 n7990 n5431 R=7.426e+00 
R7989t2105 n7990 n2106 R=1.581e+01 
R7990t3660 n7991 n3661 R=1.527e+01 
R7990t5688 n7991 n5689 R=4.018e+01 
R7990t3468 n7991 n3469 R=3.692e+00 
R7990t3183 n7991 n3184 R=2.243e+01 
R7990t1219 n7991 n1220 R=4.980e+00 
R7991t1952 n7992 n1953 R=5.615e+00 
R7991t5408 n7992 n5409 R=2.104e+01 
R7991t6051 n7992 n6052 R=3.179e+00 
R7991t6867 n7992 n6868 R=4.717e+01 
R7991t3696 n7992 n3697 R=2.622e+00 
R7992t1548 n7993 n1549 R=8.053e+01 
R7992t5350 n7993 n5351 R=7.220e+00 
R7992t6644 n7993 n6645 R=1.642e+01 
R7992t4846 n7993 n4847 R=9.464e+00 
R7993t5485 n7994 n5486 R=6.059e+00 
R7993t6461 n7994 n6462 R=6.925e+00 
R7993t4762 n7994 n4763 R=8.801e+00 
R7993t1205 n7994 n1206 R=4.632e+00 
R7993t5799 n7994 n5800 R=3.527e+01 
R7994t5062 n7995 n5063 R=4.771e+00 
R7994t4498 n7995 n4499 R=5.074e+00 
R7994t2431 n7995 n2432 R=2.236e+00 
R7995t4637 n7996 n4638 R=1.081e+01 
R7995t3505 n7996 n3506 R=3.685e+01 
R7995t6647 n7996 n6648 R=5.231e+00 
R7995t3776 n7996 n3777 R=2.905e+01 
R7996t255 n7997 n256 R=3.286e+00 
R7996t2608 n7997 n2609 R=7.011e+00 
R7996t5597 n7997 n5598 R=2.345e+01 
R7996t1761 n7997 n1762 R=9.888e+00 
R7996t7850 n7997 n7851 R=3.810e+01 
R7997t4064 n7998 n4065 R=5.928e+00 
R7997t4068 n7998 n4069 R=5.119e+00 
R7997t1509 n7998 n1510 R=1.764e+01 
R7997t4175 n7998 n4176 R=3.242e+00 
R7997t4634 n7998 n4635 R=3.047e+01 
R7998t2684 n7999 n2685 R=4.286e+00 
R7998t7289 n7999 n7290 R=2.447e+01 
R7998t917 n7999 n918 R=6.199e+00 
R7998t4581 n7999 n4582 R=9.511e+00 
R7998t7443 n7999 n7444 R=1.559e+01 
R7998t3978 n7999 n3979 R=5.890e+00 
R7998t7217 n7999 n7218 R=3.046e+01 
R7999t5474 n8000 n5475 R=1.577e+00 
R7999t6510 n8000 n6511 R=2.748e+00 
R7999t442 n8000 n443 R=1.607e+01 
R8000t927 n8001 n928 R=1.894e+01 
R8000t1658 n8001 n1659 R=3.847e+00 
R8000t1239 n8001 n1240 R=8.335e+00 
R8001t572 n8002 n573 R=6.968e+00 
R8001t1510 n8002 n1511 R=7.806e+00 
R8001t2135 n8002 n2136 R=2.192e+01 
R8001t7765 n8002 n7766 R=1.995e+01 
R8001t2723 n8002 n2724 R=6.500e+01 
R8001t749 n8002 n750 R=4.662e+00 
R8002t693 n8003 n694 R=1.365e+01 
R8002t1446 n8003 n1447 R=1.417e+01 
R8002t4010 n8003 n4011 R=8.170e+00 
R8002t1143 n8003 n1144 R=6.772e+00 
R8002t538 n8003 n539 R=1.155e+01 
R8002t5786 n8003 n5787 R=6.993e+01 
R8002t2461 n8003 n2462 R=3.729e+00 
R8003t8000 n8004 n8001 R=9.370e+01 
R8003t1151 n8004 n1152 R=1.024e+01 
R8003t5255 n8004 n5256 R=4.147e+00 
R8003t580 n8004 n581 R=6.836e+00 
R8003t1239 n8004 n1240 R=4.340e+00 
R8004t513 n8005 n514 R=1.096e+01 
R8004t7789 n8005 n7790 R=4.835e+00 
R8004t3925 n8005 n3926 R=5.608e+00 
R8004t1511 n8005 n1512 R=9.110e+00 
R8004t6631 n8005 n6632 R=4.018e+01 
R8005t4995 n8006 n4996 R=2.013e+01 
R8005t7034 n8006 n7035 R=6.789e+00 
R8005t72 n8006 n73 R=8.222e+01 
R8006t510 n8007 n511 R=4.125e+00 
R8006t1767 n8007 n1768 R=4.198e+00 
R8007t55 n8008 n56 R=5.983e+00 
R8007t5274 n8008 n5275 R=1.143e+02 
R8007t2102 n8008 n2103 R=3.044e+00 
R8007t3286 n8008 n3287 R=1.006e+01 
R8007t2453 n8008 n2454 R=3.435e+00 
R8007t7842 n8008 n7843 R=2.170e+01 
R8008t628 n8009 n629 R=2.721e+01 
R8008t4388 n8009 n4389 R=8.757e+00 
R8008t3393 n8009 n3394 R=1.092e+01 
R8008t5514 n8009 n5515 R=1.584e+01 
R8008t2875 n8009 n2876 R=9.455e+00 
R8008t6450 n8009 n6451 R=1.036e+01 
R8008t5851 n8009 n5852 R=5.818e+00 
R8009t940 n8010 n941 R=6.722e+00 
R8009t5799 n8010 n5800 R=2.361e+01 
R8009t452 n8010 n453 R=4.123e+00 
R8009t2853 n8010 n2854 R=1.918e+01 
R8009t2445 n8010 n2446 R=5.337e+00 
R8010t1859 n8011 n1860 R=2.605e+00 
R8010t2588 n8011 n2589 R=7.260e+00 
R8010t1522 n8011 n1523 R=2.104e+00 
R8010t1754 n8011 n1755 R=2.117e+01 
R8011t534 n8012 n535 R=7.243e+00 
R8011t7157 n8012 n7158 R=3.431e+00 
R8011t5761 n8012 n5762 R=1.558e+01 
R8011t85 n8012 n86 R=9.154e+00 
R8011t3177 n8012 n3178 R=2.243e+01 
R8012t4043 n8013 n4044 R=4.498e+00 
R8012t4653 n8013 n4654 R=2.104e+01 
R8012t660 n8013 n661 R=5.006e+00 
R8012t7401 n8013 n7402 R=1.055e+02 
R8012t3454 n8013 n3455 R=5.560e+00 
R8013t736 n8014 n737 R=1.674e+01 
R8013t4757 n8014 n4758 R=3.921e+00 
R8013t6724 n8014 n6725 R=2.961e+00 
R8013t1772 n8014 n1773 R=2.009e+01 
R8013t90 n8014 n91 R=5.046e+00 
R8014t1131 n8015 n1132 R=4.989e+00 
R8014t1974 n8015 n1975 R=8.254e+00 
R8014t3848 n8015 n3849 R=3.630e+02 
R8014t2652 n8015 n2653 R=3.270e+00 
R8014t2845 n8015 n2846 R=6.606e+01 
R8014t4837 n8015 n4838 R=7.279e+00 
R8015t1805 n8016 n1806 R=5.121e+00 
R8015t5205 n8016 n5206 R=1.370e+01 
R8015t653 n8016 n654 R=7.699e+00 
R8016t437 n8017 n438 R=1.200e+02 
R8016t6223 n8017 n6224 R=1.555e+00 
R8016t646 n8017 n647 R=4.337e+01 
R8016t7807 n8017 n7808 R=8.451e+00 
R8016t7008 n8017 n7009 R=3.826e+00 
R8017t177 n8018 n178 R=1.202e+01 
R8017t1042 n8018 n1043 R=2.209e+01 
R8017t6007 n8018 n6008 R=1.484e+01 
R8017t7239 n8018 n7240 R=5.791e+00 
R8017t5642 n8018 n5643 R=1.958e+01 
R8017t2977 n8018 n2978 R=9.574e+01 
R8017t7110 n8018 n7111 R=1.023e+01 
R8018t3347 n8019 n3348 R=9.612e+00 
R8018t3907 n8019 n3908 R=5.442e+00 
R8018t4987 n8019 n4988 R=1.319e+01 
R8019t526 n8020 n527 R=3.751e+00 
R8019t3795 n8020 n3796 R=3.037e+00 
R8019t4507 n8020 n4508 R=2.145e+01 
R8020t665 n8021 n666 R=3.289e+01 
R8020t1326 n8021 n1327 R=5.822e+01 
R8020t482 n8021 n483 R=2.241e+00 
R8020t7136 n8021 n7137 R=3.756e+01 
R8020t7249 n8021 n7250 R=5.131e+00 
R8020t6357 n8021 n6358 R=1.362e+01 
R8021t448 n8022 n449 R=5.558e+01 
R8021t3063 n8022 n3064 R=4.616e+00 
R8021t3686 n8022 n3687 R=6.567e+00 
R8021t3939 n8022 n3940 R=9.821e+00 
R8022t4300 n8023 n4301 R=2.747e+01 
R8022t6947 n8023 n6948 R=4.718e+00 
R8022t6985 n8023 n6986 R=3.549e+01 
R8022t7440 n8023 n7441 R=6.145e+00 
R8022t1072 n8023 n1073 R=1.732e+01 
R8022t5480 n8023 n5481 R=6.823e+00 
R8023t3942 n8024 n3943 R=7.933e+00 
R8023t4412 n8024 n4413 R=3.067e+00 
R8023t165 n8024 n166 R=1.184e+01 
R8023t308 n8024 n309 R=1.171e+01 
R8023t5983 n8024 n5984 R=1.436e+01 
R8024t208 n8025 n209 R=1.135e+01 
R8024t6211 n8025 n6212 R=1.090e+01 
R8024t124 n8025 n125 R=1.925e+01 
R8024t1506 n8025 n1507 R=1.158e+01 
R8024t2485 n8025 n2486 R=4.409e+00 
R8024t7069 n8025 n7070 R=3.160e+01 
R8024t2773 n8025 n2774 R=3.273e+00 
R8025t281 n8026 n282 R=2.287e+02 
R8025t1200 n8026 n1201 R=1.099e+01 
R8025t7273 n8026 n7274 R=9.403e+00 
R8025t351 n8026 n352 R=3.852e+00 
R8025t957 n8026 n958 R=1.223e+01 
R8025t4746 n8026 n4747 R=4.673e+00 
R8026t7395 n8027 n7396 R=4.744e+00 
R8026t6458 n8027 n6459 R=3.687e+00 
R8026t4058 n8027 n4059 R=1.574e+01 
R8026t3823 n8027 n3824 R=1.732e+01 
R8026t99 n8027 n100 R=8.901e+00 
R8027t882 n8028 n883 R=2.924e+01 
R8027t6432 n8028 n6433 R=2.564e+01 
R8027t7120 n8028 n7121 R=3.735e+01 
R8027t2540 n8028 n2541 R=9.362e+00 
R8027t2509 n8028 n2510 R=1.133e+01 
R8027t4183 n8028 n4184 R=3.756e+00 
R8027t3503 n8028 n3504 R=1.362e+01 
R8027t4120 n8028 n4121 R=7.687e+01 
R8027t6894 n8028 n6895 R=4.650e+00 
R8028t1633 n8029 n1634 R=6.060e+00 
R8028t4371 n8029 n4372 R=3.608e+01 
R8028t4601 n8029 n4602 R=1.725e+01 
R8028t2901 n8029 n2902 R=1.602e+01 
R8028t5405 n8029 n5406 R=4.995e+01 
R8028t5150 n8029 n5151 R=4.141e+00 
R8028t7628 n8029 n7629 R=2.218e+01 
R8028t2641 n8029 n2642 R=5.782e+00 
R8029t2217 n8030 n2218 R=3.318e+00 
R8029t2257 n8030 n2258 R=6.896e+00 
R8029t4386 n8030 n4387 R=5.431e+01 
R8029t5860 n8030 n5861 R=1.019e+01 
R8029t2940 n8030 n2941 R=5.016e+00 
R8029t5540 n8030 n5541 R=2.539e+01 
R8030t4001 n8031 n4002 R=5.836e+00 
R8030t7881 n8031 n7882 R=2.049e+01 
R8030t7427 n8031 n7428 R=6.010e+00 
R8030t7830 n8031 n7831 R=2.875e+01 
R8030t5870 n8031 n5871 R=8.452e+00 
R8030t7050 n8031 n7051 R=3.597e+00 
R8031t2084 n8032 n2085 R=3.582e+00 
R8031t5806 n8032 n5807 R=6.893e+00 
R8031t99 n8032 n100 R=6.296e+00 
R8031t3823 n8032 n3824 R=2.906e+01 
R8032t7420 n8033 n7421 R=1.734e+00 
R8032t7441 n8033 n7442 R=1.427e+01 
R8032t949 n8033 n950 R=1.338e+01 
R8032t2006 n8033 n2007 R=1.156e+01 
R8032t1984 n8033 n1985 R=7.922e+01 
R8033t389 n8034 n390 R=2.482e+00 
R8033t6800 n8034 n6801 R=1.149e+02 
R8033t347 n8034 n348 R=7.281e+00 
R8033t2010 n8034 n2011 R=3.638e+00 
R8033t7286 n8034 n7287 R=4.936e+00 
R8034t5743 n8035 n5744 R=1.935e+02 
R8034t6821 n8035 n6822 R=1.650e+01 
R8034t1999 n8035 n2000 R=3.164e+00 
R8034t5928 n8035 n5929 R=1.213e+01 
R8034t2027 n8035 n2028 R=8.272e+00 
R8034t536 n8035 n537 R=5.860e+00 
R8035t3928 n8036 n3929 R=8.101e+01 
R8035t7838 n8036 n7839 R=4.396e+00 
R8035t5524 n8036 n5525 R=4.601e+00 
R8035t2958 n8036 n2959 R=2.515e+01 
R8035t2673 n8036 n2674 R=8.488e+00 
R8035t5153 n8036 n5154 R=4.404e+00 
R8036t4391 n8037 n4392 R=5.069e+00 
R8036t7329 n8037 n7330 R=7.416e+00 
R8037t1707 n8038 n1708 R=3.716e+00 
R8037t587 n8038 n588 R=4.506e+00 
R8037t1137 n8038 n1138 R=3.069e+00 
R8038t3128 n8039 n3129 R=7.895e+00 
R8038t3669 n8039 n3670 R=5.142e+00 
R8039t367 n8040 n368 R=2.687e+02 
R8039t7024 n8040 n7025 R=1.018e+01 
R8039t6871 n8040 n6872 R=1.408e+01 
R8039t7538 n8040 n7539 R=2.852e+00 
R8040t1062 n8041 n1063 R=2.295e+01 
R8040t3073 n8041 n3074 R=2.672e+00 
R8040t1234 n8041 n1235 R=7.962e+01 
R8040t6447 n8041 n6448 R=6.682e+00 
R8040t4643 n8041 n4644 R=1.035e+01 
R8041t5633 n8042 n5634 R=2.433e+00 
R8041t5419 n8042 n5420 R=8.049e+00 
R8041t3935 n8042 n3936 R=2.329e+00 
R8041t6856 n8042 n6857 R=3.073e+01 
R8042t636 n8043 n637 R=7.708e+00 
R8042t1396 n8043 n1397 R=6.402e+00 
R8042t7618 n8043 n7619 R=5.059e+00 
R8042t5290 n8043 n5291 R=1.021e+02 
R8042t2853 n8043 n2854 R=6.161e+00 
R8042t796 n8043 n797 R=9.282e+00 
R8043t7987 n8044 n7988 R=4.024e+00 
R8043t7756 n8044 n7757 R=7.476e+00 
R8043t2070 n8044 n2071 R=1.351e+01 
R8043t4475 n8044 n4476 R=7.489e+00 
R8043t1425 n8044 n1426 R=1.489e+01 
R8044t6465 n8045 n6466 R=2.887e+00 
R8044t4998 n8045 n4999 R=1.074e+02 
R8044t7141 n8045 n7142 R=8.296e+00 
R8044t1246 n8045 n1247 R=9.958e+00 
R8044t2117 n8045 n2118 R=1.115e+01 
R8045t7877 n8046 n7878 R=8.865e+01 
R8045t1935 n8046 n1936 R=1.609e+01 
R8045t285 n8046 n286 R=2.113e+01 
R8045t1992 n8046 n1993 R=2.020e+01 
R8045t40 n8046 n41 R=6.322e+00 
R8046t7083 n8047 n7084 R=2.428e+03 
R8046t2353 n8047 n2354 R=3.869e+00 
R8046t5694 n8047 n5695 R=4.346e+00 
R8046t2905 n8047 n2906 R=7.023e+00 
R8047t6265 n8048 n6266 R=1.455e+01 
R8047t1261 n8048 n1262 R=8.014e+00 
R8047t4840 n8048 n4841 R=2.511e+00 
R8047t2909 n8048 n2910 R=9.653e+00 
R8047t1735 n8048 n1736 R=1.440e+01 
R8048t3592 n8049 n3593 R=6.251e+01 
R8048t5889 n8049 n5890 R=8.427e+00 
R8048t5569 n8049 n5570 R=2.470e+00 
R8048t3782 n8049 n3783 R=4.505e+01 
R8048t1255 n8049 n1256 R=4.764e+01 
R8048t1913 n8049 n1914 R=1.311e+01 
R8048t5222 n8049 n5223 R=1.124e+01 
R8049t7092 n8050 n7093 R=1.331e+01 
R8049t7308 n8050 n7309 R=2.576e+00 
R8049t4347 n8050 n4348 R=5.444e+00 
R8050t1345 n8051 n1346 R=5.900e+00 
R8050t6050 n8051 n6051 R=4.532e+00 
R8050t7448 n8051 n7449 R=2.146e+01 
R8050t725 n8051 n726 R=2.652e+01 
R8050t5964 n8051 n5965 R=6.106e+00 
R8050t4341 n8051 n4342 R=4.120e+01 
R8051t4290 n8052 n4291 R=6.912e+01 
R8051t7531 n8052 n7532 R=1.462e+01 
R8051t7913 n8052 n7914 R=3.202e+00 
R8051t5640 n8052 n5641 R=7.685e+00 
R8051t5408 n8052 n5409 R=2.863e+01 
R8051t326 n8052 n327 R=2.537e+00 
R8051t1710 n8052 n1711 R=9.914e+00 
R8052t547 n8053 n548 R=1.069e+01 
R8052t4105 n8053 n4106 R=2.695e+01 
R8052t4191 n8053 n4192 R=4.362e+00 
R8052t2456 n8053 n2457 R=5.094e+01 
R8052t1393 n8053 n1394 R=8.366e+00 
R8053t273 n8054 n274 R=7.119e+00 
R8053t3 n8054 n4 R=4.808e+00 
R8053t7844 n8054 n7845 R=3.581e+00 
R8054t723 n8055 n724 R=4.423e+00 
R8055t1334 n8056 n1335 R=1.470e+00 
R8055t2544 n8056 n2545 R=1.513e+01 
R8055t2781 n8056 n2782 R=5.197e+00 
R8055t3002 n8056 n3003 R=6.160e+00 
R8055t6503 n8056 n6504 R=6.139e+01 
R8056t3279 n8057 n3280 R=1.189e+01 
R8056t7022 n8057 n7023 R=3.715e+00 
R8056t2411 n8057 n2412 R=3.040e+01 
R8056t1731 n8057 n1732 R=9.450e+00 
R8056t6327 n8057 n6328 R=9.582e+00 
R8056t5608 n8057 n5609 R=4.349e+01 
R8057t1147 n8058 n1148 R=2.948e+00 
R8057t4125 n8058 n4126 R=6.858e+00 
R8057t2736 n8058 n2737 R=5.280e+00 
R8057t2960 n8058 n2961 R=5.251e+00 
R8057t1682 n8058 n1683 R=1.368e+01 
R8058t7832 n8059 n7833 R=7.643e+00 
R8058t77 n8059 n78 R=8.916e+00 
R8058t1424 n8059 n1425 R=5.025e+00 
R8058t7884 n8059 n7885 R=6.857e+00 
R8058t5668 n8059 n5669 R=2.752e+01 
R8059t568 n8060 n569 R=2.722e+00 
R8059t3060 n8060 n3061 R=1.037e+01 
R8059t319 n8060 n320 R=1.030e+01 
R8059t5148 n8060 n5149 R=2.835e+00 
R8059t7907 n8060 n7908 R=2.220e+01 
R8060t1708 n8061 n1 R=2.028e+01 
R8060t7222 n8061 n7223 R=4.891e+00 
R8060t4034 n8061 n4035 R=6.068e+00 
R8060t1419 n8061 n1420 R=1.065e+01 
R8060t1626 n8061 n1627 R=2.289e+00 
R8061t5115 n8062 n5116 R=2.251e+01 
R8061t7832 n8062 n7833 R=4.079e+00 
R8061t1689 n8062 n1690 R=4.779e+00 
R8061t5277 n8062 n5278 R=2.000e+01 
R8061t5832 n8062 n5833 R=7.503e+00 
R8062t4866 n8063 n4867 R=5.759e+00 
R8062t2288 n8063 n2289 R=7.231e+00 
R8062t7078 n8063 n7079 R=9.975e+00 
R8062t1609 n8063 n1610 R=5.863e+00 
R8063t1816 n8064 n1817 R=4.507e+00 
R8063t4753 n8064 n4754 R=3.381e+00 
R8063t5275 n8064 n5276 R=8.368e+01 
R8064t5863 n8065 n5864 R=4.396e+02 
R8064t6952 n8065 n6953 R=1.084e+01 
R8064t1262 n8065 n1263 R=8.528e+00 
R8064t4176 n8065 n4177 R=4.673e+00 
R8064t3410 n8065 n3411 R=2.327e+00 
R8065t2555 n8066 n2556 R=4.365e+00 
R8065t6688 n8066 n6689 R=3.229e+00 
R8066t1125 n8067 n1126 R=1.875e+00 
R8066t3053 n8067 n3054 R=1.477e+01 
R8066t4187 n8067 n4188 R=1.801e+02 
R8066t6056 n8067 n6057 R=4.296e+01 
R8066t3172 n8067 n3173 R=4.959e+02 
R8066t6858 n8067 n6859 R=2.146e+00 
R8066t2470 n8067 n2471 R=9.246e+00 
R8066t2031 n8067 n2032 R=2.942e+01 
R8067t4050 n8068 n4051 R=9.054e+00 
R8067t2146 n8068 n2147 R=9.286e+01 
R8067t5017 n8068 n5018 R=1.080e+01 
R8067t6714 n8068 n6715 R=1.907e+01 
R8067t3684 n8068 n3685 R=1.394e+01 
R8067t3016 n8068 n3017 R=1.164e+01 
R8067t954 n8068 n955 R=1.355e+01 
R8068t5877 n8069 n5878 R=8.627e+00 
R8068t5991 n8069 n5992 R=3.211e+00 
R8068t6097 n8069 n6098 R=4.362e+02 
R8068t6704 n8069 n6705 R=3.187e+00 
R8068t1959 n8069 n1960 R=1.625e+01 
R8068t7511 n8069 n7512 R=2.185e+02 
R8068t5639 n8069 n5640 R=3.083e+01 
R8069t97 n8070 n98 R=2.316e+00 
R8069t7370 n8070 n7371 R=4.606e+01 
R8069t2266 n8070 n2267 R=2.147e+00 
R8069t7330 n8070 n7331 R=8.082e+00 
R8070t3628 n8071 n3629 R=2.483e+00 
R8070t1555 n8071 n1556 R=3.545e+00 
R8070t4552 n8071 n4553 R=4.011e+01 
R8071t7400 n8072 n7401 R=1.198e+02 
R8071t5794 n8072 n5795 R=3.741e+01 
R8071t7674 n8072 n7675 R=3.515e+01 
R8071t5977 n8072 n5978 R=8.523e+00 
R8071t4588 n8072 n4589 R=2.337e+01 
R8071t2070 n8072 n2071 R=6.681e+00 
R8071t6577 n8072 n6578 R=5.949e+00 
R8072t339 n8073 n340 R=4.457e+01 
R8072t1739 n8073 n1740 R=1.752e+01 
R8072t1933 n8073 n1934 R=3.035e+00 
R8072t1834 n8073 n1835 R=6.221e+00 
R8072t3828 n8073 n3829 R=6.546e+00 
R8073t5652 n8074 n5653 R=1.837e+01 
R8073t235 n8074 n236 R=4.117e+00 
R8073t7624 n8074 n7625 R=4.501e+00 
R8073t4740 n8074 n4741 R=4.111e+00 
R8074t7454 n8075 n7455 R=4.456e+00 
R8074t4785 n8075 n4786 R=1.581e+02 
R8074t777 n8075 n778 R=1.154e+01 
R8074t7308 n8075 n7309 R=1.088e+02 
R8074t8049 n8075 n8050 R=1.569e+01 
R8075t1538 n8076 n1539 R=8.288e+01 
R8075t5259 n8076 n5260 R=6.650e+03 
R8075t6790 n8076 n6791 R=1.513e+01 
R8075t668 n8076 n669 R=4.068e+00 
R8076t4109 n8077 n4110 R=4.599e+00 
R8076t6361 n8077 n6362 R=8.386e+00 
R8076t4429 n8077 n4430 R=1.667e+01 
R8076t4863 n8077 n4864 R=6.482e+01 
R8076t4544 n8077 n4545 R=1.776e+01 
R8077t3193 n8078 n3194 R=1.290e+01 
R8077t5821 n8078 n5822 R=2.152e+01 
R8077t3126 n8078 n3127 R=2.910e+01 
R8077t6390 n8078 n6391 R=5.651e+00 
R8077t4578 n8078 n4579 R=4.289e+00 
R8078t5378 n8079 n5379 R=7.135e+00 
R8078t6948 n8079 n6949 R=4.666e+03 
R8078t4886 n8079 n4887 R=6.810e+00 
R8078t4611 n8079 n4612 R=7.448e+00 
R8078t492 n8079 n493 R=6.660e+01 
R8078t6979 n8079 n6980 R=4.477e+00 
R8079t88 n8080 n89 R=1.462e+02 
R8079t4843 n8080 n4844 R=2.332e+01 
R8079t5053 n8080 n5054 R=1.146e+01 
R8079t1658 n8080 n1659 R=2.874e+02 
R8079t4791 n8080 n4792 R=1.762e+01 
R8079t1476 n8080 n1477 R=1.787e+01 
R8079t3897 n8080 n3898 R=4.102e+00 
R8080t6379 n8081 n6380 R=9.620e+00 
R8080t7620 n8081 n7621 R=3.677e+00 
R8080t881 n8081 n882 R=1.323e+01 
R8080t3082 n8081 n3083 R=4.886e+00 
R8080t2314 n8081 n2315 R=4.489e+00 
R8081t379 n8082 n380 R=5.958e+00 
R8081t7480 n8082 n7481 R=2.330e+01 
R8081t2999 n8082 n3000 R=6.721e+00 
R8081t4306 n8082 n4307 R=4.837e+00 
R8081t2556 n8082 n2557 R=2.691e+02 
R8081t7017 n8082 n7018 R=7.982e+00 
R8081t1105 n8082 n1106 R=1.399e+01 
R8082t1496 n8083 n1497 R=4.505e+00 
R8082t7139 n8083 n7140 R=7.326e+02 
R8082t2039 n8083 n2040 R=3.940e+00 
R8083t6150 n8084 n6151 R=7.812e+00 
R8083t7813 n8084 n7814 R=6.060e+00 
R8083t5179 n8084 n5180 R=3.388e+00 
R8083t1809 n8084 n1810 R=9.208e+00 
R8083t4491 n8084 n4492 R=1.095e+01 
R8084t5741 n8085 n5742 R=1.135e+02 
R8084t7747 n8085 n7748 R=4.369e+00 
R8084t3137 n8085 n3138 R=3.976e+00 
R8084t3358 n8085 n3359 R=9.049e+00 
R8085t1450 n8086 n1451 R=4.913e+00 
R8085t3811 n8086 n3812 R=4.589e+00 
R8085t1092 n8086 n1093 R=1.139e+02 
R8085t3224 n8086 n3225 R=2.315e+01 
R8085t5699 n8086 n5700 R=4.259e+02 
R8086t436 n8087 n437 R=5.590e+01 
R8086t6296 n8087 n6297 R=3.940e+00 
R8086t3538 n8087 n3539 R=2.289e+01 
R8086t2346 n8087 n2347 R=4.868e+00 
R8086t117 n8087 n118 R=4.468e+00 
R8086t1180 n8087 n1181 R=1.245e+01 
R8086t4808 n8087 n4809 R=1.687e+02 
R8087t2779 n8088 n2780 R=8.019e+00 
R8087t3374 n8088 n3375 R=4.567e+00 
R8087t2086 n8088 n2087 R=8.741e+00 
R8087t5534 n8088 n5535 R=4.517e+00 
R8088t4260 n8089 n4261 R=1.079e+01 
R8088t899 n8089 n900 R=1.870e+01 
R8088t1888 n8089 n1889 R=1.052e+01 
R8088t4063 n8089 n4064 R=9.403e+00 
R8088t5384 n8089 n5385 R=4.419e+00 
R8089t375 n8090 n376 R=4.113e+01 
R8089t6133 n8090 n6134 R=7.325e+00 
R8089t686 n8090 n687 R=1.959e+01 
R8089t4477 n8090 n4478 R=3.645e+00 
R8089t6727 n8090 n6728 R=7.797e+00 
R8090t6769 n8091 n6770 R=1.226e+02 
R8090t6530 n8091 n6531 R=9.581e+00 
R8090t2849 n8091 n2850 R=4.492e+01 
R8090t7347 n8091 n7348 R=3.745e+00 
R8090t2013 n8091 n2014 R=9.983e+00 
R8090t6813 n8091 n6814 R=6.439e+00 
R8091t5313 n8092 n5314 R=9.561e+00 
R8091t7209 n8092 n7210 R=4.470e+00 
R8091t7441 n8092 n7442 R=4.639e+00 
R8091t7420 n8092 n7421 R=5.242e+00 
R8091t2352 n8092 n2353 R=1.770e+01 
R8092t465 n8093 n466 R=4.112e+00 
R8092t7885 n8093 n7886 R=2.377e+01 
R8092t3217 n8093 n3218 R=1.248e+02 
R8092t7378 n8093 n7379 R=7.171e+00 
R8092t6892 n8093 n6893 R=1.395e+01 
R8093t1015 n8094 n1016 R=5.232e+00 
R8093t4420 n8094 n4421 R=1.088e+01 
R8093t6968 n8094 n6969 R=1.185e+01 
R8093t4644 n8094 n4645 R=3.926e+00 
R8093t2662 n8094 n2663 R=1.482e+01 
R8093t304 n8094 n305 R=1.036e+01 
R8094t1009 n8095 n1010 R=4.324e+01 
R8094t7379 n8095 n7380 R=5.670e+00 
R8094t3832 n8095 n3833 R=2.466e+01 
R8094t5109 n8095 n5110 R=2.612e+01 
R8094t2910 n8095 n2911 R=9.517e+00 
R8095t3204 n8096 n3205 R=1.777e+02 
R8095t7463 n8096 n7464 R=1.547e+01 
R8095t2067 n8096 n2068 R=2.230e+00 
R8095t5113 n8096 n5114 R=8.136e+00 
R8095t1582 n8096 n1583 R=2.824e+00 
R8096t97 n8097 n98 R=1.044e+01 
R8096t3886 n8097 n3887 R=2.476e+00 
R8097t4139 n8098 n4140 R=1.532e+01 
R8097t5994 n8098 n5995 R=1.030e+01 
R8097t2606 n8098 n2607 R=2.528e+00 
R8098t6106 n8099 n6107 R=1.316e+01 
R8098t6981 n8099 n6982 R=9.116e+00 
R8098t6812 n8099 n6813 R=1.191e+01 
R8099t3562 n8100 n3563 R=1.563e+01 
R8099t7066 n8100 n7067 R=1.329e+01 
R8099t1230 n8100 n1231 R=1.242e+01 
R8099t5747 n8100 n5748 R=2.996e+00 
R8099t3518 n8100 n3519 R=4.585e+01 
R8100t5791 n8101 n5792 R=1.196e+01 
R8100t6795 n8101 n6796 R=4.647e+00 
R8100t6091 n8101 n6092 R=2.702e+00 
R8100t183 n8101 n184 R=1.342e+01 
R8101t6423 n8102 n6424 R=1.072e+02 
R8101t1295 n8102 n1296 R=2.750e+00 
R8101t786 n8102 n787 R=8.505e+01 
R8101t6387 n8102 n6388 R=5.264e+00 
R8101t5636 n8102 n5637 R=2.475e+00 
R8101t3768 n8102 n3769 R=2.119e+03 
R8102t1256 n8103 n1257 R=1.293e+02 
R8102t4614 n8103 n4615 R=5.316e+00 
R8102t3376 n8103 n3377 R=3.155e+02 
R8102t5177 n8103 n5178 R=4.447e+00 
R8102t1140 n8103 n1141 R=1.332e+01 
R8102t678 n8103 n679 R=1.140e+03 
R8102t1645 n8103 n1646 R=3.129e+00 
R8102t6642 n8103 n6643 R=2.696e+02 
R8103t4107 n8104 n4108 R=1.437e+01 
R8103t5684 n8104 n5685 R=1.534e+01 
R8103t410 n8104 n411 R=3.183e+01 
R8103t6024 n8104 n6025 R=4.597e+00 
R8103t5876 n8104 n5877 R=6.775e+00 
R8103t2015 n8104 n2016 R=5.906e+00 
R8104t5994 n8105 n5995 R=3.168e+01 
R8104t8097 n8105 n8098 R=1.098e+00 
R8104t2606 n8105 n2607 R=5.635e+01 
R8104t6341 n8105 n6342 R=8.649e+01 
R8104t7405 n8105 n7406 R=2.809e+00 
R8105t3218 n8106 n3219 R=1.946e+01 
R8105t5593 n8106 n5594 R=2.630e+00 
R8105t1323 n8106 n1324 R=1.886e+00 
R8105t6856 n8106 n6857 R=7.783e+01 
R8105t5189 n8106 n5190 R=5.848e+01 
R8105t6462 n8106 n6463 R=8.750e+00 
R8106t2248 n8107 n2249 R=5.566e+01 
R8106t6981 n8107 n6982 R=1.399e+01 
R8106t8098 n8107 n8099 R=3.141e+00 
R8106t1163 n8107 n1164 R=2.943e+00 
R8107t1879 n8108 n1880 R=1.446e+01 
R8107t4312 n8108 n4313 R=5.425e+00 
R8107t870 n8108 n871 R=4.805e+00 
R8107t3654 n8108 n3655 R=1.188e+01 
R8107t7182 n8108 n7183 R=6.691e+00 
R8107t1781 n8108 n1782 R=1.003e+01 
R8108t1465 n8109 n1466 R=9.002e+00 
R8108t4066 n8109 n4067 R=3.755e+00 
R8108t3708 n8109 n3709 R=2.582e+01 
R8108t682 n8109 n683 R=1.836e+00 
R8108t7531 n8109 n7532 R=4.741e+00 
R8109t989 n8110 n990 R=3.366e+02 
R8109t5140 n8110 n5141 R=9.756e+00 
R8109t6268 n8110 n6269 R=2.637e+01 
R8109t5301 n8110 n5302 R=3.624e+01 
R8109t2856 n8110 n2857 R=9.873e+00 
R8109t4802 n8110 n4803 R=4.893e+00 
R8109t1222 n8110 n1223 R=1.357e+01 
R8110t7667 n8111 n7668 R=1.255e+02 
R8110t2000 n8111 n2001 R=4.583e+00 
R8110t7408 n8111 n7409 R=3.503e+00 
R8110t7455 n8111 n7456 R=2.089e+01 
R8110t959 n8111 n960 R=2.163e+00 
R8111t128 n8112 n129 R=2.303e+01 
R8111t5181 n8112 n5182 R=1.142e+01 
R8111t4881 n8112 n4882 R=5.664e+00 
R8111t7482 n8112 n7483 R=2.867e+00 
R8112t7565 n8113 n7566 R=1.623e+01 
R8112t4210 n8113 n4211 R=4.756e+01 
R8112t2486 n8113 n2487 R=1.338e+01 
R8112t2703 n8113 n2704 R=2.243e+00 
R8113t1687 n8114 n1688 R=1.133e+02 
R8113t4436 n8114 n4437 R=2.026e+00 
R8113t866 n8114 n867 R=1.380e+01 
R8113t6929 n8114 n6930 R=1.348e+00 
R8113t2191 n8114 n2192 R=9.698e+00 
R8114t1090 n8115 n1091 R=1.003e+01 
R8114t4482 n8115 n4483 R=4.383e+01 
R8114t768 n8115 n769 R=2.695e+00 
R8114t2081 n8115 n2082 R=5.964e+00 
R8114t1967 n8115 n1968 R=1.518e+01 
R8115t4005 n8116 n4006 R=1.181e+01 
R8115t4429 n8116 n4430 R=9.101e+00 
R8115t8076 n8116 n8077 R=2.584e+00 
R8115t4863 n8116 n4864 R=3.397e+00 
R8116t1742 n8117 n1743 R=3.237e+01 
R8116t2778 n8117 n2779 R=8.674e+00 
R8116t6091 n8117 n6092 R=3.193e+01 
R8116t8100 n8117 n8101 R=6.477e+00 
R8116t6795 n8117 n6796 R=5.134e+01 
R8116t1317 n8117 n1318 R=3.052e+00 
R8116t4093 n8117 n4094 R=1.214e+01 
R8116t6578 n8117 n6579 R=2.040e+01 
R8117t655 n8118 n656 R=1.619e+00 
R8117t1675 n8118 n1676 R=3.560e+01 
R8117t7987 n8118 n7988 R=8.887e+00 
R8117t3326 n8118 n3327 R=4.710e+00 
R8117t6543 n8118 n6544 R=1.785e+01 
R8117t6313 n8118 n6314 R=1.259e+01 
R8118t3139 n8119 n3140 R=1.775e+02 
R8118t7508 n8119 n7509 R=4.040e+00 
R8118t4867 n8119 n4868 R=1.172e+01 
R8118t6525 n8119 n6526 R=2.025e+01 
R8118t6961 n8119 n6962 R=5.617e+00 
R8119t1032 n8120 n1033 R=6.698e+00 
R8119t3161 n8120 n3162 R=4.192e+00 
R8119t3703 n8120 n3704 R=3.618e+01 
R8119t2416 n8120 n2417 R=7.408e+00 
R8119t5210 n8120 n5211 R=4.737e+00 
R8119t3633 n8120 n3634 R=1.287e+02 
R8119t3882 n8120 n3883 R=2.418e+01 
R8119t4365 n8120 n4366 R=1.077e+01 
R8120t5996 n8121 n5997 R=3.000e+00 
R8120t7932 n8121 n7933 R=1.484e+01 
R8120t666 n8121 n667 R=2.318e+02 
R8120t850 n8121 n851 R=9.778e+00 
R8121t1182 n8122 n1183 R=2.159e+01 
R8121t2302 n8122 n2303 R=6.758e+00 
R8121t6305 n8122 n6306 R=1.678e+01 
R8121t7187 n8122 n7188 R=1.121e+01 
R8121t4271 n8122 n4272 R=1.171e+01 
R8121t1886 n8122 n1887 R=3.848e+01 
R8121t7121 n8122 n7122 R=8.804e+00 
R8122t7929 n8123 n7930 R=1.244e+01 
R8122t1403 n8123 n1404 R=5.322e+01 
R8122t2443 n8123 n2444 R=2.858e+01 
R8122t2991 n8123 n2992 R=4.958e+00 
R8122t2400 n8123 n2401 R=6.396e+00 
R8123t353 n8124 n354 R=1.275e+00 
R8123t2890 n8124 n2891 R=1.041e+01 
R8123t2426 n8124 n2427 R=2.145e+02 
R8123t7007 n8124 n7008 R=4.370e+00 
R8123t3690 n8124 n3691 R=1.408e+01 
R8123t3042 n8124 n3043 R=7.161e+01 
R8124t1093 n8125 n1094 R=2.378e+00 
R8124t3244 n8125 n3245 R=7.654e+00 
R8124t4577 n8125 n4578 R=2.428e+01 
R8124t6376 n8125 n6377 R=2.097e+00 
R8125t7278 n8126 n7279 R=1.404e+01 
R8125t6708 n8126 n6709 R=4.400e+00 
R8125t419 n8126 n420 R=1.266e+01 
R8125t7134 n8126 n7135 R=5.827e+00 
R8125t7311 n8126 n7312 R=1.378e+01 
R8125t7340 n8126 n7341 R=9.947e+00 
R8126t1913 n8127 n1914 R=2.976e+00 
R8126t8048 n8127 n8049 R=1.822e+01 
R8126t3377 n8127 n3378 R=2.313e+01 
R8126t2987 n8127 n2988 R=2.638e+01 
R8126t7096 n8127 n7097 R=9.438e+00 
R8126t1255 n8127 n1256 R=5.321e+00 
R8127t467 n8128 n468 R=2.182e+01 
R8127t3856 n8128 n3857 R=8.367e+00 
R8127t6650 n8128 n6651 R=6.761e+00 
R8127t7735 n8128 n7736 R=3.133e+00 
R8127t7547 n8128 n7548 R=5.037e+00 
R8127t1198 n8128 n1199 R=1.203e+02 
R8128t6309 n8129 n6310 R=2.087e+01 
R8128t7386 n8129 n7387 R=1.852e+00 
R8128t6095 n8129 n6096 R=2.400e+01 
R8128t6362 n8129 n6363 R=3.060e+00 
R8129t505 n8130 n506 R=1.096e+02 
R8129t539 n8130 n540 R=1.279e+01 
R8129t2169 n8130 n2170 R=9.779e+00 
R8129t5104 n8130 n5105 R=4.345e+01 
R8129t4080 n8130 n4081 R=7.855e+00 
R8129t1842 n8130 n1843 R=5.750e+00 
R8129t3843 n8130 n3844 R=1.382e+01 
R8130t1463 n8131 n1464 R=6.145e+01 
R8130t4825 n8131 n4826 R=2.764e+00 
R8130t7109 n8131 n7110 R=5.147e+00 
R8130t2001 n8131 n2002 R=6.593e+00 
R8131t5683 n8132 n5684 R=1.805e+01 
R8131t6634 n8132 n6635 R=5.781e+01 
R8131t1501 n8132 n1502 R=2.806e+00 
R8131t3030 n8132 n3031 R=1.305e+01 
R8131t5908 n8132 n5909 R=4.858e+00 
R8132t2843 n8133 n2844 R=1.578e+01 
R8132t7752 n8133 n7753 R=3.908e+02 
R8132t3369 n8133 n3370 R=2.599e+00 
R8132t853 n8133 n854 R=1.906e+01 
R8132t6840 n8133 n6841 R=1.196e+01 
R8133t1156 n8134 n1157 R=4.158e+00 
R8133t4488 n8134 n4489 R=1.131e+01 
R8133t6725 n8134 n6726 R=2.277e+01 
R8134t5812 n8135 n5813 R=6.849e+00 
R8134t7211 n8135 n7212 R=6.953e+00 
R8134t7074 n8135 n7075 R=4.799e+00 
R8134t7580 n8135 n7581 R=2.166e+01 
R8134t4902 n8135 n4903 R=9.384e+00 
R8135t989 n8136 n990 R=1.298e+01 
R8135t5140 n8136 n5141 R=7.098e+00 
R8135t6268 n8136 n6269 R=9.065e+00 
R8135t3225 n8136 n3226 R=2.655e+00 
R8135t1924 n8136 n1925 R=9.443e+00 
R8136t2648 n8137 n2649 R=1.315e+01 
R8136t7359 n8137 n7360 R=9.695e+00 
R8136t3448 n8137 n3449 R=1.573e+01 
R8136t4523 n8137 n4524 R=4.032e+00 
R8136t5662 n8137 n5663 R=5.065e+00 
R8137t1707 n8138 n1708 R=1.571e+01 
R8137t8037 n8138 n8038 R=6.679e+00 
R8137t3913 n8138 n3914 R=1.331e+01 
R8137t3908 n8138 n3909 R=1.098e+01 
R8137t4706 n8138 n4707 R=4.515e+00 
R8137t1137 n8138 n1138 R=2.322e+03 
R8138t1871 n8139 n1872 R=4.805e+00 
R8138t7719 n8139 n7720 R=7.015e+00 
R8138t1405 n8139 n1406 R=1.046e+01 
R8138t6261 n8139 n6262 R=3.218e+00 
R8139t331 n8140 n332 R=2.879e+01 
R8139t582 n8140 n583 R=4.909e+00 
R8139t75 n8140 n76 R=6.245e+00 
R8139t6413 n8140 n6414 R=2.826e+00 
R8140t2985 n8141 n2986 R=5.530e+00 
R8140t5444 n8141 n5445 R=6.562e+01 
R8140t7269 n8141 n7270 R=5.455e+00 
R8140t2005 n8141 n2006 R=4.583e+00 
R8140t1086 n8141 n1087 R=2.878e+01 
R8141t478 n8142 n479 R=8.609e+01 
R8141t7045 n8142 n7046 R=7.669e+01 
R8141t2213 n8142 n2214 R=4.653e+01 
R8141t1053 n8142 n1054 R=1.916e+00 
R8142t6240 n8143 n6241 R=6.748e+00 
R8142t7878 n8143 n7879 R=9.145e+00 
R8142t4756 n8143 n4757 R=1.904e+01 
R8142t3544 n8143 n3545 R=1.164e+01 
R8142t5258 n8143 n5259 R=3.528e+00 
R8143t4620 n8144 n4621 R=8.828e+00 
R8143t7928 n8144 n7929 R=1.036e+01 
R8143t2829 n8144 n2830 R=4.599e+01 
R8143t4671 n8144 n4672 R=4.012e+00 
R8144t2182 n8145 n2183 R=2.907e+02 
R8144t2235 n8145 n2236 R=3.075e+00 
R8144t3147 n8145 n3148 R=1.688e+01 
R8144t1054 n8145 n1055 R=1.267e+01 
R8144t4835 n8145 n4836 R=3.417e+01 
R8145t1534 n8146 n1535 R=3.093e+00 
R8145t7495 n8146 n7496 R=1.104e+01 
R8145t3205 n8146 n3206 R=1.526e+01 
R8145t3316 n8146 n3317 R=6.474e+00 
R8146t7624 n8147 n7625 R=9.224e+00 
R8146t4740 n8147 n4741 R=4.357e+01 
R8146t4782 n8147 n4783 R=2.636e+00 
R8146t1651 n8147 n1652 R=1.176e+01 
R8146t440 n8147 n441 R=2.197e+01 
R8147t2374 n8148 n2375 R=6.384e+00 
R8147t7234 n8148 n7235 R=8.837e+00 
R8147t6746 n8148 n6747 R=9.790e+01 
R8147t7802 n8148 n7803 R=1.791e+01 
R8147t6993 n8148 n6994 R=4.364e+00 
R8147t43 n8148 n44 R=4.362e+01 
R8147t4574 n8148 n4575 R=7.151e+00 
R8148t3379 n8149 n3380 R=5.812e+00 
R8148t5394 n8149 n5395 R=1.781e+01 
R8148t1885 n8149 n1886 R=3.312e+00 
R8148t5769 n8149 n5770 R=5.816e+00 
R8149t7216 n8150 n7217 R=7.934e+01 
R8149t7543 n8150 n7544 R=6.563e+00 
R8149t5921 n8150 n5922 R=3.077e+00 
R8149t6255 n8150 n6256 R=1.168e+01 
R8149t7855 n8150 n7856 R=4.632e+00 
R8150t1072 n8151 n1073 R=3.023e+01 
R8150t8022 n8151 n8023 R=9.021e+00 
R8150t16 n8151 n17 R=2.345e+00 
R8150t3371 n8151 n3372 R=1.376e+01 
R8150t3278 n8151 n3279 R=7.037e+00 
R8150t7440 n8151 n7441 R=1.141e+01 
R8151t2555 n8152 n2556 R=8.734e+00 
R8151t4473 n8152 n4474 R=2.667e+00 
R8151t3852 n8152 n3853 R=7.575e+00 
R8151t8065 n8152 n8066 R=5.009e+00 
R8152t1939 n8153 n1940 R=4.661e+00 
R8152t5305 n8153 n5306 R=9.988e+00 
R8152t2873 n8153 n2874 R=3.620e+01 
R8152t127 n8153 n128 R=6.307e+00 
R8152t2462 n8153 n2463 R=8.328e+00 
R8152t5426 n8153 n5427 R=1.644e+01 
R8152t7182 n8153 n7183 R=2.352e+01 
R8152t8107 n8153 n8108 R=1.541e+01 
R8152t3654 n8153 n3655 R=5.651e+01 
R8153t129 n8154 n130 R=3.899e+00 
R8153t4680 n8154 n4681 R=4.844e+00 
R8153t4003 n8154 n4004 R=3.128e+01 
R8153t5166 n8154 n5167 R=1.476e+01 
R8154t6694 n8155 n6695 R=4.976e+00 
R8154t7921 n8155 n7922 R=3.737e+00 
R8154t6273 n8155 n6274 R=8.247e+00 
R8154t3536 n8155 n3537 R=8.237e+00 
R8154t6729 n8155 n6730 R=1.072e+01 
R8154t7373 n8155 n7374 R=7.157e+01 
R8155t578 n8156 n579 R=1.654e+01 
R8155t707 n8156 n708 R=1.349e+01 
R8155t967 n8156 n968 R=1.040e+01 
R8155t7609 n8156 n7610 R=1.420e+01 
R8156t1507 n8157 n1508 R=2.784e+01 
R8156t4732 n8157 n4733 R=1.738e+01 
R8156t3465 n8157 n3466 R=2.450e+02 
R8156t2713 n8157 n2714 R=1.654e+01 
R8156t6606 n8157 n6607 R=2.348e+00 
R8157t4216 n8158 n4217 R=5.233e+00 
R8157t7219 n8158 n7220 R=1.033e+01 
R8157t562 n8158 n563 R=5.093e+00 
R8157t7201 n8158 n7202 R=2.459e+00 
R8158t3776 n8159 n3777 R=2.319e+01 
R8158t6647 n8159 n6648 R=1.717e+01 
R8158t6902 n8159 n6903 R=4.941e+00 
R8159t1133 n8160 n1134 R=3.078e+00 
R8159t7221 n8160 n7222 R=2.249e+01 
R8159t3881 n8160 n3882 R=3.646e+00 
R8159t2487 n8160 n2488 R=3.426e+01 
R8159t5660 n8160 n5661 R=2.335e+00 
R8159t7534 n8160 n7535 R=2.033e+02 
R8160t1531 n8161 n1532 R=2.491e+00 
R8160t7377 n8161 n7378 R=8.510e+00 
R8160t6661 n8161 n6662 R=1.892e+01 
R8160t2323 n8161 n2324 R=5.456e+00 
R8160t6164 n8161 n6165 R=8.456e+00 
R8161t3272 n8162 n3273 R=4.983e+02 
R8161t3838 n8162 n3839 R=3.170e+00 
R8161t1009 n8162 n1010 R=2.302e+01 
R8161t1632 n8162 n1633 R=1.642e+01 
R8161t2350 n8162 n2351 R=3.842e+00 
R8161t7 n8162 n8 R=1.047e+01 
R8161t3490 n8162 n3491 R=5.765e+00 
R8162t5073 n8163 n5074 R=1.313e+02 
R8162t6076 n8163 n6077 R=1.242e+00 
R8162t5887 n8163 n5888 R=2.860e+00 
R8162t3239 n8163 n3240 R=9.626e+00 
R8163t604 n8164 n605 R=4.295e+02 
R8163t7201 n8164 n7202 R=2.146e+02 
R8163t8157 n8164 n8158 R=1.745e+01 
R8163t562 n8164 n563 R=3.323e+00 
R8163t937 n8164 n938 R=7.359e+00 
R8163t7067 n8164 n7068 R=3.768e+00 
R8164t1005 n8165 n1006 R=8.283e+01 
R8164t5394 n8165 n5395 R=4.216e+00 
R8164t7501 n8165 n7502 R=5.816e+00 
R8164t7974 n8165 n7975 R=5.202e+01 
R8164t1785 n8165 n1786 R=8.424e+00 
R8165t3549 n8166 n3550 R=5.326e+01 
R8165t3122 n8166 n3123 R=7.926e+00 
R8165t4689 n8166 n4690 R=7.576e+00 
R8166t2633 n8167 n2634 R=4.465e+00 
R8166t7776 n8167 n7777 R=6.747e+00 
R8166t6868 n8167 n6869 R=6.001e+00 
R8166t4047 n8167 n4048 R=1.588e+01 
R8167t722 n8168 n723 R=2.742e+00 
R8167t2305 n8168 n2306 R=3.124e+00 
R8168t1660 n8169 n1661 R=3.533e+00 
R8168t7569 n8169 n7570 R=2.497e+00 
R8168t5674 n8169 n5675 R=4.802e+01 
R8168t2018 n8169 n2019 R=2.816e+01 
R8168t6901 n8169 n6902 R=7.153e+00 
R8169t3499 n8170 n3500 R=6.134e+00 
R8169t3810 n8170 n3811 R=5.076e+00 
R8169t1802 n8170 n1803 R=1.429e+01 
R8169t1932 n8170 n1933 R=4.361e+00 
R8169t3598 n8170 n3599 R=9.212e+00 
R8169t7980 n8170 n7981 R=4.571e+01 
R8170t44 n8171 n45 R=1.573e+01 
R8170t5818 n8171 n5819 R=6.611e+00 
R8170t7914 n8171 n7915 R=6.666e+00 
R8170t6998 n8171 n6999 R=7.904e+00 
R8171t3046 n8172 n3047 R=7.573e+00 
R8171t5342 n8172 n5343 R=4.537e+02 
R8171t3815 n8172 n3816 R=3.693e+00 
R8171t3761 n8172 n3762 R=1.012e+01 
R8172t8098 n8173 n8099 R=2.133e+02 
R8172t8106 n8173 n8107 R=4.692e+00 
R8172t1163 n8173 n1164 R=1.956e+01 
R8172t2306 n8173 n2307 R=6.407e+00 
R8172t5152 n8173 n5153 R=8.244e+01 
R8172t7602 n8173 n7603 R=1.928e+01 
R8172t1748 n8173 n1749 R=6.999e+00 
R8172t6812 n8173 n6813 R=1.245e+01 
R8173t6409 n8174 n6410 R=1.991e+00 
R8173t4479 n8174 n4480 R=7.839e+00 
R8173t4508 n8174 n4509 R=1.449e+01 
R8173t615 n8174 n616 R=3.092e+00 
R8174t381 n8175 n382 R=1.593e+01 
R8174t4968 n8175 n4969 R=5.322e+01 
R8174t5816 n8175 n5817 R=4.479e+00 
R8174t157 n8175 n158 R=5.133e+00 
R8174t6767 n8175 n6768 R=1.589e+00 
R8175t270 n8176 n271 R=1.118e+01 
R8175t1089 n8176 n1090 R=4.921e+01 
R8175t7038 n8176 n7039 R=4.383e+00 
R8175t4033 n8176 n4034 R=2.102e+01 
R8175t5443 n8176 n5444 R=5.503e+00 
R8176t6072 n8177 n6073 R=1.998e+02 
R8176t7586 n8177 n7587 R=6.139e+00 
R8176t1266 n8177 n1267 R=6.225e+00 
R8176t7617 n8177 n7618 R=8.669e+00 
R8176t6301 n8177 n6302 R=4.782e+00 
R8176t597 n8177 n598 R=8.765e+00 
R8177t1725 n8178 n1726 R=1.974e+01 
R8177t3785 n8178 n3786 R=1.049e+01 
R8177t1700 n8178 n1701 R=2.975e+00 
R8177t1840 n8178 n1841 R=8.851e+00 
R8177t82 n8178 n83 R=4.989e+00 
R8178t2451 n8179 n2452 R=3.893e+00 
R8178t6976 n8179 n6977 R=7.700e+02 
R8178t3306 n8179 n3307 R=1.332e+00 
R8178t7507 n8179 n7508 R=3.082e+01 
R8178t7683 n8179 n7684 R=2.251e+01 
R8179t10 n8180 n11 R=8.551e+00 
R8179t489 n8180 n490 R=2.148e+01 
R8179t5250 n8180 n5251 R=1.844e+01 
R8179t6825 n8180 n6826 R=6.651e+00 
R8179t4152 n8180 n4153 R=2.005e+01 
R8179t2524 n8180 n2525 R=4.676e+00 
R8180t5953 n8181 n5954 R=1.607e+01 
R8180t6781 n8181 n6782 R=8.480e+00 
R8180t5859 n8181 n5860 R=2.273e+01 
R8180t2886 n8181 n2887 R=1.923e+01 
R8180t7277 n8181 n7278 R=6.150e+00 
R8180t3675 n8181 n3676 R=3.140e+01 
R8181t5083 n8182 n5084 R=7.276e+00 
R8181t5491 n8182 n5492 R=1.659e+01 
R8181t1934 n8182 n1935 R=1.051e+01 
R8181t6356 n8182 n6357 R=5.403e+00 
R8181t3210 n8182 n3211 R=2.303e+01 
R8181t2220 n8182 n2221 R=4.827e+01 
R8181t570 n8182 n571 R=3.331e+01 
R8182t1193 n8183 n1194 R=1.518e+01 
R8182t5657 n8183 n5658 R=5.848e+00 
R8182t3420 n8183 n3421 R=6.708e+00 
R8182t6516 n8183 n6517 R=6.998e+00 
R8183t1624 n8184 n1625 R=1.100e+01 
R8183t5052 n8184 n5053 R=6.459e+00 
R8183t2854 n8184 n2855 R=4.321e+00 
R8183t7519 n8184 n7520 R=5.323e+00 
R8183t5881 n8184 n5882 R=1.534e+01 
R8184t2829 n8185 n2830 R=7.147e+00 
R8184t4589 n8185 n4590 R=5.588e+00 
R8184t7928 n8185 n7929 R=3.267e+00 
R8184t7196 n8185 n7197 R=7.199e+00 
R8185t5192 n8186 n5193 R=3.669e+00 
R8185t6124 n8186 n6125 R=1.001e+01 
R8185t2885 n8186 n2886 R=3.610e+01 
R8186t4653 n8187 n4654 R=3.597e+00 
R8186t6937 n8187 n6938 R=6.929e+00 
R8186t5198 n8187 n5199 R=2.318e+00 
R8186t2349 n8187 n2350 R=2.863e+01 
R8187t1779 n8188 n1 R=1.515e+01 
R8187t6966 n8188 n1 R=1.547e+01 
R8187t2095 n8188 n2096 R=5.098e+00 
R8187t2767 n8188 n2768 R=8.820e+00 
R8187t5951 n8188 n5952 R=9.171e+00 
R8187t2727 n8188 n2728 R=3.839e+00 
R8188t5057 n8189 n5058 R=5.653e+00 
R8188t3766 n8189 n3767 R=5.776e+00 
R8188t6140 n8189 n6141 R=8.096e+00 
R8188t5240 n8189 n5241 R=5.169e+00 
R8189t3440 n8190 n3441 R=2.448e+00 
R8189t4908 n8190 n4909 R=6.064e+01 
R8189t789 n8190 n790 R=4.080e+00 
R8189t3673 n8190 n3674 R=5.706e+00 
R8189t6659 n8190 n6660 R=1.412e+01 
R8190t59 n8191 n60 R=9.401e+00 
R8190t6261 n8191 n6262 R=2.219e+02 
R8190t6087 n8191 n6088 R=2.686e+01 
R8190t67 n8191 n68 R=2.885e+00 
R8190t5811 n8191 n5812 R=3.016e+01 
R8190t2452 n8191 n2453 R=3.809e+00 
R8191t927 n8192 n928 R=6.761e+00 
R8191t1658 n8192 n1659 R=1.082e+02 
R8191t8079 n8192 n8080 R=3.135e+00 
R8191t5053 n8192 n5054 R=4.672e+01 
R8191t7497 n8192 n7498 R=1.478e+01 
R8191t288 n8192 n289 R=9.029e+00 
R8192t1398 n8193 n1399 R=2.337e+00 
R8192t7170 n8193 n7171 R=3.056e+00 
R8192t3374 n8193 n3375 R=1.138e+01 
R8192t4516 n8193 n4517 R=1.634e+01 
R8193t5477 n8194 n5478 R=1.550e+01 
R8193t4058 n8194 n4059 R=4.032e+01 
R8193t3159 n8194 n3160 R=9.489e+00 
R8193t5906 n8194 n5907 R=5.736e+00 
R8193t3180 n8194 n3181 R=8.991e+00 
R8194t4094 n8195 n4095 R=4.020e+00 
R8194t5915 n8195 n5916 R=3.740e+00 
R8194t5039 n8195 n5040 R=3.715e+01 
R8194t531 n8195 n532 R=3.364e+00 
R8194t941 n8195 n942 R=5.606e+02 
R8195t394 n8196 n395 R=4.586e+00 
R8195t4092 n8196 n4093 R=4.095e+00 
R8195t2054 n8196 n2055 R=2.308e+01 
R8195t1293 n8196 n1294 R=2.370e+01 
R8195t7849 n8196 n7850 R=7.014e+00 
R8195t1743 n8196 n1744 R=7.067e+02 
R8195t3022 n8196 n3023 R=7.709e+00 
R8196t4193 n8197 n4194 R=2.881e+00 
R8196t4236 n8197 n4237 R=1.476e+01 
R8196t2471 n8197 n2472 R=1.181e+01 
R8197t8142 n8198 n8143 R=1.603e+02 
R8197t7027 n8198 n7028 R=9.361e+00 
R8197t7473 n8198 n7474 R=9.494e+00 
R8197t830 n8198 n831 R=3.832e+00 
R8197t5258 n8198 n5259 R=1.331e+01 
R8198t5366 n8199 n5367 R=9.125e+00 
R8198t6869 n8199 n6870 R=3.349e+00 
R8198t7477 n8199 n7478 R=9.034e+00 
R8198t2738 n8199 n2739 R=1.262e+01 
R8198t4157 n8199 n4158 R=4.943e+00 
R8198t5048 n8199 n5049 R=5.327e+02 
R8199t578 n8200 n579 R=1.715e+02 
R8199t8155 n8200 n8156 R=6.821e+00 
R8199t707 n8200 n708 R=3.160e+00 
R8199t6262 n8200 n6263 R=6.895e+00 
R8199t1879 n8200 n1880 R=1.064e+01 
R8200t1931 n8201 n1932 R=6.488e+00 
R8200t4733 n8201 n4734 R=4.252e+00 
R8200t4115 n8201 n4116 R=2.408e+01 
R8201t4802 n8202 n4803 R=2.751e+01 
R8201t1222 n8202 n1223 R=4.145e+00 
R8201t5884 n8202 n5885 R=4.108e+01 
R8201t2763 n8202 n2764 R=7.369e+00 
R8201t2632 n8202 n2633 R=4.491e+01 
R8201t4206 n8202 n4207 R=2.437e+01 
R8202t6597 n8203 n6598 R=5.005e+00 
R8202t5285 n8203 n5286 R=2.331e+02 
R8202t2180 n8203 n2181 R=1.836e+01 
R8202t5754 n8203 n5755 R=1.398e+01 
R8202t5996 n8203 n5997 R=1.632e+01 
R8202t8120 n8203 n8121 R=2.001e+01 
R8203t1854 n8204 n1855 R=4.533e+00 
R8203t6186 n8204 n6187 R=5.564e+00 
R8203t6596 n8204 n6597 R=3.805e+01 
R8203t3230 n8204 n3231 R=3.776e+01 
R8203t6909 n8204 n6910 R=4.396e+00 
R8203t7258 n8204 n7259 R=8.252e+00 
R8204t114 n8205 n115 R=2.415e+01 
R8204t1931 n8205 n1932 R=8.523e+01 
R8204t3734 n8205 n3735 R=1.612e+01 
R8204t918 n8205 n919 R=2.405e+00 
R8204t4115 n8205 n4116 R=2.225e+01 
R8204t8200 n8205 n8201 R=2.040e+00 
R8205t5457 n8206 n5458 R=1.846e+01 
R8205t5836 n8206 n5837 R=1.885e+00 
R8205t24 n8206 n25 R=1.688e+01 
R8205t6571 n8206 n6572 R=3.500e+00 
R8205t135 n8206 n136 R=9.679e+00 
R8206t3000 n8207 n3001 R=4.266e+01 
R8206t3560 n8207 n3561 R=7.011e+00 
R8206t831 n8207 n832 R=6.505e+00 
R8206t7318 n8207 n7319 R=2.426e+01 
R8206t4366 n8207 n4367 R=2.714e+00 
R8206t5069 n8207 n5070 R=7.626e+01 
R8206t6272 n8207 n6273 R=1.009e+02 
R8206t3526 n8207 n3527 R=7.145e+00 
R8207t5509 n8208 n5510 R=3.362e+00 
R8207t6963 n8208 n6964 R=7.770e+01 
R8207t8054 n8208 n8055 R=4.111e+02 
R8207t723 n8208 n724 R=7.132e+00 
R8207t3835 n8208 n3836 R=7.132e+00 
R8207t6020 n8208 n6021 R=1.335e+01 
R8208t298 n8209 n299 R=4.138e+00 
R8208t6418 n8209 n6419 R=5.479e+01 
R8208t2824 n8209 n2825 R=5.056e+00 
R8208t159 n8209 n160 R=6.652e+02 
R8208t4738 n8209 n4739 R=9.373e+00 
R8208t6824 n8209 n6825 R=8.716e+00 
R8209t548 n8210 n549 R=2.990e+00 
R8209t5080 n8210 n5081 R=4.189e+00 
R8209t2843 n8210 n2844 R=1.278e+02 
R8209t5458 n8210 n5459 R=2.929e+00 
R8209t6408 n8210 n6409 R=8.229e+01 
R8210t2135 n8211 n2136 R=1.406e+01 
R8210t8001 n8211 n8002 R=6.668e+00 
R8210t7765 n8211 n7766 R=5.316e+00 
R8210t7129 n8211 n7130 R=2.430e+01 
R8210t1257 n8211 n1258 R=1.152e+01 
R8210t2910 n8211 n2911 R=4.350e+00 
R8211t608 n8212 n609 R=7.130e+00 
R8211t2865 n8212 n2866 R=2.908e+01 
R8211t6831 n8212 n6832 R=8.734e+01 
R8211t3092 n8212 n3093 R=5.698e+00 
R8212t598 n8213 n599 R=2.867e+00 
R8212t5174 n8213 n5175 R=4.705e+01 
R8212t7784 n8213 n7785 R=5.045e+00 
R8212t635 n8213 n636 R=3.349e+00 
R8213t899 n8214 n900 R=1.964e+01 
R8213t6418 n8214 n6419 R=7.660e+00 
R8213t2824 n8214 n2825 R=8.706e+00 
R8213t2313 n8214 n2314 R=8.016e+00 
R8213t3140 n8214 n3141 R=4.670e+00 
R8214t2252 n8215 n2253 R=1.076e+01 
R8214t6744 n8215 n6745 R=9.588e+00 
R8214t6017 n8215 n6018 R=1.213e+01 
R8214t3273 n8215 n3274 R=1.904e+01 
R8214t7391 n8215 n7392 R=1.374e+01 
R8215t6597 n8216 n6598 R=8.705e+00 
R8215t8202 n8216 n8203 R=1.511e+01 
R8215t7612 n8216 n7613 R=2.014e+01 
R8215t7486 n8216 n7487 R=4.645e+01 
R8215t2504 n8216 n2505 R=1.151e+02 
R8216t2676 n8217 n2677 R=7.063e+00 
R8216t6377 n8217 n6378 R=2.083e+00 
R8216t240 n8217 n241 R=7.236e+00 
R8217t6934 n8218 n6935 R=2.738e+00 
R8217t7942 n8218 n7943 R=1.804e+02 
R8217t5359 n8218 n5360 R=9.005e+00 
R8217t3572 n8218 n3573 R=2.224e+00 
R8218t3147 n8219 n3148 R=4.617e+00 
R8218t8144 n8219 n8145 R=1.384e+01 
R8218t7778 n8219 n7779 R=1.057e+01 
R8218t3826 n8219 n3827 R=4.891e+00 
R8218t2235 n8219 n2236 R=1.850e+01 
R8219t4261 n8220 n4262 R=3.097e+02 
R8219t5563 n8220 n5564 R=4.023e+00 
R8219t3557 n8220 n3558 R=4.682e+00 
R8220t6000 n8221 n6001 R=2.543e+01 
R8220t6476 n8221 n6477 R=6.000e+00 
R8220t6605 n8221 n6606 R=1.042e+01 
R8220t7324 n8221 n7325 R=2.724e+00 
R8220t914 n8221 n915 R=1.082e+01 
R8220t6525 n8221 n6526 R=3.764e+01 
R8221t4174 n8222 n4175 R=6.228e+00 
R8221t7370 n8222 n7371 R=1.228e+01 
R8221t7866 n8222 n7867 R=6.546e+00 
R8221t2677 n8222 n2678 R=8.803e+00 
R8221t3758 n8222 n3759 R=5.567e+00 
R8222t2033 n8223 n2034 R=2.285e+00 
R8222t5607 n8223 n5608 R=1.040e+01 
R8222t2870 n8223 n2871 R=9.084e+00 
R8222t2142 n8223 n2143 R=5.464e+01 
R8222t5549 n8223 n5550 R=6.398e+00 
R8222t1962 n8223 n1963 R=2.038e+01 
R8223t5106 n8224 n5107 R=3.076e+00 
R8223t5470 n8224 n5471 R=9.963e+00 
R8223t775 n8224 n776 R=1.881e+02 
R8223t7156 n8224 n7157 R=3.327e+00 
R8224t4345 n8225 n4346 R=3.771e+02 
R8224t2357 n8225 n2358 R=5.312e+00 
R8224t1467 n8225 n1468 R=1.515e+01 
R8224t1002 n8225 n1003 R=3.295e+00 
R8225t4232 n8226 n4233 R=1.823e+00 
R8225t478 n8226 n479 R=7.888e+00 
R8225t8141 n8226 n8142 R=1.243e+00 
R8226t1376 n8227 n1377 R=1.812e+01 
R8226t4919 n8227 n1 R=3.591e+01 
R8226t2859 n8227 n2860 R=1.492e+01 
R8226t4480 n8227 n4481 R=1.164e+01 
R8226t5613 n8227 n5614 R=3.283e+00 
R8226t6174 n8227 n1 R=2.867e+00 
R8227t3810 n8228 n3811 R=7.599e+00 
R8227t7992 n8228 n7993 R=9.085e+00 
R8227t4846 n8228 n4847 R=4.158e+00 
R8227t5621 n8228 n5622 R=5.174e+01 
R8227t7585 n8228 n7586 R=6.975e+00 
R8228t374 n8229 n375 R=1.309e+01 
R8228t6818 n8229 n6819 R=6.509e+00 
R8228t2490 n8229 n2491 R=8.726e+00 
R8228t5343 n8229 n5344 R=4.634e+00 
R8228t7818 n8229 n7819 R=8.281e+00 
R8228t6501 n8229 n6502 R=1.246e+02 
R8229t6265 n8230 n6266 R=9.700e+00 
R8229t5926 n8230 n5927 R=8.560e+00 
R8229t7535 n8230 n7536 R=2.063e+00 
R8229t1735 n8230 n1736 R=2.729e+01 
R8230t5271 n8231 n5272 R=2.444e+01 
R8230t1421 n8231 n1422 R=2.785e+01 
R8230t5163 n8231 n5164 R=4.827e+00 
R8230t761 n8231 n762 R=8.432e+00 
R8230t3006 n8231 n3007 R=1.078e+01 
R8231t3202 n8232 n3203 R=2.377e+01 
R8231t7433 n8232 n7434 R=3.703e+00 
R8231t4045 n8232 n4046 R=4.732e+00 
R8231t6984 n8232 n6985 R=3.291e+00 
R8231t4301 n8232 n4302 R=3.170e+01 
R8232t1230 n8233 n1231 R=4.039e+02 
R8232t3562 n8233 n3563 R=8.233e+00 
R8232t8099 n8233 n8100 R=2.108e+00 
R8233t3121 n8234 n3122 R=5.311e+00 
R8233t6350 n8234 n6351 R=6.286e+00 
R8233t6670 n8234 n6671 R=6.281e+00 
R8233t7770 n8234 n7771 R=3.122e+01 
R8233t5971 n8234 n5972 R=6.217e+00 
R8233t5979 n8234 n5980 R=1.067e+01 
R8234t2987 n8235 n2988 R=3.609e+00 
R8234t3377 n8235 n3378 R=1.060e+01 
R8234t8126 n8235 n8127 R=9.727e+00 
R8235t2815 n8236 n2816 R=6.782e+00 
R8235t6598 n8236 n6599 R=8.213e+00 
R8235t2580 n8236 n2581 R=1.576e+01 
R8235t345 n8236 n346 R=8.075e+00 
R8235t1288 n8236 n1289 R=5.719e+00 
R8236t5633 n8237 n5634 R=9.049e+00 
R8236t8041 n8237 n8042 R=4.517e+01 
R8236t5292 n8237 n5293 R=6.096e+00 
R8236t7846 n8237 n7847 R=3.787e+00 
R8236t2904 n8237 n2905 R=2.079e+01 
R8236t6856 n8237 n6857 R=5.551e+00 
R8237t3183 n8238 n3184 R=1.963e+00 
R8237t7990 n8238 n7991 R=4.882e+01 
R8237t2317 n8238 n2318 R=9.540e+00 
R8237t6962 n8238 n6963 R=4.446e+00 
R8237t6794 n8238 n6795 R=2.984e+02 
R8237t1219 n8238 n1220 R=5.846e+00 
R8238t6738 n8239 n6739 R=6.330e+01 
R8238t27 n8239 n28 R=3.670e+00 
R8238t5036 n8239 n5037 R=6.660e+00 
R8239t6018 n8240 n6019 R=2.719e+01 
R8239t3338 n8240 n3339 R=5.684e+01 
R8239t7798 n8240 n7799 R=4.754e+00 
R8239t3867 n8240 n3868 R=9.339e+00 
R8240t544 n8241 n545 R=1.218e+01 
R8240t7588 n8241 n7589 R=1.201e+01 
R8240t2888 n8241 n2889 R=7.295e+01 
R8240t7371 n8241 n7372 R=4.036e+00 
R8240t4630 n8241 n4631 R=9.084e+00 
R8240t7102 n8241 n7103 R=7.825e+00 
R8241t2787 n8242 n2788 R=2.796e+01 
R8241t7739 n8242 n7740 R=1.513e+01 
R8241t825 n8242 n826 R=1.080e+01 
R8241t3369 n8242 n3370 R=1.029e+01 
R8241t7752 n8242 n7753 R=5.633e+00 
R8241t3138 n8242 n3139 R=9.471e+00 
R8241t7180 n8242 n7181 R=3.811e+00 
R8242t2008 n8243 n2009 R=2.398e+01 
R8242t7106 n8243 n7107 R=4.907e+01 
R8242t5744 n8243 n5745 R=1.707e+00 
R8242t6515 n8243 n6516 R=1.372e+01 
R8242t6061 n8243 n6062 R=2.484e+00 
R8243t3110 n8244 n3111 R=2.635e+00 
R8243t7658 n8244 n7659 R=6.358e+00 
R8243t2534 n8244 n2535 R=7.646e+01 
R8243t103 n8244 n104 R=2.455e+00 
R8243t5865 n8244 n5866 R=1.194e+01 
R8243t3714 n8244 n3715 R=4.179e+01 
R8244t5352 n8245 n5353 R=2.594e+01 
R8244t5898 n8245 n5899 R=1.850e+01 
R8244t5070 n8245 n5071 R=5.224e+00 
R8244t5838 n8245 n5839 R=6.338e+00 
R8244t7145 n8245 n7146 R=6.165e+01 
R8244t1156 n8245 n1157 R=5.521e+00 
R8244t8133 n8245 n8134 R=6.618e+00 
R8244t6725 n8245 n6726 R=1.933e+01 
R8245t352 n8246 n353 R=2.728e+00 
R8245t1301 n8246 n1302 R=8.424e+00 
R8245t1476 n8246 n1477 R=4.326e+01 
R8245t3926 n8246 n3927 R=2.717e+00 
R8245t3897 n8246 n3898 R=1.641e+02 
R8245t7794 n8246 n7795 R=2.048e+02 
R8245t5897 n8246 n5898 R=6.990e+01 
R8246t6336 n8247 n6337 R=4.223e+00 
R8246t7845 n8247 n7846 R=1.950e+01 
R8246t6126 n8247 n6127 R=2.629e+01 
R8246t560 n8247 n561 R=3.964e+00 
R8246t6764 n8247 n6765 R=9.211e+00 
R8247t3243 n8248 n3244 R=7.516e+00 
R8247t4899 n8248 n4900 R=4.331e+00 
R8247t2716 n8248 n2717 R=1.738e+01 
R8247t431 n8248 n432 R=2.652e+00 
R8248t857 n8249 n858 R=7.977e+00 
R8248t6737 n8249 n6738 R=2.725e+01 
R8248t3785 n8249 n3786 R=8.387e+00 
R8248t737 n8249 n738 R=9.957e+00 
R8248t969 n8249 n970 R=1.289e+01 
R8248t2447 n8249 n2448 R=7.780e+01 
R8248t5121 n8249 n5122 R=4.123e+00 
R8248t5536 n8249 n5537 R=1.386e+02 
R8248t1231 n8249 n1232 R=5.898e+01 
R8249t5770 n8250 n5771 R=2.262e+01 
R8249t7556 n8250 n7557 R=4.399e+00 
R8249t1690 n8250 n1691 R=3.042e+00 
R8249t7599 n8250 n7600 R=1.626e+01 
R8249t150 n8250 n151 R=6.029e+00 
R8250t7461 n8251 n7462 R=3.128e+01 
R8250t710 n8251 n711 R=5.266e+00 
R8250t4687 n8251 n4688 R=8.556e+00 
R8250t150 n8251 n151 R=5.067e+00 
R8250t7599 n8251 n7600 R=1.448e+01 
R8250t3446 n8251 n3447 R=3.870e+00 
R8251t4819 n8252 n4820 R=1.901e+00 
R8251t7064 n8252 n7065 R=3.276e+01 
R8251t1587 n8252 n1588 R=6.402e+00 
R8251t1981 n8252 n1982 R=2.380e+00 
R8252t209 n8253 n210 R=1.628e+01 
R8252t843 n8253 n844 R=6.925e+00 
R8252t2986 n8253 n2987 R=7.208e+00 
R8253t6425 n8254 n6426 R=4.256e+00 
R8253t5414 n8254 n5415 R=2.938e+00 
R8253t1747 n8254 n1748 R=2.551e+01 
R8253t3615 n8254 n3616 R=1.443e+01 
R8254t1178 n8255 n1179 R=2.023e+00 
R8254t4195 n8255 n4196 R=3.612e+00 
R8254t1227 n8255 n1228 R=9.710e+00 
R8254t2074 n8255 n2075 R=1.345e+01 
R8255t5212 n8256 n5213 R=9.652e+00 
R8255t5669 n8256 n5670 R=3.292e+00 
R8255t1711 n8256 n1712 R=4.311e+01 
R8255t3922 n8256 n3923 R=4.913e+00 
R8255t672 n8256 n673 R=7.247e+00 
R8256t6877 n8257 n6878 R=1.650e+01 
R8256t7461 n8257 n7462 R=5.153e+01 
R8256t1226 n8257 n1227 R=3.602e+00 
R8256t705 n8257 n706 R=2.016e+01 
R8256t3964 n8257 n3965 R=3.454e+00 
R8256t5628 n8257 n5629 R=4.329e+00 
R8257t6910 n8258 n6911 R=1.481e+01 
R8257t7818 n8258 n7819 R=1.606e+02 
R8257t7312 n8258 n7313 R=8.220e+00 
R8257t913 n8258 n914 R=6.441e+00 
R8257t5114 n8258 n5115 R=6.202e+00 
R8257t6501 n8258 n6502 R=2.271e+00 
R8258t2649 n8259 n2650 R=8.486e+00 
R8258t7695 n8259 n7696 R=8.531e+00 
R8258t684 n8259 n685 R=3.820e+00 
R8259t4053 n8260 n4054 R=1.363e+01 
R8259t5403 n8260 n5404 R=2.580e+01 
R8259t841 n8260 n842 R=1.382e+01 
R8259t2368 n8260 n2369 R=5.480e+00 
R8259t6633 n8260 n6634 R=1.226e+01 
R8259t5592 n8260 n5593 R=1.005e+01 
R8260t3242 n8261 n3243 R=1.962e+01 
R8260t4566 n8261 n4567 R=3.960e+00 
R8260t7374 n8261 n7375 R=4.528e+00 
R8260t4390 n8261 n4391 R=1.158e+01 
R8261t2025 n8262 n2026 R=6.302e+01 
R8261t6354 n8262 n6355 R=2.924e+00 
R8261t6963 n8262 n6964 R=5.202e+01 
R8261t8054 n8262 n8055 R=2.092e+01 
R8262t3517 n8263 n3518 R=1.105e+02 
R8262t4463 n8263 n4464 R=5.481e+01 
R8262t75 n8263 n76 R=6.365e+00 
R8262t582 n8263 n583 R=1.665e+01 
R8262t6800 n8263 n6801 R=4.977e+00 
R8262t7286 n8263 n7287 R=1.049e+01 
R8262t563 n8263 n564 R=9.110e+00 
R8262t3763 n8263 n3764 R=6.628e+00 
R8262t1984 n8263 n1985 R=3.832e+01 
R8263t3543 n8264 n3544 R=1.512e+01 
R8263t4820 n8264 n4821 R=4.612e+00 
R8263t1558 n8264 n1559 R=3.775e+00 
R8263t265 n8264 n266 R=1.397e+01 
R8263t6218 n8264 n6219 R=8.083e+00 
R8263t3375 n8264 n3376 R=2.985e+01 
R8264t7892 n8265 n7893 R=4.243e+00 
R8264t4396 n8265 n4397 R=6.864e+00 
R8264t6782 n8265 n6783 R=3.027e+01 
R8264t7539 n8265 n7540 R=1.780e+00 
R8265t290 n8266 n291 R=6.821e+00 
R8265t1164 n8266 n1165 R=4.522e+00 
R8265t6730 n8266 n6731 R=8.433e+00 
R8266t2110 n8267 n2111 R=1.275e+02 
R8266t7504 n8267 n7505 R=7.014e+00 
R8266t5827 n8267 n5828 R=2.481e+01 
R8266t215 n8267 n216 R=2.477e+01 
R8266t1780 n8267 n1781 R=2.584e+01 
R8266t4145 n8267 n4146 R=6.367e+00 
R8266t3752 n8267 n3753 R=1.168e+02 
R8266t1246 n8267 n1247 R=4.479e+00 
R8267t1955 n8268 n1956 R=9.003e+00 
R8267t5062 n8268 n5063 R=1.670e+01 
R8267t5216 n8268 n5217 R=3.249e+00 
R8267t3126 n8268 n3127 R=4.504e+00 
R8267t2431 n8268 n2432 R=1.977e+01 
R8267t7994 n8268 n7995 R=1.392e+01 
R8268t5088 n8269 n5089 R=1.386e+01 
R8268t6991 n8269 n6992 R=2.263e+00 
R8268t1057 n8269 n1058 R=1.189e+01 
R8269t1956 n8270 n1957 R=6.902e+00 
R8269t7742 n8270 n7743 R=4.077e+01 
R8269t4186 n8270 n4187 R=2.780e+01 
R8269t6021 n8270 n6022 R=4.474e+00 
R8269t5685 n8270 n5686 R=5.978e+00 
R8269t858 n8270 n859 R=4.845e+01 
R8269t2409 n8270 n2410 R=3.833e+00 
R8270t4145 n8271 n4146 R=7.867e+00 
R8270t4536 n8271 n4537 R=2.261e+01 
R8270t3509 n8271 n3510 R=8.419e+00 
R8270t5100 n8271 n5101 R=9.449e+00 
R8270t3752 n8271 n3753 R=9.686e+00 
R8270t8266 n8271 n8267 R=6.216e+00 
R8271t3630 n8272 n3631 R=2.025e+00 
R8271t3486 n8272 n3487 R=1.014e+01 
R8271t5120 n8272 n5121 R=2.233e+01 
R8272t2784 n8273 n2785 R=7.243e+00 
R8272t3873 n8273 n3874 R=9.281e+00 
R8272t4005 n8273 n4006 R=2.356e+01 
R8272t4429 n8273 n4430 R=4.958e+00 
R8272t1619 n8273 n1620 R=3.165e+01 
R8272t4150 n8273 n4151 R=9.224e+00 
R8272t5372 n8273 n5373 R=6.862e+00 
R8273t2280 n8274 n2281 R=6.168e+01 
R8273t2109 n8274 n2110 R=3.674e+00 
R8273t7411 n8274 n7412 R=4.266e+00 
R8273t5067 n8274 n5068 R=1.088e+01 
R8274t301 n8275 n302 R=2.469e+00 
R8274t7595 n8275 n7596 R=4.596e+00 
R8274t6901 n8275 n6902 R=1.258e+01 
R8274t706 n8275 n707 R=1.288e+01 
R8274t7416 n8275 n7417 R=5.384e+01 
R8275t7290 n8276 n7291 R=1.171e+02 
R8275t4143 n8276 n4144 R=2.076e+01 
R8275t7953 n8276 n7954 R=1.272e+01 
R8275t996 n8276 n997 R=2.495e+00 
R8276t4745 n8277 n4746 R=2.781e+02 
R8276t5834 n8277 n5835 R=2.994e+00 
R8276t6526 n8277 n6527 R=5.332e+01 
R8276t6748 n8277 n6749 R=2.968e+00 
R8276t6162 n8277 n6163 R=6.891e+00 
R8276t6941 n8277 n6942 R=2.077e+01 
R8276t2059 n8277 n2060 R=1.079e+01 
R8277t482 n8278 n483 R=6.934e+00 
R8277t8020 n8278 n8021 R=4.906e+01 
R8277t7136 n8278 n7137 R=7.508e+00 
R8277t5880 n8278 n5881 R=7.464e+00 
R8277t6411 n8278 n6412 R=8.359e+00 
R8278t1678 n8279 n1679 R=4.771e+00 
R8278t3979 n8279 n3980 R=8.039e+00 
R8278t6248 n8279 n6249 R=2.364e+02 
R8279t3754 n8280 n3755 R=2.881e+01 
R8279t2711 n8280 n2712 R=8.822e+01 
R8279t1162 n8280 n1163 R=3.064e+01 
R8279t3194 n8280 n3195 R=3.301e+01 
R8279t5776 n8280 n5777 R=1.744e+00 
R8280t4184 n8281 n4185 R=2.722e+00 
R8280t6710 n8281 n6711 R=4.199e+01 
R8280t7575 n8281 n7576 R=8.739e+00 
R8280t3191 n8281 n3192 R=4.315e+00 
R8281t2894 n8282 n2895 R=1.085e+01 
R8281t7715 n8282 n7716 R=4.475e+00 
R8281t6293 n8282 n6294 R=3.138e+00 
R8282t109 n8283 n110 R=2.994e+00 
R8282t2423 n8283 n2424 R=1.262e+02 
R8282t4069 n8283 n4070 R=2.216e+00 
R8282t4986 n8283 n4987 R=9.571e+00 
R8282t7277 n8283 n7278 R=3.758e+01 
R8282t3675 n8283 n3676 R=5.492e+00 
R8283t4387 n8284 n4388 R=9.255e+00 
R8283t7951 n8284 n7952 R=1.276e+02 
R8283t7684 n8284 n7685 R=1.386e+01 
R8283t1959 n8284 n1960 R=1.190e+01 
R8283t8068 n8284 n8069 R=9.175e+00 
R8283t7511 n8284 n7512 R=2.488e+00 
R8283t2635 n8284 n2636 R=1.088e+01 
R8284t7146 n8285 n7147 R=2.018e+00 
R8284t7492 n8285 n7493 R=5.962e+01 
R8284t672 n8285 n673 R=1.470e+01 
R8284t3922 n8285 n3923 R=3.129e+00 
R8284t5820 n8285 n5821 R=8.958e+00 
R8285t7905 n8286 n7906 R=4.072e+00 
R8285t3385 n8286 n3386 R=1.881e+02 
R8286t3257 n8287 n3258 R=1.820e+01 
R8286t1152 n8287 n1153 R=4.099e+00 
R8286t6673 n8287 n6674 R=5.913e+00 
R8287t864 n8288 n865 R=1.769e+01 
R8287t7059 n8288 n7060 R=3.230e+01 
R8287t7795 n8288 n7796 R=3.176e+00 
R8287t5808 n8288 n5809 R=2.024e+01 
R8287t4978 n8288 n4979 R=3.431e+00 
R8287t2251 n8288 n2252 R=2.066e+01 
R8287t284 n8288 n285 R=3.679e+01 
R8288t1021 n8289 n1022 R=1.274e+01 
R8288t1192 n8289 n1193 R=3.011e+02 
R8288t4983 n8289 n4984 R=3.192e+00 
R8288t5339 n8289 n5340 R=5.487e+00 
R8288t4086 n8289 n4087 R=4.528e+00 
R8289t2875 n8290 n2876 R=3.173e+00 
R8289t5514 n8290 n5515 R=1.004e+01 
R8289t629 n8290 n630 R=5.713e+00 
R8289t4585 n8290 n4586 R=7.418e+00 
R8290t1548 n8291 n1549 R=4.095e+00 
R8290t7992 n8291 n7993 R=3.139e+01 
R8290t6441 n8291 n6442 R=1.459e+01 
R8290t4497 n8291 n4498 R=5.848e+00 
R8290t5350 n8291 n5351 R=2.471e+00 
R8291t4586 n8292 n4587 R=6.400e+00 
R8291t7307 n8292 n7308 R=2.520e+01 
R8291t1774 n8292 n1775 R=3.771e+00 
R8291t1637 n8292 n1638 R=1.844e+01 
R8291t1200 n8292 n1201 R=2.881e+01 
R8291t2708 n8292 n2709 R=2.191e+00 
R8292t2815 n8293 n2816 R=2.749e+00 
R8292t3974 n8293 n3975 R=4.572e+01 
R8292t5051 n8293 n5052 R=4.062e+00 
R8292t698 n8293 n699 R=3.104e+01 
R8293t6228 n8294 n6229 R=3.140e+00 
R8293t6835 n8294 n6836 R=2.456e+01 
R8293t2618 n8294 n2619 R=6.644e+00 
R8294t1339 n8295 n1340 R=5.390e+00 
R8294t7223 n8295 n7224 R=6.881e+00 
R8294t27 n8295 n28 R=1.102e+02 
R8294t8238 n8295 n8239 R=4.500e+00 
R8294t2839 n8295 n2840 R=5.339e+00 
R8295t1148 n8296 n1149 R=2.018e+01 
R8295t4705 n8296 n4706 R=7.003e+01 
R8295t6512 n8296 n6513 R=5.453e+00 
R8295t5439 n8296 n5440 R=1.567e+01 
R8295t6924 n8296 n6925 R=8.052e+00 
R8295t3971 n8296 n3972 R=4.803e+01 
R8295t720 n8296 n721 R=8.899e+00 
R8295t2111 n8296 n2112 R=2.287e+01 
R8296t2382 n8297 n2383 R=2.339e+01 
R8296t7981 n8297 n7982 R=5.411e+00 
R8296t2068 n8297 n2069 R=5.817e+01 
R8296t1303 n8297 n1304 R=9.457e+01 
R8296t2219 n8297 n2220 R=1.759e+02 
R8297t1778 n8298 n1779 R=2.762e+01 
R8297t7410 n8298 n7411 R=1.036e+01 
R8298t588 n8299 n589 R=2.819e+00 
R8298t2490 n8299 n2491 R=1.377e+01 
R8298t7447 n8299 n7448 R=6.162e+00 
R8298t7489 n8299 n7490 R=1.628e+01 
R8298t4672 n8299 n4673 R=7.063e+00 
R8298t4667 n8299 n4668 R=4.324e+01 
R8299t1652 n8300 n1653 R=5.028e+00 
R8299t4220 n8300 n4221 R=1.191e+01 
R8299t4792 n8300 n4793 R=2.328e+01 
R8299t2570 n8300 n2571 R=5.335e+01 
R8300t6086 n8301 n6087 R=4.431e+00 
R8300t2617 n8301 n2618 R=8.485e+00 
R8300t3915 n8301 n3916 R=3.349e+00 
R8300t3975 n8301 n3976 R=1.869e+01 
R8300t6505 n8301 n6506 R=1.139e+01 
R8301t2590 n8302 n2591 R=2.303e+00 
R8301t1058 n8302 n1059 R=8.053e+00 
R8301t5050 n8302 n5051 R=1.112e+01 
R8301t5903 n8302 n5904 R=1.189e+01 
R8302t6301 n8303 n6302 R=2.955e+00 
R8302t6638 n8303 n6639 R=5.739e+00 
R8302t8176 n8303 n8177 R=1.981e+01 
R8302t597 n8303 n598 R=2.364e+02 
R8302t3581 n8303 n3582 R=1.052e+02 
R8302t5507 n8303 n5508 R=2.982e+00 
R8303t578 n8304 n579 R=2.998e+00 
R8303t6618 n8304 n6619 R=2.002e+01 
R8303t8155 n8304 n8156 R=4.555e+00 
R8303t7609 n8304 n7610 R=3.661e+00 
R8304t2668 n8305 n2669 R=5.218e+00 
R8304t6370 n8305 n6371 R=1.704e+01 
R8304t405 n8305 n406 R=4.311e+00 
R8304t7792 n8305 n7793 R=5.707e+00 
R8304t1065 n8305 n1066 R=2.363e+01 
R8304t4920 n8305 n4921 R=8.456e+00 
R8305t5125 n8306 n5126 R=4.272e+00 
R8305t6198 n8306 n6199 R=1.667e+01 
R8305t6399 n8306 n6400 R=2.306e+00 
R8305t307 n8306 n308 R=3.478e+00 
R8306t3350 n8307 n3351 R=3.063e+01 
R8306t4182 n8307 n4183 R=3.325e+00 
R8306t5612 n8307 n5613 R=1.351e+01 
R8306t3996 n8307 n3997 R=2.874e+00 
R8306t7179 n8307 n7180 R=7.691e+00 
R8307t1050 n8308 n1051 R=6.603e+00 
R8307t4270 n8308 n4271 R=5.670e+00 
R8307t2658 n8308 n2659 R=5.612e+00 
R8307t5520 n8308 n5521 R=4.816e+00 
R8307t4903 n8308 n4904 R=2.004e+01 
R8308t2436 n8309 n2437 R=4.525e+01 
R8308t6034 n8309 n6035 R=7.947e+00 
R8308t6482 n8309 n6483 R=5.887e+00 
R8308t5157 n8309 n5158 R=4.534e+00 
R8309t2486 n8310 n2487 R=3.701e+00 
R8309t4210 n8310 n4211 R=2.396e+01 
R8309t5067 n8310 n5068 R=7.393e+00 
R8309t8273 n8310 n8274 R=3.218e+00 
R8309t2280 n8310 n2281 R=1.212e+01 
R8310t4132 n8311 n4133 R=2.558e+01 
R8310t4389 n8311 n4390 R=8.288e+01 
R8310t3162 n8311 n3163 R=3.586e+00 
R8310t2004 n8311 n2005 R=1.497e+01 
R8310t1429 n8311 n1430 R=1.848e+00 
R8310t7451 n8311 n7452 R=3.200e+01 
R8311t1067 n8312 n1068 R=2.577e+01 
R8311t3753 n8312 n3754 R=2.466e+00 
R8311t7598 n8312 n7599 R=8.286e+00 
R8311t2484 n8312 n2485 R=1.734e+01 
R8311t6026 n8312 n6027 R=2.204e+01 
R8312t4117 n8313 n4118 R=5.906e+00 
R8312t7218 n8313 n7219 R=4.963e+01 
R8312t4279 n8313 n4280 R=8.848e+00 
R8312t5021 n8313 n5022 R=1.015e+02 
R8312t2806 n8313 n2807 R=4.718e+00 
R8312t2193 n8313 n2194 R=8.291e+00 
R8312t6522 n8313 n6523 R=2.057e+01 
R8313t8297 n8314 n8298 R=3.913e+01 
R8313t937 n8314 n938 R=7.260e+00 
R8313t562 n8314 n563 R=9.266e+00 
R8313t3941 n8314 n3942 R=6.079e+00 
R8313t7410 n8314 n7411 R=3.455e+00 
R8314t6260 n8315 n6261 R=7.105e+00 
R8314t7627 n8315 n7628 R=2.959e+00 
R8314t122 n8315 n123 R=6.701e+00 
R8314t3794 n8315 n3795 R=6.030e+00 
R8315t784 n8316 n785 R=6.970e+01 
R8315t2922 n8316 n2923 R=3.303e+00 
R8315t4134 n8316 n4135 R=5.780e+01 
R8315t146 n8316 n147 R=7.110e+00 
R8315t3762 n8316 n3763 R=8.498e+00 
R8316t1761 n8317 n1762 R=3.688e+00 
R8316t7880 n8317 n7881 R=4.509e+00 
R8316t7996 n8317 n7997 R=5.771e+00 
R8316t5891 n8317 n5892 R=8.459e+00 
R8316t6953 n8317 n6954 R=3.718e+01 
R8317t6302 n8318 n6303 R=4.812e+00 
R8317t2339 n8318 n2340 R=2.345e+01 
R8317t1119 n8318 n1120 R=8.663e+00 
R8318t383 n8319 n384 R=1.103e+01 
R8318t558 n8319 n559 R=4.376e+00 
R8318t5774 n8319 n5775 R=6.352e+01 
R8318t6276 n8319 n6277 R=3.191e+00 
R8319t931 n8320 n932 R=2.938e+00 
R8319t7404 n8320 n7405 R=1.613e+01 
R8319t135 n8320 n136 R=9.558e+00 
R8319t6571 n8320 n6572 R=1.546e+01 
R8319t3548 n8320 n3549 R=2.117e+01 
R8319t5459 n8320 n5460 R=5.462e+00 
R8320t3307 n8321 n3308 R=2.225e+01 
R8320t7175 n8321 n7176 R=2.883e+00 
R8320t1717 n8321 n1718 R=1.705e+01 
R8320t4230 n8321 n4231 R=7.684e+00 
R8320t4207 n8321 n4208 R=1.659e+01 
R8320t453 n8321 n454 R=6.711e+00 
R8321t6268 n8322 n6269 R=3.782e+00 
R8321t8135 n8322 n8136 R=1.064e+01 
R8321t7766 n8322 n7767 R=2.987e+00 
R8322t1300 n8323 n1301 R=6.033e+00 
R8322t6322 n8323 n6323 R=4.994e+00 
R8322t1409 n8323 n1410 R=1.785e+01 
R8322t1443 n8323 n1444 R=4.921e+00 
R8322t1210 n8323 n1211 R=1.252e+01 
R8323t1163 n8324 n1164 R=1.792e+01 
R8323t2248 n8324 n2249 R=8.410e+00 
R8323t2335 n8324 n2336 R=1.799e+01 
R8323t2683 n8324 n2684 R=3.183e+01 
R8323t5925 n8324 n5926 R=3.835e+00 
R8323t6026 n8324 n6027 R=6.365e+00 
R8324t1014 n8325 n1015 R=4.017e+00 
R8324t5118 n8325 n5119 R=7.075e+00 
R8324t7973 n8325 n7974 R=7.589e+00 
R8324t2064 n8325 n2065 R=3.966e+00 
R8325t2390 n8326 n2391 R=7.499e+00 
R8325t556 n8326 n557 R=1.833e+01 
R8325t7439 n8326 n7440 R=2.076e+01 
R8325t3539 n8326 n3540 R=7.848e+01 
R8325t4980 n8326 n4981 R=1.203e+02 
R8325t7423 n8326 n7424 R=8.438e+00 
R8325t6956 n8326 n6957 R=5.216e+00 
R8326t8175 n8327 n8176 R=8.900e+00 
R8326t3631 n8327 n3632 R=1.799e+02 
R8326t5328 n8327 n5329 R=3.835e+00 
R8326t2920 n8327 n2921 R=1.527e+01 
R8326t5443 n8327 n5444 R=6.837e+00 
R8327t6406 n8328 n6407 R=1.221e+01 
R8327t7036 n8328 n7037 R=1.477e+01 
R8327t2226 n8328 n2227 R=6.775e+00 
R8327t7518 n8328 n7519 R=5.566e+00 
R8327t2591 n8328 n2592 R=1.858e+02 
R8327t4768 n8328 n4769 R=4.566e+00 
R8327t3923 n8328 n3924 R=1.685e+02 
R8328t6089 n8329 n6090 R=1.869e+01 
R8328t7123 n8329 n7124 R=3.499e+00 
R8329t3880 n8330 n3881 R=7.205e+00 
R8329t4500 n8330 n4501 R=5.429e+00 
R8329t3862 n8330 n3863 R=8.327e+00 
R8329t6719 n8330 n6720 R=1.239e+01 
R8329t4125 n8330 n4126 R=4.414e+00 
R8330t202 n8331 n203 R=5.208e+00 
R8330t2986 n8331 n2987 R=1.144e+01 
R8330t8252 n8331 n8253 R=2.768e+00 
R8331t1742 n8332 n1743 R=2.572e+00 
R8331t2778 n8332 n2779 R=4.500e+00 
R8331t1224 n8332 n1225 R=4.975e+00 
R8332t936 n8333 n937 R=1.550e+02 
R8332t4348 n8333 n4349 R=3.787e+00 
R8332t1882 n8333 n1883 R=3.482e+00 
R8332t5864 n8333 n5865 R=6.101e+00 
R8332t2761 n8333 n2762 R=1.941e+01 
R8332t4254 n8333 n4255 R=5.525e+00 
R8333t2898 n8334 n2899 R=2.646e+01 
R8333t3190 n8334 n3191 R=9.497e+01 
R8333t6659 n8334 n6660 R=2.433e+01 
R8333t2329 n8334 n2330 R=4.043e+00 
R8333t7443 n8334 n7444 R=8.816e+01 
R8333t3626 n8334 n3627 R=5.898e+00 
R8333t3174 n8334 n3175 R=4.677e+00 
R8333t342 n8334 n343 R=6.823e+00 
R8334t6518 n8335 n6519 R=5.267e+01 
R8334t7943 n8335 n7944 R=1.346e+00 
R8334t2780 n8335 n2781 R=1.907e+01 
R8334t2844 n8335 n2845 R=1.934e+00 
R8334t3297 n8335 n3298 R=1.867e+01 
R8334t7139 n8335 n7140 R=3.048e+01 
R8335t3156 n1 n3157 R=9.385e+00 
R8336t5604 n8337 n5605 R=1.489e+01 
R8336t6959 n8337 n6960 R=5.657e+00 
R8336t7372 n8337 n7373 R=1.404e+01 
R8336t2696 n8337 n2697 R=6.672e+00 
R8336t450 n8337 n451 R=9.577e+01 
R8336t5035 n8337 n5036 R=1.516e+01 
R8336t6343 n8337 n6344 R=1.393e+01 
R8337t1816 n8338 n1817 R=3.342e+01 
R8337t6436 n8338 n6437 R=9.171e+00 
R8337t1660 n8338 n1661 R=3.271e+01 
R8337t7569 n8338 n7570 R=1.839e+00 
R8337t8063 n8338 n8064 R=4.159e+00 
R8338t352 n8339 n353 R=7.903e+00 
R8338t1301 n8339 n1302 R=1.980e+01 
R8338t8018 n8339 n8019 R=7.296e+00 
R8338t3907 n8339 n3908 R=4.724e+00 
R8338t2917 n8339 n2918 R=2.045e+02 
R8338t3265 n8339 n3266 R=1.430e+01 
R8338t4631 n8339 n4632 R=1.051e+01 
R8339t7321 n8340 n7322 R=2.737e+00 
R8339t439 n8340 n440 R=6.802e+01 
R8340t3046 n8341 n3047 R=8.449e+00 
R8340t5749 n8341 n5750 R=1.196e+01 
R8340t452 n8341 n453 R=6.923e+00 
R8340t5290 n8341 n5291 R=1.296e+01 
R8340t5342 n8341 n5343 R=7.424e+00 
R8340t8171 n8341 n8172 R=5.495e+00 
R8341t693 n8342 n694 R=4.116e+01 
R8341t4010 n8342 n4011 R=4.288e+01 
R8341t1023 n8342 n1024 R=8.862e+00 
R8341t965 n8342 n966 R=7.827e+01 
R8341t3962 n8342 n3963 R=9.838e+00 
R8341t4620 n8342 n4621 R=7.549e+00 
R8341t8143 n8342 n8144 R=4.780e+00 
R8341t659 n8342 n660 R=4.021e+00 
R8342t4557 n8343 n4558 R=6.466e+00 
R8342t6092 n8343 n6093 R=6.845e+00 
R8342t1384 n8343 n1385 R=2.395e+01 
R8342t2085 n8343 n2086 R=2.054e+01 
R8342t6097 n8343 n6098 R=5.543e+00 
R8343t5832 n8344 n5833 R=4.328e+00 
R8343t7207 n8344 n7208 R=1.198e+01 
R8343t7819 n8344 n7820 R=2.907e+01 
R8343t7205 n8344 n7206 R=7.332e+00 
R8343t1030 n8344 n1031 R=6.821e+00 
R8343t1433 n8344 n1434 R=1.828e+01 
R8344t2663 n8345 n2664 R=7.322e+00 
R8344t6657 n8345 n6658 R=1.418e+02 
R8344t2326 n8345 n2327 R=9.081e+00 
R8344t4518 n8345 n4519 R=2.372e+00 
R8344t4119 n8345 n4120 R=1.313e+01 
R8344t1004 n8345 n1005 R=7.994e+00 
R8345t6699 n8346 n6700 R=1.438e+00 
R8345t6763 n8346 n6764 R=6.387e+00 
R8345t3358 n8346 n3359 R=1.331e+01 
R8345t37 n8346 n38 R=5.539e+00 
R8346t1045 n8347 n1046 R=1.785e+00 
R8346t7246 n8347 n7247 R=2.439e+01 
R8346t7323 n8347 n7324 R=2.097e+01 
R8346t7383 n8347 n7384 R=2.469e+00 
R8346t2295 n8347 n2296 R=1.144e+01 
R8347t5376 n8348 n5377 R=8.075e+00 
R8347t1333 n8348 n1334 R=1.561e+01 
R8347t2759 n8348 n2760 R=1.520e+01 
R8347t6266 n8348 n6267 R=6.504e+00 
R8347t3051 n8348 n3052 R=9.419e+00 
R8348t6479 n8349 n6480 R=1.007e+01 
R8348t6535 n8349 n6536 R=4.234e+01 
R8348t5943 n8349 n5944 R=5.139e+00 
R8348t2372 n8349 n2373 R=3.054e+00 
R8348t1359 n8349 n1360 R=5.151e+00 
R8349t825 n8350 n826 R=5.374e+00 
R8349t7815 n8350 n7816 R=2.871e+00 
R8349t7739 n8350 n7740 R=3.073e+00 
R8349t5382 n8350 n5383 R=4.350e+01 
R8350t7325 n8351 n7326 R=3.748e+01 
R8350t1187 n8351 n1188 R=5.569e+00 
R8350t5656 n8351 n5657 R=8.281e+00 
R8350t6379 n8351 n6380 R=2.072e+01 
R8350t6511 n8351 n6512 R=6.151e+00 
R8351t2969 n8352 n2970 R=2.726e+00 
R8351t4143 n8352 n4144 R=4.709e+00 
R8351t4857 n8352 n4858 R=2.716e+01 
R8351t5418 n8352 n5419 R=2.351e+00 
R8352t618 n8353 n619 R=9.149e+00 
R8352t3372 n8353 n3373 R=8.445e+01 
R8352t2014 n8353 n2015 R=5.737e+00 
R8352t6876 n8353 n6877 R=1.312e+01 
R8352t1653 n8353 n1654 R=4.331e+00 
R8352t7931 n8353 n7932 R=5.519e+00 
R8353t936 n8354 n937 R=9.193e+00 
R8353t2445 n8354 n2446 R=1.344e+01 
R8353t1882 n8354 n1883 R=6.738e+00 
R8353t5864 n8354 n5865 R=2.755e+01 
R8353t5775 n8354 n5776 R=7.140e+00 
R8353t4062 n8354 n4063 R=1.248e+01 
R8353t8009 n8354 n8010 R=1.830e+01 
R8354t6699 n8355 n6700 R=6.393e+02 
R8354t6923 n8355 n6924 R=3.563e+00 
R8354t2511 n8355 n2512 R=3.284e+00 
R8354t6763 n8355 n6764 R=2.136e+00 
R8354t8345 n8355 n8346 R=1.443e+02 
R8355t7156 n8356 n7157 R=1.212e+01 
R8355t7215 n8356 n7216 R=5.089e+01 
R8355t3624 n8356 n3625 R=2.158e+00 
R8355t5784 n8356 n5785 R=3.036e+01 
R8355t134 n8356 n135 R=5.870e+01 
R8356t3669 n8357 n3670 R=7.105e+00 
R8356t8038 n8357 n8039 R=1.421e+01 
R8356t6883 n8357 n6884 R=1.026e+01 
R8356t198 n8357 n199 R=1.031e+02 
R8356t4779 n8357 n4780 R=2.973e+00 
R8357t5345 n8358 n5346 R=3.514e+00 
R8357t4890 n8358 n4891 R=3.022e+00 
R8357t4771 n8358 n4772 R=2.088e+01 
R8358t1321 n8359 n1322 R=3.146e+00 
R8358t4209 n8359 n4210 R=2.041e+01 
R8358t7360 n8359 n7361 R=2.771e+01 
R8358t5099 n8359 n5100 R=4.882e+00 
R8358t5732 n8359 n5733 R=8.188e+00 
R8358t3630 n8359 n3631 R=4.127e+01 
R8358t8271 n8359 n8272 R=1.036e+01 
R8359t970 n8360 n971 R=1.887e+01 
R8359t5535 n8360 n5536 R=9.142e+00 
R8359t2455 n8360 n2456 R=3.651e+01 
R8359t6498 n8360 n6499 R=2.982e+01 
R8359t4418 n8360 n4419 R=1.538e+01 
R8359t4243 n8360 n4244 R=4.416e+00 
R8359t5843 n8360 n5844 R=5.461e+00 
R8359t5923 n8360 n5924 R=3.775e+01 
R8360t4299 n8361 n4300 R=3.756e+01 
R8360t4661 n8361 n4662 R=7.558e+00 
R8360t1358 n8361 n1359 R=4.817e+00 
R8360t2837 n8361 n2838 R=1.255e+01 
R8360t1280 n8361 n1281 R=8.785e+00 
R8360t6397 n8361 n6398 R=3.662e+00 
R8361t160 n8362 n161 R=1.869e+01 
R8361t6362 n8362 n6363 R=6.214e+00 
R8361t8128 n8362 n8129 R=1.600e+01 
R8361t6095 n8362 n6096 R=8.330e+00 
R8361t2495 n8362 n2496 R=4.271e+01 
R8361t3293 n8362 n3294 R=8.882e+00 
R8361t4617 n8362 n4618 R=3.425e+00 
R8362t4807 n8363 n1 R=5.965e+00 
R8362t7710 n8363 n7711 R=7.030e+00 
R8362t3989 n8363 n3990 R=3.197e+00 
R8362t3236 n8363 n3237 R=3.543e+01 
R8362t4975 n8363 n4976 R=9.886e+00 
R8362t1322 n8363 n1 R=7.103e+00 
R8363t4003 n8364 n4004 R=1.038e+01 
R8363t8153 n8364 n8154 R=3.585e+00 
R8363t4680 n8364 n4681 R=3.119e+01 
R8363t2851 n8364 n2852 R=7.982e+00 
R8363t1777 n8364 n1778 R=7.357e+00 
R8363t176 n8364 n177 R=5.245e+00 
R8364t1391 n8365 n1392 R=1.033e+01 
R8364t7983 n8365 n7984 R=2.619e+00 
R8364t6599 n8365 n6600 R=4.268e+00 
R8364t7064 n8365 n7065 R=1.451e+02 
R8364t3136 n8365 n3137 R=7.325e+00 
R8364t7890 n8365 n7891 R=4.034e+01 
R8365t1141 n8366 n1142 R=7.008e+01 
R8365t7989 n8366 n7990 R=2.274e+00 
R8365t694 n8366 n695 R=2.364e+01 
R8365t6705 n8366 n6706 R=5.144e+00 
R8365t6508 n8366 n6509 R=9.173e+01 
R8365t1820 n8366 n1821 R=2.928e+00 
R8366t1946 n8367 n1947 R=5.671e+00 
R8366t7784 n8367 n7785 R=5.647e+00 
R8366t2640 n8367 n2641 R=2.786e+01 
R8367t1145 n8368 n1146 R=3.951e+00 
R8367t4332 n8368 n4333 R=6.655e+00 
R8367t4363 n8368 n4364 R=1.516e+01 
R8367t6413 n8368 n6414 R=1.646e+01 
R8367t8139 n8368 n8140 R=1.388e+01 
R8368t3391 n8369 n3392 R=6.559e+00 
R8368t5773 n8369 n5774 R=4.073e+00 
R8369t1679 n8370 n1680 R=1.076e+01 
R8369t7128 n8370 n7129 R=2.271e+00 
R8369t2367 n8370 n2368 R=1.127e+01 
R8370t2604 n8371 n2605 R=6.537e+00 
R8370t2744 n8371 n2745 R=2.061e+01 
R8370t141 n8371 n142 R=7.433e+00 
R8370t3649 n8371 n3650 R=1.643e+01 
R8370t6842 n8371 n6843 R=1.391e+01 
R8370t3432 n8371 n3433 R=1.732e+01 
R8370t3260 n8371 n3261 R=1.226e+01 
R8371t233 n8372 n234 R=1.107e+01 
R8371t2155 n8372 n2156 R=3.304e+00 
R8371t3242 n8372 n3243 R=4.932e+00 
R8372t7152 n8373 n7153 R=1.293e+02 
R8372t4637 n8373 n4638 R=7.534e+00 
R8372t7095 n8373 n7096 R=4.319e+00 
R8373t1363 n8374 n1364 R=3.257e+00 
R8373t4819 n8374 n4820 R=9.863e+01 
R8373t1587 n8374 n1588 R=6.572e+00 
R8373t7523 n8374 n7524 R=1.432e+01 
R8373t5702 n8374 n5703 R=3.495e+01 
R8373t567 n8374 n568 R=3.453e+00 
R8373t5914 n8374 n5915 R=1.677e+02 
R8373t3248 n8374 n3249 R=4.407e+01 
R8374t1080 n8375 n1081 R=3.491e+00 
R8374t3007 n8375 n3008 R=9.089e+01 
R8374t4928 n8375 n4929 R=7.566e+01 
R8374t3063 n8375 n3064 R=2.061e+00 
R8374t7282 n8375 n7283 R=3.735e+00 
R8375t3283 n8376 n3284 R=9.209e+00 
R8375t4927 n8376 n4928 R=8.374e+00 
R8375t6019 n8376 n6020 R=1.172e+01 
R8375t2622 n8376 n2623 R=3.957e+00 
R8375t1139 n8376 n1140 R=1.467e+02 
R8376t4496 n8377 n4497 R=6.157e+00 
R8376t7627 n8377 n7628 R=1.857e+01 
R8376t3736 n8377 n3737 R=7.984e+00 
R8376t5011 n8377 n5012 R=4.881e+00 
R8377t499 n8378 n500 R=4.358e+00 
R8377t2274 n8378 n2275 R=5.236e+00 
R8377t2230 n8378 n2231 R=1.121e+01 
R8377t6254 n8378 n6255 R=2.740e+00 
R8377t4826 n8378 n4827 R=3.347e+01 
R8377t1702 n8378 n1703 R=1.234e+03 
R8378t6134 n8379 n6135 R=1.467e+01 
R8378t4075 n8379 n4076 R=7.504e+00 
R8378t3120 n8379 n3121 R=3.565e+01 
R8378t2909 n8379 n2910 R=6.186e+00 
R8378t4313 n8379 n4314 R=1.867e+02 
R8378t7047 n8379 n7048 R=5.019e+00 
R8378t1770 n8379 n1771 R=2.847e+01 
R8379t6829 n8380 n6830 R=4.872e+00 
R8379t7430 n8380 n7431 R=5.773e+00 
R8379t1120 n8380 n1121 R=3.364e+00 
R8380t5175 n8381 n5176 R=1.739e+01 
R8380t3485 n8381 n3486 R=3.740e+00 
R8380t7678 n8381 n7679 R=4.052e+00 
R8380t4740 n8381 n4741 R=1.675e+01 
R8380t2958 n8381 n2959 R=9.314e+00 
R8380t4335 n8381 n4336 R=5.470e+01 
R8381t1296 n8382 n1297 R=8.788e+00 
R8381t4489 n8382 n4490 R=5.071e+00 
R8381t4114 n8382 n4115 R=5.751e+00 
R8381t1144 n8382 n1145 R=5.394e+01 
R8381t136 n8382 n137 R=7.891e+00 
R8381t6524 n8382 n6525 R=1.120e+01 
R8381t5235 n8382 n5236 R=1.707e+01 
R8382t1647 n8383 n1648 R=1.777e+01 
R8382t7716 n8383 n7717 R=4.814e+00 
R8382t3051 n8383 n3052 R=5.591e+00 
R8382t8347 n8383 n8348 R=3.466e+01 
R8382t6266 n8383 n6267 R=2.525e+00 
R8383t5536 n8384 n5537 R=2.638e+00 
R8383t6449 n8384 n6450 R=1.141e+01 
R8383t5121 n8384 n5122 R=6.969e+00 
R8384t4506 n8385 n4507 R=2.943e+00 
R8384t7831 n8385 n7832 R=1.657e+01 
R8384t2515 n8385 n2516 R=3.830e+00 
R8385t3431 n8386 n3432 R=1.813e+02 
R8385t3884 n8386 n3885 R=1.917e+01 
R8385t2386 n8386 n2387 R=1.005e+01 
R8385t434 n8386 n435 R=3.092e+00 
R8385t7647 n8386 n7648 R=1.119e+02 
R8385t4204 n8386 n4205 R=2.450e+00 
R8385t5161 n8386 n5162 R=2.858e+01 
R8385t5159 n8386 n5160 R=1.636e+01 
R8386t8074 n8387 n8075 R=3.666e+00 
R8386t3768 n8387 n3769 R=3.321e+00 
R8387t6074 n8388 n6075 R=7.230e+00 
R8387t7552 n8388 n7553 R=5.287e+01 
R8387t5056 n8388 n5057 R=5.187e+00 
R8387t6531 n8388 n6532 R=5.972e+00 
R8387t1471 n8388 n1472 R=3.993e+01 
R8387t6134 n8388 n6135 R=3.104e+01 
R8387t5201 n8388 n5202 R=1.898e+01 
R8387t1469 n8388 n1470 R=4.144e+00 
R8388t2832 n8389 n2833 R=3.128e+00 
R8388t6614 n8389 n6615 R=6.013e+00 
R8388t2775 n8389 n2776 R=5.293e+01 
R8388t5955 n8389 n5956 R=6.073e+00 
R8388t6590 n8389 n6591 R=3.286e+00 
R8389t299 n8390 n300 R=4.362e+00 
R8389t7731 n8390 n7732 R=1.202e+01 
R8389t1193 n8390 n1194 R=2.273e+00 
R8389t4727 n8390 n4728 R=1.276e+01 
R8390t5857 n8391 n5858 R=4.160e+00 
R8390t3690 n8391 n3691 R=7.799e+00 
R8390t142 n8391 n143 R=6.981e+00 
R8391t3243 n8392 n3244 R=3.722e+00 
R8391t4899 n8392 n4900 R=5.843e+00 
R8391t1012 n8392 n1013 R=1.198e+01 
R8391t3733 n8392 n3734 R=4.861e+01 
R8391t422 n8392 n423 R=3.679e+00 
R8391t7350 n8392 n7351 R=1.402e+01 
R8392t6858 n8393 n6859 R=5.197e+00 
R8392t5878 n8393 n5879 R=3.345e+00 
R8392t3779 n8393 n3780 R=1.352e+01 
R8393t5419 n8394 n5420 R=6.044e+00 
R8393t1228 n8394 n1229 R=3.360e+01 
R8393t4747 n8394 n4748 R=3.985e+00 
R8394t5553 n8395 n5554 R=8.932e+00 
R8394t7868 n8395 n7869 R=3.252e+00 
R8394t572 n8395 n573 R=1.043e+01 
R8394t5930 n8395 n5931 R=9.779e+00 
R8394t4337 n8395 n4338 R=6.153e+00 
R8394t6118 n8395 n6119 R=5.376e+01 
R8395t4274 n8396 n4275 R=4.263e+00 
R8395t6288 n8396 n6289 R=3.992e+00 
R8395t7958 n8396 n7959 R=1.120e+01 
R8396t7070 n8397 n7071 R=1.163e+01 
R8396t7024 n8397 n7025 R=1.688e+01 
R8396t8039 n8397 n8040 R=3.191e+00 
R8396t6871 n8397 n6872 R=2.440e+01 
R8396t1998 n8397 n1999 R=6.148e+00 
R8397t3273 n8398 n3274 R=2.687e+01 
R8397t8214 n8398 n8215 R=7.507e+02 
R8397t4492 n8398 n4493 R=4.196e+00 
R8397t7629 n8398 n7630 R=3.939e+02 
R8397t2242 n8398 n2243 R=3.721e+00 
R8398t2704 n8399 n2705 R=3.686e+00 
R8398t6287 n8399 n6288 R=4.983e+01 
R8398t458 n8399 n459 R=9.246e+00 
R8398t3658 n8399 n3659 R=1.391e+01 
R8398t2885 n8399 n2886 R=6.386e+00 
R8399t6401 n8400 n6402 R=3.707e+00 
R8399t6450 n8400 n6451 R=4.911e+01 
R8399t8008 n8400 n8009 R=1.509e+01 
R8399t2875 n8400 n2876 R=3.287e+00 
R8399t7745 n8400 n7746 R=7.868e+00 
R8400t6963 n8401 n6964 R=3.279e+00 
R8400t8261 n8401 n8262 R=1.518e+01 
R8400t8207 n8401 n8208 R=5.714e+00 
R8400t8054 n8401 n8055 R=2.335e+00 
R8401t3661 n8402 n3662 R=8.197e+00 
R8401t5481 n8402 n5482 R=5.808e+00 
R8401t6301 n8402 n6302 R=1.223e+01 
R8401t6638 n8402 n6639 R=4.568e+00 
R8402t3621 n8403 n3622 R=4.190e+00 
R8402t4039 n8403 n4040 R=3.866e+00 
R8402t6443 n8403 n6444 R=2.554e+01 
R8403t5554 n8404 n5555 R=5.880e+00 
R8403t1941 n8404 n1942 R=4.536e+01 
R8403t4329 n8404 n4330 R=2.140e+01 
R8404t5197 n8405 n5198 R=3.098e+01 
R8404t6310 n8405 n6311 R=3.440e+00 
R8404t2035 n8405 n2036 R=1.075e+01 
R8404t7057 n8405 n7058 R=5.855e+00 
R8404t1923 n8405 n1924 R=7.009e+00 
R8404t3385 n8405 n3386 R=1.915e+02 
R8404t4635 n8405 n4636 R=6.382e+00 
R8405t63 n8406 n64 R=2.577e+01 
R8405t6936 n8406 n6937 R=4.600e+00 
R8405t1499 n8406 n1500 R=6.190e+00 
R8405t1176 n8406 n1177 R=7.697e+00 
R8405t2177 n8406 n2178 R=7.392e+00 
R8406t917 n8407 n918 R=6.814e+00 
R8406t3673 n8407 n3674 R=3.821e+00 
R8406t4581 n8407 n4582 R=9.646e+01 
R8406t2329 n8407 n2330 R=2.525e+00 
R8406t6659 n8407 n6660 R=9.330e+00 
R8407t1678 n8408 n1679 R=1.065e+01 
R8407t8278 n8408 n8279 R=7.420e+00 
R8407t6248 n8408 n6249 R=6.137e+00 
R8407t5640 n8408 n5641 R=9.584e+00 
R8407t7913 n8408 n7914 R=1.155e+01 
R8407t6722 n8408 n6723 R=7.133e+00 
R8408t466 n8409 n467 R=3.972e+01 
R8408t5765 n8409 n5766 R=2.068e+00 
R8408t1393 n8409 n1394 R=3.045e+01 
R8408t2456 n8409 n2457 R=2.594e+00 
R8409t137 n8410 n138 R=1.364e+01 
R8409t6942 n8410 n6943 R=1.595e+01 
R8409t4628 n8410 n4629 R=3.261e+01 
R8409t7257 n8410 n7258 R=1.249e+01 
R8410t1285 n8411 n1286 R=4.166e+00 
R8410t6426 n8411 n6427 R=9.424e+00 
R8410t7461 n8411 n7462 R=5.108e+00 
R8410t8250 n8411 n8251 R=6.458e+02 
R8410t3446 n8411 n3447 R=3.553e+00 
R8411t2835 n8412 n2836 R=1.268e+01 
R8411t2575 n8412 n2576 R=3.039e+00 
R8411t4147 n8412 n4148 R=1.388e+01 
R8411t3903 n8412 n3904 R=2.784e+01 
R8412t3085 n8413 n3086 R=4.159e+00 
R8412t2592 n8413 n2593 R=3.573e+00 
R8412t953 n8413 n954 R=1.321e+02 
R8412t7076 n8413 n7077 R=4.322e+00 
R8412t2259 n8413 n2260 R=6.131e+01 
R8413t5928 n8414 n5929 R=5.031e+00 
R8413t6438 n8414 n6439 R=9.099e+00 
R8413t8034 n8414 n8035 R=1.753e+01 
R8413t1999 n8414 n2000 R=5.080e+00 
R8413t1214 n8414 n1215 R=8.830e+00 
R8414t1871 n8415 n1872 R=1.063e+01 
R8414t8138 n8415 n8139 R=1.263e+01 
R8414t6261 n8415 n6262 R=5.799e+01 
R8414t2452 n8415 n2453 R=1.875e+01 
R8414t6919 n8415 n6920 R=6.180e+00 
R8414t238 n8415 n239 R=1.101e+01 
R8414t1101 n8415 n1102 R=3.694e+00 
R8415t4964 n8416 n4965 R=1.339e+01 
R8415t7116 n8416 n7117 R=4.984e+00 
R8415t1478 n8416 n1479 R=1.336e+01 
R8415t1850 n8416 n1851 R=2.208e+01 
R8415t3807 n8416 n3808 R=7.755e+00 
R8415t6210 n8416 n6211 R=4.660e+00 
R8416t4117 n8417 n4118 R=3.990e+00 
R8416t8312 n8417 n8313 R=1.250e+01 
R8416t6522 n8417 n6523 R=4.680e+00 
R8416t1561 n8417 n1562 R=1.212e+01 
R8417t5325 n8418 n5326 R=3.509e+00 
R8417t3106 n8418 n3107 R=2.207e+01 
R8417t3009 n8418 n3010 R=2.417e+00 
R8417t4416 n8418 n4417 R=2.756e+01 
R8418t31 n8419 n32 R=1.183e+01 
R8418t3915 n8419 n3916 R=1.093e+01 
R8418t2098 n8419 n2099 R=5.734e+00 
R8418t271 n8419 n272 R=7.892e+00 
R8418t580 n8419 n581 R=5.961e+00 
R8418t589 n8419 n590 R=5.315e+00 
R8419t2527 n8420 n2528 R=4.233e+03 
R8419t3925 n8420 n3926 R=8.715e+00 
R8419t1511 n8420 n1512 R=2.414e+02 
R8419t4133 n8420 n4134 R=1.818e+01 
R8419t2681 n8420 n2682 R=7.151e+00 
R8419t5727 n8420 n5728 R=7.591e+00 
R8419t5212 n8420 n5213 R=6.479e+00 
R8420t6207 n8421 n6208 R=5.830e+00 
R8420t5837 n8421 n5838 R=9.598e+00 
R8420t5495 n8421 n5496 R=1.263e+01 
R8420t4511 n8421 n4512 R=4.968e+01 
R8420t1720 n8421 n1721 R=2.346e+01 
R8421t1987 n8422 n1988 R=5.254e+00 
R8421t6461 n8422 n6462 R=6.388e+01 
R8421t2445 n8422 n2446 R=1.139e+01 
R8421t940 n8422 n941 R=2.301e+00 
R8421t5799 n8422 n5800 R=7.335e+02 
R8421t7993 n8422 n7994 R=4.528e+00 
R8422t5169 n8423 n5170 R=3.230e+01 
R8422t5756 n8423 n5757 R=7.378e+00 
R8422t7215 n8423 n7216 R=7.538e+00 
R8422t7156 n8423 n7157 R=1.547e+02 
R8422t8223 n8423 n8224 R=8.454e+00 
R8422t5106 n8423 n5107 R=1.212e+01 
R8422t5410 n8423 n5411 R=5.268e+00 
R8423t555 n8424 n556 R=1.742e+01 
R8423t6086 n8424 n6087 R=1.257e+01 
R8423t5236 n8424 n5237 R=4.363e+00 
R8423t3397 n8424 n3398 R=1.673e+01 
R8423t2617 n8424 n2618 R=6.303e+00 
R8423t8300 n8424 n8301 R=6.580e+00 
R8424t6420 n8425 n6421 R=5.721e+01 
R8424t8061 n8425 n8062 R=1.524e+01 
R8424t5115 n8425 n5116 R=6.865e+00 
R8424t2161 n8425 n2162 R=6.620e+01 
R8424t1311 n8425 n1312 R=4.679e+00 
R8425t4126 n8426 n4127 R=5.180e+01 
R8425t7345 n8426 n7346 R=7.412e+00 
R8425t1431 n8426 n1432 R=2.899e+00 
R8425t4248 n8426 n4249 R=5.027e+01 
R8425t5972 n8426 n5973 R=3.205e+00 
R8426t1005 n8427 n1006 R=4.340e+00 
R8426t1785 n8427 n1786 R=2.886e+01 
R8426t2950 n8427 n2951 R=1.021e+02 
R8426t321 n8427 n322 R=3.893e+00 
R8426t319 n8427 n320 R=3.440e+00 
R8427t7662 n8428 n1 R=6.672e+00 
R8427t2063 n8428 n1 R=1.595e+01 
R8427t3638 n8428 n3639 R=4.786e+01 
R8427t5455 n8428 n5456 R=1.753e+01 
R8427t6368 n8428 n6369 R=1.220e+01 
R8427t2395 n8428 n1 R=6.797e+00 
R8428t542 n8429 n543 R=8.996e+00 
R8428t1081 n8429 n1082 R=2.103e+02 
R8428t5239 n8429 n5240 R=2.009e+00 
R8428t3422 n8429 n3423 R=3.235e+01 
R8428t7137 n8429 n7138 R=2.575e+00 
R8428t3415 n8429 n3416 R=7.520e+00 
R8429t5561 n8430 n5562 R=1.415e+01 
R8429t1851 n8430 n1852 R=1.095e+01 
R8429t3650 n8430 n3651 R=1.287e+02 
R8429t4956 n8430 n4957 R=2.077e+00 
R8429t3596 n8430 n3597 R=1.134e+01 
R8429t5131 n8430 n5132 R=1.395e+02 
R8430t3279 n8431 n3280 R=5.275e+01 
R8430t5465 n8431 n5466 R=1.704e+01 
R8430t2399 n8431 n2400 R=5.211e+00 
R8430t5093 n8431 n5094 R=4.780e+00 
R8431t6194 n8432 n6195 R=4.581e+00 
R8431t7841 n8432 n7842 R=6.118e+00 
R8431t6449 n8432 n6450 R=7.600e+00 
R8431t1382 n8432 n1383 R=1.905e+01 
R8431t808 n8432 n809 R=1.316e+01 
R8432t2004 n8433 n2005 R=3.761e+00 
R8432t8310 n8433 n8311 R=2.518e+01 
R8432t3011 n8433 n3012 R=9.617e+00 
R8432t471 n8433 n472 R=9.665e+00 
R8432t3162 n8433 n3163 R=3.899e+00 
R8433t7950 n8434 n7951 R=3.097e+00 
R8433t4442 n8434 n4443 R=4.695e+00 
R8433t54 n8434 n55 R=2.934e+01 
R8434t1972 n8435 n1973 R=7.463e+00 
R8434t2136 n8435 n2137 R=1.545e+01 
R8434t2208 n8435 n2209 R=1.808e+01 
R8434t5762 n8435 n5763 R=8.445e+00 
R8434t901 n8435 n902 R=7.269e+00 
R8434t3254 n8435 n3255 R=7.116e+00 
R8434t3251 n8435 n3252 R=1.147e+01 
R8435t2754 n8436 n2755 R=2.690e+00 
R8435t3655 n8436 n3656 R=1.081e+01 
R8435t5574 n8436 n5575 R=2.232e+01 
R8435t7349 n8436 n7350 R=3.301e+00 
R8435t2163 n8436 n2164 R=1.185e+01 
R8436t2277 n8437 n2278 R=1.743e+01 
R8436t6903 n8437 n6904 R=3.813e+00 
R8436t7727 n8437 n7728 R=4.129e+00 
R8436t893 n8437 n894 R=8.441e+00 
R8436t7209 n8437 n7210 R=6.615e+01 
R8436t5313 n8437 n5314 R=5.928e+00 
R8437t192 n8438 n193 R=2.197e+01 
R8437t3570 n8438 n3571 R=6.997e+00 
R8437t6950 n8438 n6951 R=2.680e+01 
R8437t5057 n8438 n5058 R=3.157e+01 
R8437t8188 n8438 n8189 R=1.038e+01 
R8437t5240 n8438 n5241 R=7.634e+00 
R8437t3139 n8438 n3140 R=3.125e+03 
R8437t6961 n8438 n6962 R=1.457e+01 
R8438t7077 n8439 n7078 R=3.948e+00 
R8438t5285 n8439 n5286 R=4.256e+00 
R8438t8202 n8439 n8203 R=1.552e+01 
R8439t5753 n8440 n5754 R=7.159e+01 
R8439t6337 n8440 n6338 R=2.058e+00 
R8439t7350 n8440 n7351 R=3.076e+00 
R8439t3015 n8440 n3016 R=5.360e+01 
R8439t5733 n8440 n5734 R=6.849e+00 
R8440t1117 n8441 n1118 R=6.962e+00 
R8440t7471 n8441 n7472 R=3.131e+01 
R8440t6874 n8441 n6875 R=3.092e+01 
R8440t2246 n8441 n2247 R=4.496e+00 
R8440t7570 n8441 n7571 R=8.114e+00 
R8440t7764 n8441 n7765 R=1.134e+01 
R8440t5427 n8441 n5428 R=2.415e+01 
R8441t4535 n8442 n4536 R=4.368e+00 
R8441t1474 n8442 n1475 R=1.382e+01 
R8441t6276 n8442 n6277 R=4.505e+01 
R8441t8318 n8442 n8319 R=5.492e+00 
R8441t5774 n8442 n5775 R=2.569e+01 
R8442t964 n8443 n965 R=2.455e+00 
R8442t1836 n8443 n1837 R=5.480e+00 
R8442t3216 n8443 n3217 R=6.095e+00 
R8442t7230 n8443 n7231 R=1.252e+02 
R8442t5976 n8443 n5977 R=1.459e+01 
R8443t6930 n8444 n6931 R=5.374e+01 
R8443t760 n8444 n761 R=9.250e+00 
R8443t6900 n8444 n6901 R=1.161e+02 
R8443t2695 n8444 n2696 R=1.111e+01 
R8443t2317 n8444 n2318 R=2.874e+01 
R8443t6962 n8444 n6963 R=3.976e+00 
R8443t5797 n8444 n5798 R=2.395e+02 
R8443t974 n8444 n975 R=4.215e+00 
R8444t1 n8445 n2 R=4.949e+00 
R8444t6319 n8445 n6320 R=2.602e+01 
R8444t7938 n8445 n1 R=4.204e+00 
R8444t5602 n8445 n1 R=1.059e+01 
R8444t3796 n8445 n3797 R=3.901e+00 
R8444t1650 n8445 n1651 R=5.969e+01 
R8445t5354 n8446 n5355 R=5.547e+00 
R8445t218 n8446 n219 R=4.285e+00 
R8445t7247 n8446 n7248 R=1.022e+01 
R8446t1547 n8447 n1548 R=4.586e+00 
R8446t6671 n8447 n6672 R=5.293e+00 
R8446t6262 n8447 n6263 R=1.075e+01 
R8447t1016 n8448 n1017 R=7.726e+00 
R8447t2725 n8448 n2726 R=3.216e+00 
R8447t3489 n8448 n3490 R=2.845e+01 
R8447t4549 n8448 n4550 R=1.889e+01 
R8447t6299 n8448 n6300 R=2.808e+01 
R8448t4724 n8449 n4725 R=2.021e+01 
R8448t5995 n8449 n5996 R=4.357e+00 
R8448t2173 n8449 n2174 R=8.831e+00 
R8449t1632 n8450 n1633 R=3.806e+00 
R8449t5949 n8450 n5950 R=1.062e+01 
R8449t2769 n8450 n2770 R=1.420e+01 
R8449t8094 n8450 n8095 R=2.257e+01 
R8449t1009 n8450 n1010 R=2.722e+00 
R8449t8161 n8450 n8162 R=1.163e+02 
R8450t5650 n8451 n5651 R=1.021e+01 
R8450t6858 n8451 n6859 R=6.111e+00 
R8450t8392 n8451 n8393 R=5.711e+00 
R8450t3779 n8451 n3780 R=4.054e+00 
R8450t1580 n8451 n1581 R=6.373e+01 
R8451t2680 n8452 n2681 R=2.126e+01 
R8451t5669 n8452 n5670 R=2.046e+01 
R8451t3373 n8452 n3374 R=6.473e+00 
R8451t3036 n8452 n3037 R=6.330e+00 
R8451t1158 n8452 n1159 R=1.364e+01 
R8451t12 n8452 n13 R=9.540e+00 
R8452t2990 n8453 n2991 R=1.535e+01 
R8452t5020 n8453 n5021 R=3.254e+00 
R8452t5063 n8453 n5064 R=7.846e+00 
R8452t7709 n8453 n7710 R=7.422e+00 
R8452t1399 n8453 n1400 R=7.117e+00 
R8453t2037 n8454 n2038 R=1.944e+01 
R8453t2171 n8454 n2172 R=3.781e+00 
R8453t2577 n8454 n2578 R=2.803e+02 
R8453t1662 n8454 n1663 R=3.086e+00 
R8453t3042 n8454 n3043 R=2.289e+01 
R8453t3685 n8454 n3686 R=6.573e+00 
R8454t2224 n8455 n2225 R=3.033e+00 
R8454t2065 n8455 n2066 R=3.402e+01 
R8454t3019 n8455 n3020 R=1.061e+01 
R8454t4490 n8455 n4491 R=1.626e+02 
R8454t612 n8455 n613 R=9.237e+00 
R8454t6274 n8455 n6275 R=3.102e+02 
R8454t2079 n8455 n2080 R=2.700e+00 
R8455t812 n8456 n813 R=1.586e+01 
R8455t2332 n8456 n2333 R=4.879e+00 
R8455t1693 n8456 n1694 R=4.025e+00 
R8455t7585 n8456 n7586 R=7.265e+01 
R8455t5621 n8456 n5622 R=2.461e+00 
R8456t2939 n8457 n2940 R=2.525e+00 
R8456t1256 n8457 n1257 R=1.564e+01 
R8456t3376 n8457 n3377 R=9.389e+00 
R8456t2945 n8457 n2946 R=1.280e+01 
R8457t2411 n8458 n2412 R=1.428e+02 
R8457t6576 n8458 n6577 R=3.106e+00 
R8457t2746 n8458 n2747 R=1.878e+02 
R8457t3662 n8458 n3663 R=3.216e+00 
R8457t359 n8458 n360 R=2.635e+02 
R8457t2880 n8458 n2881 R=9.127e+00 
R8457t5031 n8458 n5032 R=5.017e+01 
R8457t4282 n8458 n4283 R=1.161e+01 
R8457t3921 n8458 n3922 R=2.082e+01 
R8458t7459 n8459 n7460 R=7.225e+00 
R8458t7817 n8459 n7818 R=4.617e+00 
R8458t4684 n8459 n4685 R=1.247e+01 
R8458t3100 n8459 n3101 R=5.431e+00 
R8458t2353 n8459 n2354 R=1.797e+02 
R8458t5694 n8459 n5695 R=1.452e+01 
R8458t6459 n8459 n6460 R=1.850e+01 
R8459t2188 n8460 n2189 R=2.610e+00 
R8459t3652 n8460 n3653 R=2.104e+01 
R8459t7435 n8460 n7436 R=2.924e+00 
R8459t3953 n8460 n3954 R=2.357e+01 
R8460t50 n8461 n51 R=2.445e+00 
R8460t4421 n8461 n4422 R=2.145e+01 
R8460t4386 n8461 n4387 R=6.433e+00 
R8460t7706 n8461 n7707 R=5.270e+00 
R8460t5545 n8461 n5546 R=1.537e+01 
R8460t757 n8461 n758 R=1.953e+01 
R8461t1215 n8462 n1216 R=6.162e+00 
R8461t2896 n8462 n2897 R=2.742e+00 
R8461t7557 n8462 n7558 R=4.096e+00 
R8461t1272 n8462 n1273 R=1.046e+01 
R8462t4269 n8463 n4270 R=2.212e+01 
R8462t5927 n8463 n5928 R=1.895e+01 
R8462t5937 n8463 n5938 R=4.793e+00 
R8462t3469 n8463 n3470 R=3.207e+01 
R8462t5012 n8463 n5013 R=1.370e+01 
R8462t2911 n8463 n2912 R=5.555e+00 
R8462t3555 n8463 n3556 R=1.403e+01 
R8462t358 n8463 n359 R=7.776e+01 
R8462t5127 n8463 n5128 R=6.041e+00 
R8463t1911 n8464 n1912 R=1.539e+01 
R8463t6532 n8464 n6533 R=4.416e+00 
R8463t37 n8464 n38 R=5.792e+00 
R8464t2892 n8465 n2893 R=4.386e+00 
R8464t3277 n8465 n3278 R=3.313e+00 
R8464t7663 n8465 n7664 R=2.503e+02 
R8464t5795 n8465 n5796 R=8.409e+00 
R8464t2464 n8465 n2465 R=4.242e+00 
R8465t5812 n8466 n5813 R=4.464e+00 
R8465t8134 n8466 n8135 R=1.381e+01 
R8465t4902 n8466 n4903 R=2.404e+00 
R8465t7792 n8466 n7793 R=1.283e+02 
R8465t1065 n8466 n1066 R=3.760e+00 
R8465t1803 n8466 n1804 R=3.705e+02 
R8466t95 n8467 n96 R=1.956e+01 
R8466t699 n8467 n700 R=2.844e+01 
R8466t5624 n8467 n5625 R=1.464e+01 
R8466t5778 n8467 n5779 R=1.538e+02 
R8466t2913 n8467 n2914 R=2.808e+00 
R8466t5466 n8467 n5467 R=2.999e+00 
R8467t45 n8468 n46 R=4.874e+00 
R8467t2951 n8468 n2952 R=2.297e+01 
R8467t2888 n8468 n2889 R=6.828e+00 
R8467t4142 n8468 n4143 R=1.071e+01 
R8467t3457 n8468 n3458 R=4.291e+00 
R8468t2322 n8469 n2323 R=7.627e+00 
R8468t6880 n8469 n6881 R=4.142e+00 
R8468t7011 n8469 n7012 R=9.777e+00 
R8468t364 n8469 n365 R=3.305e+00 
R8468t6005 n8469 n6006 R=3.724e+03 
R8469t547 n8470 n548 R=6.001e+00 
R8469t8052 n8470 n8053 R=3.462e+00 
R8469t1467 n8470 n1468 R=7.250e+00 
R8469t1415 n8470 n1416 R=4.250e+01 
R8469t4105 n8470 n4106 R=4.269e+00 
R8470t3327 n8471 n3328 R=2.256e+01 
R8470t7005 n8471 n7006 R=3.324e+00 
R8470t1547 n8471 n1548 R=9.769e+00 
R8470t8446 n8471 n8447 R=8.914e+00 
R8470t6262 n8471 n6263 R=4.991e+00 
R8470t870 n8471 n871 R=5.218e+01 
R8471t2949 n8472 n2950 R=6.729e+00 
R8471t6010 n8472 n6011 R=9.385e+00 
R8471t7199 n8472 n7200 R=1.133e+01 
R8471t4287 n8472 n4288 R=1.820e+01 
R8471t1250 n8472 n1251 R=3.038e+01 
R8471t1515 n8472 n1516 R=3.404e+00 
R8472t6323 n8473 n6324 R=6.310e+00 
R8472t6456 n8473 n6457 R=1.930e+01 
R8472t430 n8473 n431 R=2.877e+00 
R8472t1448 n8473 n1449 R=8.670e+01 
R8472t7890 n8473 n7891 R=4.108e+00 
R8473t2336 n8474 n2337 R=7.848e+01 
R8473t3309 n8474 n3310 R=1.415e+01 
R8473t349 n8474 n350 R=6.464e+00 
R8473t7605 n8474 n7606 R=3.694e+01 
R8473t3986 n8474 n3987 R=5.330e+00 
R8473t140 n8474 n141 R=3.854e+00 
R8473t6627 n8474 n6628 R=2.181e+01 
R8474t4518 n8475 n4519 R=6.352e+00 
R8474t7581 n8475 n7582 R=5.427e+01 
R8474t8344 n8475 n8345 R=3.395e+01 
R8474t2326 n8475 n2327 R=3.872e+00 
R8474t2831 n8475 n2832 R=8.604e+00 
R8474t7131 n8475 n7132 R=3.162e+00 
R8475t2025 n8476 n2026 R=5.823e+00 
R8475t5195 n8476 n5196 R=4.793e+01 
R8475t691 n8476 n692 R=5.285e+00 
R8475t5233 n8476 n5234 R=1.651e+01 
R8475t6619 n8476 n6620 R=4.525e+00 
R8475t6354 n8476 n6355 R=5.278e+00 
R8475t8261 n8476 n8262 R=1.185e+02 
R8476t5256 n8477 n5257 R=1.521e+01 
R8476t6136 n8477 n6137 R=1.920e+01 
R8476t2029 n8477 n2030 R=5.535e+00 
R8477t5699 n8478 n5700 R=2.668e+00 
R8477t8085 n8478 n8086 R=3.261e+00 
R8477t3224 n8478 n3225 R=1.376e+01 
R8478t5208 n8479 n5209 R=2.463e+00 
R8478t5745 n8479 n5746 R=5.958e+00 
R8478t194 n8479 n195 R=6.306e+00 
R8479t544 n8480 n545 R=5.656e+00 
R8479t4180 n8480 n4181 R=6.178e+00 
R8479t1953 n8480 n1954 R=5.905e+00 
R8479t5698 n8480 n5699 R=1.242e+01 
R8479t4142 n8480 n4143 R=2.723e+02 
R8479t2888 n8480 n2889 R=6.810e+00 
R8480t1910 n8481 n1911 R=6.899e+00 
R8480t7716 n8481 n7717 R=8.876e+00 
R8480t2639 n8481 n2640 R=1.551e+01 
R8480t1794 n8481 n1795 R=6.612e+00 
R8480t7962 n8481 n7963 R=1.193e+01 
R8480t535 n8481 n536 R=3.422e+01 
R8481t2606 n8482 n2607 R=1.743e+01 
R8481t4139 n8482 n4140 R=2.586e+00 
R8481t1040 n8482 n1041 R=6.142e+00 
R8481t2435 n8482 n2436 R=1.849e+01 
R8481t5755 n8482 n5756 R=5.030e+00 
R8481t4842 n8482 n4843 R=6.693e+00 
R8482t826 n8483 n827 R=1.298e+02 
R8482t6137 n8483 n6138 R=6.429e+00 
R8482t2508 n8483 n2509 R=1.848e+00 
R8482t4856 n8483 n4857 R=2.404e+01 
R8482t1353 n8483 n1354 R=3.221e+00 
R8483t4677 n8484 n4678 R=4.502e+01 
R8483t5346 n8484 n5347 R=2.728e+00 
R8483t7538 n8484 n7539 R=4.421e+01 
R8483t8039 n8484 n8040 R=8.794e+00 
R8483t367 n8484 n368 R=8.840e+02 
R8483t6667 n8484 n6668 R=2.698e+00 
R8483t3409 n8484 n3410 R=7.582e+01 
R8483t7276 n8484 n7277 R=1.382e+01 
R8483t5938 n8484 n5939 R=5.548e+01 
R8484t4344 n8485 n4345 R=3.788e+01 
R8484t6774 n8485 n6775 R=4.969e+00 
R8484t6247 n8485 n6248 R=6.397e+00 
R8484t5337 n8485 n5338 R=4.208e+00 
R8484t1915 n8485 n1916 R=1.692e+01 
R8485t883 n8486 n884 R=1.959e+01 
R8485t3535 n8486 n3536 R=8.081e+00 
R8485t6806 n8486 n6807 R=2.720e+00 
R8485t1815 n8486 n1816 R=1.297e+01 
R8485t3256 n8486 n3257 R=5.322e+00 
R8486t89 n8487 n90 R=1.181e+01 
R8486t3416 n8487 n3417 R=2.576e+00 
R8486t6995 n8487 n6996 R=5.398e+01 
R8486t154 n8487 n155 R=1.391e+01 
R8487t1536 n8488 n1537 R=8.892e+00 
R8487t5622 n8488 n5623 R=1.179e+01 
R8487t4645 n8488 n4646 R=2.873e+01 
R8487t7717 n8488 n7718 R=3.160e+00 
R8487t4604 n8488 n4605 R=8.829e+00 
R8487t7245 n8488 n7246 R=6.919e+00 
R8488t2821 n8489 n2822 R=1.041e+01 
R8488t3902 n8489 n3903 R=7.467e+00 
R8488t3933 n8489 n3934 R=1.250e+01 
R8488t5445 n8489 n5446 R=3.011e+01 
R8488t2593 n8489 n2594 R=3.905e+00 
R8488t1280 n8489 n1281 R=2.343e+01 
R8488t6397 n8489 n6398 R=9.315e+00 
R8489t929 n8490 n930 R=3.561e+00 
R8489t3141 n8490 n3142 R=2.740e+01 
R8489t3861 n8490 n3862 R=3.978e+00 
R8489t835 n8490 n836 R=7.877e+00 
R8489t7193 n8490 n7194 R=1.515e+01 
R8489t3045 n8490 n3046 R=1.306e+01 
R8490t211 n8491 n212 R=3.565e+00 
R8490t808 n8491 n809 R=4.207e+01 
R8490t7841 n8491 n7842 R=4.460e+00 
R8490t1868 n8491 n1869 R=1.280e+01 
R8490t366 n8491 n367 R=5.588e+00 
R8490t2818 n8491 n2819 R=6.876e+01 
R8491t1707 n8492 n1708 R=1.318e+01 
R8491t6551 n8492 n6552 R=3.292e+00 
R8491t6188 n8492 n6189 R=1.104e+01 
R8491t4262 n8492 n4263 R=8.427e+00 
R8491t587 n8492 n588 R=3.294e+01 
R8492t3624 n8493 n3625 R=8.338e+00 
R8492t5784 n8493 n5785 R=2.932e+00 
R8492t4164 n8493 n4165 R=5.114e+00 
R8492t2624 n8493 n2625 R=5.795e+00 
R8493t2648 n8494 n2649 R=3.621e+01 
R8493t6778 n8494 n6779 R=5.034e+00 
R8493t3024 n8494 n3025 R=2.444e+01 
R8493t6243 n8494 n6244 R=1.129e+01 
R8493t6039 n8494 n6040 R=5.280e+00 
R8493t5042 n8494 n5043 R=4.889e+00 
R8494t2547 n8495 n2548 R=6.265e+00 
R8494t3911 n8495 n3912 R=7.137e+00 
R8494t2178 n8495 n2179 R=4.832e+00 
R8494t5967 n8495 n5968 R=1.271e+01 
R8494t3551 n8495 n3552 R=4.766e+00 
R8494t3073 n8495 n3074 R=3.167e+01 
R8495t1933 n8496 n1934 R=8.511e+00 
R8495t6166 n8496 n6167 R=1.757e+01 
R8495t6565 n8496 n6566 R=5.641e+00 
R8495t5098 n8496 n5099 R=7.537e+00 
R8495t1739 n8496 n1740 R=7.141e+00 
R8496t6577 n8497 n6578 R=1.064e+01 
R8496t8071 n8497 n8072 R=3.468e+00 
R8496t7400 n8497 n7401 R=2.491e+00 
R8496t5449 n8497 n5450 R=1.877e+02 
R8497t5000 n8498 n5001 R=9.811e+01 
R8497t6055 n8498 n6056 R=3.987e+01 
R8497t6348 n8498 n6349 R=3.154e+00 
R8497t1489 n8498 n1490 R=1.647e+01 
R8497t6326 n8498 n6327 R=4.812e+00 
R8497t7593 n8498 n7594 R=2.519e+01 
R8497t6529 n8498 n6530 R=5.047e+00 
R8498t4213 n8499 n4214 R=1.573e+00 
R8498t4675 n8499 n4676 R=4.050e+01 
R8498t6601 n8499 n6602 R=3.063e+00 
R8498t1672 n8499 n1673 R=8.346e+00 
R8498t3163 n8499 n3164 R=3.196e+01 
R8498t2271 n8499 n2272 R=8.268e+01 
R8499t5787 n1 n5788 R=1.176e+01 
R8499t1787 n1 n1788 R=6.388e+00 
R8500t5141 n8501 n5142 R=9.996e+00 
R8500t2927 n8501 n2928 R=8.791e+01 
R8500t510 n8501 n511 R=9.173e+00 
R8500t8006 n8501 n8007 R=3.299e+00 
R8500t1767 n8501 n1768 R=2.269e+02 
R8500t3043 n8501 n3044 R=4.590e+00 
R8501t5046 n8502 n5047 R=3.726e+00 
R8501t6757 n8502 n6758 R=1.382e+02 
R8501t3149 n8502 n3150 R=3.729e+00 
R8501t4469 n8502 n4470 R=8.524e+00 
R8502t1679 n8503 n1680 R=8.965e+00 
R8502t5805 n8503 n5806 R=3.645e+00 
R8502t2367 n8503 n2368 R=4.536e+00 
R8502t8369 n8503 n8370 R=5.884e+00 
R8503t3193 n8504 n3194 R=6.827e+00 
R8503t1422 n8504 n1423 R=3.862e+00 
R8504t4552 n8505 n4553 R=8.381e+00 
R8504t5237 n8505 n5238 R=1.760e+01 
R8504t7129 n8505 n7130 R=5.002e+00 
R8505t5745 n8506 n5746 R=1.461e+01 
R8505t6480 n8506 n6481 R=3.423e+00 
R8505t8478 n8506 n8479 R=2.628e+01 
R8505t5208 n8506 n5209 R=7.928e+00 
R8505t4030 n8506 n4031 R=1.394e+01 
R8505t6245 n8506 n6246 R=2.041e+01 
R8505t1244 n8506 n1245 R=5.736e+01 
R8505t1606 n8506 n1607 R=7.399e+00 
R8506t4948 n8507 n4949 R=4.746e+00 
R8506t5961 n8507 n5962 R=2.715e+01 
R8506t6259 n8507 n6260 R=3.586e+01 
R8506t5098 n8507 n5099 R=3.454e+00 
R8506t8495 n8507 n8496 R=3.037e+01 
R8506t6565 n8507 n6566 R=7.122e+00 
R8506t2403 n8507 n2404 R=8.096e+01 
R8507t2523 n8508 n2524 R=4.949e+00 
R8507t199 n8508 n200 R=4.842e+00 
R8507t1253 n8508 n1254 R=1.231e+01 
R8507t804 n8508 n805 R=1.118e+01 
R8508t3992 n8509 n3993 R=5.891e+00 
R8508t4300 n8509 n4301 R=6.583e+01 
R8508t1217 n8509 n1218 R=1.523e+02 
R8508t3801 n8509 n3802 R=7.592e+00 
R8508t7675 n8509 n7676 R=3.718e+00 
R8508t4505 n8509 n4506 R=2.678e+01 
R8509t5135 n8510 n5136 R=8.391e+00 
R8509t5774 n8510 n5775 R=9.399e+00 
R8509t558 n8510 n559 R=3.240e+00 
R8509t2291 n8510 n2292 R=1.010e+01 
R8509t476 n8510 n477 R=6.204e+00 
R8510t1228 n8511 n1229 R=1.313e+01 
R8510t8393 n8511 n8394 R=4.170e+00 
R8510t3688 n8511 n3689 R=2.856e+01 
R8510t2519 n8511 n2520 R=4.680e+00 
R8511t8017 n8512 n8018 R=5.762e+00 
R8511t1412 n8512 n1413 R=4.368e+01 
R8511t2308 n8512 n2309 R=7.238e+00 
R8511t3708 n8512 n3709 R=4.981e+01 
R8511t2977 n8512 n2978 R=1.218e+01 
R8512t1955 n8513 n1956 R=1.429e+01 
R8512t5216 n8513 n5217 R=7.699e+00 
R8512t4464 n8513 n4465 R=4.635e+00 
R8512t2221 n8513 n2222 R=4.728e+01 
R8512t3808 n8513 n3809 R=2.431e+00 
R8513t5956 n8514 n5957 R=1.174e+01 
R8513t6905 n8514 n6906 R=7.924e+00 
R8513t420 n8514 n421 R=8.093e+00 
R8513t2852 n8514 n2853 R=5.783e+00 
R8513t7054 n8514 n7055 R=7.179e+00 
R8514t4604 n8515 n4605 R=4.030e+01 
R8514t571 n8515 n572 R=3.360e+00 
R8514t5676 n8515 n5677 R=8.033e+00 
R8514t7380 n8515 n7381 R=2.973e+00 
R8515t8476 n8516 n8477 R=6.798e+00 
R8515t2029 n8516 n2030 R=3.000e+01 
R8515t6726 n8516 n6727 R=4.411e+02 
R8515t5626 n8516 n5627 R=5.702e+00 
R8516t5532 n8517 n5533 R=7.822e+00 
R8516t5720 n8517 n5721 R=1.827e+02 
R8516t6375 n8517 n6376 R=1.097e+01 
R8516t6604 n8517 n6605 R=8.080e+00 
R8517t3234 n8518 n3235 R=2.450e+01 
R8517t7267 n8518 n7268 R=3.351e+01 
R8517t2835 n8518 n2836 R=1.811e+00 
R8517t8411 n8518 n8412 R=1.165e+01 
R8517t2575 n8518 n2576 R=2.036e+01 
R8517t6304 n8518 n6305 R=2.341e+00 
R8518t5535 n8519 n5536 R=6.615e+00 
R8518t2455 n8519 n2456 R=3.180e+00 
R8518t212 n8519 n213 R=1.106e+01 
R8519t3228 n8520 n3229 R=2.798e+00 
R8519t3995 n8520 n3996 R=5.274e+01 
R8519t5089 n8520 n5090 R=5.463e+00 
R8519t2150 n8520 n2151 R=6.396e+00 
R8519t4028 n8520 n4029 R=5.224e+00 
R8520t7885 n8521 n7886 R=1.133e+01 
R8520t1855 n8521 n1856 R=3.621e+00 
R8520t6399 n8521 n6400 R=2.105e+01 
R8520t8305 n8521 n8306 R=5.164e+03 
R8520t307 n8521 n308 R=5.606e+01 
R8520t7172 n8521 n7173 R=4.733e+00 
R8520t3217 n8521 n3218 R=4.814e+00 
R8521t180 n8522 n181 R=4.544e+00 
R8521t7281 n8522 n7282 R=1.887e+02 
R8521t2341 n8522 n2342 R=5.925e+00 
R8521t6346 n8522 n6347 R=1.758e+01 
R8521t6320 n8522 n6321 R=2.985e+01 
R8521t4027 n8522 n4028 R=2.426e+01 
R8521t5347 n8522 n5348 R=4.775e+00 
R8522t7566 n8523 n7567 R=1.614e+01 
R8522t1556 n8523 n1557 R=2.786e+00 
R8523t7138 n8524 n7139 R=2.690e+01 
R8523t4362 n8524 n4363 R=5.420e+01 
R8523t3342 n8524 n3343 R=2.686e+00 
R8524t2419 n8525 n2420 R=6.789e+00 
R8524t2699 n8525 n2700 R=2.591e+01 
R8524t5529 n8525 n5530 R=8.866e+00 
R8524t5045 n8525 n5046 R=1.497e+01 
R8524t3590 n8525 n3591 R=2.138e+01 
R8525t1385 n8526 n1386 R=2.451e+01 
R8525t2599 n8526 n2600 R=4.979e+00 
R8525t4303 n8526 n4304 R=6.331e+00 
R8525t2041 n8526 n2042 R=4.571e+01 
R8525t6053 n8526 n6054 R=2.161e+01 
R8525t4281 n8526 n4282 R=6.794e+00 
R8525t7385 n8526 n7386 R=3.934e+00 
R8526t3298 n8527 n3299 R=1.212e+01 
R8526t5454 n8527 n5455 R=2.325e+01 
R8526t3222 n8527 n3223 R=7.302e+00 
R8526t5168 n8527 n5169 R=2.435e+01 
R8526t7482 n8527 n7483 R=1.200e+01 
R8526t8111 n8527 n8112 R=7.249e+00 
R8526t4881 n8527 n4882 R=8.736e+00 
R8527t1566 n8528 n1567 R=1.165e+01 
R8527t4129 n8528 n4130 R=3.639e+00 
R8527t2372 n8528 n2373 R=5.280e+01 
R8527t1359 n8528 n1360 R=1.582e+01 
R8527t2730 n8528 n2731 R=6.794e+00 
R8528t4198 n8529 n4199 R=1.483e+01 
R8528t6113 n8529 n6114 R=2.906e+01 
R8528t5804 n8529 n5805 R=1.253e+01 
R8528t1906 n8529 n1907 R=9.978e+03 
R8528t5114 n8529 n5115 R=2.624e+00 
R8528t6818 n8529 n6819 R=2.820e+01 
R8528t7854 n8529 n7855 R=1.613e+01 
R8528t593 n8529 n594 R=1.812e+01 
R8528t2720 n8529 n2721 R=1.055e+01 
R8529t1342 n8530 n1343 R=4.777e+00 
R8529t3438 n8530 n3439 R=8.825e+00 
R8529t4979 n8530 n4980 R=2.937e+01 
R8529t7399 n8530 n7400 R=1.418e+01 
R8529t3360 n8530 n3361 R=2.942e+00 
R8530t2970 n8531 n2971 R=3.871e+02 
R8530t7344 n8531 n7345 R=4.284e+00 
R8530t837 n8531 n838 R=7.068e+00 
R8530t1070 n8531 n1071 R=2.856e+01 
R8530t537 n8531 n538 R=6.496e+00 
R8530t3098 n8531 n3099 R=7.377e+00 
R8531t4347 n8532 n4348 R=6.010e+00 
R8531t7308 n8532 n7309 R=5.493e+00 
R8531t777 n8532 n778 R=1.111e+01 
R8531t1509 n8532 n1510 R=5.528e+01 
R8531t1417 n8532 n1418 R=1.182e+01 
R8531t2204 n8532 n2205 R=3.833e+00 
R8531t3142 n8532 n3143 R=1.464e+01 
R8531t3157 n8532 n3158 R=1.207e+02 
R8532t2348 n8533 n2349 R=5.425e+01 
R8532t3263 n8533 n3264 R=1.019e+01 
R8532t2611 n8533 n2612 R=1.097e+01 
R8532t4871 n8533 n4872 R=9.773e+00 
R8532t5026 n8533 n5027 R=2.074e+01 
R8532t3354 n8533 n3355 R=8.035e+00 
R8532t513 n8533 n514 R=3.823e+00 
R8533t735 n8534 n736 R=1.101e+01 
R8533t6486 n8534 n6487 R=1.043e+01 
R8533t2916 n8534 n2917 R=1.996e+01 
R8533t8253 n8534 n8254 R=1.996e+01 
R8533t5414 n8534 n5415 R=8.531e+01 
R8533t3974 n8534 n3975 R=6.006e+00 
R8533t7418 n8534 n7419 R=1.582e+01 
R8534t2051 n8535 n2052 R=7.602e+00 
R8534t3269 n8535 n3270 R=1.116e+01 
R8534t529 n8535 n530 R=4.190e+00 
R8534t3592 n8535 n3593 R=1.383e+01 
R8534t5958 n8535 n5959 R=4.807e+00 
R8535t684 n8536 n685 R=1.625e+01 
R8535t5985 n8536 n5986 R=8.133e+00 
R8535t6264 n8536 n6265 R=1.965e+01 
R8535t7939 n8536 n7940 R=5.020e+00 
R8535t2849 n8536 n2850 R=6.275e+00 
R8535t6530 n8536 n6531 R=3.852e+01 
R8535t7695 n8536 n7696 R=3.899e+00 
R8536t3773 n8537 n3774 R=6.048e+00 
R8536t7783 n8537 n7784 R=1.005e+01 
R8536t5060 n8537 n5061 R=8.167e+00 
R8536t5014 n8537 n5015 R=1.819e+01 
R8536t8295 n8537 n8296 R=1.359e+01 
R8536t5439 n8537 n5440 R=3.458e+01 
R8536t6359 n8537 n6360 R=7.999e+00 
R8537t686 n8538 n687 R=4.101e+00 
R8537t8089 n8538 n8090 R=6.986e+00 
R8537t3747 n8538 n3748 R=4.323e+00 
R8537t4971 n8538 n4972 R=6.749e+00 
R8537t4477 n8538 n4478 R=2.900e+01 
R8538t1895 n8539 n1896 R=1.454e+00 
R8538t4683 n8539 n4684 R=5.687e+01 
R8538t5819 n8539 n5820 R=7.036e+00 
R8538t7008 n8539 n7009 R=3.800e+00 
R8538t8016 n8539 n8017 R=1.185e+01 
R8538t437 n8539 n438 R=1.411e+02 
R8539t3052 n8540 n3053 R=4.515e+00 
R8539t7295 n8540 n7296 R=3.595e+00 
R8539t6333 n8540 n6334 R=2.514e+01 
R8540t24 n8541 n25 R=1.544e+00 
R8540t4190 n8541 n4191 R=4.324e+00 
R8541t5261 n8542 n5262 R=2.286e+01 
R8541t5378 n8542 n5379 R=1.084e+01 
R8541t4944 n8542 n4945 R=2.504e+00 
R8541t6123 n8542 n6124 R=2.139e+03 
R8541t1745 n8542 n1746 R=4.439e+01 
R8541t4886 n8542 n4887 R=2.405e+00 
R8541t8078 n8542 n8079 R=1.615e+01 
R8542t152 n8543 n153 R=2.285e+01 
R8542t6851 n8543 n6852 R=1.185e+01 
R8542t6060 n8543 n6061 R=3.955e+00 
R8542t4841 n8543 n4842 R=1.574e+01 
R8542t2365 n8543 n2366 R=1.955e+01 
R8542t4579 n8543 n4580 R=1.748e+01 
R8542t5516 n8543 n5517 R=3.055e+00 
R8543t261 n8544 n262 R=1.060e+01 
R8543t1535 n8544 n1536 R=6.270e+00 
R8543t7626 n8544 n7627 R=2.210e+01 
R8543t1738 n8544 n1739 R=7.530e+00 
R8543t1914 n8544 n1915 R=8.318e+00 
R8543t1497 n8544 n1498 R=4.599e+00 
R8544t1234 n8545 n1235 R=7.098e+00 
R8544t8040 n8545 n8041 R=4.821e+00 
R8544t1828 n8545 n1829 R=3.143e+00 
R8544t2087 n8545 n2088 R=2.328e+01 
R8544t6447 n8545 n6448 R=6.503e+00 
R8545t1996 n8546 n1 R=5.575e+00 
R8545t6469 n8546 n1 R=1.442e+01 
R8545t8499 n8546 n1 R=6.341e+00 
R8545t1787 n8546 n1788 R=2.430e+01 
R8545t5330 n8546 n5331 R=4.281e+00 
R8546t827 n8547 n828 R=8.846e+01 
R8546t3625 n8547 n3626 R=2.316e+00 
R8546t6176 n8547 n6177 R=1.255e+01 
R8546t3691 n8547 n3692 R=2.520e+00 
R8546t6127 n8547 n6128 R=1.574e+01 
R8547t3824 n8548 n3825 R=1.836e+01 
R8547t4698 n8548 n4699 R=5.799e+00 
R8547t3818 n8548 n3819 R=3.796e+00 
R8547t5181 n8548 n5182 R=4.019e+00 
R8547t4881 n8548 n4882 R=1.878e+01 
R8548t8165 n8549 n8166 R=1.556e+01 
R8548t2574 n8549 n2575 R=4.338e+00 
R8549t5168 n8550 n5169 R=9.455e+00 
R8549t8526 n8550 n8527 R=1.169e+01 
R8549t3222 n8550 n3223 R=6.100e+00 
R8549t1435 n8550 n1436 R=1.634e+01 
R8549t3189 n8550 n3190 R=1.098e+01 
R8549t4991 n8550 n4992 R=6.031e+00 
R8550t3188 n8551 n3189 R=8.286e+00 
R8550t5605 n8551 n5606 R=2.316e+00 
R8550t4890 n8551 n4891 R=3.514e+02 
R8550t8357 n8551 n8358 R=1.343e+01 
R8550t4771 n8551 n4772 R=8.581e+00 
R8551t950 n8552 n951 R=6.582e+00 
R8551t559 n8552 n560 R=1.942e+01 
R8551t5538 n8552 n5539 R=7.391e+00 
R8552t6998 n8553 n6999 R=9.995e+00 
R8552t4444 n8553 n4445 R=1.790e+01 
R8552t4998 n8553 n4999 R=4.693e+00 
R8552t7141 n8553 n7142 R=2.196e+01 
R8552t7914 n8553 n7915 R=1.068e+01 
R8552t8170 n8553 n8171 R=3.039e+00 
R8553t980 n8554 n981 R=1.375e+02 
R8553t1074 n8554 n1075 R=5.285e+00 
R8553t3103 n8554 n3104 R=2.686e+01 
R8553t3899 n8554 n3900 R=1.052e+01 
R8553t993 n8554 n994 R=9.994e+00 
R8554t7176 n1 n7177 R=1.813e+01 
R8554t3366 n1 n3367 R=5.321e+00 
R8554t3455 n1 n3456 R=3.674e+01 
R8555t2425 n8556 n2426 R=4.573e+01 
R8555t7944 n8556 n7945 R=8.752e+00 
R8555t3999 n8556 n4000 R=5.657e+00 
R8555t2119 n8556 n2120 R=5.103e+00 
R8555t6237 n8556 n6238 R=2.082e+02 
R8555t4769 n8556 n4770 R=8.821e+00 
R8556t4205 n8557 n4206 R=3.007e+00 
R8556t363 n8557 n364 R=3.752e+01 
R8556t2870 n8557 n2871 R=7.846e+00 
R8556t2033 n8557 n2034 R=1.199e+01 
R8556t3604 n8557 n3605 R=1.157e+01 
R8557t1126 n8558 n1127 R=1.435e+01 
R8557t8260 n8558 n8261 R=5.102e+00 
R8557t7374 n8558 n7375 R=1.944e+01 
R8558t1551 n8559 n1552 R=3.125e+00 
R8558t1806 n8559 n1807 R=2.253e+01 
R8558t367 n8559 n368 R=3.602e+01 
R8558t7109 n8559 n7110 R=1.853e+01 
R8558t2003 n8559 n2004 R=6.792e+00 
R8558t4143 n8559 n4144 R=1.703e+01 
R8558t3885 n8559 n3886 R=3.473e+00 
R8559t4781 n8560 n4782 R=8.078e+01 
R8559t7029 n8560 n7030 R=5.637e+00 
R8559t5634 n8560 n5635 R=2.923e+01 
R8559t5371 n8560 n5372 R=3.267e+00 
R8559t6147 n8560 n6148 R=4.046e+00 
R8559t1719 n8560 n1720 R=1.429e+01 
R8560t4646 n8561 n4647 R=2.969e+02 
R8560t5547 n8561 n5548 R=3.008e+01 
R8560t2939 n8561 n2940 R=3.115e+01 
R8560t8456 n8561 n8457 R=3.432e+00 
R8560t1256 n8561 n1257 R=6.820e+01 
R8560t4016 n8561 n4017 R=5.111e+00 
R8560t1873 n8561 n1874 R=1.254e+01 
R8560t6222 n8561 n6223 R=5.005e+01 
R8560t6799 n8561 n6800 R=9.308e+01 
R8561t3211 n8562 n3212 R=4.787e+01 
R8561t4977 n8562 n4978 R=8.522e+00 
R8561t6386 n8562 n6387 R=4.018e+00 
R8561t3148 n8562 n3149 R=5.898e+00 
R8561t1066 n8562 n1067 R=8.831e+00 
R8561t1845 n8562 n1846 R=9.531e+00 
R8562t854 n8563 n855 R=3.124e+01 
R8562t8202 n8563 n8203 R=1.326e+01 
R8562t8215 n8563 n8216 R=5.757e+01 
R8562t2959 n8563 n2960 R=4.842e+00 
R8563t1946 n8564 n1947 R=5.700e+00 
R8563t2270 n8564 n2271 R=1.939e+01 
R8563t519 n8564 n520 R=5.231e+01 
R8563t5023 n8564 n5024 R=3.066e+00 
R8563t5355 n8564 n5356 R=8.206e+00 
R8563t2642 n8564 n2643 R=2.491e+01 
R8563t5949 n8564 n5950 R=1.901e+01 
R8564t4039 n8565 n4040 R=2.540e+01 
R8564t5294 n8565 n5295 R=3.381e+00 
R8564t1810 n8565 n1811 R=5.571e+00 
R8564t6515 n8565 n6516 R=2.580e+01 
R8564t6061 n8565 n6062 R=1.764e+01 
R8564t4603 n8565 n4604 R=5.572e+00 
R8564t6643 n8565 n6644 R=1.184e+03 
R8565t642 n8566 n643 R=7.481e+00 
R8565t5162 n8566 n5163 R=5.558e+01 
R8565t1499 n8566 n1500 R=3.506e+00 
R8565t8405 n8566 n8406 R=1.871e+01 
R8565t1176 n8566 n1177 R=8.907e+01 
R8565t881 n8566 n882 R=2.886e+00 
R8565t3082 n8566 n3083 R=2.167e+01 
R8566t2891 n8567 n2892 R=1.357e+01 
R8566t4882 n8567 n4883 R=2.512e+01 
R8566t715 n8567 n716 R=6.990e+00 
R8566t4707 n8567 n4708 R=4.343e+00 
R8566t6838 n8567 n6839 R=5.426e+02 
R8566t7021 n8567 n7022 R=6.121e+00 
R8566t6236 n8567 n6237 R=5.414e+00 
R8567t2203 n8568 n2204 R=4.475e+00 
R8567t6771 n8568 n6772 R=1.130e+03 
R8567t2654 n8568 n2655 R=4.757e+00 
R8567t5563 n8568 n5564 R=4.899e+01 
R8567t5120 n8568 n5121 R=1.871e+00 
R8567t8271 n8568 n8272 R=8.853e+01 
R8567t3630 n8568 n3631 R=3.311e+01 
R8568t4531 n8569 n4532 R=1.384e+02 
R8568t7843 n8569 n7844 R=2.844e+00 
R8568t450 n8569 n451 R=1.951e+01 
R8568t2696 n8569 n2697 R=1.465e+01 
R8568t7982 n8569 n7983 R=8.360e+00 
R8568t7697 n8569 n7698 R=8.767e+00 
R8568t2205 n8569 n2206 R=4.701e+01 
R8569t2202 n8570 n2203 R=5.186e+00 
R8569t7237 n8570 n7238 R=4.350e+00 
R8569t1926 n8570 n1927 R=1.603e+01 
R8569t651 n8570 n652 R=2.106e+01 
R8569t7229 n8570 n7230 R=3.675e+00 
R8570t1398 n8571 n1399 R=8.659e+00 
R8570t3541 n8571 n3542 R=2.969e+01 
R8570t8192 n8571 n8193 R=1.011e+01 
R8570t3374 n8571 n3375 R=1.294e+01 
R8570t2779 n8571 n2780 R=4.799e+00 
R8570t3559 n8571 n3560 R=4.281e+01 
R8571t3381 n8572 n3382 R=3.636e+00 
R8571t4672 n8572 n4673 R=1.173e+01 
R8571t5986 n8572 n5987 R=9.142e+00 
R8571t7489 n8572 n7490 R=1.765e+00 
R8571t8298 n8572 n8299 R=1.725e+01 
R8572t356 n8573 n357 R=4.328e+01 
R8572t5134 n8573 n5135 R=4.746e+00 
R8572t6234 n8573 n6235 R=5.422e+00 
R8572t7074 n8573 n7075 R=9.992e+00 
R8572t4293 n8573 n4294 R=5.309e+00 
R8573t3040 n8574 n3041 R=1.370e+01 
R8573t3262 n8574 n3263 R=7.481e+00 
R8573t7497 n8574 n7498 R=1.088e+02 
R8573t288 n8574 n289 R=1.883e+01 
R8573t1928 n8574 n1929 R=5.742e+00 
R8573t5590 n8574 n5591 R=2.689e+01 
R8573t337 n8574 n338 R=3.710e+01 
R8573t6657 n8574 n6658 R=5.892e+01 
R8573t1306 n8574 n1307 R=1.066e+01 
R8573t4035 n8574 n4036 R=6.596e+00 
R8574t4397 n8575 n4398 R=1.780e+01 
R8574t6159 n8575 n6160 R=3.124e+00 
R8574t333 n8575 n334 R=1.518e+01 
R8574t3148 n8575 n3149 R=5.900e+00 
R8574t6843 n8575 n6844 R=6.813e+00 
R8575t4697 n8576 n4698 R=4.618e+00 
R8575t6665 n8576 n6666 R=4.907e+00 
R8575t2925 n8576 n2926 R=3.673e+01 
R8575t3800 n8576 n3801 R=1.020e+02 
R8575t6443 n8576 n6444 R=3.816e+00 
R8575t8402 n8576 n8403 R=1.255e+02 
R8575t3621 n8576 n3622 R=1.399e+01 
R8576t2234 n8577 n2235 R=1.947e+00 
R8576t6499 n8577 n6500 R=2.506e+04 
R8576t2130 n8577 n2131 R=7.237e+00 
R8576t3825 n8577 n3826 R=4.697e+00 
R8576t4660 n8577 n4661 R=5.678e+00 
R8577t4546 n8578 n4547 R=1.877e+01 
R8577t7885 n8578 n7886 R=5.256e+01 
R8577t5687 n8578 n5688 R=2.763e+00 
R8577t5891 n8578 n5892 R=1.510e+01 
R8577t2120 n8578 n2121 R=1.953e+01 
R8577t1741 n8578 n1742 R=2.286e+01 
R8577t5751 n8578 n5752 R=3.292e+01 
R8577t5913 n8578 n5914 R=1.332e+01 
R8577t1855 n8578 n1856 R=1.395e+01 
R8577t8520 n8578 n8521 R=2.266e+01 
R8578t6381 n8579 n6382 R=5.960e+00 
R8578t6779 n8579 n6780 R=6.972e+01 
R8578t1361 n8579 n1362 R=3.950e+00 
R8578t7580 n8579 n7581 R=1.168e+02 
R8579t2783 n8580 n2784 R=2.695e+01 
R8579t2932 n8580 n2933 R=1.338e+01 
R8579t3995 n8580 n3996 R=4.219e+00 
R8579t6621 n8580 n6622 R=5.319e+02 
R8579t3676 n8580 n3677 R=5.093e+01 
R8579t7978 n8580 n7979 R=4.786e+00 
R8579t4990 n8580 n4991 R=1.519e+02 
R8580t1402 n8581 n1403 R=1.936e+01 
R8580t3123 n8581 n3124 R=4.731e+00 
R8580t5741 n8581 n5742 R=1.160e+01 
R8580t1342 n8581 n1343 R=5.521e+01 
R8580t8529 n8581 n8530 R=2.113e+01 
R8581t1342 n8582 n1343 R=3.971e+00 
R8581t5741 n8582 n5742 R=2.838e+00 
R8581t2342 n8582 n2343 R=7.248e+00 
R8582t3371 n8583 n3372 R=3.533e+02 
R8582t3278 n8583 n3279 R=4.762e+00 
R8582t7440 n8583 n7441 R=5.434e+01 
R8582t7103 n8583 n7104 R=6.287e+01 
R8582t5551 n8583 n5552 R=1.185e+02 
R8583t2891 n8584 n2892 R=3.343e+00 
R8583t4882 n8584 n4883 R=2.828e+00 
R8583t7597 n8584 n7598 R=8.277e+00 
R8583t1160 n8584 n1161 R=9.567e+01 
R8583t2324 n8584 n2325 R=1.040e+01 
R8584t3982 n8585 n3983 R=2.223e+01 
R8584t5744 n8585 n5745 R=1.220e+01 
R8584t8242 n8585 n8243 R=1.780e+01 
R8584t6515 n8585 n6516 R=5.116e+00 
R8584t5357 n8585 n5358 R=9.892e+00 
R8584t2787 n8585 n2788 R=1.130e+01 
R8584t3749 n8585 n3750 R=1.140e+01 
R8585t985 n8586 n986 R=3.498e+01 
R8585t6701 n8586 n6702 R=1.717e+00 
R8585t2016 n8586 n2017 R=3.330e+01 
R8585t1589 n8586 n1590 R=6.908e+00 
R8585t4806 n8586 n4807 R=6.053e+00 
R8586t392 n8587 n393 R=5.439e+00 
R8586t6536 n8587 n6537 R=2.676e+01 
R8586t1365 n8587 n1366 R=2.808e+00 
R8587t3329 n8588 n3330 R=6.062e+00 
R8587t7351 n8588 n7352 R=4.928e+00 
R8587t1087 n8588 n1088 R=2.371e+01 
R8587t5488 n8588 n5489 R=7.817e+00 
R8587t1134 n8588 n1135 R=1.448e+01 
R8587t116 n8588 n117 R=1.650e+02 
R8587t4575 n8588 n4576 R=5.179e+00 
R8588t2600 n8589 n2601 R=5.972e+00 
R8588t3421 n8589 n3422 R=1.361e+01 
R8588t3585 n8589 n3586 R=4.251e+00 
R8588t1541 n8589 n1542 R=2.508e+01 
R8589t5367 n8590 n5368 R=4.869e+00 
R8589t5671 n8590 n5672 R=4.753e+00 
R8589t2906 n8590 n2907 R=2.064e+01 
R8589t877 n8590 n878 R=3.628e+00 
R8589t5905 n8590 n5906 R=1.887e+01 
R8590t2049 n8591 n2050 R=1.793e+01 
R8590t7099 n8591 n7100 R=2.687e+00 
R8590t1190 n8591 n1191 R=1.002e+01 
R8590t7108 n8591 n7109 R=4.876e+00 
R8590t6990 n8591 n6991 R=8.926e+00 
R8591t4014 n8592 n4015 R=8.571e+00 
R8591t7967 n8592 n7968 R=2.854e+02 
R8591t6406 n8592 n6407 R=5.254e+00 
R8591t7036 n8592 n7037 R=8.656e+00 
R8591t1693 n8592 n1694 R=9.654e+01 
R8591t1802 n8592 n1803 R=9.071e+00 
R8592t6401 n8593 n6402 R=4.254e+00 
R8592t8399 n8593 n8400 R=1.468e+01 
R8592t7745 n8593 n7746 R=9.120e+00 
R8593t463 n8594 n464 R=4.339e+01 
R8593t2004 n8594 n2005 R=8.745e+00 
R8593t4929 n8594 n4930 R=8.937e+00 
R8593t275 n8594 n276 R=9.273e+00 
R8593t1909 n8594 n1910 R=1.764e+01 
R8593t3793 n8594 n3794 R=6.425e+00 
R8594t502 n8595 n503 R=1.372e+00 
R8594t2398 n8595 n2399 R=1.774e+01 
R8594t1158 n8595 n1159 R=5.769e+00 
R8594t2210 n8595 n2211 R=4.682e+00 
R8594t4181 n8595 n4182 R=1.761e+01 
R8595t3725 n8596 n3726 R=1.373e+01 
R8595t7754 n8596 n7755 R=7.804e+00 
R8595t926 n8596 n927 R=3.701e+00 
R8595t6182 n8596 n6183 R=1.138e+02 
R8595t1790 n8596 n1791 R=7.093e+00 
R8596t1729 n8597 n1730 R=1.277e+01 
R8596t3373 n8597 n3374 R=3.483e+00 
R8596t2210 n8597 n2211 R=6.934e+02 
R8596t4181 n8597 n4182 R=3.293e+01 
R8597t4475 n8598 n4476 R=4.275e+00 
R8597t6577 n8598 n6578 R=5.587e+00 
R8597t3326 n8598 n3327 R=2.247e+01 
R8597t2565 n8598 n2566 R=3.873e+01 
R8597t1468 n8598 n1469 R=2.418e+00 
R8598t3588 n8599 n3589 R=2.513e+01 
R8598t4949 n8599 n4950 R=2.130e+02 
R8598t3864 n8599 n3865 R=3.037e+00 
R8598t687 n8599 n688 R=2.542e+01 
R8598t2942 n8599 n2943 R=7.044e+01 
R8598t7128 n8599 n7129 R=3.765e+01 
R8598t8369 n8599 n8370 R=5.962e+00 
R8598t2367 n8599 n2368 R=1.016e+01 
R8598t7012 n8599 n7013 R=8.608e+00 
R8599t2721 n8600 n2722 R=1.403e+01 
R8599t6425 n8600 n6426 R=1.054e+01 
R8599t2916 n8600 n2917 R=6.279e+00 
R8599t8533 n8600 n8534 R=2.327e+00 
R8599t8253 n8600 n8254 R=4.214e+00 
R8600t1692 n8601 n1693 R=4.731e+00 
R8600t7657 n8601 n7658 R=3.729e+01 
R8600t7964 n8601 n7965 R=3.539e+01 
R8600t4335 n8601 n4336 R=7.878e+00 
R8601t5231 n8602 n5232 R=8.939e+00 
R8601t5283 n8602 n5284 R=4.110e+01 
R8601t1559 n8602 n1560 R=4.509e+00 
R8601t4787 n8602 n4788 R=1.308e+01 
R8601t2996 n8602 n2997 R=2.795e+00 
R8601t5169 n8602 n5170 R=1.040e+02 
R8602t6691 n1 n6692 R=7.720e+00 
R8602t5442 n1 n5443 R=4.081e+00 
R8603t5900 n8604 n5901 R=6.694e+00 
R8603t7292 n8604 n7293 R=6.198e+00 
R8603t7968 n8604 n7969 R=6.612e+00 
R8603t4417 n8604 n4418 R=1.053e+02 
R8603t5782 n8604 n5783 R=4.299e+00 
R8603t5267 n8604 n5268 R=6.266e+01 
R8604t8448 n8605 n8449 R=6.170e+00 
R8604t5995 n8605 n5996 R=1.079e+01 
R8604t6232 n8605 n6233 R=1.067e+01 
R8604t7635 n8605 n7636 R=2.855e+00 
R8605t3316 n8606 n3317 R=8.833e+00 
R8605t7495 n8606 n7496 R=7.017e+00 
R8605t2819 n8606 n2820 R=6.380e+01 
R8605t4121 n8606 n4122 R=7.038e+00 
R8605t1196 n8606 n1197 R=1.269e+01 
R8605t5701 n8606 n5702 R=4.987e+00 
R8605t5482 n8606 n5483 R=6.164e+00 
R8606t3532 n8607 n3533 R=9.225e+01 
R8606t7285 n8607 n7286 R=3.852e+01 
R8606t6513 n8607 n6514 R=1.679e+01 
R8606t4752 n8607 n4753 R=3.872e+00 
R8606t556 n8607 n557 R=5.053e+00 
R8607t7518 n8608 n7519 R=2.238e+00 
R8607t8327 n8608 n8328 R=2.024e+01 
R8607t2591 n8608 n2592 R=4.311e+00 
R8607t4625 n8608 n4626 R=1.095e+01 
R8607t1808 n8608 n1809 R=4.188e+01 
R8608t405 n8609 n406 R=2.665e+00 
R8608t4017 n8609 n4018 R=1.324e+01 
R8608t7792 n8609 n7793 R=3.336e+01 
R8608t7689 n8609 n7690 R=6.384e+00 
R8608t4726 n8609 n4727 R=7.972e+00 
R8609t3115 n8610 n3116 R=7.696e+00 
R8609t6697 n8610 n6698 R=2.940e+01 
R8609t3700 n8610 n3701 R=1.139e+01 
R8609t6615 n8610 n6616 R=7.768e+00 
R8609t1801 n8610 n1802 R=2.554e+00 
R8609t2183 n8610 n2184 R=9.259e+00 
R8610t1167 n8611 n1168 R=4.673e+00 
R8610t5194 n8611 n5195 R=2.366e+00 
R8610t4303 n8611 n4304 R=1.488e+01 
R8610t2467 n8611 n2468 R=5.446e+00 
R8611t289 n8612 n290 R=4.125e+00 
R8611t4787 n8612 n4788 R=1.287e+02 
R8611t3781 n8612 n3782 R=5.396e+00 
R8611t5828 n8612 n5829 R=9.280e+00 
R8611t7193 n8612 n7194 R=6.018e+01 
R8611t3045 n8612 n3046 R=3.268e+01 
R8611t2650 n8612 n2651 R=2.042e+01 
R8612t1670 n8613 n1671 R=4.354e+00 
R8612t6342 n8613 n1 R=4.660e+00 
R8612t3389 n8613 n1 R=1.633e+01 
R8612t2247 n8613 n2248 R=1.208e+01 
R8613t1399 n8614 n1400 R=3.073e+00 
R8613t2531 n8614 n2532 R=3.854e+00 
R8613t1730 n8614 n1731 R=6.960e+00 
R8614t6599 n8615 n6600 R=6.837e+00 
R8614t7947 n8615 n7948 R=1.063e+01 
R8614t7064 n8615 n7065 R=2.710e+00 
R8614t4819 n8615 n4820 R=1.068e+01 
R8615t6731 n8616 n6732 R=2.095e+03 
R8615t6834 n8616 n6835 R=4.418e+01 
R8615t5538 n8616 n5539 R=3.087e+00 
R8615t8551 n8616 n8552 R=1.243e+01 
R8615t950 n8616 n951 R=6.499e+00 
R8615t6297 n8616 n6298 R=2.773e+00 
R8616t2570 n8617 n2571 R=4.178e+00 
R8616t8299 n8617 n8300 R=4.988e+00 
R8616t5295 n8617 n5296 R=2.076e+01 
R8616t3239 n8617 n3240 R=1.961e+01 
R8616t573 n8617 n574 R=7.888e+00 
R8616t4792 n8617 n4793 R=7.479e+00 
R8617t653 n8618 n654 R=3.099e+00 
R8617t867 n8618 n868 R=2.749e+00 
R8618t3199 n8619 n3200 R=9.596e+00 
R8618t6089 n8619 n6090 R=4.036e+01 
R8618t4219 n8619 n4220 R=4.325e+00 
R8618t4655 n8619 n4656 R=9.795e+00 
R8618t4180 n8619 n4181 R=1.515e+01 
R8618t4591 n8619 n4592 R=7.708e+00 
R8619t2726 n8620 n2727 R=1.297e+01 
R8619t7467 n8620 n7468 R=7.491e+00 
R8619t6013 n8620 n6014 R=5.467e+00 
R8619t352 n8620 n353 R=1.921e+02 
R8619t1476 n8620 n1477 R=8.562e+00 
R8619t4791 n8620 n4792 R=4.374e+01 
R8619t852 n8620 n853 R=3.199e+00 
R8620t2826 n8621 n2827 R=1.541e+01 
R8620t5327 n8621 n5328 R=8.259e+00 
R8620t4310 n8621 n4311 R=7.186e+00 
R8620t7548 n8621 n7549 R=1.023e+01 
R8620t5117 n8621 n5118 R=8.505e+00 
R8621t2959 n8622 n2960 R=2.716e+00 
R8621t8562 n8622 n8563 R=7.224e+00 
R8621t8215 n8622 n8216 R=2.228e+00 
R8621t2504 n8622 n2505 R=6.047e+00 
R8622t2952 n8623 n2953 R=2.087e+00 
R8622t4991 n8623 n4992 R=6.933e+00 
R8622t3732 n8623 n3733 R=1.531e+01 
R8622t752 n8623 n753 R=7.491e+00 
R8622t1867 n8623 n1868 R=2.279e+01 
R8623t6930 n8624 n6931 R=8.917e+01 
R8623t8443 n8624 n8444 R=7.445e+00 
R8623t760 n8624 n761 R=4.223e+00 
R8623t4097 n8624 n4098 R=1.370e+01 
R8623t4605 n8624 n4606 R=7.110e+00 
R8623t5829 n8624 n5830 R=5.798e+00 
R8624t2317 n8625 n2318 R=2.470e+02 
R8624t7781 n8625 n7782 R=3.991e+00 
R8624t4695 n8625 n4696 R=6.882e+00 
R8624t3721 n8625 n3722 R=2.300e+00 
R8625t2885 n8626 n2886 R=5.761e+00 
R8625t8398 n8626 n8399 R=5.139e+00 
R8625t2558 n8626 n2559 R=8.573e+00 
R8625t3658 n8626 n3659 R=1.661e+01 
R8626t348 n8627 n349 R=9.914e+00 
R8626t3473 n8627 n3474 R=2.899e+00 
R8626t7160 n8627 n7161 R=1.678e+01 
R8626t3957 n8627 n3958 R=2.996e+02 
R8627t1014 n8628 n1015 R=1.510e+01 
R8627t2064 n8628 n2065 R=6.021e+00 
R8627t3359 n8628 n3360 R=1.761e+01 
R8627t2206 n8628 n2207 R=5.398e+00 
R8627t6544 n8628 n6545 R=1.480e+01 
R8627t6829 n8628 n6830 R=4.432e+00 
R8627t6088 n8628 n6089 R=7.540e+01 
R8628t1283 n8629 n1284 R=9.610e+00 
R8628t3506 n8629 n3507 R=5.141e+00 
R8628t6103 n8629 n6104 R=5.131e+00 
R8628t3085 n8629 n3086 R=1.137e+01 
R8628t8412 n8629 n8413 R=8.108e+00 
R8628t2592 n8629 n2593 R=5.306e+01 
R8629t3315 n8630 n3316 R=1.216e+01 
R8629t6983 n8630 n6984 R=5.736e+00 
R8629t7172 n8630 n7173 R=6.475e+00 
R8629t8520 n8630 n8521 R=1.212e+02 
R8629t3217 n8630 n3218 R=1.068e+01 
R8629t2330 n8630 n2331 R=3.525e+01 
R8630t10 n8631 n11 R=1.335e+01 
R8630t4570 n8631 n4571 R=9.760e+00 
R8630t4465 n8631 n4466 R=6.860e+00 
R8630t5088 n8631 n5089 R=6.883e+00 
R8630t8268 n8631 n8269 R=2.699e+00 
R8630t6991 n8631 n6992 R=1.052e+01 
R8631t2569 n8632 n2570 R=4.069e+00 
R8631t4168 n8632 n4169 R=4.716e+00 
R8631t354 n8632 n355 R=4.229e+01 
R8631t5875 n8632 n5876 R=7.413e+00 
R8631t5700 n8632 n5701 R=6.482e+01 
R8632t4135 n8633 n4136 R=3.532e+00 
R8632t5292 n8633 n5293 R=2.167e+01 
R8632t5633 n8633 n5634 R=2.903e+00 
R8632t5419 n8633 n5420 R=2.611e+02 
R8632t8393 n8633 n8394 R=4.848e+01 
R8632t4747 n8633 n4748 R=2.838e+01 
R8632t6589 n8633 n6590 R=5.262e+00 
R8633t4046 n8634 n4047 R=9.308e+01 
R8633t5822 n8634 n5823 R=1.011e+01 
R8633t6212 n8634 n6213 R=2.290e+00 
R8633t5016 n8634 n5017 R=4.919e+02 
R8633t930 n8634 n931 R=2.831e+00 
R8634t4947 n8635 n4948 R=9.219e+01 
R8634t5256 n8635 n5257 R=3.009e+00 
R8634t6832 n8635 n6833 R=4.806e+00 
R8634t5598 n8635 n5599 R=3.301e+00 
R8635t3904 n8636 n3905 R=4.358e+01 
R8635t4925 n8636 n4926 R=6.258e+00 
R8635t4859 n8636 n4860 R=1.050e+01 
R8635t709 n8636 n710 R=1.995e+01 
R8635t2145 n8636 n2146 R=1.644e+01 
R8636t3629 n8637 n3630 R=1.021e+01 
R8636t5299 n8637 n5300 R=5.008e+00 
R8636t5511 n8637 n5512 R=1.210e+01 
R8637t2137 n8638 n2138 R=1.099e+01 
R8637t6931 n8638 n6932 R=2.068e+01 
R8637t4171 n8638 n4172 R=3.522e+00 
R8638t4606 n8639 n4607 R=6.943e+00 
R8638t850 n8639 n851 R=1.335e+01 
R8638t3960 n8639 n3961 R=4.336e+00 
R8639t1398 n8640 n1399 R=8.764e+01 
R8639t3541 n8640 n3542 R=3.934e+01 
R8639t7170 n8640 n7171 R=7.499e+00 
R8639t4225 n8640 n4226 R=1.594e+02 
R8639t205 n8640 n206 R=6.040e+00 
R8639t5304 n8640 n5305 R=4.969e+00 
R8639t2893 n8640 n2894 R=3.321e+00 
R8640t8175 n8641 n8176 R=1.506e+01 
R8640t6068 n8641 n6069 R=3.184e+00 
R8640t3631 n8641 n3632 R=1.885e+01 
R8640t8326 n8641 n8327 R=3.506e+00 
R8641t4107 n8642 n4108 R=6.127e+00 
R8641t5684 n8642 n5685 R=5.207e+00 
R8641t6121 n8642 n6122 R=1.774e+01 
R8641t3529 n8642 n3530 R=2.591e+01 
R8641t3215 n8642 n3216 R=5.054e+00 
R8641t7565 n8642 n7566 R=1.188e+01 
R8641t2560 n8642 n2561 R=1.368e+01 
R8642t2748 n8643 n2749 R=1.006e+01 
R8642t5988 n8643 n5989 R=5.014e+00 
R8643t665 n8644 n666 R=1.941e+00 
R8643t8020 n8644 n8021 R=7.664e+00 
R8643t6357 n8644 n6358 R=4.500e+00 
R8644t305 n8645 n306 R=9.411e+00 
R8644t6651 n8645 n6652 R=2.041e+01 
R8644t2472 n8645 n2473 R=4.433e+00 
R8644t488 n8645 n489 R=1.764e+01 
R8644t1090 n8645 n1091 R=1.877e+01 
R8644t5469 n8645 n5470 R=1.513e+00 
R8645t4583 n8646 n4584 R=1.892e+01 
R8645t4777 n8646 n4778 R=4.310e+00 
R8645t3109 n8646 n3110 R=6.615e+00 
R8645t5327 n8646 n5328 R=5.148e+00 
R8645t4310 n8646 n4311 R=5.423e+00 
R8646t724 n8647 n725 R=2.631e+01 
R8646t595 n8647 n596 R=3.186e+00 
R8646t57 n8647 n58 R=8.770e+00 
R8646t1694 n8647 n1695 R=4.844e+01 
R8646t1433 n8647 n1434 R=3.262e+01 
R8647t1778 n8648 n1779 R=2.519e+00 
R8647t8297 n8648 n8298 R=3.519e+00 
R8647t3282 n8648 n3283 R=2.095e+01 
R8647t937 n8648 n938 R=1.780e+01 
R8647t8313 n8648 n8314 R=7.148e+00 
R8648t1659 n8649 n1660 R=5.804e+00 
R8648t4604 n8649 n4605 R=1.349e+02 
R8648t8514 n8649 n8515 R=5.753e+01 
R8648t7380 n8649 n7381 R=6.932e+00 
R8648t7714 n8649 n7715 R=1.644e+01 
R8648t3780 n8649 n3781 R=1.073e+01 
R8648t6783 n8649 n6784 R=1.658e+01 
R8648t6693 n8649 n6694 R=6.815e+00 
R8648t4624 n8649 n4625 R=1.027e+01 
R8649t3652 n8650 n3653 R=4.163e+00 
R8649t7115 n8650 n7116 R=4.592e+00 
R8649t5311 n8650 n5312 R=2.076e+01 
R8649t1070 n8650 n1071 R=1.141e+01 
R8649t837 n8650 n838 R=1.288e+01 
R8650t2580 n8651 n2581 R=3.391e+00 
R8650t2815 n8651 n2816 R=1.629e+01 
R8650t698 n8651 n699 R=4.982e+01 
R8650t8292 n8651 n8293 R=2.780e+00 
R8651t5201 n8652 n5202 R=2.682e+00 
R8651t6134 n8652 n6135 R=4.123e+00 
R8651t7563 n8652 n7564 R=6.786e+01 
R8651t4075 n8652 n4076 R=6.334e+00 
R8651t8378 n8652 n8379 R=8.043e+00 
R8652t3133 n8653 n3134 R=2.860e+01 
R8652t1259 n8653 n1260 R=3.178e+00 
R8652t6073 n8653 n6074 R=7.824e+00 
R8653t620 n8654 n621 R=1.337e+01 
R8653t7946 n8654 n7947 R=1.767e+01 
R8653t6098 n8654 n6099 R=5.643e+00 
R8653t2401 n8654 n2402 R=1.691e+01 
R8653t266 n8654 n267 R=4.909e+00 
R8654t1008 n8655 n1009 R=4.276e+00 
R8654t1895 n8655 n1896 R=1.535e+01 
R8654t3165 n8655 n3166 R=1.461e+01 
R8654t6197 n8655 n6198 R=6.662e+00 
R8654t4154 n8655 n4155 R=7.944e+00 
R8654t437 n8655 n438 R=1.883e+01 
R8655t4053 n8656 n4054 R=1.287e+01 
R8655t4649 n8656 n4650 R=3.484e+00 
R8655t4120 n8656 n4121 R=6.629e+01 
R8655t3809 n8656 n3810 R=1.122e+01 
R8655t5403 n8656 n5404 R=3.463e+00 
R8655t8259 n8656 n8260 R=6.771e+00 
R8656t2630 n8657 n2631 R=1.569e+01 
R8656t2742 n8657 n2743 R=3.454e+01 
R8656t1490 n8657 n1491 R=1.197e+02 
R8656t1593 n8657 n1594 R=1.953e+01 
R8656t5895 n8657 n5896 R=1.457e+01 
R8656t1667 n8657 n1668 R=3.230e+01 
R8656t1106 n8657 n1107 R=2.898e+00 
R8656t4278 n8657 n4279 R=2.137e+02 
R8657t7657 n8658 n7658 R=5.604e+00 
R8657t8600 n8658 n8601 R=1.197e+01 
R8657t4335 n8658 n4336 R=4.159e+00 
R8657t8380 n8658 n8381 R=4.381e+01 
R8657t5175 n8658 n5176 R=3.719e+00 
R8657t1524 n8658 n1525 R=1.135e+01 
R8657t5767 n8658 n5768 R=5.363e+01 
R8658t2414 n8659 n2415 R=5.956e+00 
R8658t1936 n8659 n1937 R=4.930e+00 
R8658t2392 n8659 n2393 R=6.600e+00 
R8658t3076 n8659 n3077 R=1.398e+01 
R8658t3859 n8659 n3860 R=2.150e+01 
R8659t2361 n8660 n2362 R=6.719e+00 
R8659t4492 n8660 n4493 R=1.454e+03 
R8659t8397 n8660 n8398 R=1.223e+01 
R8659t3273 n8660 n3274 R=2.096e+00 
R8659t4799 n8660 n4800 R=3.926e+01 
R8660t3305 n8661 n3306 R=1.338e+01 
R8660t3426 n8661 n3427 R=1.974e+00 
R8660t7429 n8661 n7430 R=6.931e+01 
R8660t5794 n8661 n5795 R=2.650e+01 
R8660t7674 n8661 n7675 R=3.991e+00 
R8660t5977 n8661 n5978 R=4.524e+01 
R8660t6549 n8661 n6550 R=7.008e+00 
R8661t4470 n8662 n4471 R=2.331e+01 
R8661t6028 n8662 n6029 R=7.171e+00 
R8661t6780 n8662 n6781 R=1.985e+01 
R8661t5157 n8662 n5158 R=8.266e+00 
R8661t8308 n8662 n8309 R=1.637e+01 
R8661t6482 n8662 n6483 R=8.055e+00 
R8661t3244 n8662 n3245 R=1.105e+01 
R8661t3552 n8662 n3553 R=6.285e+01 
R8662t5321 n8663 n5322 R=4.307e+00 
R8662t7331 n8663 n7332 R=9.839e+00 
R8662t183 n8663 n184 R=5.704e+00 
R8662t2516 n8663 n2517 R=4.235e+01 
R8662t7122 n8663 n7123 R=2.445e+00 
R8662t6980 n8663 n6981 R=1.160e+02 
R8663t2371 n8664 n2372 R=1.872e+01 
R8663t4761 n8664 n4762 R=1.221e+01 
R8663t1671 n8664 n1672 R=3.683e+00 
R8663t7734 n8664 n7735 R=2.986e+01 
R8663t6366 n8664 n6367 R=4.766e+00 
R8663t2011 n8664 n2012 R=9.201e+00 
R8664t83 n8665 n84 R=1.128e+01 
R8664t1451 n8665 n1452 R=1.315e+01 
R8664t1567 n8665 n1568 R=7.263e+00 
R8664t1056 n8665 n1057 R=5.726e+00 
R8664t1218 n8665 n1219 R=6.258e+00 
R8665t8403 n8666 n8404 R=3.024e+00 
R8665t5554 n8666 n5555 R=7.126e+00 
R8665t2228 n8666 n2229 R=1.457e+01 
R8665t3955 n8666 n3956 R=3.458e+00 
R8665t1111 n8666 n1112 R=2.855e+01 
R8666t7155 n8667 n7156 R=1.067e+01 
R8666t520 n8667 n521 R=5.109e+00 
R8666t7148 n8667 n7149 R=6.681e+00 
R8667t424 n8668 n425 R=2.104e+00 
R8667t6331 n8668 n6332 R=3.425e+01 
R8667t5230 n8668 n5231 R=2.992e+00 
R8667t4735 n8668 n4736 R=3.388e+00 
R8668t4682 n8669 n4683 R=3.422e+00 
R8669t2197 n8670 n2198 R=1.695e+02 
R8669t6433 n8670 n6434 R=4.997e+00 
R8669t5644 n8670 n5645 R=1.684e+01 
R8669t2671 n8670 n2672 R=7.260e+00 
R8669t3180 n8670 n3181 R=2.395e+00 
R8669t7169 n8670 n7170 R=1.887e+01 
R8670t3557 n8671 n3558 R=2.827e+01 
R8670t8219 n8671 n8220 R=1.137e+01 
R8670t2430 n8671 n2431 R=5.073e+00 
R8670t5010 n8671 n5011 R=6.492e+01 
R8670t3106 n8671 n3107 R=1.040e+01 
R8670t3009 n8671 n3010 R=3.153e+01 
R8670t3606 n8671 n3607 R=4.722e+00 
R8671t352 n8672 n353 R=1.810e+01 
R8671t6013 n8672 n6014 R=5.687e+00 
R8671t8338 n8672 n8339 R=1.271e+01 
R8671t8018 n8672 n8019 R=2.566e+00 
R8671t4987 n8672 n4988 R=6.199e+00 
R8672t6280 n8673 n6281 R=4.026e+01 
R8672t8348 n8673 n8349 R=1.322e+03 
R8672t5943 n8673 n5944 R=4.024e+01 
R8672t5796 n8673 n5797 R=7.935e+00 
R8672t1487 n8673 n1488 R=8.870e+00 
R8672t6391 n8673 n6392 R=5.962e+00 
R8673t7667 n8674 n7668 R=5.431e+00 
R8673t8110 n8674 n8111 R=1.166e+02 
R8673t711 n8674 n712 R=1.112e+01 
R8673t6489 n8674 n6490 R=2.046e+01 
R8673t350 n8674 n351 R=3.322e+00 
R8673t2000 n8674 n2001 R=6.804e+00 
R8674t3040 n8675 n3041 R=1.166e+01 
R8674t5247 n8675 n5248 R=2.203e+00 
R8674t4538 n8675 n4539 R=6.986e+00 
R8674t2855 n8675 n2856 R=3.610e+01 
R8674t4593 n8675 n4594 R=2.397e+00 
R8675t6878 n8676 n6879 R=8.996e+00 
R8675t7477 n8676 n7478 R=3.557e+00 
R8675t2738 n8676 n2739 R=1.271e+01 
R8675t3356 n8676 n3357 R=3.412e+01 
R8675t106 n8676 n107 R=4.798e+01 
R8675t2292 n8676 n2293 R=3.059e+00 
R8676t7883 n8677 n7884 R=3.965e+01 
R8676t5904 n8677 n5905 R=2.685e+00 
R8676t7010 n8677 n7011 R=9.719e+00 
R8676t3961 n8677 n3962 R=4.394e+00 
R8677t1946 n8678 n1947 R=7.426e+00 
R8677t8366 n8678 n8367 R=3.352e+00 
R8677t2640 n8678 n2641 R=1.541e+01 
R8677t2769 n8678 n2770 R=3.859e+00 
R8677t5949 n8678 n5950 R=8.027e+00 
R8678t3020 n8679 n3021 R=1.757e+01 
R8678t5341 n8679 n5342 R=8.329e+00 
R8678t1113 n8679 n1114 R=5.844e+01 
R8678t5174 n8679 n5175 R=3.837e+00 
R8678t635 n8679 n636 R=6.330e+00 
R8678t2370 n8679 n2371 R=9.272e+00 
R8678t4613 n8679 n4614 R=1.407e+02 
R8678t800 n8679 n801 R=6.928e+00 
R8679t4454 n1 n4455 R=1.200e+01 
R8679t6293 n1 n6294 R=1.682e+01 
R8679t8281 n1 n8282 R=4.234e+01 
R8679t4042 n1 n4043 R=5.437e+00 
R8680t1484 n8681 n1 R=1.015e+01 
R8680t6041 n8681 n1 R=1.443e+02 
R8680t1383 n8681 n1384 R=3.803e+00 
R8680t7844 n8681 n7845 R=4.823e+01 
R8680t6646 n8681 n1 R=2.463e+00 
R8681t2558 n8682 n2559 R=5.430e+00 
R8681t8185 n8682 n8186 R=3.902e+00 
R8681t2885 n8682 n2886 R=5.009e+01 
R8681t8625 n8682 n8626 R=6.725e+00 
R8682t3651 n8683 n3652 R=1.453e+01 
R8682t4351 n8683 n4352 R=1.758e+01 
R8682t4976 n8683 n4977 R=1.034e+01 
R8682t1076 n8683 n1077 R=9.018e+00 
R8682t4079 n8683 n4080 R=1.735e+01 
R8682t2844 n8683 n2845 R=1.920e+01 
R8682t3297 n8683 n3298 R=5.329e+00 
R8683t970 n8684 n971 R=1.074e+01 
R8683t2237 n8684 n2238 R=3.418e+00 
R8683t484 n8684 n485 R=2.489e+01 
R8683t8518 n8684 n8519 R=1.547e+01 
R8683t5535 n8684 n5536 R=5.612e+00 
R8684t2266 n8685 n2267 R=2.300e+00 
R8684t7370 n8685 n7371 R=3.372e+01 
R8684t5790 n8685 n5791 R=8.222e+01 
R8684t5136 n8685 n5137 R=1.253e+01 
R8684t8395 n8685 n8396 R=1.453e+01 
R8684t4274 n8685 n4275 R=2.335e+01 
R8685t3757 n8686 n3758 R=3.035e+00 
R8685t2448 n8686 n2449 R=3.200e+01 
R8685t7044 n8686 n7045 R=1.086e+01 
R8685t77 n8686 n78 R=3.467e+01 
R8685t584 n8686 n585 R=4.610e+00 
R8686t3143 n8687 n3144 R=1.322e+01 
R8686t3330 n8687 n3331 R=3.648e+01 
R8686t1428 n8687 n1429 R=5.389e+00 
R8686t5384 n8687 n5385 R=1.960e+01 
R8686t8088 n8687 n8089 R=1.087e+01 
R8686t4260 n8687 n4261 R=7.531e+00 
R8687t3723 n8688 n3724 R=3.595e+01 
R8687t7528 n8688 n7529 R=4.827e+00 
R8687t2038 n8688 n2039 R=3.025e+00 
R8687t6713 n8688 n6714 R=9.953e+00 
R8687t1408 n8688 n1409 R=4.211e+00 
R8688t6170 n8689 n6171 R=9.208e+01 
R8688t7162 n8689 n7163 R=1.126e+01 
R8688t2410 n8689 n2411 R=4.677e+00 
R8688t4013 n8689 n4014 R=5.273e+00 
R8688t6867 n8689 n6868 R=5.670e+00 
R8688t6931 n8689 n6932 R=9.593e+01 
R8688t6822 n8689 n6823 R=5.939e+02 
R8688t6747 n8689 n6748 R=1.508e+02 
R8689t5018 n8690 n5019 R=3.887e+01 
R8689t7731 n8690 n7732 R=6.815e+00 
R8689t1193 n8690 n1194 R=4.586e+00 
R8689t1120 n8690 n1121 R=2.304e+00 
R8690t6289 n8691 n6290 R=1.713e+01 
R8690t7413 n8691 n7414 R=2.414e+01 
R8690t3266 n8691 n3267 R=2.906e+00 
R8690t1867 n8691 n1868 R=8.103e+00 
R8690t6417 n8691 n6418 R=3.925e+00 
R8691t5468 n8692 n5469 R=2.420e+01 
R8691t7854 n8692 n7855 R=3.522e+00 
R8691t8528 n8692 n8529 R=9.168e+02 
R8691t593 n8692 n594 R=2.276e+00 
R8691t4209 n8692 n4210 R=3.246e+00 
R8692t2040 n8693 n2041 R=9.029e+00 
R8692t2656 n8693 n2657 R=2.191e+01 
R8692t6913 n8693 n6914 R=2.633e+01 
R8692t5666 n8693 n5667 R=8.367e+00 
R8692t6203 n8693 n6204 R=9.690e+00 
R8693t1300 n8694 n1301 R=5.157e+00 
R8693t8322 n8694 n8323 R=8.488e+00 
R8693t6322 n8694 n6323 R=2.409e+01 
R8693t6338 n8694 n6339 R=1.197e+01 
R8693t3865 n8694 n3866 R=3.041e+00 
R8693t6238 n8694 n6239 R=9.386e+00 
R8693t1330 n8694 n1331 R=1.872e+02 
R8694t3724 n8695 n3725 R=4.101e+00 
R8694t5286 n8695 n5287 R=4.966e+00 
R8694t801 n8695 n802 R=1.190e+01 
R8694t2253 n8695 n2254 R=8.978e+00 
R8695t2633 n8696 n2634 R=1.726e+01 
R8695t8166 n8696 n8167 R=6.150e+00 
R8695t4047 n8696 n4048 R=4.280e+00 
R8695t5498 n8696 n5499 R=8.065e+00 
R8695t4128 n8696 n4129 R=5.031e+00 
R8695t1513 n8696 n1514 R=1.092e+01 
R8696t1989 n8697 n1990 R=1.043e+01 
R8696t6224 n8697 n6225 R=2.849e+00 
R8696t2432 n8697 n2433 R=1.615e+01 
R8696t2194 n8697 n2195 R=3.506e+00 
R8696t3840 n8697 n3841 R=2.637e+01 
R8697t5309 n8698 n5310 R=4.670e+00 
R8697t4244 n8698 n4245 R=1.962e+01 
R8697t3390 n8698 n3391 R=5.017e+01 
R8697t5293 n8698 n5294 R=4.138e+00 
R8697t6884 n8698 n6885 R=1.364e+01 
R8698t982 n8699 n983 R=7.183e+00 
R8698t3364 n8699 n3365 R=9.197e+00 
R8698t7144 n8699 n7145 R=6.505e+00 
R8698t7527 n8699 n7528 R=3.386e+00 
R8698t3953 n8699 n3954 R=3.897e+01 
R8698t7435 n8699 n7436 R=5.806e+00 
R8699t8277 n8700 n8278 R=4.092e+00 
R8699t482 n8700 n483 R=6.549e+00 
R8699t1326 n8700 n1327 R=3.773e+00 
R8699t993 n8700 n994 R=4.068e+01 
R8699t3711 n8700 n3712 R=1.694e+01 
R8699t2413 n8700 n2414 R=1.617e+02 
R8700t1193 n8701 n1194 R=4.642e+00 
R8700t8689 n8701 n8690 R=8.423e+00 
R8700t8182 n8701 n8183 R=1.466e+01 
R8700t5657 n8701 n5658 R=1.664e+01 
R8700t3114 n8701 n3115 R=2.983e+01 
R8700t5107 n8701 n5108 R=4.773e+00 
R8700t6829 n8701 n6830 R=5.352e+01 
R8700t8379 n8701 n8380 R=3.806e+01 
R8700t1120 n8701 n1121 R=5.359e+01 
R8701t4119 n8702 n4120 R=2.506e+01 
R8701t6045 n8702 n6046 R=3.929e+01 
R8701t5247 n8702 n5248 R=1.504e+00 
R8701t4538 n8702 n4539 R=3.098e+01 
R8701t1532 n8702 n1533 R=2.024e+00 
R8701t2420 n8702 n2421 R=4.440e+01 
R8702t1792 n8703 n1793 R=1.188e+01 
R8702t5931 n8703 n5932 R=1.030e+01 
R8702t1444 n8703 n1445 R=1.546e+01 
R8702t2454 n8703 n2455 R=5.126e+01 
R8702t4217 n8703 n4218 R=3.961e+00 
R8703t413 n8704 n414 R=2.831e+00 
R8703t3691 n8704 n3692 R=1.167e+01 
R8703t1573 n8704 n1574 R=1.664e+01 
R8703t190 n8704 n191 R=1.055e+01 
R8703t5769 n8704 n5770 R=1.721e+01 
R8704t7539 n8705 n7540 R=4.346e+00 
R8704t1262 n8705 n1263 R=6.656e+01 
R8704t6782 n8705 n6783 R=2.424e+00 
R8705t2159 n8706 n2160 R=1.111e+01 
R8705t3929 n8706 n3930 R=3.043e+00 
R8705t2733 n8706 n2734 R=2.251e+00 
R8705t5165 n8706 n5166 R=6.643e+00 
R8705t451 n8706 n452 R=3.194e+01 
R8706t3132 n8707 n3133 R=3.294e+00 
R8706t5833 n8707 n5834 R=1.763e+01 
R8706t38 n8707 n39 R=6.444e+00 
R8707t2260 n8708 n2261 R=1.841e+01 
R8707t4535 n8708 n4536 R=1.300e+01 
R8707t739 n8708 n740 R=1.195e+01 
R8707t5654 n8708 n5655 R=9.638e+00 
R8707t1474 n8708 n1475 R=2.966e+01 
R8707t8441 n8708 n8442 R=3.290e+00 
R8708t3548 n8709 n3549 R=4.713e+00 
R8708t7889 n8709 n7890 R=4.381e+00 
R8708t6571 n8709 n6572 R=7.505e+01 
R8708t8205 n8709 n8206 R=2.470e+01 
R8708t24 n8709 n25 R=8.588e+01 
R8708t8540 n8709 n8541 R=2.934e+00 
R8708t4190 n8709 n4191 R=2.238e+01 
R8709t2099 n8710 n2100 R=7.265e+00 
R8709t5821 n8710 n5822 R=4.014e+00 
R8709t6485 n8710 n6486 R=6.557e+00 
R8709t5111 n8710 n5112 R=2.691e+00 
R8710t885 n8711 n886 R=1.458e+01 
R8710t4280 n8711 n4281 R=1.473e+01 
R8710t1923 n8711 n1924 R=4.173e+00 
R8710t2012 n8711 n2013 R=2.519e+00 
R8711t744 n8712 n745 R=3.145e+00 
R8711t2194 n8712 n2195 R=3.930e+01 
R8711t5058 n8712 n5059 R=3.314e+01 
R8711t6525 n8712 n6526 R=5.672e+00 
R8711t8220 n8712 n8221 R=9.361e+00 
R8711t6000 n8712 n6001 R=9.073e+00 
R8711t2928 n8712 n2929 R=6.792e+00 
R8712t2382 n8713 n2383 R=5.151e+01 
R8712t8296 n8713 n8297 R=2.685e+00 
R8712t7981 n8713 n7982 R=5.876e+00 
R8712t2794 n8713 n2795 R=5.559e+00 
R8713t722 n8714 n723 R=1.364e+01 
R8713t5532 n8714 n5533 R=5.813e+01 
R8713t8516 n8714 n8517 R=8.271e+00 
R8713t6604 n8714 n6605 R=2.509e+00 
R8713t4177 n8714 n4178 R=7.716e+01 
R8713t2305 n8714 n2306 R=1.173e+01 
R8713t8167 n8714 n8168 R=6.287e+00 
R8714t2135 n8715 n2136 R=1.055e+01 
R8714t7432 n8715 n7433 R=1.318e+01 
R8714t8210 n8715 n8211 R=1.295e+01 
R8714t2910 n8715 n2911 R=5.338e+00 
R8714t8094 n8715 n8095 R=1.701e+01 
R8714t1009 n8715 n1010 R=2.659e+00 
R8715t4932 n8716 n4933 R=9.696e+00 
R8715t6084 n8716 n6085 R=6.730e+00 
R8715t5029 n8716 n5030 R=6.804e+00 
R8715t4218 n8716 n4219 R=8.966e+00 
R8715t5572 n8716 n5573 R=4.247e+00 
R8716t58 n8717 n59 R=1.102e+01 
R8716t6669 n8717 n6670 R=1.784e+02 
R8716t5497 n8717 n5498 R=2.625e+00 
R8716t456 n8717 n457 R=7.925e+00 
R8716t1970 n8717 n1971 R=3.447e+00 
R8717t2799 n8718 n2800 R=6.972e+01 
R8717t7246 n8718 n7247 R=5.168e+00 
R8717t7323 n8718 n7324 R=6.451e+02 
R8717t3485 n8718 n3486 R=1.011e+01 
R8717t8380 n8718 n8381 R=1.424e+01 
R8717t7678 n8718 n7679 R=7.640e+00 
R8717t4782 n8718 n4783 R=6.209e+00 
R8717t1651 n8718 n1652 R=1.820e+01 
R8718t867 n8719 n868 R=4.579e+00 
R8718t54 n8719 n55 R=5.110e+01 
R8718t8433 n8719 n8434 R=4.630e+00 
R8718t4442 n8719 n4443 R=4.323e+00 
R8718t7161 n8719 n7162 R=1.127e+01 
R8718t653 n8719 n654 R=3.913e+01 
R8718t8617 n8719 n8618 R=7.683e+00 
R8719t6420 n8720 n6421 R=1.772e+01 
R8719t2899 n8720 n2900 R=4.558e+00 
R8719t5832 n8720 n5833 R=3.711e+01 
R8719t8061 n8720 n8062 R=1.904e+01 
R8719t8424 n8720 n8425 R=2.690e+00 
R8720t4411 n8721 n4412 R=9.039e+00 
R8720t7899 n8721 n7900 R=1.477e+01 
R8720t7381 n8721 n7382 R=6.893e+01 
R8720t6557 n8721 n6558 R=2.440e+00 
R8721t5879 n8722 n5880 R=8.072e+01 
R8721t6814 n8722 n6815 R=4.786e+00 
R8721t7403 n8722 n7404 R=1.269e+01 
R8721t2228 n8722 n2229 R=4.030e+00 
R8721t3955 n8722 n3956 R=5.121e+00 
R8721t7510 n8722 n7511 R=9.797e+00 
R8722t1892 n8723 n1893 R=8.713e+00 
R8722t2525 n8723 n2526 R=3.446e+00 
R8722t83 n8723 n84 R=4.889e+01 
R8722t8664 n8723 n8665 R=1.040e+01 
R8722t1218 n8723 n1219 R=7.687e+00 
R8723t992 n8724 n993 R=5.416e+00 
R8723t1018 n8724 n1019 R=5.405e+02 
R8723t5556 n8724 n5557 R=7.590e+00 
R8723t6970 n8724 n6971 R=1.109e+01 
R8723t3178 n8724 n3179 R=5.151e+00 
R8723t754 n8724 n755 R=1.754e+01 
R8723t5896 n8724 n5897 R=9.314e+01 
R8723t1035 n8724 n1036 R=9.786e+00 
R8723t1370 n8724 n1371 R=2.172e+01 
R8723t5970 n8724 n5971 R=1.216e+02 
R8724t2369 n8725 n2370 R=5.385e+01 
R8724t6108 n8725 n6109 R=6.949e+01 
R8724t112 n8725 n113 R=2.032e+02 
R8724t5856 n8725 n5857 R=1.222e+01 
R8724t6653 n8725 n6654 R=5.696e+00 
R8724t2028 n8725 n2029 R=3.098e+02 
R8724t3666 n8725 n3667 R=2.785e+00 
R8725t4924 n8726 n4925 R=5.997e+00 
R8725t3510 n8726 n3511 R=2.648e+01 
R8725t591 n8726 n592 R=6.285e+00 
R8725t1867 n8726 n1868 R=3.286e+02 
R8725t6417 n8726 n6418 R=3.984e+00 
R8726t4255 n8727 n4256 R=3.416e+00 
R8726t6369 n8727 n6370 R=4.420e+02 
R8726t427 n8727 n428 R=1.846e+01 
R8726t7720 n8727 n7721 R=3.515e+00 
R8726t3067 n8727 n3068 R=1.436e+01 
R8726t6777 n8727 n6778 R=3.455e+02 
R8726t1793 n8727 n1794 R=1.541e+01 
R8727t2743 n8728 n2744 R=1.581e+01 
R8727t7852 n8728 n7853 R=1.274e+01 
R8727t9 n8728 n10 R=8.166e+00 
R8727t7299 n8728 n7300 R=2.966e+01 
R8727t7488 n8728 n7489 R=2.449e+00 
R8728t175 n8729 n176 R=8.601e+00 
R8728t4606 n8729 n4607 R=7.788e+00 
R8728t751 n8729 n752 R=1.811e+01 
R8729t3585 n8730 n3586 R=7.945e+01 
R8729t8588 n8730 n8589 R=4.038e+00 
R8729t7088 n8730 n7089 R=8.922e+00 
R8729t3459 n8730 n3460 R=1.501e+01 
R8729t5999 n8730 n6000 R=1.432e+01 
R8729t1541 n8730 n1542 R=2.200e+01 
R8730t1788 n8731 n1789 R=2.419e+00 
R8730t7753 n8731 n7754 R=1.838e+00 
R8730t3311 n8731 n3312 R=1.212e+01 
R8730t6584 n8731 n6585 R=8.394e+00 
R8730t6340 n8731 n6341 R=6.694e+01 
R8731t2322 n8732 n2323 R=6.771e+00 
R8731t5263 n8732 n5264 R=1.409e+01 
R8731t822 n8732 n823 R=1.638e+01 
R8731t6574 n8732 n6575 R=4.697e+00 
R8731t3204 n8732 n3205 R=2.557e+01 
R8731t227 n8732 n228 R=3.114e+00 
R8732t3379 n8733 n3380 R=1.899e+01 
R8732t5394 n8733 n5395 R=5.722e+00 
R8732t8164 n8733 n8165 R=5.817e+00 
R8733t4934 n8734 n4935 R=8.165e+02 
R8733t6513 n8734 n6514 R=1.420e+01 
R8733t1966 n8734 n1967 R=6.072e+00 
R8733t5711 n8734 n5712 R=8.544e+00 
R8734t2776 n8735 n2777 R=4.127e+00 
R8734t3680 n8735 n3681 R=3.268e+01 
R8735t4234 n8736 n4235 R=3.241e+00 
R8735t7693 n8736 n7694 R=4.459e+00 
R8735t2661 n8736 n2662 R=6.700e+01 
R8735t5817 n8736 n5818 R=1.079e+01 
R8736t3632 n8737 n3633 R=2.013e+00 
R8736t4768 n8737 n4769 R=9.526e+00 
R8736t3022 n8737 n3023 R=2.650e+00 
R8737t7077 n8738 n7078 R=4.302e+00 
R8737t6886 n8738 n6887 R=8.562e+00 
R8737t2533 n8738 n2534 R=1.434e+02 
R8737t81 n8738 n82 R=3.912e+00 
R8737t5285 n8738 n5286 R=8.208e+00 
R8738t809 n8739 n810 R=1.679e+02 
R8738t1837 n8739 n1838 R=5.507e+00 
R8738t4147 n8739 n4148 R=7.675e+00 
R8738t3949 n8739 n3950 R=5.827e+00 
R8739t968 n8740 n969 R=9.201e+00 
R8739t7901 n8740 n7902 R=7.982e+00 
R8739t2865 n8740 n2866 R=5.524e+00 
R8739t6831 n8740 n6832 R=1.489e+01 
R8739t632 n8740 n633 R=5.898e+00 
R8740t32 n8741 n33 R=2.159e+00 
R8740t2163 n8741 n2164 R=6.313e+00 
R8740t3868 n8741 n3869 R=1.939e+02 
R8740t3093 n8741 n3094 R=2.021e+00 
R8741t4759 n8742 n4760 R=2.547e+00 
R8741t5352 n8742 n5353 R=1.591e+01 
R8741t3927 n8742 n3928 R=7.940e+00 
R8741t895 n8742 n896 R=3.910e+01 
R8741t4628 n8742 n4629 R=9.402e+01 
R8741t8409 n8742 n8410 R=2.160e+00 
R8741t7257 n8742 n7258 R=3.268e+01 
R8741t1763 n8742 n1764 R=3.105e+01 
R8741t2792 n8742 n2793 R=7.206e+01 
R8742t5112 n8743 n5113 R=5.211e+00 
R8742t7967 n8743 n7968 R=3.557e+00 
R8743t1406 n8744 n1407 R=5.794e+00 
R8743t3391 n8744 n3392 R=1.436e+01 
R8743t8368 n8744 n8369 R=5.261e+00 
R8743t5773 n8744 n5774 R=1.351e+01 
R8743t6042 n8744 n6043 R=7.910e+00 
R8743t7339 n8744 n7340 R=6.685e+00 
R8744t3083 n8745 n3084 R=3.630e+01 
R8744t5830 n8745 n5831 R=3.652e+00 
R8744t7236 n8745 n7237 R=1.769e+01 
R8744t6891 n8745 n6892 R=5.159e+00 
R8744t1242 n8745 n1243 R=1.037e+01 
R8744t2808 n8745 n2809 R=4.457e+00 
R8745t2776 n8746 n2777 R=4.270e+01 
R8745t8734 n8746 n8735 R=1.004e+01 
R8745t7871 n8746 n7872 R=2.835e+00 
R8745t4026 n8746 n4027 R=3.874e+00 
R8746t997 n8747 n998 R=3.443e+01 
R8746t7908 n8747 n7909 R=3.196e+00 
R8746t7827 n8747 n7828 R=9.506e+00 
R8746t2839 n8747 n2840 R=3.875e+00 
R8746t8294 n8747 n8295 R=3.683e+02 
R8746t8238 n8747 n8239 R=5.699e+00 
R8746t5036 n8747 n5037 R=9.290e+02 
R8747t3754 n8748 n3755 R=3.524e+00 
R8747t8279 n8748 n8280 R=4.041e+01 
R8747t2711 n8748 n2712 R=5.034e+00 
R8747t5456 n8748 n5457 R=1.595e+01 
R8747t3172 n8748 n3173 R=5.841e+00 
R8748t2953 n8749 n2954 R=2.581e+01 
R8748t7631 n8749 n7632 R=5.246e+00 
R8748t2245 n8749 n2246 R=2.849e+01 
R8748t6156 n8749 n6157 R=1.385e+01 
R8748t239 n8749 n240 R=5.549e+00 
R8748t3748 n8749 n3749 R=1.136e+01 
R8749t650 n8750 n651 R=4.168e+00 
R8749t6172 n8750 n6173 R=1.114e+01 
R8749t1705 n8750 n1706 R=9.122e+00 
R8749t4476 n8750 n4477 R=5.537e+01 
R8749t3839 n8750 n3840 R=5.360e+00 
R8750t2955 n8751 n2956 R=3.600e+01 
R8750t6467 n8751 n6468 R=5.577e+01 
R8750t7483 n8751 n7484 R=6.401e+00 
R8750t4076 n8751 n4077 R=2.475e+00 
R8750t6441 n8751 n6442 R=2.587e+01 
R8750t4497 n8751 n4498 R=4.533e+00 
R8750t3109 n8751 n3110 R=3.028e+01 
R8751t3810 n8752 n3811 R=1.641e+01 
R8751t7992 n8752 n7993 R=1.377e+01 
R8751t1548 n8752 n1549 R=2.053e+01 
R8751t3894 n8752 n3895 R=3.172e+00 
R8751t1211 n8752 n1212 R=1.173e+01 
R8751t7980 n8752 n7981 R=3.185e+01 
R8751t8169 n8752 n8170 R=6.206e+02 
R8752t6018 n8753 n6019 R=1.515e+01 
R8752t8239 n8753 n8240 R=3.367e+00 
R8752t1284 n8753 n1285 R=4.019e+00 
R8752t2428 n8753 n2429 R=1.236e+01 
R8752t3338 n8753 n3339 R=1.108e+01 
R8753t273 n8754 n274 R=4.268e+00 
R8753t8053 n8754 n8054 R=9.118e+00 
R8753t7844 n8754 n7845 R=1.257e+01 
R8753t4880 n8754 n4881 R=1.403e+01 
R8753t1655 n8754 n1656 R=5.243e+01 
R8754t386 n8755 n387 R=1.047e+01 
R8754t3124 n8755 n3125 R=8.841e+00 
R8754t2724 n8755 n2725 R=7.516e+00 
R8754t4142 n8755 n4143 R=1.540e+01 
R8754t5698 n8755 n5699 R=3.320e+00 
R8755t5597 n8756 n5598 R=3.770e+00 
R8755t5687 n8756 n5688 R=3.376e+00 
R8755t7996 n8756 n7997 R=2.480e+01 
R8755t8316 n8756 n8317 R=4.130e+01 
R8755t5891 n8756 n5892 R=3.594e+00 
R8755t8577 n8756 n8578 R=6.017e+02 
R8756t6401 n8757 n6402 R=1.749e+01 
R8756t8592 n8757 n8593 R=3.847e+00 
R8756t3399 n8757 n3400 R=6.620e+00 
R8756t3179 n8757 n3180 R=2.132e+01 
R8756t6575 n8757 n6576 R=2.302e+00 
R8756t7745 n8757 n7746 R=2.197e+01 
R8757t431 n8758 n432 R=3.572e+00 
R8757t8247 n8758 n8248 R=1.931e+01 
R8757t2716 n8758 n2717 R=2.032e+01 
R8757t1250 n8758 n1251 R=5.414e+01 
R8757t1515 n8758 n1516 R=3.151e+00 
R8757t6010 n8758 n6011 R=9.480e+00 
R8757t3554 n8758 n3555 R=1.721e+01 
R8757t3015 n8758 n3016 R=7.808e+01 
R8758t272 n8759 n273 R=1.685e+01 
R8758t5804 n8759 n5805 R=3.623e+00 
R8758t3116 n8759 n3117 R=7.259e+00 
R8758t4824 n8759 n4825 R=1.985e+02 
R8758t1950 n8759 n1951 R=3.828e+00 
R8758t7559 n8759 n7560 R=1.096e+01 
R8759t4629 n8760 n4630 R=9.874e+00 
R8759t7530 n8760 n7531 R=5.523e+01 
R8759t6006 n8760 n6007 R=3.625e+00 
R8759t719 n8760 n720 R=3.458e+00 
R8759t2576 n8760 n2577 R=1.776e+02 
R8759t2333 n8760 n2334 R=6.604e+00 
R8760t617 n8761 n618 R=6.562e+00 
R8760t5623 n8761 n5624 R=6.943e+00 
R8760t7973 n8761 n7974 R=8.111e+00 
R8760t6400 n8761 n6401 R=4.845e+00 
R8761t8214 n8762 n8215 R=4.295e+00 
R8761t8397 n8762 n8398 R=3.743e+00 
R8761t6017 n8762 n6018 R=1.062e+01 
R8761t2242 n8762 n2243 R=7.771e+01 
R8762t577 n8763 n578 R=9.262e+00 
R8762t3041 n8763 n3042 R=3.349e+00 
R8762t991 n8763 n992 R=7.185e+01 
R8762t4573 n8763 n4574 R=3.285e+00 
R8762t3433 n8763 n3434 R=3.377e+03 
R8763t908 n8764 n909 R=1.467e+02 
R8763t3616 n8764 n3617 R=4.674e+00 
R8763t7842 n8764 n7843 R=7.638e+00 
R8763t6195 n8764 n6196 R=1.617e+01 
R8763t2930 n8764 n2931 R=2.926e+00 
R8764t1007 n8765 n1008 R=4.639e+00 
R8764t3619 n8765 n3620 R=2.638e+00 
R8764t5013 n8765 n5014 R=3.006e+01 
R8764t1449 n8765 n1450 R=5.350e+00 
R8764t3807 n8765 n3808 R=1.000e+02 
R8764t3813 n8765 n3814 R=3.105e+01 
R8765t2315 n8766 n2316 R=7.804e+00 
R8765t3720 n8766 n3721 R=7.582e+00 
R8765t6570 n8766 n6571 R=6.214e+01 
R8765t5611 n8766 n5612 R=6.380e+00 
R8765t7483 n8766 n7484 R=6.844e+00 
R8765t5187 n8766 n5188 R=6.139e+00 
R8766t7327 n8767 n7328 R=2.811e+00 
R8766t2968 n8767 n2969 R=1.034e+01 
R8766t4565 n8767 n4566 R=2.485e+00 
R8767t816 n8768 n817 R=9.892e+01 
R8767t4055 n8768 n4056 R=3.376e+00 
R8767t607 n8768 n608 R=8.495e+00 
R8767t3084 n8768 n3085 R=1.965e+02 
R8767t4671 n8768 n4672 R=3.772e+00 
R8767t8143 n8768 n8144 R=8.909e+00 
R8767t8341 n8768 n8342 R=7.689e+01 
R8767t659 n8768 n660 R=8.168e+01 
R8768t4316 n8769 n4317 R=4.403e+00 
R8768t4933 n8769 n4934 R=1.675e+02 
R8768t7896 n8769 n7897 R=9.478e+00 
R8768t7687 n8769 n7688 R=5.894e+00 
R8768t4242 n8769 n4243 R=2.570e+00 
R8769t141 n8770 n142 R=7.127e+00 
R8769t7690 n8770 n7691 R=3.379e+00 
R8769t4394 n8770 n4395 R=1.578e+01 
R8770t3402 n8771 n3403 R=2.425e+00 
R8770t6019 n8771 n6020 R=3.985e+00 
R8770t6107 n8771 n6108 R=3.087e+00 
R8771t7941 n8772 n7942 R=8.314e+00 
R8771t5376 n8772 n5377 R=7.687e+00 
R8771t8347 n8772 n8348 R=5.216e+00 
R8771t1333 n8772 n1334 R=5.581e+00 
R8771t7123 n8772 n7124 R=1.209e+02 
R8771t8328 n8772 n8329 R=6.807e+01 
R8772t5002 n8773 n5003 R=4.154e+00 
R8772t5831 n8773 n5832 R=1.295e+01 
R8772t2555 n8773 n2556 R=7.837e+01 
R8772t8151 n8773 n8152 R=2.577e+01 
R8772t4473 n8773 n4474 R=2.195e+01 
R8772t133 n8773 n134 R=1.116e+01 
R8772t445 n8773 n446 R=3.945e+00 
R8772t7767 n8773 n7768 R=1.647e+01 
R8772t5717 n8773 n5718 R=2.618e+01 
R8772t1858 n8773 n1859 R=3.074e+03 
R8773t1090 n8774 n1091 R=3.788e+01 
R8773t488 n8774 n489 R=6.284e+00 
R8773t6898 n8774 n6899 R=8.291e+00 
R8774t8017 n8775 n8018 R=2.661e+01 
R8774t8511 n8775 n8512 R=3.541e+00 
R8774t1412 n8775 n1413 R=4.183e+00 
R8774t6142 n8775 n6143 R=1.145e+01 
R8774t7110 n8775 n7111 R=4.315e+00 
R8775t5460 n8776 n5461 R=7.789e+00 
R8775t4679 n8776 n4680 R=9.125e+00 
R8775t6218 n8776 n6219 R=3.362e+00 
R8776t6577 n8777 n6578 R=1.005e+02 
R8776t8496 n8777 n8497 R=7.308e+00 
R8776t5449 n8777 n5450 R=6.617e+00 
R8776t1116 n8777 n1117 R=6.615e+00 
R8776t1468 n8777 n1469 R=2.603e+00 
R8777t439 n8778 n440 R=7.071e+00 
R8777t1635 n8778 n1636 R=2.049e+01 
R8777t8339 n8778 n8340 R=1.926e+01 
R8777t2661 n8778 n2662 R=2.972e+00 
R8777t4234 n8778 n4235 R=1.452e+02 
R8777t1617 n8778 n1618 R=4.110e+00 
R8778t728 n8779 n729 R=1.319e+01 
R8778t1563 n8779 n1564 R=5.344e+00 
R8778t7298 n8779 n7299 R=1.318e+01 
R8778t7975 n8779 n7976 R=2.103e+01 
R8778t2152 n8779 n2153 R=4.601e+00 
R8778t1493 n8779 n1494 R=6.669e+00 
R8779t115 n8780 n116 R=3.777e+01 
R8779t5338 n8780 n5339 R=2.948e+00 
R8779t11 n8780 n12 R=4.264e+00 
R8779t4420 n8780 n4421 R=1.768e+01 
R8779t1819 n8780 n1820 R=3.185e+00 
R8779t2755 n8780 n2756 R=6.692e+01 
R8780t449 n8781 n450 R=2.554e+01 
R8780t2436 n8781 n2437 R=4.175e+00 
R8780t2285 n8781 n2286 R=1.208e+01 
R8780t3816 n8781 n3817 R=9.727e+00 
R8780t2482 n8781 n2483 R=6.146e+00 
R8780t2715 n8781 n2716 R=9.439e+00 
R8781t7327 n8782 n7328 R=1.533e+01 
R8781t8766 n8782 n8767 R=7.870e+00 
R8781t4565 n8782 n4566 R=8.628e+01 
R8781t2393 n8782 n2394 R=9.054e+00 
R8781t532 n8782 n533 R=6.135e+00 
R8782t3453 n8783 n3454 R=8.654e+00 
R8782t3739 n8783 n3740 R=1.066e+01 
R8782t4001 n8783 n4002 R=1.153e+01 
R8782t726 n8783 n727 R=1.059e+02 
R8782t2990 n8783 n2991 R=5.470e+00 
R8782t7734 n8783 n7735 R=1.755e+01 
R8782t1671 n8783 n1672 R=5.164e+00 
R8783t3374 n8784 n3375 R=7.738e+00 
R8783t8087 n8784 n8088 R=4.107e+01 
R8783t5534 n8784 n5535 R=5.080e+00 
R8783t5680 n8784 n5681 R=1.839e+01 
R8783t6546 n8784 n6547 R=5.578e+00 
R8783t3276 n8784 n3277 R=5.656e+00 
R8784t4794 n8785 n4795 R=3.269e+01 
R8784t4946 n8785 n4947 R=2.120e+01 
R8784t4600 n8785 n4601 R=5.058e+00 
R8784t7912 n8785 n7913 R=5.713e+00 
R8784t6307 n8785 n6308 R=3.941e+00 
R8784t5092 n8785 n5093 R=1.009e+01 
R8785t734 n8786 n735 R=3.045e+00 
R8785t5770 n8786 n5771 R=5.221e+01 
R8785t5833 n8786 n5834 R=4.465e+02 
R8785t7306 n8786 n7307 R=3.015e+00 
R8785t6182 n8786 n6183 R=6.917e+00 
R8786t8000 n8787 n8001 R=2.045e+00 
R8786t8003 n8787 n8004 R=1.875e+01 
R8786t1151 n8787 n1152 R=2.620e+00 
R8786t6040 n8787 n6041 R=2.918e+04 
R8786t1928 n8787 n1929 R=2.041e+02 
R8786t927 n8787 n928 R=6.694e+01 
R8787t2200 n8788 n2201 R=1.815e+01 
R8787t2347 n8788 n2348 R=7.628e+00 
R8787t7091 n8788 n7092 R=4.643e+00 
R8787t3163 n8788 n3164 R=4.996e+00 
R8787t6324 n8788 n6325 R=1.368e+01 
R8787t6078 n8788 n6079 R=6.917e+00 
R8788t3000 n8789 n3001 R=4.646e+00 
R8788t5841 n8789 n5842 R=2.483e+00 
R8788t831 n8789 n832 R=4.187e+00 
R8789t73 n8790 n74 R=3.650e+00 
R8789t5814 n8790 n5815 R=1.065e+01 
R8789t1475 n8790 n1476 R=4.605e+00 
R8789t3481 n8790 n3482 R=1.191e+02 
R8789t6053 n8790 n6054 R=1.452e+01 
R8790t5736 n8791 n5737 R=1.882e+01 
R8790t7653 n8791 n7654 R=5.630e+00 
R8790t4952 n8791 n4953 R=6.823e+00 
R8790t7690 n8791 n7691 R=9.260e+00 
R8790t8769 n8791 n8770 R=1.500e+01 
R8790t4394 n8791 n4395 R=7.213e+00 
R8791t6090 n8792 n6091 R=1.056e+01 
R8791t4385 n8792 n1 R=1.528e+01 
R8791t5396 n8792 n5397 R=1.106e+01 
R8791t6345 n8792 n6346 R=1.985e+00 
R8792t1678 n8793 n1679 R=8.963e+00 
R8792t8278 n8793 n8279 R=1.489e+01 
R8792t3979 n8793 n3980 R=2.856e+00 
R8792t3235 n8793 n3236 R=9.662e+00 
R8792t3814 n8793 n3815 R=1.634e+01 
R8793t1972 n8794 n1973 R=2.554e+01 
R8793t5725 n8794 n5726 R=2.655e+00 
R8793t5181 n8794 n5182 R=9.751e+00 
R8794t854 n8795 n855 R=1.634e+01 
R8794t4179 n8795 n4180 R=7.223e+00 
R8794t8562 n8795 n8563 R=2.684e+00 
R8794t8202 n8795 n8203 R=3.733e+02 
R8794t8120 n8795 n8121 R=3.659e+00 
R8794t2543 n8795 n2544 R=1.492e+01 
R8795t6680 n8796 n6681 R=3.537e+00 
R8795t7742 n8796 n7743 R=3.852e+00 
R8795t3639 n8796 n3640 R=7.560e+00 
R8795t6906 n8796 n6907 R=2.211e+02 
R8795t5262 n8796 n5263 R=8.168e+00 
R8796t1470 n8797 n1471 R=1.231e+01 
R8796t3049 n8797 n3050 R=6.284e+00 
R8796t5551 n8797 n5552 R=6.732e+00 
R8796t8582 n8797 n8583 R=3.236e+00 
R8796t3371 n8797 n3372 R=9.112e+00 
R8797t4208 n8798 n4209 R=3.607e+00 
R8797t7020 n8798 n7021 R=4.558e+00 
R8797t5937 n8798 n5938 R=5.149e+01 
R8797t3469 n8798 n3470 R=1.943e+01 
R8797t7478 n8798 n7479 R=4.284e+00 
R8797t4043 n8798 n4044 R=2.048e+01 
R8798t4263 n8799 n4264 R=5.260e+00 
R8798t164 n8799 n165 R=4.431e+00 
R8798t2359 n8799 n2360 R=2.801e+01 
R8799t1957 n8800 n1958 R=1.686e+01 
R8799t4048 n8800 n4049 R=5.480e+00 
R8799t3059 n8800 n3060 R=5.842e+00 
R8799t6502 n8800 n6503 R=1.398e+01 
R8799t4809 n8800 n4810 R=4.250e+00 
R8799t4978 n8800 n4979 R=1.549e+01 
R8799t2785 n8800 n2786 R=2.973e+01 
R8800t3973 n8801 n3974 R=1.021e+01 
R8800t4557 n8801 n4558 R=1.166e+02 
R8800t4096 n8801 n4097 R=7.317e+00 
R8800t2191 n8801 n2192 R=8.226e+00 
R8800t6092 n8801 n6093 R=5.650e+00 
R8800t8342 n8801 n8343 R=4.644e+00 
R8801t1690 n8802 n1691 R=4.889e+02 
R8801t1790 n8802 n1791 R=8.970e+00 
R8801t2151 n8802 n2152 R=8.719e+00 
R8801t2800 n8802 n2801 R=2.418e+02 
R8802t2893 n8803 n2894 R=2.840e+00 
R8802t5304 n8803 n5305 R=1.411e+01 
R8802t6837 n8803 n6838 R=2.231e+01 
R8802t7597 n8803 n7598 R=4.492e+00 
R8802t3777 n8803 n3778 R=9.183e+01 
R8803t5857 n8804 n5858 R=7.350e+00 
R8803t7165 n8804 n7166 R=8.442e+00 
R8803t182 n8804 n183 R=6.064e+01 
R8803t2822 n8804 n2823 R=1.425e+01 
R8803t142 n8804 n143 R=5.947e+00 
R8804t1494 n8805 n1495 R=3.167e+01 
R8804t4546 n8805 n4547 R=2.236e+00 
R8804t8577 n8805 n8578 R=6.185e+01 
R8804t5687 n8805 n5688 R=1.014e+01 
R8804t5597 n8805 n5598 R=4.256e+00 
R8804t2174 n8805 n2175 R=1.086e+01 
R8805t1372 n8806 n1373 R=8.731e+00 
R8805t5422 n8806 n5423 R=8.927e+00 
R8805t2954 n8806 n2955 R=7.517e+00 
R8805t2709 n8806 n2710 R=1.042e+01 
R8805t71 n8806 n72 R=2.514e+00 
R8806t235 n8807 n236 R=3.631e+01 
R8806t2104 n8807 n2105 R=3.562e+00 
R8806t6207 n8807 n6208 R=7.239e+00 
R8806t8420 n8807 n8421 R=4.337e+00 
R8806t1720 n8807 n1721 R=5.301e+00 
R8807t4456 n8808 n4457 R=7.652e+00 
R8807t7548 n8808 n7549 R=1.886e+01 
R8807t4284 n8808 n4285 R=4.923e+00 
R8807t5117 n8808 n5118 R=8.855e+00 
R8808t2649 n8809 n2650 R=9.470e+00 
R8808t7663 n8809 n7664 R=2.902e+00 
R8808t3277 n8809 n3278 R=1.513e+01 
R8808t3481 n8809 n3482 R=1.412e+01 
R8808t684 n8809 n685 R=1.414e+02 
R8808t8258 n8809 n8259 R=1.676e+01 
R8809t2932 n8810 n2933 R=3.898e+00 
R8809t7214 n8810 n7215 R=6.713e+00 
R8809t1764 n8810 n1765 R=7.119e+00 
R8809t4990 n8810 n4991 R=1.877e+03 
R8809t8579 n8810 n8580 R=3.705e+00 
R8810t1130 n8811 n1131 R=1.815e+01 
R8810t2359 n8811 n2360 R=5.436e+00 
R8810t7925 n8811 n7926 R=3.205e+00 
R8810t5589 n8811 n5590 R=1.699e+01 
R8810t5361 n8811 n5362 R=4.521e+00 
R8810t7472 n8811 n7473 R=1.392e+01 
R8811t2770 n8812 n2771 R=1.735e+01 
R8811t3069 n8812 n3070 R=1.518e+02 
R8811t7145 n8812 n7146 R=4.899e+02 
R8811t1786 n8812 n1787 R=6.858e+00 
R8811t7920 n8812 n7921 R=1.214e+01 
R8811t3101 n8812 n3102 R=5.586e+00 
R8811t1030 n8812 n1031 R=2.314e+01 
R8811t3799 n8812 n3800 R=3.858e+00 
R8812t4637 n8813 n4638 R=2.659e+01 
R8812t7995 n8813 n7996 R=7.649e+00 
R8812t3505 n8813 n3506 R=4.203e+00 
R8812t7095 n8813 n7096 R=1.541e+01 
R8812t8372 n8813 n8373 R=6.659e+00 
R8813t4345 n8814 n4346 R=6.473e+00 
R8813t5693 n8814 n5694 R=4.648e+00 
R8813t3899 n8814 n3900 R=3.463e+01 
R8813t7960 n8814 n7961 R=3.650e+00 
R8813t1002 n8814 n1003 R=4.221e+01 
R8813t8224 n8814 n8225 R=8.095e+00 
R8814t4528 n8815 n4529 R=6.593e+00 
R8814t6302 n8815 n6303 R=4.773e+00 
R8814t8317 n8815 n8318 R=1.412e+01 
R8814t1119 n8815 n1120 R=9.692e+00 
R8814t2500 n8815 n2501 R=7.695e+00 
R8815t3380 n8816 n3381 R=4.011e+00 
R8815t6170 n8816 n6171 R=4.038e+01 
R8815t2398 n8816 n2399 R=6.567e+01 
R8815t12 n8816 n13 R=1.239e+01 
R8815t3005 n8816 n3006 R=6.608e+00 
R8816t1407 n8817 n1408 R=1.039e+00 
R8816t3415 n8817 n3416 R=7.480e+01 
R8816t3715 n8817 n3716 R=6.975e+02 
R8816t1313 n8817 n1314 R=2.898e+00 
R8816t7468 n8817 n7469 R=5.713e+00 
R8817t1639 n8818 n1640 R=5.281e+00 
R8817t7287 n8818 n7288 R=1.364e+01 
R8817t3389 n8818 n1 R=2.416e+01 
R8817t2964 n8818 n2965 R=3.916e+00 
R8817t3924 n8818 n3925 R=1.673e+01 
R8817t4969 n8818 n4970 R=9.055e+00 
R8818t836 n8819 n837 R=3.716e+00 
R8818t890 n8819 n891 R=3.081e+00 
R8818t7608 n8819 n7609 R=3.317e+01 
R8819t1386 n8820 n1387 R=1.028e+01 
R8819t6420 n8820 n6421 R=2.586e+01 
R8819t6427 n8820 n6428 R=8.602e+00 
R8819t833 n8820 n834 R=6.862e+00 
R8819t2899 n8820 n2900 R=1.181e+01 
R8819t8719 n8820 n8720 R=4.701e+00 
R8820t3814 n8821 n3815 R=1.366e+01 
R8820t5362 n8821 n5363 R=3.428e+00 
R8820t8792 n8821 n8793 R=3.719e+00 
R8820t3235 n8821 n3236 R=6.536e+00 
R8820t741 n8821 n742 R=1.702e+01 
R8821t5693 n8822 n5694 R=5.522e+00 
R8821t8813 n8822 n8814 R=1.334e+01 
R8821t747 n8822 n748 R=1.514e+01 
R8821t3103 n8822 n3104 R=6.485e+00 
R8821t3899 n8822 n3900 R=4.154e+00 
R8822t5261 n8823 n5262 R=2.280e+00 
R8822t5900 n8823 n5901 R=8.789e+00 
R8822t8603 n8823 n8604 R=2.122e+01 
R8822t5267 n8823 n5268 R=1.633e+00 
R8823t4434 n8824 n4435 R=8.661e+00 
R8823t5559 n8824 n5560 R=1.177e+01 
R8823t2119 n8824 n2120 R=7.549e+00 
R8823t8555 n8824 n8556 R=6.308e+00 
R8823t3999 n8824 n4000 R=4.047e+01 
R8823t2989 n8824 n2990 R=6.228e+00 
R8823t7604 n8824 n7605 R=1.284e+01 
R8824t4101 n8825 n4102 R=5.325e+00 
R8824t5068 n8825 n5069 R=1.382e+01 
R8824t1274 n8825 n1275 R=9.009e+00 
R8824t5792 n8825 n5793 R=2.269e+01 
R8825t7501 n8826 n7502 R=2.356e+01 
R8825t369 n8826 n370 R=4.506e+01 
R8825t1573 n8826 n1574 R=7.180e+01 
R8825t190 n8826 n191 R=1.336e+01 
R8825t3379 n8826 n3380 R=4.328e+00 
R8825t8732 n8826 n8733 R=4.743e+00 
R8825t8164 n8826 n8165 R=2.660e+01 
R8826t4539 n8827 n4540 R=4.785e+01 
R8826t4233 n8827 n4234 R=2.030e+01 
R8826t6388 n8827 n6389 R=8.737e+00 
R8827t8775 n8828 n8776 R=1.322e+01 
R8827t2376 n8828 n2377 R=3.528e+00 
R8827t3335 n8828 n3336 R=7.040e+00 
R8827t7355 n8828 n7356 R=1.527e+01 
R8827t265 n8828 n266 R=1.325e+01 
R8827t6218 n8828 n6219 R=4.506e+01 
R8828t1514 n8829 n1515 R=2.615e+00 
R8828t3199 n8829 n3200 R=3.786e+00 
R8828t6286 n8829 n6287 R=8.111e+00 
R8828t4219 n8829 n4220 R=1.176e+02 
R8828t8618 n8829 n8619 R=7.465e+00 
R8829t2620 n8830 n2621 R=1.407e+00 
R8829t4876 n8830 n4877 R=1.683e+02 
R8829t6674 n8830 n6675 R=5.234e+00 
R8829t7898 n8830 n7899 R=3.177e+00 
R8829t3577 n8830 n3578 R=5.249e+01 
R8830t7323 n8831 n7324 R=5.461e+00 
R8830t7383 n8831 n7384 R=5.181e+00 
R8830t3485 n8831 n3486 R=1.164e+01 
R8830t5175 n8831 n5176 R=4.281e+00 
R8830t43 n8831 n44 R=2.665e+01 
R8831t8622 n8832 n8623 R=1.215e+02 
R8831t4991 n8832 n4992 R=1.661e+01 
R8831t8549 n8832 n8550 R=6.309e+00 
R8831t5168 n8832 n5169 R=3.278e+01 
R8831t7895 n8832 n7896 R=3.975e+00 
R8831t6884 n8832 n6885 R=2.532e+01 
R8831t3266 n8832 n3267 R=2.938e+01 
R8832t314 n8833 n315 R=5.992e+00 
R8832t4611 n8833 n4612 R=1.749e+01 
R8832t903 n8833 n904 R=1.422e+01 
R8832t4359 n8833 n4360 R=1.963e+01 
R8832t8330 n8833 n8331 R=1.022e+01 
R8832t2986 n8833 n2987 R=1.860e+01 
R8833t28 n8834 n29 R=5.649e+02 
R8833t6611 n8834 n6612 R=1.365e+01 
R8833t8653 n8834 n8654 R=5.851e+00 
R8833t266 n8834 n267 R=6.483e+00 
R8834t198 n8835 n199 R=6.727e+01 
R8834t743 n8835 n744 R=7.055e+00 
R8834t3960 n8835 n3961 R=2.182e+01 
R8834t8638 n8835 n8639 R=6.406e+00 
R8834t850 n8835 n851 R=8.000e+00 
R8834t666 n8835 n667 R=5.693e+01 
R8835t5118 n8836 n5119 R=3.731e+01 
R8835t1014 n8836 n1015 R=2.773e+00 
R8835t3359 n8836 n3360 R=3.364e+01 
R8835t5840 n8836 n5841 R=3.356e+00 
R8836t421 n8837 n422 R=1.248e+01 
R8836t5066 n8837 n5067 R=3.416e+00 
R8836t616 n8837 n617 R=3.341e+01 
R8836t7498 n8837 n7499 R=1.173e+01 
R8836t4405 n8837 n4406 R=1.046e+01 
R8836t6532 n8837 n6533 R=3.922e+00 
R8837t8173 n8838 n8174 R=9.934e+00 
R8837t6409 n8838 n6410 R=2.841e+01 
R8837t5360 n8838 n5361 R=2.898e+02 
R8837t5402 n8838 n5403 R=9.151e+00 
R8837t6872 n8838 n6873 R=6.262e+00 
R8837t4051 n8838 n4052 R=4.937e+00 
R8838t3375 n8839 n3376 R=1.799e+00 
R8838t8263 n8839 n8264 R=3.359e+01 
R8838t6218 n8839 n6219 R=1.449e+01 
R8838t5145 n8839 n5146 R=2.398e+01 
R8838t4500 n8839 n4501 R=9.989e+00 
R8838t2984 n8839 n2985 R=4.053e+00 
R8838t3259 n8839 n3260 R=3.755e+01 
R8839t2057 n8840 n2058 R=1.376e+01 
R8839t5387 n8840 n5388 R=2.852e+01 
R8839t5713 n8840 n5714 R=3.984e+00 
R8839t66 n8840 n67 R=8.715e+01 
R8839t3192 n8840 n3193 R=2.303e+01 
R8839t5476 n8840 n5477 R=4.704e+00 
R8840t4368 n8841 n4369 R=8.603e+00 
R8840t5072 n8841 n5073 R=2.373e+01 
R8840t7112 n8841 n7113 R=7.237e+01 
R8840t6032 n8841 n6033 R=3.150e+00 
R8840t5479 n8841 n5480 R=6.586e+00 
R8840t5303 n8841 n5304 R=5.437e+00 
R8841t2743 n8842 n2744 R=4.695e+00 
R8841t8727 n8842 n8728 R=4.697e+00 
R8841t9 n8842 n10 R=1.075e+01 
R8841t7561 n8842 n7562 R=1.118e+01 
R8841t1826 n8842 n1827 R=7.543e+00 
R8841t2437 n8842 n2438 R=3.761e+01 
R8842t5708 n1 n5709 R=1.006e+01 
R8842t6158 n1 n6159 R=5.004e+00 
R8842t327 n1 n328 R=1.110e+01 
R8843t323 n8844 n324 R=5.556e+01 
R8843t3342 n8844 n3343 R=1.760e+01 
R8843t7166 n8844 n7167 R=3.622e+01 
R8843t7089 n8844 n7090 R=1.542e+01 
R8843t3890 n8844 n3891 R=3.072e+00 
R8843t4362 n8844 n4363 R=1.631e+01 
R8843t8523 n8844 n8524 R=4.689e+00 
R8844t3343 n8845 n3344 R=2.088e+01 
R8844t5105 n8845 n5106 R=3.821e+00 
R8844t3771 n8845 n3772 R=1.108e+01 
R8844t871 n8845 n872 R=5.339e+00 
R8844t5208 n8845 n5209 R=9.731e+00 
R8845t4902 n8846 n4903 R=2.669e+00 
R8845t7792 n8846 n7793 R=2.109e+01 
R8845t3334 n8846 n3335 R=4.479e+00 
R8845t6832 n8846 n6833 R=1.625e+01 
R8845t2862 n8846 n2863 R=6.084e+00 
R8846t1914 n8847 n1915 R=1.731e+01 
R8846t3607 n8847 n3608 R=3.775e+00 
R8846t3715 n8847 n3716 R=6.837e+00 
R8846t5221 n8847 n5222 R=5.611e+02 
R8846t1108 n8847 n1109 R=7.039e+00 
R8846t1738 n8847 n1739 R=5.252e+00 
R8847t8142 n8848 n8143 R=1.046e+01 
R8847t8197 n8848 n8198 R=3.564e+00 
R8847t6240 n8848 n6241 R=9.172e+00 
R8847t4898 n8848 n4899 R=8.236e+00 
R8847t7027 n8848 n7028 R=1.013e+01 
R8848t167 n8849 n168 R=8.684e+00 
R8848t4547 n8849 n4548 R=3.926e+00 
R8848t3579 n8849 n3580 R=1.528e+01 
R8848t392 n8849 n393 R=2.252e+02 
R8848t8586 n8849 n8587 R=2.364e+00 
R8848t6536 n8849 n6537 R=1.017e+01 
R8849t4442 n8850 n4443 R=7.577e+00 
R8849t8433 n8850 n8434 R=4.525e+01 
R8849t7950 n8850 n7951 R=1.965e+01 
R8849t6492 n8850 n6493 R=7.638e+00 
R8849t414 n8850 n415 R=1.922e+01 
R8849t5122 n8850 n5123 R=1.091e+01 
R8849t7309 n8850 n7310 R=8.198e+00 
R8849t7161 n8850 n7162 R=2.217e+01 
R8850t5532 n8851 n5533 R=3.086e+01 
R8850t8516 n8851 n8517 R=1.890e+00 
R8850t5720 n8851 n5721 R=2.829e+00 
R8850t2999 n8851 n3000 R=3.233e+01 
R8850t7480 n8851 n7481 R=6.106e+00 
R8851t598 n8852 n599 R=1.654e+01 
R8851t4328 n8852 n4329 R=9.957e+00 
R8851t2270 n8852 n2271 R=1.408e+01 
R8851t1946 n8852 n1947 R=4.242e+01 
R8851t8366 n8852 n8367 R=1.110e+01 
R8851t7784 n8852 n7785 R=5.443e+00 
R8852t692 n8853 n1 R=7.641e+00 
R8852t1161 n8853 n1162 R=7.587e+00 
R8852t2900 n8853 n1 R=1.899e+02 
R8852t7416 n8853 n7417 R=5.032e+00 
R8852t8274 n8853 n8275 R=7.665e+00 
R8852t706 n8853 n707 R=4.612e+00 
R8853t3826 n8854 n3827 R=4.812e+01 
R8853t8218 n8854 n8219 R=6.339e+00 
R8853t7900 n8854 n7901 R=3.925e+01 
R8853t4037 n8854 n4038 R=5.088e+00 
R8853t4505 n8854 n4506 R=1.707e+01 
R8853t3992 n8854 n3993 R=5.641e+00 
R8853t7778 n8854 n7779 R=4.633e+00 
R8854t4921 n8855 n4922 R=2.525e+01 
R8854t1114 n8855 n1115 R=1.172e+01 
R8854t7342 n8855 n7343 R=1.701e+01 
R8854t7606 n8855 n7607 R=3.622e+00 
R8854t3947 n8855 n3948 R=2.343e+01 
R8854t2154 n8855 n2155 R=4.552e+01 
R8854t7204 n8855 n7205 R=1.076e+01 
R8855t6206 n8856 n6207 R=1.207e+01 
R8855t4291 n8856 n4292 R=5.148e+00 
R8855t815 n8856 n816 R=7.113e+00 
R8855t5460 n8856 n5461 R=5.125e+00 
R8856t8285 n8857 n8286 R=1.665e+00 
R8856t3385 n8857 n3386 R=1.040e+01 
R8856t4280 n8857 n4281 R=9.382e+00 
R8856t3909 n8857 n3910 R=3.921e+00 
R8856t7296 n8857 n7297 R=3.402e+01 
R8857t2004 n8858 n2005 R=7.382e+00 
R8857t8432 n8858 n8433 R=4.890e+01 
R8857t3011 n8858 n3012 R=2.571e+00 
R8857t1475 n8858 n1476 R=2.290e+01 
R8857t3793 n8858 n3794 R=1.353e+01 
R8857t8593 n8858 n8594 R=3.854e+00 
R8858t1276 n8859 n1277 R=3.938e+01 
R8858t2601 n8859 n2602 R=4.384e+00 
R8858t5880 n8859 n5881 R=1.292e+01 
R8858t3295 n8859 n3296 R=3.736e+00 
R8858t2716 n8859 n2717 R=6.485e+00 
R8858t6911 n8859 n6912 R=9.516e+00 
R8859t7642 n8860 n7643 R=2.483e+00 
R8859t6141 n8860 n6142 R=3.889e+01 
R8859t7612 n8860 n7613 R=8.806e+00 
R8859t3176 n8860 n3177 R=5.030e+00 
R8859t4789 n8860 n4790 R=1.709e+01 
R8860t499 n8861 n500 R=5.443e+01 
R8860t7970 n8861 n7971 R=1.091e+01 
R8860t1169 n8861 n1170 R=2.153e+00 
R8860t6168 n8861 n6169 R=6.359e+01 
R8860t2698 n8861 n2699 R=3.891e+02 
R8860t2669 n8861 n2670 R=3.899e+00 
R8860t5893 n8861 n5894 R=6.068e+00 
R8861t1632 n8862 n1633 R=7.508e+00 
R8861t8449 n8862 n8450 R=2.619e+01 
R8861t5949 n8862 n5950 R=2.681e+00 
R8861t8563 n8862 n8564 R=1.013e+01 
R8861t2642 n8862 n2643 R=9.131e+00 
R8861t2350 n8862 n2351 R=1.032e+01 
R8862t4083 n8863 n4084 R=2.313e+00 
R8862t5256 n8863 n5257 R=6.149e+00 
R8862t1958 n8863 n1959 R=1.748e+01 
R8862t6136 n8863 n6137 R=3.393e+01 
R8862t8476 n8863 n8477 R=2.800e+00 
R8863t2607 n8864 n2608 R=6.486e+00 
R8863t4426 n8864 n4427 R=3.595e+00 
R8863t4488 n8864 n4489 R=1.383e+01 
R8863t8133 n8864 n8134 R=2.838e+00 
R8863t6725 n8864 n6726 R=1.915e+02 
R8863t1599 n8864 n1600 R=2.064e+01 
R8864t6741 n8865 n6742 R=3.108e+00 
R8864t1935 n8865 n1936 R=4.045e+00 
R8864t8045 n8865 n8046 R=7.688e+00 
R8864t285 n8865 n286 R=1.633e+01 
R8865t3313 n8866 n3314 R=8.864e+00 
R8865t6059 n8866 n6060 R=7.817e+00 
R8865t662 n8866 n663 R=6.052e+00 
R8865t284 n8866 n285 R=2.137e+02 
R8865t3430 n8866 n3431 R=4.420e+00 
R8865t7051 n8866 n7052 R=7.170e+01 
R8865t1554 n8866 n1555 R=1.000e+01 
R8866t3925 n8867 n3926 R=3.246e+02 
R8866t8004 n8867 n8005 R=7.903e+00 
R8866t2887 n8867 n2888 R=5.447e+00 
R8866t2549 n8867 n2550 R=1.291e+01 
R8866t2137 n8867 n2138 R=1.272e+01 
R8866t3354 n8867 n3355 R=5.283e+00 
R8866t513 n8867 n514 R=1.714e+01 
R8867t5351 n8868 n5352 R=6.200e+00 
R8867t6474 n8868 n6475 R=1.829e+01 
R8867t7837 n8868 n7838 R=2.336e+01 
R8867t1826 n8868 n1827 R=8.078e+00 
R8867t7786 n8868 n7787 R=1.050e+01 
R8867t4674 n8868 n4675 R=1.439e+01 
R8867t3876 n8868 n3877 R=5.361e+00 
R8868t6222 n8869 n6223 R=2.023e+00 
R8868t8560 n8869 n8561 R=1.109e+01 
R8868t2193 n8869 n2194 R=8.236e+00 
R8868t4095 n8869 n4096 R=3.462e+00 
R8868t6799 n8869 n6800 R=1.486e+01 
R8869t5327 n8870 n5328 R=7.604e+00 
R8869t5465 n8870 n5466 R=3.574e+00 
R8869t3109 n8870 n3110 R=1.510e+02 
R8869t4514 n8870 n4515 R=2.047e+00 
R8869t2399 n8870 n2400 R=6.341e+00 
R8870t2826 n8871 n2827 R=2.525e+00 
R8870t8620 n8871 n8621 R=1.537e+01 
R8870t814 n8871 n815 R=1.057e+01 
R8870t6576 n8871 n6577 R=2.747e+02 
R8870t3921 n8871 n3922 R=7.842e+00 
R8870t5117 n8871 n5118 R=4.628e+01 
R8871t3251 n8872 n3252 R=8.956e+00 
R8871t5725 n8872 n5726 R=1.626e+01 
R8871t3390 n8872 n3391 R=3.052e+00 
R8871t5293 n8872 n5294 R=1.212e+02 
R8871t4324 n8872 n4325 R=1.083e+01 
R8871t7040 n8872 n7041 R=3.980e+00 
R8871t128 n8872 n129 R=4.449e+01 
R8872t723 n8873 n724 R=4.433e+00 
R8872t2025 n8873 n2026 R=1.692e+01 
R8872t8054 n8873 n8055 R=5.677e+00 
R8872t8261 n8873 n8262 R=2.627e+00 
R8873t2414 n8874 n2415 R=8.125e+00 
R8873t8658 n8874 n8659 R=1.376e+01 
R8873t5825 n8874 n5826 R=7.964e+00 
R8873t1291 n8874 n1292 R=2.504e+01 
R8873t3859 n8874 n3860 R=5.353e+00 
R8874t1462 n8875 n1463 R=9.966e+01 
R8874t7582 n8875 n7583 R=2.906e+00 
R8874t3985 n8875 n3986 R=1.627e+01 
R8874t7318 n8875 n7319 R=5.071e+00 
R8874t4366 n8875 n4367 R=3.319e+00 
R8875t4834 n8876 n4835 R=1.851e+00 
R8876t7092 n8877 n7093 R=2.369e+00 
R8876t8049 n8877 n8050 R=1.332e+01 
R8876t8074 n8877 n8075 R=2.572e+01 
R8876t8386 n8877 n8387 R=3.755e+00 
R8876t3768 n8877 n3769 R=1.875e+01 
R8876t8101 n8877 n8102 R=2.092e+01 
R8876t6423 n8877 n6424 R=2.673e+01 
R8876t3157 n8877 n3158 R=3.458e+01 
R8877t2020 n8878 n2021 R=1.085e+01 
R8877t3005 n8878 n3006 R=3.669e+00 
R8877t8637 n8878 n8638 R=5.933e+00 
R8877t6931 n8878 n6932 R=2.306e+01 
R8877t6822 n8878 n6823 R=1.160e+01 
R8878t588 n8879 n589 R=6.622e+01 
R8878t4667 n8879 n4668 R=4.932e+00 
R8878t6235 n8879 n6236 R=2.468e+00 
R8878t7818 n8879 n7819 R=1.026e+01 
R8878t5343 n8879 n5344 R=5.603e+00 
R8879t2118 n8880 n2119 R=5.481e+00 
R8879t4958 n8880 n4959 R=7.110e+01 
R8879t440 n8880 n441 R=6.493e+00 
R8879t7873 n8880 n7874 R=4.858e+01 
R8879t1249 n8880 n1250 R=1.808e+01 
R8879t4166 n8880 n4167 R=2.761e+00 
R8880t2685 n8881 n2686 R=1.444e+01 
R8880t7227 n8881 n7228 R=1.608e+01 
R8880t2545 n8881 n2546 R=4.222e+00 
R8880t4113 n8881 n4114 R=4.429e+00 
R8880t2657 n8881 n2658 R=2.212e+01 
R8880t7893 n8881 n7894 R=9.010e+00 
R8881t206 n8882 n207 R=1.425e+01 
R8881t2489 n8882 n2490 R=1.481e+01 
R8881t2488 n8882 n2489 R=4.252e+01 
R8881t5753 n8882 n5754 R=2.300e+01 
R8881t1022 n8882 n1023 R=4.889e+00 
R8882t2579 n8883 n2580 R=2.541e+00 
R8882t6786 n8883 n6787 R=3.005e+00 
R8882t4507 n8883 n4508 R=6.188e+00 
R8882t8019 n8883 n8020 R=1.358e+01 
R8882t526 n8883 n527 R=6.485e+01 
R8883t2390 n8884 n2391 R=2.515e+00 
R8883t6458 n8884 n6459 R=6.179e+00 
R8883t8026 n8884 n8027 R=1.506e+01 
R8883t4058 n8884 n4059 R=3.371e+00 
R8884t1717 n8885 n1718 R=3.201e+00 
R8884t4230 n8885 n4231 R=2.633e+01 
R8884t2207 n8885 n2208 R=5.221e+00 
R8884t1347 n8885 n1348 R=6.148e+00 
R8884t1319 n8885 n1320 R=9.639e+00 
R8885t4637 n8886 n4638 R=2.253e+01 
R8885t6896 n8886 n6897 R=1.332e+02 
R8885t8372 n8886 n8373 R=2.806e+00 
R8885t7152 n8886 n7153 R=8.026e+01 
R8885t7403 n8886 n7404 R=2.949e+00 
R8885t2228 n8886 n2229 R=1.310e+01 
R8885t3077 n8886 n3078 R=1.886e+01 
R8885t3701 n8886 n3702 R=2.003e+01 
R8886t5112 n8887 n5113 R=5.255e+01 
R8886t8742 n8887 n8743 R=1.948e+00 
R8886t1496 n8887 n1497 R=2.081e+01 
R8886t8082 n8887 n8083 R=2.839e+00 
R8886t2039 n8887 n2040 R=6.248e+01 
R8887t626 n8888 n627 R=1.045e+01 
R8887t1684 n8888 n1685 R=4.565e+00 
R8887t3574 n8888 n3575 R=1.164e+01 
R8887t3744 n8888 n3745 R=1.884e+01 
R8888t5883 n8889 n5884 R=1.923e+01 
R8888t4011 n8889 n4012 R=5.846e+01 
R8888t1676 n8889 n1677 R=3.287e+02 
R8888t1657 n8889 n1658 R=1.905e+00 
R8888t7338 n8889 n7339 R=2.349e+01 
R8888t2139 n8889 n2140 R=5.134e+00 
R8889t1451 n8890 n1452 R=4.507e+00 
R8889t6864 n8890 n6865 R=2.965e+00 
R8889t2480 n8890 n2481 R=1.011e+01 
R8889t2638 n8890 n2639 R=3.337e+01 
R8889t6917 n8890 n6918 R=4.986e+01 
R8890t1392 n8891 n1393 R=5.232e+01 
R8890t4499 n8891 n4500 R=1.335e+01 
R8890t3227 n8891 n3228 R=1.235e+01 
R8890t3569 n8891 n3570 R=2.408e+02 
R8890t5497 n8891 n5498 R=6.292e+00 
R8890t456 n8891 n457 R=6.961e+00 
R8890t2275 n8891 n2276 R=1.864e+01 
R8891t1115 n8892 n1116 R=4.431e+00 
R8891t1150 n8892 n1151 R=7.138e+00 
R8891t2996 n8892 n2997 R=1.736e+01 
R8891t5169 n8892 n5170 R=3.861e+00 
R8891t5756 n8892 n5757 R=1.469e+01 
R8892t1269 n8893 n1270 R=3.566e+00 
R8892t2794 n8893 n2795 R=8.292e+00 
R8892t8712 n8893 n8713 R=3.266e+00 
R8892t7981 n8893 n7982 R=2.612e+01 
R8893t5650 n8894 n5651 R=2.259e+00 
R8893t8450 n8894 n8451 R=2.518e+00 
R8893t1580 n8894 n1581 R=3.932e+00 
R8894t5299 n8895 n5300 R=6.835e+00 
R8894t256 n8895 n257 R=5.846e+00 
R8894t2412 n8895 n2413 R=5.399e+00 
R8895t914 n8896 n915 R=8.034e+00 
R8895t1938 n8896 n1939 R=1.606e+02 
R8895t764 n8896 n765 R=1.696e+01 
R8895t671 n8896 n672 R=6.744e+00 
R8895t5660 n8896 n5661 R=1.889e+01 
R8895t2528 n8896 n2529 R=3.186e+00 
R8896t3968 n8897 n3969 R=2.421e+00 
R8896t4451 n8897 n4452 R=7.102e+01 
R8896t5544 n8897 n5545 R=5.827e+00 
R8896t4804 n8897 n4805 R=2.833e+00 
R8897t5369 n8898 n5370 R=7.333e+00 
R8897t7293 n8898 n7294 R=2.324e+01 
R8897t7283 n8898 n7284 R=3.883e+00 
R8897t2250 n8898 n2251 R=1.427e+01 
R8897t7489 n8898 n7490 R=8.914e+00 
R8897t5986 n8898 n5987 R=1.196e+01 
R8897t2351 n8898 n2352 R=1.605e+01 
R8898t927 n8899 n928 R=2.348e+00 
R8898t8786 n8899 n8787 R=1.298e+01 
R8898t8191 n8899 n8192 R=1.213e+01 
R8898t288 n8899 n289 R=1.068e+01 
R8898t1928 n8899 n1929 R=3.458e+00 
R8899t6305 n8900 n6306 R=3.460e+00 
R8899t8121 n8900 n8122 R=1.990e+01 
R8899t2415 n8900 n2416 R=2.377e+01 
R8899t6854 n8900 n6855 R=8.902e+00 
R8899t5348 n8900 n5349 R=4.448e+01 
R8899t4868 n8900 n4869 R=4.498e+00 
R8899t2722 n8900 n2723 R=2.493e+02 
R8899t2302 n8900 n2303 R=7.864e+00 
R8900t585 n8901 n586 R=1.978e+01 
R8900t3312 n8901 n3313 R=8.806e+01 
R8900t2752 n8901 n2753 R=3.874e+00 
R8900t794 n8901 n795 R=5.646e+00 
R8900t1784 n8901 n1785 R=2.831e+01 
R8900t6706 n8901 n6707 R=2.143e+00 
R8901t4995 n8902 n4996 R=3.019e+01 
R8901t8005 n8902 n8006 R=3.640e+00 
R8901t123 n8902 n124 R=2.967e+00 
R8901t1767 n8902 n1768 R=8.020e+00 
R8902t6006 n8903 n6007 R=6.404e+00 
R8902t1223 n8903 n1224 R=8.814e+00 
R8902t478 n8903 n479 R=1.080e+01 
R8902t3386 n8903 n3387 R=7.390e+01 
R8902t6055 n8903 n6056 R=5.950e+00 
R8902t1517 n8903 n1518 R=6.770e+00 
R8903t7066 n8904 n7067 R=2.657e+00 
R8903t8099 n8904 n8100 R=9.144e+01 
R8903t3518 n8904 n3519 R=4.114e+00 
R8903t3515 n8904 n3516 R=6.523e+00 
R8903t5034 n8904 n5035 R=1.125e+01 
R8903t118 n8904 n119 R=1.640e+01 
R8904t5818 n8905 n5819 R=7.028e+01 
R8904t8170 n8905 n8171 R=8.929e+01 
R8904t6998 n8905 n6999 R=1.664e+00 
R8904t3207 n8905 n3208 R=7.090e+01 
R8904t1588 n8905 n1589 R=8.226e+00 
R8904t2809 n8905 n2810 R=2.540e+00 
R8905t4927 n8906 n4928 R=4.112e+01 
R8905t8375 n8906 n8376 R=4.709e+00 
R8905t5246 n8906 n5247 R=2.216e+00 
R8905t1139 n8906 n1140 R=3.559e+00 
R8906t2278 n8907 n2279 R=4.068e+00 
R8906t5388 n8907 n5389 R=1.160e+02 
R8906t2508 n8907 n2509 R=4.697e+00 
R8906t3596 n8907 n3597 R=8.557e+00 
R8906t1170 n8907 n1171 R=5.024e+00 
R8907t5915 n8908 n5916 R=1.963e+01 
R8907t6150 n8908 n6151 R=2.336e+00 
R8907t2719 n8908 n2720 R=3.419e+00 
R8907t2233 n8908 n2234 R=4.478e+00 
R8908t1549 n8909 n1550 R=3.548e+00 
R8908t2111 n8909 n2112 R=1.522e+01 
R8908t7634 n8909 n7635 R=6.211e+00 
R8908t7245 n8909 n7246 R=1.579e+01 
R8908t802 n8909 n803 R=3.234e+00 
R8909t1269 n8910 n1270 R=6.632e+00 
R8909t3460 n8910 n3461 R=7.216e+00 
R8909t6315 n8910 n6316 R=1.140e+01 
R8909t214 n8910 n215 R=1.538e+01 
R8909t1556 n8910 n1557 R=7.007e+00 
R8910t5118 n8911 n5119 R=7.686e+01 
R8910t8835 n8911 n8836 R=4.056e+00 
R8910t5840 n8911 n5841 R=1.035e+01 
R8910t3512 n8911 n3513 R=1.777e+01 
R8910t557 n8911 n558 R=2.887e+00 
R8911t3886 n8912 n3887 R=4.227e+02 
R8911t8096 n8912 n8097 R=4.087e+00 
R8911t3618 n8912 n3619 R=5.166e+00 
R8911t4067 n8912 n4068 R=8.682e+01 
R8911t7330 n8912 n7331 R=8.026e+00 
R8911t97 n8912 n98 R=1.339e+01 
R8912t695 n8913 n696 R=1.207e+02 
R8912t1372 n8913 n1373 R=2.313e+01 
R8912t4067 n8913 n4068 R=1.221e+01 
R8912t3827 n8913 n3828 R=7.922e+00 
R8912t748 n8913 n749 R=5.719e+00 
R8912t7436 n8913 n7437 R=1.534e+02 
R8912t3428 n8913 n3429 R=3.815e+00 
R8913t1351 n8914 n1352 R=3.270e+00 
R8913t5191 n8914 n5192 R=9.302e+00 
R8913t25 n8914 n26 R=8.209e+00 
R8913t6335 n8914 n6336 R=1.671e+01 
R8913t4309 n8914 n4310 R=3.599e+00 
R8914t3024 n8915 n3025 R=4.294e+00 
R8914t7183 n8915 n7184 R=2.446e+00 
R8914t2514 n8915 n2515 R=1.372e+01 
R8914t2019 n8915 n2020 R=7.765e+01 
R8914t4709 n8915 n4710 R=4.967e+00 
R8915t6265 n8916 n6266 R=2.760e+00 
R8915t8229 n8916 n8230 R=9.131e+00 
R8915t8047 n8916 n8048 R=9.336e+00 
R8915t1735 n8916 n1736 R=4.735e+00 
R8916t260 n8917 n261 R=2.275e+01 
R8916t4236 n8917 n4237 R=8.952e+00 
R8916t7257 n8917 n7258 R=2.981e+00 
R8916t2471 n8917 n2472 R=1.979e+01 
R8916t8196 n8917 n8197 R=1.840e+00 
R8917t3057 n8918 n3058 R=4.028e+00 
R8917t5730 n8918 n5731 R=1.603e+01 
R8917t2680 n8918 n2681 R=5.523e+00 
R8917t3373 n8918 n3374 R=1.992e+01 
R8917t8596 n8918 n8597 R=1.329e+01 
R8917t1729 n8918 n1730 R=1.124e+01 
R8918t4479 n8919 n4480 R=7.717e+00 
R8918t6099 n8919 n6100 R=1.567e+01 
R8918t4508 n8919 n4509 R=1.190e+01 
R8918t5551 n8919 n5552 R=5.290e+01 
R8918t8582 n8919 n8583 R=2.309e+00 
R8918t7103 n8919 n7104 R=3.999e+00 
R8919t1706 n8920 n1707 R=9.415e+00 
R8919t5057 n8920 n5058 R=3.400e+00 
R8919t8437 n8920 n8438 R=7.501e+00 
R8919t6950 n8920 n6951 R=3.233e+00 
R8920t4186 n8921 n4187 R=5.932e+00 
R8920t5018 n8921 n5019 R=8.444e+00 
R8920t3994 n8921 n3995 R=3.946e+00 
R8920t1029 n8921 n1030 R=1.553e+01 
R8920t3844 n8921 n3845 R=4.737e+01 
R8920t1925 n8921 n1926 R=6.298e+02 
R8920t1776 n8921 n1777 R=1.703e+01 
R8920t7430 n8921 n7431 R=2.749e+01 
R8920t1120 n8921 n1121 R=1.175e+01 
R8921t4827 n8922 n4828 R=4.664e+00 
R8921t1706 n8922 n1707 R=1.006e+01 
R8921t6802 n8922 n6803 R=9.570e+00 
R8921t1769 n8922 n1770 R=1.079e+01 
R8921t848 n8922 n849 R=1.351e+01 
R8921t7105 n8922 n7106 R=6.705e+01 
R8922t6068 n8923 n6069 R=5.568e+00 
R8922t8640 n8923 n8641 R=4.298e+01 
R8922t4592 n8923 n4593 R=9.606e+00 
R8922t514 n8923 n515 R=2.970e+00 
R8923t3594 n8924 n3595 R=3.237e+00 
R8923t544 n8924 n545 R=3.011e+01 
R8923t4591 n8924 n4592 R=8.526e+00 
R8923t6089 n8924 n6090 R=1.164e+01 
R8923t8328 n8924 n8329 R=7.168e+00 
R8924t3862 n8925 n3863 R=2.585e+00 
R8924t8329 n8925 n8330 R=1.618e+01 
R8924t6719 n8925 n6720 R=4.839e+01 
R8924t2026 n8925 n2027 R=1.950e+01 
R8924t6477 n8925 n6478 R=1.110e+01 
R8924t5145 n8925 n5146 R=6.581e+00 
R8924t4500 n8925 n4501 R=1.710e+01 
R8925t4880 n1 n4881 R=4.463e+00 
R8925t8753 n1 n8754 R=5.165e+00 
R8925t7844 n1 n7845 R=1.962e+01 
R8925t8680 n1 n8681 R=1.089e+01 
R8926t2775 n8927 n2776 R=2.222e+00 
R8926t5849 n8927 n5850 R=2.609e+01 
R8926t3576 n8927 n3577 R=2.063e+01 
R8926t2482 n8927 n2483 R=3.465e+00 
R8926t4509 n8927 n4510 R=1.933e+01 
R8926t5955 n8927 n5956 R=1.665e+01 
R8927t1071 n8928 n1072 R=3.467e+00 
R8927t5141 n8928 n5142 R=4.425e+01 
R8927t2927 n8928 n2928 R=2.198e+00 
R8927t2967 n8928 n2968 R=7.912e+00 
R8927t2477 n8928 n2478 R=2.464e+01 
R8928t1803 n8929 n1804 R=1.063e+01 
R8928t3920 n8929 n3921 R=2.696e+00 
R8928t4265 n8929 n4266 R=7.008e+00 
R8928t5146 n8929 n5147 R=3.551e+01 
R8928t4025 n8929 n4026 R=2.623e+01 
R8928t4920 n8929 n4921 R=5.915e+00 
R8928t1065 n8929 n1066 R=4.286e+02 
R8929t1067 n8930 n1068 R=7.516e+00 
R8929t8311 n8930 n8312 R=3.169e+02 
R8929t4140 n8930 n4141 R=1.616e+01 
R8929t1918 n8930 n1919 R=3.957e+00 
R8929t503 n8930 n504 R=5.678e+00 
R8930t1350 n8931 n1351 R=3.442e+00 
R8930t5246 n8931 n5247 R=4.334e+00 
R8930t1307 n8931 n1308 R=1.079e+01 
R8930t3824 n8931 n3825 R=8.923e+00 
R8930t3818 n8931 n3819 R=3.174e+01 
R8931t6022 n8932 n6023 R=5.493e+00 
R8931t2377 n8932 n2378 R=4.164e+00 
R8931t708 n8932 n709 R=5.538e+00 
R8932t899 n8933 n900 R=2.946e+00 
R8932t8213 n8933 n8214 R=4.955e+00 
R8932t3140 n8933 n3141 R=1.659e+01 
R8932t1888 n8933 n1889 R=1.357e+01 
R8932t8088 n8933 n8089 R=8.319e+00 
R8933t5665 n8934 n5666 R=2.690e+00 
R8933t5706 n8934 n5707 R=2.379e+00 
R8933t618 n8934 n619 R=3.203e+00 
R8934t1990 n8935 n1991 R=1.864e+00 
R8934t2839 n8935 n2840 R=1.438e+01 
R8934t6696 n8935 n6697 R=8.770e+00 
R8934t7393 n8935 n7394 R=8.850e+00 
R8934t2933 n8935 n2934 R=5.368e+00 
R8935t5263 n8936 n5264 R=4.921e+00 
R8935t5508 n8936 n5509 R=9.743e+00 
R8935t1762 n8936 n1763 R=3.038e+00 
R8935t227 n8936 n228 R=5.294e+00 
R8936t1523 n8937 n1524 R=3.757e+00 
R8936t5610 n8937 n5611 R=5.463e+00 
R8936t7268 n8937 n7269 R=5.996e+00 
R8937t290 n8938 n291 R=2.204e+01 
R8937t308 n8938 n309 R=3.866e+00 
R8937t5983 n8938 n5984 R=9.370e+00 
R8937t8265 n8938 n8266 R=7.646e+00 
R8938t7167 n8939 n7168 R=2.338e+00 
R8938t3702 n8939 n3703 R=1.501e+01 
R8938t7670 n8939 n7671 R=1.187e+01 
R8938t6629 n8939 n6630 R=2.741e+01 
R8938t287 n8939 n288 R=5.099e+00 
R8939t2429 n8940 n2430 R=2.906e+01 
R8939t4874 n8940 n4875 R=6.707e+01 
R8939t7630 n8940 n7631 R=4.019e+00 
R8939t6975 n8940 n6976 R=1.229e+01 
R8939t3567 n8940 n3568 R=5.112e+00 
R8939t296 n8940 n297 R=4.185e+00 
R8940t5558 n8941 n5559 R=5.299e+00 
R8940t5791 n8941 n5792 R=9.765e+00 
R8940t8100 n8941 n8101 R=3.838e+01 
R8940t183 n8941 n184 R=7.097e+00 
R8940t738 n8941 n739 R=6.342e+00 
R8940t1281 n8941 n1282 R=5.160e+00 
R8941t4947 n8942 n4948 R=1.941e+00 
R8941t8634 n8942 n8635 R=8.866e+00 
R8941t5598 n8942 n5599 R=3.700e+00 
R8941t5530 n8942 n5531 R=1.088e+01 
R8942t4067 n8943 n4068 R=4.365e+01 
R8942t8912 n8943 n8913 R=3.607e+01 
R8942t8911 n8943 n8912 R=3.270e+00 
R8942t7330 n8943 n7331 R=1.939e+01 
R8942t381 n8943 n382 R=9.904e+00 
R8942t7300 n8943 n7301 R=2.939e+01 
R8942t6244 n8943 n6245 R=2.695e+01 
R8942t3827 n8943 n3828 R=2.019e+00 
R8943t7501 n8944 n7502 R=3.007e+00 
R8943t8825 n8944 n8826 R=4.001e+00 
R8943t369 n8944 n370 R=2.397e+00 
R8943t5280 n8944 n5281 R=5.966e+02 
R8943t7974 n8944 n7975 R=3.768e+01 
R8944t2524 n8945 n2525 R=8.923e+00 
R8944t3984 n8945 n3985 R=3.434e+00 
R8944t109 n8945 n110 R=5.720e+00 
R8944t4152 n8945 n4153 R=4.840e+00 
R8944t8179 n8945 n8180 R=9.816e+00 
R8945t2492 n8946 n2493 R=1.125e+01 
R8945t6838 n8946 n6839 R=3.500e+00 
R8945t8566 n8946 n8567 R=4.010e+01 
R8945t4707 n8946 n4708 R=1.870e+01 
R8945t7382 n8946 n7383 R=1.888e+00 
R8946t7031 n8947 n7032 R=1.457e+01 
R8946t6316 n8947 n6317 R=3.831e+00 
R8947t202 n8948 n203 R=5.606e+01 
R8947t8330 n8948 n8331 R=9.256e+00 
R8947t8832 n8948 n8833 R=4.551e+00 
R8947t4359 n8948 n4360 R=7.066e+01 
R8947t3646 n8948 n3647 R=6.617e+00 
R8947t191 n8948 n192 R=8.489e+00 
R8947t2647 n8948 n2648 R=6.175e+00 
R8948t4332 n8949 n4333 R=1.351e+01 
R8948t8367 n8949 n8368 R=6.729e+00 
R8948t8139 n8949 n8140 R=2.722e+01 
R8948t75 n8949 n76 R=2.844e+00 
R8948t4463 n8949 n4464 R=1.667e+01 
R8948t3731 n8949 n3732 R=6.245e+00 
R8948t3797 n8949 n3798 R=6.177e+02 
R8949t276 n8950 n277 R=4.513e+00 
R8949t3992 n8950 n3993 R=8.038e+00 
R8949t8508 n8950 n8509 R=5.423e+00 
R8949t4300 n8950 n4301 R=1.239e+01 
R8950t3591 n8951 n3592 R=8.981e+00 
R8950t7342 n8951 n7343 R=2.628e+01 
R8950t7626 n8951 n7627 R=1.040e+01 
R8950t4943 n8951 n4944 R=1.084e+01 
R8950t2186 n8951 n2187 R=7.829e+00 
R8950t3714 n8951 n3715 R=1.424e+01 
R8950t5546 n8951 n5547 R=7.938e+00 
R8951t4263 n8952 n4264 R=3.133e+02 
R8951t8798 n8952 n8799 R=6.608e+00 
R8951t146 n8952 n147 R=3.411e+00 
R8951t3762 n8952 n3763 R=1.409e+01 
R8951t6046 n8952 n6047 R=5.360e+00 
R8952t1428 n8953 n1429 R=6.059e+00 
R8952t8686 n8953 n8687 R=8.237e+00 
R8952t2017 n8953 n2018 R=1.317e+01 
R8952t2213 n8953 n2214 R=1.023e+01 
R8952t5384 n8953 n5385 R=5.879e+00 
R8953t5325 n8954 n5326 R=2.843e+00 
R8953t7532 n8954 n7533 R=1.026e+01 
R8953t8417 n8954 n8418 R=1.231e+01 
R8953t4416 n8954 n4417 R=6.877e+00 
R8953t3620 n8954 n3621 R=4.969e+00 
R8954t4648 n8955 n4649 R=6.724e+00 
R8954t5550 n8955 n5551 R=7.775e+00 
R8954t1321 n8955 n1322 R=1.318e+01 
R8954t8358 n8955 n8359 R=3.420e+01 
R8954t8271 n8955 n8272 R=6.622e+00 
R8954t3486 n8955 n3487 R=3.472e+00 
R8954t7010 n8955 n7011 R=5.349e+01 
R8955t765 n8956 n766 R=1.546e+01 
R8955t1808 n8956 n1809 R=4.764e+00 
R8955t8607 n8956 n8608 R=9.303e+00 
R8955t4625 n8956 n4626 R=6.905e+00 
R8955t4006 n8956 n4007 R=9.460e+00 
R8956t5613 n8957 n5614 R=8.490e+01 
R8956t7367 n8957 n7368 R=7.063e+00 
R8956t5951 n8957 n5952 R=3.061e+00 
R8956t2727 n8957 n2728 R=2.075e+00 
R8957t7747 n8958 n7748 R=1.705e+00 
R8957t5086 n8958 n5087 R=1.272e+01 
R8957t3468 n8958 n3469 R=1.526e+01 
R8958t966 n8959 n967 R=3.949e+01 
R8958t3290 n8959 n3291 R=7.251e+00 
R8958t5780 n8959 n5781 R=9.910e+00 
R8958t6327 n8959 n6328 R=7.360e+00 
R8958t1731 n8959 n1732 R=4.522e+00 
R8959t2318 n8960 n2319 R=6.252e+01 
R8959t6788 n8960 n6789 R=5.647e+00 
R8959t7598 n8960 n7599 R=1.289e+01 
R8959t8311 n8960 n8312 R=3.746e+00 
R8959t8929 n8960 n8930 R=6.389e+00 
R8959t4140 n8960 n4141 R=4.347e+01 
R8960t2361 n8961 n2362 R=2.054e+00 
R8960t4972 n8961 n4973 R=1.190e+01 
R8960t4532 n8961 n4533 R=6.370e+01 
R8960t3133 n8961 n3134 R=3.084e+00 
R8961t6435 n8962 n6436 R=1.925e+01 
R8961t6532 n8962 n6533 R=6.580e+01 
R8961t8463 n8962 n8464 R=5.928e+00 
R8961t1911 n8962 n1912 R=3.073e+00 
R8961t3468 n8962 n3469 R=1.688e+01 
R8961t3660 n8962 n3661 R=5.640e+00 
R8962t3463 n8963 n3464 R=6.097e+00 
R8962t6883 n8963 n6884 R=1.888e+01 
R8962t8356 n8963 n8357 R=2.256e+01 
R8962t198 n8963 n199 R=1.290e+01 
R8962t3960 n8963 n3961 R=5.053e+00 
R8962t8638 n8963 n8639 R=1.341e+01 
R8962t4606 n8963 n4607 R=2.167e+01 
R8962t8728 n8963 n8729 R=5.745e+00 
R8962t175 n8963 n176 R=5.851e+01 
R8963t1722 n8964 n1723 R=7.465e+00 
R8963t3321 n8964 n3322 R=2.464e+01 
R8963t4215 n8964 n4216 R=6.358e+00 
R8963t6554 n8964 n6555 R=1.023e+01 
R8963t5048 n8964 n5049 R=1.003e+01 
R8963t3134 n8964 n3135 R=1.831e+01 
R8963t7734 n8964 n7735 R=4.230e+00 
R8964t376 n8965 n377 R=6.734e+00 
R8964t1464 n8965 n1465 R=3.217e+00 
R8964t701 n8965 n702 R=7.113e+01 
R8964t1920 n8965 n1921 R=2.502e+00 
R8964t3789 n8965 n3790 R=1.020e+01 
R8965t2272 n8966 n2273 R=7.158e+00 
R8965t3599 n8966 n3600 R=2.522e+00 
R8965t5014 n8966 n5015 R=8.018e+01 
R8965t1391 n8966 n1392 R=1.023e+01 
R8966t4898 n8967 n4899 R=7.231e+00 
R8966t6240 n8967 n6241 R=2.723e+01 
R8966t84 n8967 n85 R=1.210e+01 
R8966t5959 n8967 n5960 R=1.598e+01 
R8966t5619 n8967 n5620 R=2.024e+02 
R8966t1612 n8967 n1613 R=5.151e+00 
R8966t573 n8967 n574 R=6.518e+00 
R8966t1818 n8967 n1819 R=3.199e+02 
R8967t781 n8968 n782 R=9.040e+00 
R8967t4341 n8968 n4342 R=2.029e+02 
R8967t8050 n8968 n8051 R=6.324e+00 
R8967t5964 n8968 n5965 R=4.327e+00 
R8967t1445 n8968 n1446 R=6.058e+01 
R8967t4021 n8968 n4022 R=4.420e+00 
R8967t402 n8968 n403 R=1.282e+01 
R8968t2137 n8969 n2138 R=1.177e+02 
R8968t8866 n8969 n8867 R=1.139e+01 
R8968t2549 n8969 n2550 R=5.282e+00 
R8968t3005 n8969 n3006 R=1.973e+02 
R8968t8877 n8969 n8878 R=1.158e+01 
R8968t8637 n8969 n8638 R=3.768e+00 
R8969t1723 n8970 n1724 R=5.072e+00 
R8969t6226 n8970 n6227 R=2.341e+00 
R8969t6908 n8970 n6909 R=8.097e+00 
R8970t649 n8971 n650 R=1.789e+01 
R8970t3545 n8971 n3546 R=5.340e+00 
R8970t5848 n8971 n5849 R=3.675e+00 
R8970t1171 n8971 n1172 R=2.585e+00 
R8971t3027 n8972 n3028 R=1.722e+01 
R8971t4085 n8972 n4086 R=2.772e+00 
R8971t2289 n8972 n2290 R=9.558e+00 
R8971t8557 n8972 n8558 R=2.901e+02 
R8971t1126 n8972 n1127 R=6.259e+00 
R8972t461 n8973 n462 R=6.288e+00 
R8972t2918 n8973 n2919 R=4.108e+00 
R8972t2114 n8973 n2115 R=1.069e+01 
R8972t475 n8973 n476 R=5.266e+00 
R8972t3759 n8973 n3760 R=5.991e+01 
R8973t2398 n8974 n2399 R=2.361e+00 
R8973t4700 n8974 n4701 R=1.311e+01 
R8973t6572 n8974 n6573 R=3.044e+00 
R8973t4071 n8974 n4072 R=5.771e+01 
R8973t3380 n8974 n3381 R=1.122e+01 
R8973t8815 n8974 n8816 R=1.509e+01 
R8974t2021 n8975 n2022 R=3.922e+00 
R8974t4840 n8975 n4841 R=5.630e+01 
R8974t6027 n8975 n6028 R=3.381e+00 
R8974t5401 n8975 n5402 R=6.562e+00 
R8975t5424 n8976 n5425 R=1.991e+00 
R8975t6938 n8976 n6939 R=1.994e+02 
R8975t3387 n8976 n3388 R=4.818e+01 
R8975t5461 n8976 n5462 R=2.653e+00 
R8975t2137 n8976 n2138 R=8.134e+00 
R8976t2198 n8977 n1 R=9.323e+00 
R8976t6191 n8977 n6192 R=5.533e+00 
R8976t278 n8977 n1 R=1.161e+01 
R8976t6966 n8977 n1 R=5.906e+00 
R8976t8187 n8977 n8188 R=1.211e+02 
R8976t2095 n8977 n2096 R=3.964e+00 
R8977t1642 n8978 n1643 R=2.046e+00 
R8977t7117 n8978 n7118 R=8.127e+00 
R8977t796 n8978 n797 R=3.362e+00 
R8977t527 n8978 n528 R=3.301e+01 
R8978t1530 n8979 n1531 R=9.481e+00 
R8978t7636 n8979 n7637 R=1.755e+01 
R8978t137 n8979 n138 R=1.064e+03 
R8978t8409 n8979 n8410 R=3.155e+00 
R8978t7257 n8979 n7258 R=1.893e+02 
R8978t2471 n8979 n2472 R=2.579e+00 
R8978t787 n8979 n788 R=1.112e+01 
R8979t7070 n8980 n7071 R=3.978e+01 
R8979t8396 n8980 n8397 R=5.325e+00 
R8979t1998 n8980 n1999 R=6.037e+00 
R8979t6871 n8980 n6872 R=6.763e+00 
R8979t4231 n8980 n4232 R=2.092e+01 
R8979t6111 n8980 n6112 R=1.980e+00 
R8980t722 n8981 n723 R=2.794e+01 
R8980t2305 n8981 n2306 R=6.859e+00 
R8980t4711 n8981 n4712 R=7.470e+00 
R8980t4990 n8981 n4991 R=4.296e+00 
R8980t2756 n8981 n2757 R=1.228e+01 
R8980t4796 n8981 n4797 R=7.555e+00 
R8980t5532 n8981 n5533 R=1.073e+01 
R8981t4339 n8982 n4340 R=5.481e+00 
R8981t7042 n8982 n7043 R=3.157e+00 
R8981t424 n8982 n425 R=2.403e+00 
R8981t6331 n8982 n6332 R=4.829e+01 
R8981t1752 n8982 n1753 R=4.860e+01 
R8982t966 n8983 n967 R=4.641e+00 
R8982t3290 n8983 n3291 R=4.055e+00 
R8982t2746 n8983 n2747 R=1.230e+03 
R8982t3333 n8983 n3334 R=3.194e+00 
R8982t4739 n8983 n4740 R=8.045e+00 
R8983t4413 n8984 n4414 R=2.934e+01 
R8983t6412 n8984 n6413 R=9.846e+01 
R8983t2427 n8984 n2428 R=2.318e+00 
R8983t7299 n8984 n7300 R=7.366e+00 
R8983t9 n8984 n10 R=1.934e+01 
R8983t7786 n8984 n7787 R=2.757e+00 
R8984t554 n8985 n555 R=1.078e+01 
R8984t2426 n8985 n2427 R=2.538e+00 
R8984t8123 n8985 n8124 R=2.929e+01 
R8984t7007 n8985 n7008 R=3.360e+00 
R8984t2822 n8985 n2823 R=9.160e+00 
R8985t7328 n8986 n7329 R=1.820e+01 
R8985t7554 n8986 n7555 R=2.084e+00 
R8985t327 n8986 n328 R=1.621e+00 
R8985t2080 n8986 n2081 R=6.787e+00 
R8986t1148 n8987 n1149 R=5.314e+00 
R8986t7977 n8987 n7978 R=7.237e+00 
R8986t4393 n8987 n4394 R=9.828e+00 
R8986t579 n8987 n580 R=9.523e+00 
R8986t7634 n8987 n7635 R=7.400e+00 
R8987t3395 n8988 n3396 R=1.367e+01 
R8987t6076 n8988 n6077 R=1.164e+02 
R8987t4441 n8988 n4442 R=7.400e+00 
R8987t1351 n8988 n1352 R=1.265e+01 
R8987t8913 n8988 n8914 R=5.524e+01 
R8987t4309 n8988 n4310 R=2.264e+01 
R8987t2115 n8988 n2116 R=4.505e+00 
R8987t5757 n8988 n5758 R=9.496e+00 
R8987t5887 n8988 n5888 R=1.217e+01 
R8988t5136 n8989 n5137 R=2.548e+00 
R8988t8684 n8989 n8685 R=5.904e+00 
R8988t8395 n8989 n8396 R=5.160e+00 
R8988t6288 n8989 n6289 R=1.618e+01 
R8989t1759 n8990 n1760 R=1.265e+01 
R8989t4632 n8990 n4633 R=1.161e+01 
R8989t1654 n8990 n1655 R=2.321e+00 
R8989t4152 n8990 n4153 R=1.950e+01 
R8989t6825 n8990 n6826 R=8.975e+01 
R8989t2375 n8990 n2376 R=2.729e+00 
R8990t5576 n8991 n5577 R=2.621e+01 
R8990t7055 n8991 n7056 R=4.404e+00 
R8990t6730 n8991 n6731 R=1.031e+01 
R8990t8265 n8991 n8266 R=5.862e+00 
R8990t8937 n8991 n8938 R=5.100e+00 
R8991t1440 n8992 n1441 R=9.951e+00 
R8991t3406 n8992 n3407 R=4.510e+00 
R8991t2583 n8992 n2584 R=8.593e+00 
R8991t516 n8992 n517 R=2.349e+01 
R8991t5226 n8992 n5227 R=2.197e+01 
R8991t1013 n8992 n1014 R=7.243e+00 
R8991t5160 n8992 n5161 R=4.220e+02 
R8991t4116 n8992 n4117 R=1.794e+01 
R8992t2782 n8993 n2783 R=3.871e+00 
R8992t7594 n8993 n7595 R=4.555e+00 
R8992t5362 n8993 n5363 R=1.483e+01 
R8992t741 n8993 n742 R=1.460e+00 
R8992t4439 n8993 n4440 R=3.702e+01 
R8993t2672 n8994 n2673 R=2.992e+01 
R8993t5561 n8994 n5562 R=3.874e+00 
R8993t8429 n8994 n8430 R=3.418e+00 
R8993t5131 n8994 n5132 R=3.532e+00 
R8994t4445 n8995 n4446 R=6.286e+00 
R8994t5474 n8995 n5475 R=2.532e+02 
R8994t107 n8995 n108 R=2.836e+01 
R8994t2627 n8995 n2628 R=6.239e+00 
R8994t2090 n8995 n2091 R=8.802e+00 
R8994t7107 n8995 n7108 R=1.736e+01 
R8994t6510 n8995 n6511 R=2.870e+01 
R8994t7999 n8995 n8000 R=7.995e+00 
R8995t4563 n8996 n4564 R=2.300e+00 
R8995t6524 n8996 n6525 R=6.948e+01 
R8995t2077 n8996 n2078 R=2.259e+00 
R8995t3495 n8996 n3496 R=1.676e+01 
R8995t5517 n8996 n5518 R=6.490e+00 
R8996t5748 n8997 n5749 R=1.563e+01 
R8996t508 n8997 n509 R=2.920e+00 
R8997t263 n8998 n264 R=2.300e+01 
R8997t5049 n8998 n5050 R=5.682e+00 
R8997t3212 n8998 n3213 R=6.770e+00 
R8997t7658 n8998 n7659 R=1.305e+01 
R8997t2534 n8998 n2535 R=6.568e+00 
R8997t3589 n8998 n3590 R=9.876e+00 
R8998t6289 n8999 n6290 R=1.567e+01 
R8998t7240 n8999 n7241 R=3.484e+01 
R8998t7080 n8999 n7081 R=5.837e+00 
R8998t4266 n8999 n4267 R=3.252e+00 
R8998t4924 n8999 n4925 R=4.461e+01 
R8998t8725 n8999 n8726 R=1.853e+01 
R8998t6417 n8999 n6418 R=8.940e+00 
R8999t2040 n9000 n2041 R=7.270e+00 
R8999t6203 n9000 n6204 R=4.288e+00 
R8999t2358 n9000 n2359 R=3.307e+00 
R8999t2873 n9000 n2874 R=8.887e+00 
R9000t1003 n9001 n1004 R=2.877e+00 
R9000t5735 n9001 n5736 R=1.774e+01 
R9000t443 n9001 n444 R=2.208e+01 
R9000t49 n9001 n50 R=5.142e+00 
R9000t5667 n9001 n5668 R=6.242e+00 
R9000t2665 n9001 n2666 R=2.907e+01 
R9001t688 n9002 n689 R=2.714e+01 
R9001t4921 n9002 n4922 R=5.513e+00 
R9001t8854 n9002 n8855 R=7.441e+00 
R9001t1114 n9002 n1115 R=4.544e+00 
R9001t3591 n9002 n3592 R=5.632e+01 
R9001t999 n9002 n1000 R=7.145e+00 
R9002t306 n9003 n307 R=1.883e+01 
R9002t2026 n9003 n2027 R=7.621e+00 
R9002t6477 n9003 n6478 R=4.475e+01 
R9002t2979 n9003 n2980 R=2.405e+00 
R9002t1807 n9003 n1808 R=9.881e+00 
R9002t6555 n9003 n6556 R=5.487e+00 
R9003t1540 n9004 n1541 R=5.031e+01 
R9003t5704 n9004 n5705 R=2.160e+00 
R9003t7843 n9004 n7844 R=1.009e+01 
R9003t8568 n9004 n8569 R=1.033e+01 
R9003t450 n9004 n451 R=8.581e+00 
R9003t6216 n9004 n6217 R=7.320e+00 
R9004t2749 n9005 n2750 R=2.538e+00 
R9004t4995 n9005 n4996 R=6.483e+00 
R9004t510 n9005 n511 R=1.227e+01 
R9005t4180 n9006 n4181 R=6.585e+01 
R9005t8618 n9006 n8619 R=4.338e+01 
R9005t4655 n9006 n4656 R=4.684e+00 
R9005t979 n9006 n980 R=4.584e+00 
R9005t860 n9006 n861 R=1.031e+02 
R9005t386 n9006 n387 R=1.061e+02 
R9005t5719 n9006 n5720 R=4.209e+00 
R9005t1953 n9006 n1954 R=4.945e+00 
R9006t622 n9007 n623 R=3.200e+00 
R9006t7478 n9007 n7479 R=2.441e+01 
R9006t8797 n9007 n8798 R=1.450e+01 
R9006t4043 n9007 n4044 R=2.967e+01 
R9006t8012 n9007 n8013 R=5.700e+00 
R9006t4653 n9007 n4654 R=1.220e+01 
R9006t8186 n9007 n8187 R=1.136e+01 
R9006t2349 n9007 n2350 R=3.348e+01 
R9007t1220 n9008 n1221 R=6.191e+00 
R9007t5453 n9008 n5454 R=5.967e+01 
R9007t2080 n9008 n2081 R=3.718e+00 
R9007t7701 n9008 n7702 R=6.256e+00 
R9008t1875 n9009 n1876 R=4.845e+00 
R9008t4597 n9009 n4598 R=2.060e+01 
R9008t2907 n9009 n2908 R=8.063e+01 
R9008t2767 n9009 n2768 R=2.636e+00 
R9008t8187 n9009 n8188 R=8.563e+01 
R9008t5951 n9009 n5952 R=1.392e+01 
R9009t1452 n9010 n1453 R=3.026e+01 
R9009t3629 n9010 n3630 R=6.933e+00 
R9009t196 n9010 n197 R=1.215e+01 
R9009t5849 n9010 n5850 R=7.244e+00 
R9009t1159 n9010 n1160 R=5.722e+00 
R9009t7919 n9010 n7920 R=9.492e+00 
R9010t5074 n9011 n5075 R=3.218e+01 
R9010t6139 n9011 n6140 R=3.286e+00 
R9010t159 n9011 n160 R=8.640e+01 
R9010t601 n9011 n602 R=1.009e+01 
R9010t2564 n9011 n2565 R=2.856e+00 
R9010t6033 n9011 n6034 R=1.495e+01 
R9011t7157 n9012 n7158 R=2.238e+02 
R9011t8011 n9012 n8012 R=5.269e+00 
R9011t1370 n9012 n1371 R=2.037e+01 
R9011t7696 n9012 n7697 R=3.238e+00 
R9011t5896 n9012 n5897 R=5.751e+00 
R9011t5761 n9012 n5762 R=4.941e+00 
R9012t2327 n9013 n2328 R=2.551e+01 
R9012t2495 n9013 n2496 R=8.097e+00 
R9012t7375 n9013 n7376 R=3.765e+00 
R9012t5113 n9013 n5114 R=1.810e+01 
R9012t1582 n9013 n1583 R=1.344e+01 
R9012t3934 n9013 n3935 R=9.892e+01 
R9012t7631 n9013 n7632 R=7.369e+01 
R9012t8748 n9013 n8749 R=5.965e+00 
R9012t3748 n9013 n3749 R=2.530e+01 
R9013t4232 n9014 n4233 R=3.706e+00 
R9013t8225 n9014 n8226 R=3.383e+01 
R9013t7481 n9014 n7482 R=5.337e+00 
R9013t7660 n9014 n7661 R=6.378e+01 
R9013t3883 n9014 n3884 R=5.332e+01 
R9013t7035 n9014 n7036 R=3.775e+00 
R9013t6982 n9014 n6983 R=1.397e+01 
R9013t2213 n9014 n2214 R=2.161e+01 
R9013t8141 n9014 n8142 R=1.482e+02 
R9014t1560 n9015 n1561 R=5.801e+00 
R9014t3072 n9015 n3073 R=1.179e+01 
R9014t4019 n9015 n4020 R=7.980e+00 
R9014t5024 n9015 n5025 R=5.534e+00 
R9015t1447 n9016 n1448 R=1.754e+01 
R9015t6365 n9016 n6366 R=3.075e+00 
R9015t1521 n9016 n1522 R=8.095e+00 
R9015t4146 n9016 n4147 R=6.396e+00 
R9016t13 n9017 n14 R=2.423e+01 
R9016t673 n9017 n674 R=1.744e+01 
R9016t4554 n9017 n4555 R=9.052e+02 
R9016t652 n9017 n653 R=3.188e+00 
R9016t1109 n9017 n1110 R=1.269e+01 
R9017t3672 n9018 n3673 R=1.364e+01 
R9017t6472 n9018 n6473 R=2.414e+01 
R9017t3837 n9018 n3838 R=2.853e+00 
R9017t5110 n9018 n5111 R=1.116e+01 
R9017t6595 n9018 n6596 R=1.019e+01 
R9017t108 n9018 n109 R=4.601e+00 
R9018t1650 n9019 n1651 R=2.676e+01 
R9018t7490 n9019 n7491 R=1.075e+01 
R9018t5490 n9019 n5491 R=2.027e+00 
R9018t4362 n9019 n4363 R=1.467e+02 
R9018t2595 n9019 n2596 R=1.184e+01 
R9018t6002 n9019 n6003 R=2.599e+00 
R9019t1355 n9020 n1356 R=6.511e+00 
R9019t6958 n9020 n6959 R=7.325e+00 
R9019t5308 n9020 n5309 R=5.602e+00 
R9019t2752 n9020 n2753 R=7.005e+01 
R9019t3151 n9020 n3152 R=7.451e+00 
R9019t6060 n9020 n6061 R=7.103e+00 
R9019t4841 n9020 n4842 R=2.628e+01 
R9020t2551 n9021 n2552 R=1.219e+01 
R9020t6545 n9021 n6546 R=3.618e+00 
R9020t6769 n9021 n6770 R=2.502e+00 
R9020t8090 n9021 n8091 R=5.986e+00 
R9020t6813 n9021 n6814 R=1.333e+01 
R9021t1086 n9022 n1087 R=4.826e+00 
R9021t3407 n9022 n3408 R=4.076e+00 
R9021t1254 n9022 n1255 R=1.131e+01 
R9021t7356 n9022 n7357 R=1.046e+01 
R9021t1024 n9022 n1025 R=1.591e+01 
R9022t2393 n9023 n2394 R=6.228e+01 
R9022t8781 n9023 n8782 R=5.820e+00 
R9022t680 n9023 n681 R=1.294e+01 
R9022t3997 n9023 n3998 R=1.340e+01 
R9022t5466 n9023 n5467 R=3.628e+01 
R9022t532 n9023 n533 R=4.960e+00 
R9023t5652 n9024 n5653 R=2.903e+00 
R9023t8073 n9024 n8074 R=4.905e+01 
R9023t2673 n9024 n2674 R=1.967e+01 
R9023t2958 n9024 n2959 R=2.776e+00 
R9023t4740 n9024 n4741 R=1.416e+01 
R9024t335 n9025 n336 R=3.392e+00 
R9024t7564 n9025 n7565 R=3.109e+00 
R9024t1172 n9025 n1173 R=7.884e+00 
R9024t4165 n9025 n4166 R=8.548e+00 
R9025t1765 n9026 n1766 R=2.858e+01 
R9025t2167 n9026 n2168 R=5.932e+00 
R9025t2450 n9026 n2451 R=4.056e+00 
R9025t824 n9026 n825 R=1.303e+01 
R9025t1601 n9026 n1602 R=2.680e+01 
R9025t4008 n9026 n4009 R=3.617e+01 
R9026t716 n9027 n717 R=4.468e+01 
R9026t7387 n9027 n7388 R=7.220e+00 
R9026t994 n9027 n995 R=1.679e+02 
R9026t2983 n9027 n2984 R=2.821e+00 
R9026t1194 n9027 n1195 R=1.466e+01 
R9026t1525 n9027 n1526 R=2.940e+00 
R9027t2272 n9028 n2273 R=5.136e+00 
R9027t7303 n9028 n7304 R=2.198e+02 
R9027t1442 n9028 n1443 R=4.709e+00 
R9028t1876 n9029 n1877 R=2.730e+02 
R9028t6519 n9029 n6520 R=6.261e+00 
R9028t2855 n9029 n2856 R=9.594e+00 
R9028t7681 n9029 n7682 R=3.213e+00 
R9028t1038 n9029 n1039 R=1.263e+01 
R9029t1905 n9030 n1906 R=5.452e+02 
R9029t4551 n9030 n4552 R=2.266e+00 
R9029t2166 n9030 n2167 R=5.958e+01 
R9029t5697 n9030 n5698 R=3.695e+00 
R9029t2058 n9030 n2059 R=1.813e+01 
R9030t5510 n9031 n5511 R=9.570e+00 
R9030t5784 n9031 n5785 R=4.707e+01 
R9030t368 n9031 n369 R=4.392e+00 
R9030t2325 n9031 n2326 R=8.856e+00 
R9030t2934 n9031 n2935 R=1.299e+01 
R9030t134 n9031 n135 R=7.198e+00 
R9030t8355 n9031 n8356 R=9.220e+01 
R9031t1778 n9032 n1779 R=1.581e+02 
R9031t8297 n9032 n8298 R=6.320e+00 
R9031t2493 n9032 n2494 R=5.042e+00 
R9031t140 n9032 n141 R=9.460e+01 
R9031t3986 n9032 n3987 R=5.584e+00 
R9031t4545 n9032 n4546 R=5.456e+01 
R9031t3173 n9032 n3174 R=2.545e+01 
R9031t7410 n9032 n7411 R=3.802e+00 
R9032t7139 n9033 n7140 R=1.048e+01 
R9032t8082 n9033 n8083 R=7.650e+00 
R9032t8334 n9033 n8335 R=1.962e+01 
R9032t3297 n9033 n3298 R=8.531e+00 
R9032t4351 n9033 n4352 R=9.386e+00 
R9032t1075 n9033 n1076 R=1.424e+01 
R9032t1066 n9033 n1067 R=4.012e+01 
R9032t1845 n9033 n1846 R=7.069e+00 
R9032t1496 n9033 n1497 R=5.287e+01 
R9033t3084 n9034 n3085 R=2.782e+00 
R9033t8767 n9034 n8768 R=1.462e+01 
R9033t2073 n9034 n2074 R=1.030e+01 
R9033t7936 n9034 n7937 R=1.314e+01 
R9033t3668 n9034 n3669 R=1.872e+01 
R9033t2946 n9034 n2947 R=7.844e+00 
R9033t2829 n9034 n2830 R=1.663e+01 
R9033t4671 n9034 n4672 R=2.350e+01 
R9034t6911 n9035 n6912 R=9.590e+00 
R9034t37 n9035 n38 R=1.901e+01 
R9034t6699 n9035 n6700 R=1.923e+00 
R9034t4287 n9035 n4288 R=7.571e+00 
R9034t1250 n9035 n1251 R=5.345e+00 
R9035t8178 n9036 n8179 R=6.719e+00 
R9035t7683 n9036 n7684 R=6.100e+00 
R9035t6424 n9036 n6425 R=2.893e+00 
R9035t3550 n9036 n3551 R=1.101e+01 
R9036t2926 n9037 n2927 R=3.268e+01 
R9036t7343 n9037 n7344 R=4.821e+00 
R9036t5401 n9037 n5402 R=1.867e+01 
R9036t2303 n9037 n2304 R=6.583e+01 
R9036t3444 n9037 n3445 R=2.018e+01 
R9036t6132 n9037 n6133 R=2.362e+01 
R9036t6495 n9037 n6496 R=3.424e+00 
R9037t1994 n9038 n1995 R=1.260e+01 
R9037t4455 n9038 n4456 R=1.556e+01 
R9037t7402 n9038 n7403 R=1.657e+01 
R9037t6640 n9038 n6641 R=1.976e+01 
R9037t4201 n9038 n4202 R=2.732e+00 
R9037t4916 n9038 n4917 R=3.390e+00 
R9038t4033 n9039 n4034 R=2.291e+00 
R9038t8175 n9039 n8176 R=6.214e+01 
R9038t8640 n9039 n8641 R=1.177e+01 
R9038t8922 n9039 n8923 R=3.735e+00 
R9038t514 n9039 n515 R=3.575e+01 
R9038t6850 n9039 n6851 R=7.738e+01 
R9038t3665 n9039 n3666 R=9.990e+00 
R9039t4423 n9040 n4424 R=7.504e+00 
R9039t5614 n9040 n5615 R=9.942e+00 
R9039t2567 n9040 n2568 R=7.302e+00 
R9039t444 n9040 n445 R=5.008e+00 
R9039t4812 n9040 n4813 R=3.616e+00 
R9039t1083 n9040 n1084 R=6.791e+01 
R9040t3132 n9041 n3133 R=1.060e+02 
R9040t6202 n9041 n6203 R=2.028e+00 
R9040t5349 n9041 n5350 R=1.192e+01 
R9040t7958 n9041 n7959 R=2.129e+00 
R9040t38 n9041 n39 R=2.500e+01 
R9040t8706 n9041 n8707 R=5.128e+01 
R9041t5441 n9042 n5442 R=1.774e+00 
R9041t6204 n9042 n6205 R=1.378e+04 
R9042t230 n9043 n231 R=3.995e+01 
R9042t1415 n9043 n1416 R=4.245e+00 
R9042t1421 n9043 n1422 R=6.534e+01 
R9042t2840 n9043 n2841 R=3.588e+00 
R9042t2947 n9043 n2948 R=9.352e+00 
R9042t5000 n9043 n5001 R=1.121e+01 
R9043t2574 n9044 n2575 R=1.218e+01 
R9043t8548 n9044 n8549 R=3.852e+00 
R9043t4089 n9044 n4090 R=8.353e+00 
R9043t7616 n9044 n7617 R=3.050e+00 
R9043t4689 n9044 n4690 R=4.032e+01 
R9044t6154 n9045 n6155 R=1.531e+01 
R9044t6984 n9045 n6985 R=1.209e+01 
R9044t703 n9045 n704 R=1.338e+01 
R9044t1857 n9045 n1858 R=9.746e+00 
R9044t6853 n9045 n6854 R=6.098e+00 
R9044t4045 n9045 n4046 R=1.409e+01 
R9045t3331 n9046 n3332 R=8.466e+00 
R9045t4821 n9046 n4822 R=1.547e+01 
R9045t3867 n9046 n3868 R=7.058e+01 
R9045t8239 n9046 n8240 R=4.985e+00 
R9045t7798 n9046 n7799 R=1.696e+01 
R9045t5344 n9046 n5345 R=7.463e+00 
R9045t6560 n9046 n6561 R=4.585e+00 
R9046t3751 n9047 n3752 R=5.294e+00 
R9046t7713 n9047 n7714 R=2.698e+00 
R9046t949 n9047 n950 R=1.202e+01 
R9046t8032 n9047 n8033 R=2.645e+01 
R9046t7441 n9047 n7442 R=4.413e+00 
R9047t3493 n9048 n3494 R=3.001e+00 
R9047t4004 n9048 n4005 R=3.741e+00 
R9047t4963 n9048 n4964 R=3.805e+00 
R9048t6374 n9049 n6375 R=6.962e+00 
R9048t8894 n9049 n8895 R=6.694e+00 
R9048t2412 n9049 n2413 R=5.910e+00 
R9048t5786 n9049 n5787 R=5.950e+00 
R9049t663 n9050 n664 R=1.696e+01 
R9049t3201 n9050 n3202 R=2.978e+00 
R9049t6190 n9050 n6191 R=1.137e+01 
R9049t8826 n9050 n8827 R=6.665e+00 
R9049t6388 n9050 n6389 R=1.393e+01 
R9049t1135 n9050 n1136 R=2.762e+01 
R9050t6723 n9051 n6724 R=1.336e+01 
R9050t6768 n9051 n6769 R=6.308e+00 
R9050t4414 n9051 n4415 R=1.283e+01 
R9050t6706 n9051 n6707 R=5.971e+00 
R9050t8900 n9051 n8901 R=8.203e+01 
R9050t1784 n9051 n1785 R=2.970e+00 
R9051t2318 n9052 n2319 R=5.825e+00 
R9051t8959 n9052 n8960 R=4.189e+00 
R9051t1245 n9052 n1246 R=2.561e+01 
R9051t3857 n9052 n3858 R=2.791e+00 
R9051t6788 n9052 n6789 R=2.831e+01 
R9052t206 n9053 n207 R=8.179e+00 
R9052t8881 n9053 n8882 R=6.444e+00 
R9052t2489 n9053 n2490 R=4.590e+00 
R9052t102 n9053 n103 R=1.044e+01 
R9052t5108 n9053 n5109 R=1.274e+01 
R9052t842 n9053 n843 R=2.459e+01 
R9053t590 n9054 n591 R=2.891e+01 
R9053t4822 n9054 n4823 R=1.609e+02 
R9053t7126 n9054 n7127 R=2.712e+00 
R9053t6925 n9054 n6926 R=4.251e+00 
R9053t1358 n9054 n1359 R=1.337e+01 
R9053t4661 n9054 n4662 R=3.280e+00 
R9054t3230 n9055 n3231 R=5.249e+00 
R9054t6451 n9055 n6452 R=1.772e+01 
R9054t6909 n9055 n6910 R=8.472e+00 
R9054t6558 n9055 n6559 R=4.911e+00 
R9054t1440 n9055 n1441 R=4.266e+00 
R9055t1366 n9056 n1367 R=3.144e+00 
R9055t5436 n9056 n5437 R=2.231e+01 
R9055t5245 n9056 n5246 R=1.789e+01 
R9055t2164 n9056 n2165 R=6.214e+00 
R9055t1181 n9056 n1182 R=6.871e+00 
R9055t3235 n9056 n3236 R=5.536e+00 
R9056t257 n9057 n258 R=1.748e+01 
R9056t6468 n9057 n6469 R=2.941e+01 
R9056t1949 n9057 n1950 R=3.017e+01 
R9056t3006 n9057 n3007 R=5.879e+00 
R9056t8230 n9057 n8231 R=8.203e+00 
R9056t761 n9057 n762 R=5.422e+00 
R9057t1063 n9058 n1064 R=3.192e+01 
R9057t4356 n9058 n4357 R=4.614e+00 
R9057t7095 n9058 n7096 R=3.220e+00 
R9057t8372 n9058 n8373 R=2.649e+01 
R9057t7152 n9058 n7153 R=1.565e+01 
R9058t8393 n9059 n8394 R=1.339e+01 
R9058t8510 n9059 n8511 R=6.332e+00 
R9058t5419 n9059 n5420 R=5.336e+00 
R9058t2857 n9059 n2858 R=1.230e+01 
R9058t4491 n9059 n4492 R=6.601e+00 
R9058t1809 n9059 n1810 R=1.789e+01 
R9058t3688 n9059 n3689 R=3.054e+01 
R9059t714 n9060 n715 R=7.983e+00 
R9059t3756 n9060 n3757 R=6.170e+00 
R9059t2515 n9060 n2516 R=1.890e+01 
R9059t8384 n9060 n8385 R=6.083e+00 
R9059t4506 n9060 n4507 R=1.586e+02 
R9059t7496 n9060 n7497 R=1.946e+01 
R9059t1308 n9060 n1309 R=2.499e+01 
R9059t731 n9060 n732 R=1.025e+01 
R9060t701 n9061 n702 R=1.555e+02 
R9060t2739 n9061 n2740 R=2.161e+00 
R9060t3831 n9061 n3832 R=5.824e+00 
R9061t743 n9062 n744 R=1.758e+01 
R9061t8834 n9062 n8835 R=4.272e+00 
R9061t666 n9062 n667 R=3.897e+00 
R9061t6677 n9062 n6678 R=3.411e+00 
R9061t7959 n9062 n7960 R=7.341e+01 
R9062t8173 n9063 n8174 R=7.891e+01 
R9062t8837 n9063 n8838 R=7.156e+00 
R9062t4051 n9063 n4052 R=8.232e+00 
R9062t3049 n9063 n3050 R=7.411e+00 
R9062t5551 n9063 n5552 R=8.032e+00 
R9062t4508 n9063 n4509 R=1.199e+02 
R9062t615 n9063 n616 R=3.557e+00 
R9063t6110 n9064 n6111 R=4.028e+00 
R9063t4205 n9064 n4206 R=1.013e+01 
R9063t4470 n9064 n4471 R=7.517e+00 
R9063t8661 n9064 n8662 R=5.751e+00 
R9063t6780 n9064 n6781 R=6.732e+01 
R9063t4911 n9064 n4912 R=7.085e+00 
R9064t5979 n9065 n5980 R=1.965e+01 
R9064t6350 n9065 n6351 R=7.976e+00 
R9064t3679 n9065 n3680 R=1.106e+01 
R9064t7469 n9065 n7470 R=1.301e+01 
R9064t2238 n9065 n2239 R=1.343e+01 
R9064t6625 n9065 n6626 R=4.677e+00 
R9064t1423 n9065 n1424 R=6.471e+01 
R9064t7093 n9065 n7094 R=4.793e+00 
R9065t1363 n9066 n1364 R=5.765e+00 
R9065t7947 n9066 n7948 R=7.424e+00 
R9065t8614 n9066 n8615 R=6.720e+00 
R9065t4819 n9066 n4820 R=3.058e+00 
R9066t5805 n9067 n5806 R=3.857e+00 
R9066t6600 n9067 n6601 R=1.164e+01 
R9066t1619 n9067 n1620 R=3.572e+00 
R9066t4150 n9067 n4151 R=4.335e+00 
R9067t2242 n9068 n2243 R=1.339e+01 
R9067t8761 n9068 n8762 R=3.563e+00 
R9067t6017 n9068 n6018 R=1.221e+01 
R9067t3774 n9068 n3775 R=6.904e+00 
R9067t7091 n9068 n7092 R=4.375e+00 
R9068t3674 n9069 n3675 R=9.744e+00 
R9068t4220 n9069 n4221 R=3.951e+00 
R9068t6797 n9069 n6798 R=1.607e+01 
R9068t5289 n9069 n5290 R=4.679e+00 
R9068t1337 n9069 n1338 R=8.106e+00 
R9069t2182 n9070 n2183 R=4.018e+00 
R9069t8144 n9070 n8145 R=3.748e+00 
R9069t4835 n9070 n4836 R=3.902e+01 
R9069t6470 n9070 n6471 R=3.787e+00 
R9069t3542 n9070 n3543 R=1.365e+01 
R9069t2123 n9070 n2124 R=9.058e+01 
R9069t2584 n9070 n2585 R=1.336e+02 
R9070t3652 n9071 n3653 R=8.589e+00 
R9070t8649 n9071 n8650 R=8.769e+00 
R9070t7452 n9071 n7453 R=4.588e+00 
R9070t1305 n9071 n1306 R=1.365e+01 
R9070t7694 n9071 n7695 R=9.944e+00 
R9070t1569 n9071 n1570 R=3.319e+01 
R9070t837 n9071 n838 R=1.289e+01 
R9071t3604 n9072 n3605 R=5.751e+00 
R9071t6110 n9072 n6111 R=4.052e+00 
R9071t8556 n9072 n8557 R=7.407e+00 
R9071t4205 n9072 n4206 R=1.626e+01 
R9071t9063 n9072 n9064 R=4.138e+01 
R9072t885 n9073 n886 R=2.533e+01 
R9072t5389 n9073 n5390 R=1.391e+01 
R9072t3096 n9073 n3097 R=2.761e+00 
R9072t6063 n9073 n6064 R=3.373e+01 
R9072t3324 n9073 n3325 R=3.663e+00 
R9072t7862 n9073 n7863 R=1.253e+01 
R9073t2563 n9074 n2564 R=6.003e+00 
R9073t5382 n9074 n5383 R=6.554e+00 
R9073t8349 n9074 n8350 R=1.025e+02 
R9073t7815 n9074 n7816 R=4.368e+00 
R9073t5777 n9074 n5778 R=1.699e+01 
R9073t1656 n9074 n1657 R=7.090e+00 
R9074t5789 n9075 n5790 R=6.624e+01 
R9074t6384 n9075 n6385 R=5.330e+00 
R9074t2196 n9075 n2197 R=4.293e+00 
R9074t6789 n9075 n6790 R=6.100e+00 
R9074t4769 n9075 n4770 R=4.092e+01 
R9075t7039 n9076 n7040 R=2.071e+01 
R9075t7757 n9076 n7758 R=1.977e+01 
R9075t7050 n9076 n7051 R=2.885e+00 
R9075t5870 n9076 n5871 R=7.576e+00 
R9076t5699 n9077 n5700 R=8.800e+01 
R9076t8477 n9077 n8478 R=4.779e+00 
R9076t3224 n9077 n3225 R=5.102e+00 
R9076t1144 n9077 n1145 R=4.123e+00 
R9076t6742 n9077 n6743 R=5.280e+00 
R9077t1693 n9078 n1694 R=3.626e+01 
R9077t8591 n9078 n8592 R=2.152e+00 
R9077t3499 n9078 n3500 R=2.552e+00 
R9077t8169 n9078 n8170 R=3.370e+01 
R9077t1802 n9078 n1803 R=8.636e+00 
R9078t384 n9079 n385 R=4.897e+00 
R9078t2330 n9079 n2331 R=4.179e+00 
R9078t8629 n9079 n8630 R=2.724e+00 
R9079t2758 n9080 n2759 R=4.816e+00 
R9079t7867 n9080 n7868 R=8.086e+01 
R9079t4409 n9080 n4410 R=4.026e+00 
R9079t7704 n9080 n7705 R=7.425e+01 
R9079t2925 n9080 n2926 R=1.065e+01 
R9079t2304 n9080 n2305 R=2.642e+00 
R9080t1552 n9081 n1553 R=7.534e+00 
R9080t5345 n9081 n5346 R=8.813e+00 
R9080t3325 n9081 n3326 R=8.389e+00 
R9080t5291 n9081 n5292 R=1.701e+01 
R9080t3847 n9081 n3848 R=7.369e+00 
R9080t4890 n9081 n4891 R=5.671e+01 
R9080t8357 n9081 n8358 R=1.012e+01 
R9081t5435 n1 n5436 R=2.855e+00 
R9081t7361 n1 n7362 R=2.776e+01 
R9081t6691 n1 n6692 R=1.760e+01 
R9081t5393 n1 n5394 R=1.454e+01 
R9082t2215 n9083 n2216 R=4.762e+00 
R9082t5413 n9083 n5414 R=3.585e+00 
R9082t1756 n9083 n1757 R=1.550e+00 
R9082t6688 n9083 n6689 R=3.645e+01 
R9082t7723 n9083 n7724 R=1.056e+02 
R9083t8109 n9084 n8110 R=5.063e+01 
R9083t7766 n9084 n7767 R=3.417e+00 
R9083t7244 n9084 n7245 R=4.088e+01 
R9083t5301 n9084 n5302 R=3.775e+00 
R9084t272 n9085 n273 R=2.435e+01 
R9084t5586 n9085 n5587 R=3.618e+00 
R9084t584 n9085 n585 R=8.959e+00 
R9084t8685 n9085 n8686 R=6.146e+00 
R9084t3757 n9085 n3758 R=2.367e+01 
R9084t787 n9085 n788 R=1.245e+01 
R9084t7851 n9085 n7852 R=2.235e+01 
R9085t209 n9086 n210 R=5.978e+00 
R9085t7614 n9086 n7615 R=7.318e+00 
R9085t6749 n9086 n6750 R=7.953e+00 
R9085t2432 n9086 n2433 R=7.674e+00 
R9085t6885 n9086 n6886 R=1.115e+01 
R9086t1303 n9087 n1304 R=2.047e+01 
R9086t4562 n9087 n4563 R=6.980e+00 
R9086t5771 n9087 n5772 R=4.062e+00 
R9086t2219 n9087 n2220 R=1.758e+01 
R9086t8296 n9087 n8297 R=1.218e+00 
R9087t6473 n9088 n6474 R=3.001e+00 
R9087t7051 n9088 n7052 R=1.277e+01 
R9087t6426 n9088 n6427 R=6.222e+00 
R9087t4342 n9088 n4343 R=4.074e+00 
R9087t7059 n9088 n7060 R=9.673e+00 
R9087t864 n9088 n865 R=3.279e+01 
R9088t3115 n9089 n3116 R=1.334e+01 
R9088t5946 n9089 n5947 R=3.896e+00 
R9088t5970 n9089 n5971 R=1.267e+03 
R9088t3192 n9089 n3193 R=4.583e+01 
R9088t8839 n9089 n8840 R=2.819e+00 
R9088t66 n9089 n67 R=8.295e+00 
R9089t1695 n9090 n1696 R=1.466e+01 
R9089t6241 n9090 n6242 R=7.279e+00 
R9089t4072 n9090 n4073 R=2.327e+00 
R9089t1041 n9090 n1042 R=6.651e+01 
R9089t5366 n9090 n5367 R=3.382e+00 
R9090t2388 n9091 n2389 R=9.250e+00 
R9090t6149 n9091 n6150 R=4.553e+00 
R9090t6472 n9091 n6473 R=3.922e+00 
R9090t3837 n9091 n3838 R=6.161e+00 
R9090t818 n9091 n819 R=4.001e+01 
R9091t3320 n9092 n3321 R=8.427e+00 
R9091t7041 n9092 n7042 R=5.209e+00 
R9091t3622 n9092 n3623 R=3.367e+00 
R9091t6689 n9092 n6690 R=8.814e+00 
R9092t1653 n9093 n1654 R=1.113e+01 
R9092t6142 n9093 n6143 R=5.292e+00 
R9092t7110 n9093 n7111 R=6.728e+00 
R9092t2537 n9093 n2538 R=7.156e+00 
R9092t3991 n9093 n3992 R=6.050e+00 
R9093t217 n9094 n218 R=2.366e+00 
R9093t2263 n9094 n2264 R=6.523e+00 
R9093t1634 n9094 n1635 R=1.510e+02 
R9093t7381 n9094 n7382 R=3.090e+01 
R9093t8720 n9094 n8721 R=1.053e+01 
R9093t1543 n9094 n1544 R=2.028e+01 
R9093t2401 n9094 n2402 R=3.811e+01 
R9093t6098 n9094 n6099 R=2.362e+02 
R9094t779 n9095 n780 R=1.953e+01 
R9094t4217 n9095 n4218 R=1.085e+01 
R9094t8702 n9095 n8703 R=4.982e+00 
R9094t1792 n9095 n1793 R=2.808e+00 
R9095t3821 n9096 n3822 R=6.384e+01 
R9095t4308 n9096 n4309 R=2.330e+00 
R9095t4396 n9096 n4397 R=6.184e+00 
R9095t8264 n9096 n8265 R=6.354e+01 
R9095t6782 n9096 n6783 R=9.003e+02 
R9095t7768 n9096 n7769 R=3.297e+01 
R9095t6957 n9096 n6958 R=1.502e+00 
R9095t5655 n9096 n5656 R=1.624e+01 
R9096t1686 n9097 n1687 R=5.138e+00 
R9096t3392 n9097 n3393 R=8.819e+00 
R9096t5989 n9097 n5990 R=3.273e+01 
R9096t2031 n9097 n2032 R=6.853e+00 
R9096t4211 n9097 n4212 R=2.588e+02 
R9096t7916 n9097 n7917 R=4.076e+00 
R9096t4513 n9097 n4514 R=1.062e+02 
R9096t7800 n9097 n7801 R=1.676e+01 
R9097t7624 n9098 n7625 R=6.609e+00 
R9097t8146 n9098 n8147 R=3.087e+00 
R9097t440 n9098 n441 R=5.975e+00 
R9097t7873 n9098 n7874 R=3.503e+00 
R9098t2876 n9099 n2877 R=5.538e+01 
R9098t6682 n9099 n6683 R=2.970e+01 
R9098t7639 n9099 n7640 R=1.700e+00 
R9098t5243 n9099 n1 R=2.979e+01 
R9098t7197 n9099 n7198 R=3.641e+00 
R9098t7799 n9099 n7800 R=6.073e+00 
R9099t2761 n9100 n2762 R=4.689e+00 
R9099t4450 n9100 n4451 R=1.369e+01 
R9099t8275 n9100 n8276 R=1.661e+01 
R9099t7290 n9100 n7291 R=5.237e+00 
R9099t1312 n9100 n1313 R=3.254e+02 
R9099t220 n9100 n221 R=1.960e+01 
R9100t4061 n9101 n4062 R=5.187e+00 
R9100t6952 n9101 n6953 R=8.847e+00 
R9100t7768 n9101 n7769 R=9.612e+00 
R9100t4401 n9101 n4402 R=6.058e+00 
R9100t4021 n9101 n4022 R=4.879e+00 
R9101t8036 n9102 n8037 R=2.795e+00 
R9101t1047 n9102 n1048 R=4.509e+01 
R9101t3341 n9102 n3342 R=1.612e+00 
R9102t5736 n9103 n5737 R=5.622e+00 
R9102t7653 n9103 n7654 R=4.149e+00 
R9102t7685 n9103 n7686 R=9.636e+01 
R9102t8875 n9103 n8876 R=1.922e+00 
R9102t5082 n9103 n5083 R=3.686e+01 
R9102t3320 n9103 n3321 R=1.752e+01 
R9103t568 n9104 n569 R=7.058e+00 
R9103t3060 n9104 n3061 R=1.593e+01 
R9103t3616 n9104 n3617 R=3.023e+00 
R9103t7907 n9104 n7908 R=1.281e+01 
R9103t8059 n9104 n8060 R=1.256e+01 
R9104t1475 n9105 n1476 R=1.215e+01 
R9104t8789 n9105 n8790 R=4.878e+00 
R9104t8857 n9105 n8858 R=1.550e+02 
R9104t3793 n9105 n3794 R=2.361e+00 
R9104t1909 n9105 n1910 R=5.932e+01 
R9104t2892 n9105 n2893 R=2.257e+01 
R9104t3277 n9105 n3278 R=8.908e+00 
R9104t3481 n9105 n3482 R=1.853e+01 
R9105t2361 n9106 n2362 R=1.031e+03 
R9105t8960 n9106 n8961 R=5.294e+00 
R9105t3133 n9106 n3134 R=4.437e+00 
R9105t8652 n9106 n8653 R=5.821e+00 
R9105t6073 n9106 n6074 R=4.582e+01 
R9105t4799 n9106 n4800 R=3.335e+00 
R9105t8659 n9106 n8660 R=5.988e+02 
R9106t4003 n9107 n4004 R=1.952e+01 
R9106t4167 n9107 n4168 R=6.083e+00 
R9106t756 n9107 n757 R=1.532e+01 
R9106t384 n9107 n385 R=3.008e+00 
R9106t9078 n9107 n9079 R=9.276e+01 
R9106t2330 n9107 n2331 R=1.879e+01 
R9106t5166 n9107 n5167 R=6.659e+00 
R9106t8153 n9107 n8154 R=2.391e+01 
R9107t3441 n9108 n3442 R=2.061e+00 
R9107t6805 n9108 n6806 R=2.139e+01 
R9107t4278 n9108 n4279 R=8.182e+00 
R9107t8656 n9108 n8657 R=3.522e+00 
R9107t2630 n9108 n2631 R=1.335e+01 
R9108t3580 n9109 n3581 R=9.399e+01 
R9108t7490 n9109 n7491 R=4.738e+00 
R9108t1252 n9109 n1253 R=1.768e+00 
R9108t5370 n9109 n5371 R=5.780e+01 
R9108t2595 n9109 n2596 R=3.503e+01 
R9108t6002 n9109 n6003 R=2.244e+00 
R9109t375 n9110 n376 R=3.373e+00 
R9109t6133 n9110 n6134 R=1.232e+01 
R9109t6803 n9110 n6804 R=4.736e+02 
R9109t1055 n9110 n1056 R=2.618e+00 
R9109t7399 n9110 n7400 R=6.493e+00 
R9110t1058 n9111 n1059 R=2.718e+00 
R9110t8301 n9111 n8302 R=2.817e+01 
R9110t1329 n9111 n1330 R=7.283e+00 
R9110t6992 n9111 n6993 R=4.133e+00 
R9110t5050 n9111 n5051 R=6.629e+00 
R9111t308 n9112 n309 R=2.072e+00 
R9111t5922 n9112 n5923 R=1.033e+01 
R9111t8023 n9112 n8024 R=1.355e+01 
R9111t165 n9112 n166 R=1.647e+00 
R9112t3257 n9113 n3258 R=4.271e+00 
R9112t6891 n9113 n6892 R=1.148e+01 
R9112t1103 n9113 n1104 R=2.809e+00 
R9112t7491 n9113 n7492 R=1.332e+01 
R9112t1152 n9113 n1153 R=4.429e+00 
R9113t1796 n9114 n1797 R=3.028e+00 
R9113t3726 n9114 n3727 R=1.292e+01 
R9113t7779 n9114 n7780 R=5.945e+00 
R9113t6014 n9114 n6015 R=1.141e+01 
R9113t2639 n9114 n2640 R=6.588e+00 
R9113t6496 n9114 n6497 R=4.269e+01 
R9114t4742 n9115 n4743 R=6.555e+00 
R9114t7837 n9115 n7838 R=5.546e+00 
R9114t5351 n9115 n5352 R=1.320e+01 
R9114t6474 n9115 n6475 R=4.993e+00 
R9114t6075 n9115 n6076 R=2.642e+02 
R9114t479 n9115 n480 R=4.410e+00 
R9115t1302 n9116 n1303 R=2.587e+00 
R9115t2405 n9116 n2406 R=6.462e+00 
R9115t2836 n9116 n2837 R=6.635e+01 
R9115t3791 n9116 n3792 R=3.259e+00 
R9115t3131 n9116 n3132 R=1.588e+01 
R9116t3391 n9117 n3392 R=6.386e+01 
R9116t4374 n9117 n4375 R=8.941e+00 
R9116t5773 n9117 n5774 R=6.073e+00 
R9116t8368 n9117 n8369 R=7.021e+00 
R9117t3159 n9118 n3160 R=3.411e+00 
R9117t5510 n9118 n5511 R=6.913e+02 
R9117t8193 n9118 n8194 R=9.785e+00 
R9117t4058 n9118 n4059 R=1.799e+01 
R9117t2390 n9118 n2391 R=7.344e+02 
R9117t3047 n9118 n3048 R=4.878e+00 
R9117t4164 n9118 n4165 R=6.007e+00 
R9117t8492 n9118 n8493 R=3.110e+01 
R9117t5784 n9118 n5785 R=5.796e+01 
R9118t2043 n9119 n2044 R=1.974e+01 
R9118t4009 n9119 n4010 R=8.931e+00 
R9118t1270 n9119 n1271 R=3.502e+00 
R9118t4798 n9119 n4799 R=1.655e+01 
R9118t902 n9119 n903 R=1.048e+01 
R9118t6257 n9119 n6258 R=8.139e+00 
R9119t1375 n9120 n1376 R=1.526e+01 
R9119t6656 n9120 n6657 R=3.357e+01 
R9119t7238 n9120 n7239 R=1.899e+01 
R9119t5939 n9120 n5940 R=7.570e+00 
R9119t5868 n9120 n5869 R=6.760e+00 
R9120t6374 n9121 n6375 R=6.823e+00 
R9120t9048 n9121 n9049 R=6.149e+00 
R9120t7919 n9121 n7920 R=2.266e+01 
R9120t3629 n9121 n3630 R=4.943e+01 
R9120t8636 n9121 n8637 R=3.845e+00 
R9120t5299 n9121 n5300 R=2.442e+01 
R9120t8894 n9121 n8895 R=3.143e+01 
R9121t1470 n9122 n1471 R=6.609e+00 
R9121t5158 n9122 n5159 R=1.255e+01 
R9121t6198 n9122 n6199 R=1.031e+01 
R9121t16 n9122 n17 R=2.342e+01 
R9121t3371 n9122 n3372 R=4.185e+00 
R9122t4449 n9123 n4450 R=4.224e+01 
R9122t7252 n9123 n7253 R=1.202e+01 
R9122t3681 n9123 n3682 R=5.177e+00 
R9122t1110 n9123 n1111 R=4.349e+00 
R9122t4082 n9123 n4083 R=2.173e+01 
R9122t4355 n9123 n4356 R=4.786e+00 
R9123t360 n9124 n361 R=1.382e+01 
R9123t3164 n9124 n3165 R=6.116e+00 
R9123t7785 n9124 n7786 R=1.316e+01 
R9123t6567 n9124 n6568 R=3.463e+00 
R9123t2529 n9124 n2530 R=2.644e+01 
R9123t2681 n9124 n2682 R=5.451e+00 
R9124t230 n9125 n231 R=6.005e+00 
R9124t3153 n9125 n3154 R=7.786e+00 
R9124t204 n9125 n205 R=9.419e+00 
R9124t3519 n9125 n3520 R=3.966e+00 
R9124t1415 n9125 n1416 R=2.462e+01 
R9125t4255 n9126 n4256 R=9.607e+00 
R9125t5279 n9126 n5280 R=7.095e+00 
R9125t2189 n9126 n2190 R=9.441e+00 
R9125t2072 n9126 n2073 R=7.416e+00 
R9125t6369 n9126 n6370 R=6.980e+00 
R9125t8726 n9126 n8727 R=1.383e+01 
R9126t3380 n9127 n3381 R=2.169e+02 
R9126t6170 n9127 n6171 R=4.139e+01 
R9126t7003 n9127 n7004 R=6.767e+01 
R9126t7571 n9127 n7572 R=8.443e+00 
R9126t4905 n9127 n4906 R=7.930e+00 
R9126t2536 n9127 n2537 R=4.395e+00 
R9126t7000 n9127 n7001 R=2.632e+01 
R9126t253 n9127 n254 R=1.387e+01 
R9126t1410 n9127 n1411 R=1.912e+00 
R9127t5016 n9128 n5017 R=4.886e+00 
R9127t8633 n9128 n8634 R=1.231e+01 
R9127t4365 n9128 n4366 R=4.564e+00 
R9127t3882 n9128 n3883 R=1.011e+01 
R9127t2833 n9128 n2834 R=8.794e+00 
R9127t930 n9128 n931 R=1.471e+01 
R9128t2351 n9129 n2352 R=3.165e+01 
R9128t7293 n9129 n7294 R=7.217e+01 
R9128t3657 n9129 n3658 R=3.377e+00 
R9128t6348 n9129 n6349 R=8.501e+02 
R9128t1887 n9129 n1888 R=3.316e+00 
R9129t1269 n9130 n1270 R=4.208e+01 
R9129t8909 n9130 n8910 R=1.508e+01 
R9129t3460 n9130 n3461 R=1.011e+01 
R9129t6988 n9130 n6989 R=4.193e+00 
R9129t2068 n9130 n2069 R=7.886e+00 
R9129t7981 n9130 n7982 R=1.259e+01 
R9129t8892 n9130 n8893 R=1.076e+01 
R9130t6108 n9131 n6109 R=1.641e+00 
R9130t7195 n9131 n7196 R=4.165e+00 
R9130t3666 n9131 n3667 R=1.660e+01 
R9130t3496 n9131 n3497 R=3.606e+00 
R9131t554 n9132 n555 R=1.063e+01 
R9131t7872 n9132 n7873 R=8.046e+00 
R9131t182 n9132 n183 R=3.717e+00 
R9131t8803 n9132 n8804 R=5.880e+00 
R9131t2822 n9132 n2823 R=7.342e+00 
R9132t2498 n9133 n2499 R=1.631e+01 
R9132t6103 n9133 n6104 R=4.128e+00 
R9132t2169 n9133 n2170 R=1.166e+01 
R9132t8129 n9133 n8130 R=3.055e+00 
R9132t5104 n9133 n5105 R=1.708e+01 
R9132t4988 n9133 n4989 R=1.598e+01 
R9133t6377 n9134 n6378 R=1.506e+01 
R9133t8216 n9134 n8217 R=1.446e+01 
R9133t2806 n9134 n2807 R=3.515e+01 
R9133t5021 n9134 n5022 R=3.923e+00 
R9133t4279 n9134 n4280 R=1.893e+01 
R9133t2380 n9134 n2381 R=5.383e+00 
R9133t240 n9134 n241 R=5.563e+00 
R9134t300 n9135 n301 R=7.696e+00 
R9134t4415 n9135 n4416 R=3.759e+00 
R9134t3189 n9135 n3190 R=1.058e+01 
R9134t6460 n9135 n6461 R=4.673e+00 
R9135t4904 n9136 n4905 R=8.663e+00 
R9135t7474 n9136 n7475 R=2.960e+01 
R9135t2933 n9136 n2934 R=9.600e+00 
R9135t6875 n9136 n6876 R=2.148e+00 
R9135t7524 n9136 n7525 R=1.574e+01 
R9135t7492 n9136 n7493 R=5.842e+00 
R9136t650 n9137 n651 R=8.233e+00 
R9136t3839 n9137 n3840 R=3.212e+01 
R9136t203 n9137 n204 R=6.688e+00 
R9136t7985 n9137 n7986 R=3.615e+00 
R9137t4472 n1 n4473 R=1.490e+01 
R9137t4224 n1 n4225 R=4.347e+01 
R9137t7639 n1 n7640 R=9.866e+01 
R9137t9098 n1 n9099 R=2.383e+01 
R9138t632 n9139 n633 R=7.799e+00 
R9138t4788 n9139 n4789 R=4.502e+00 
R9138t508 n9139 n509 R=5.869e+01 
R9138t6831 n9139 n6832 R=4.008e+00 
R9139t3471 n9140 n3472 R=1.877e+00 
R9139t6100 n9140 n6101 R=8.035e+00 
R9139t7650 n9140 n7651 R=1.039e+01 
R9139t5659 n9140 n5660 R=4.074e+00 
R9139t2312 n9140 n2313 R=6.425e+01 
R9140t4431 n9141 n4432 R=5.798e+00 
R9140t703 n9141 n704 R=3.277e+00 
R9140t9044 n9141 n9045 R=1.079e+01 
R9140t1857 n9141 n1858 R=1.006e+01 
R9140t3427 n9141 n3428 R=1.544e+01 
R9141t4844 n9142 n4845 R=2.233e+01 
R9141t5729 n9142 n5730 R=3.121e+01 
R9141t4686 n9142 n4687 R=4.526e+00 
R9141t527 n9142 n528 R=5.390e+00 
R9141t8977 n9142 n8978 R=2.062e+01 
R9141t1642 n9142 n1643 R=1.974e+01 
R9141t6208 n9142 n6209 R=4.350e+00 
R9142t8720 n9143 n8721 R=5.008e+00 
R9142t9093 n9143 n9094 R=3.256e+00 
R9142t1543 n9143 n1544 R=4.819e+00 
R9142t7899 n9143 n7900 R=5.485e+00 
R9143t1312 n9144 n1313 R=1.253e+01 
R9143t2776 n9144 n2777 R=2.812e+00 
R9143t3680 n9144 n3681 R=1.335e+01 
R9143t8734 n9144 n8735 R=8.736e+00 
R9144t2378 n9145 n2379 R=3.421e+00 
R9144t2967 n9145 n2968 R=2.713e+01 
R9144t3497 n9145 n3498 R=7.523e+00 
R9144t6439 n9145 n6440 R=8.620e+00 
R9144t3784 n9145 n3785 R=2.825e+00 
R9145t3550 n9146 n3551 R=9.127e+00 
R9145t6151 n9146 n6152 R=3.464e+01 
R9145t9035 n9146 n9036 R=5.317e+00 
R9145t8178 n9146 n8179 R=8.344e+02 
R9145t7507 n9146 n7508 R=2.720e+00 
R9145t2209 n9146 n2210 R=5.892e+00 
R9146t4696 n9147 n4697 R=3.348e+00 
R9146t5381 n9147 n5382 R=1.533e+01 
R9146t1656 n9147 n1657 R=1.528e+01 
R9146t5777 n9147 n5778 R=3.989e+00 
R9146t6840 n9147 n6841 R=8.815e+00 
R9147t2560 n9148 n2561 R=4.257e+00 
R9147t7565 n9148 n7566 R=2.647e+01 
R9147t1577 n9148 n1578 R=6.149e+00 
R9147t5282 n9148 n5283 R=2.248e+01 
R9147t4210 n9148 n4211 R=3.467e+01 
R9147t8112 n9148 n8113 R=1.506e+00 
R9148t577 n9149 n578 R=5.106e+00 
R9148t8762 n9149 n8763 R=1.207e+01 
R9148t1989 n9149 n1990 R=3.985e+00 
R9148t873 n9149 n874 R=2.832e+01 
R9148t1601 n9149 n1602 R=6.975e+00 
R9148t3433 n9149 n3434 R=3.227e+00 
R9149t1614 n9150 n1615 R=3.004e+01 
R9149t4259 n9150 n4260 R=6.037e+00 
R9149t4707 n9150 n4708 R=6.849e+01 
R9149t715 n9150 n716 R=4.550e+00 
R9149t2891 n9150 n2892 R=1.723e+01 
R9149t7597 n9150 n7598 R=2.183e+01 
R9149t8802 n9150 n8803 R=6.377e+00 
R9149t6837 n9150 n6838 R=2.677e+01 
R9149t2861 n9150 n2862 R=1.286e+01 
R9150t7039 n9151 n7040 R=2.044e+01 
R9150t9075 n9151 n9076 R=2.218e+00 
R9150t6429 n9151 n6430 R=1.004e+01 
R9150t6861 n9151 n6862 R=1.683e+01 
R9150t1528 n9151 n1529 R=6.058e+00 
R9150t7757 n9151 n7758 R=1.479e+01 
R9151t7718 n9152 n7719 R=3.673e+00 
R9151t7882 n9152 n7883 R=3.420e+00 
R9152t2563 n9153 n2564 R=4.672e+00 
R9152t6058 n9153 n6059 R=3.572e+00 
R9152t3683 n9153 n3684 R=2.271e+00 
R9153t5086 n9154 n5087 R=3.990e+00 
R9153t8957 n9154 n8958 R=8.466e+00 
R9153t4433 n9154 n4434 R=8.837e+00 
R9153t7836 n9154 n7837 R=7.106e+01 
R9153t6226 n9154 n6227 R=3.222e+01 
R9153t8969 n9154 n8970 R=2.279e+01 
R9153t6908 n9154 n6909 R=3.186e+00 
R9153t3468 n9154 n3469 R=1.313e+01 
R9154t4453 n9155 n4454 R=1.730e+01 
R9154t7728 n9155 n7729 R=4.374e+00 
R9154t5574 n9155 n5575 R=8.051e+00 
R9154t7349 n9155 n7350 R=7.292e+00 
R9155t4502 n9156 n4503 R=3.875e+00 
R9155t5221 n9156 n5222 R=9.736e+00 
R9155t2383 n9156 n2384 R=4.620e+00 
R9155t999 n9156 n1000 R=4.521e+01 
R9155t9001 n9156 n9002 R=9.938e+00 
R9155t3591 n9156 n3592 R=9.580e+00 
R9156t1615 n9157 n1616 R=4.196e+01 
R9156t6809 n9157 n6810 R=5.119e+00 
R9156t3877 n9157 n3878 R=1.146e+01 
R9156t5499 n9157 n5500 R=1.743e+01 
R9156t5718 n9157 n5719 R=3.575e+01 
R9156t1869 n9157 n1870 R=5.134e+00 
R9156t1472 n9157 n1473 R=3.508e+00 
R9157t698 n9158 n699 R=1.029e+01 
R9157t1595 n9158 n1596 R=2.620e+01 
R9157t8650 n9158 n8651 R=4.238e+00 
R9157t2580 n9158 n2581 R=2.449e+01 
R9157t2961 n9158 n2962 R=1.323e+01 
R9157t2002 n9158 n2003 R=7.173e+00 
R9157t4136 n9158 n4137 R=6.894e+00 
R9157t1485 n9158 n1486 R=1.766e+01 
R9158t1815 n9159 n1816 R=9.162e+00 
R9158t3579 n9159 n3580 R=5.977e+00 
R9159t1420 n9160 n1421 R=1.904e+00 
R9159t634 n9160 n635 R=8.967e+00 
R9159t3368 n9160 n3369 R=3.528e+00 
R9159t2700 n9160 n2701 R=1.344e+01 
R9160t1899 n9161 n1900 R=7.915e+00 
R9160t5183 n9161 n5184 R=1.076e+01 
R9160t4240 n9161 n4241 R=1.402e+01 
R9160t5530 n9161 n5531 R=3.885e+00 
R9160t4947 n9161 n4948 R=5.067e+00 
R9161t1332 n9162 n1333 R=4.212e+00 
R9161t3274 n9162 n3275 R=7.471e+00 
R9161t3970 n9162 n3971 R=7.089e+00 
R9161t5496 n9162 n5497 R=1.210e+01 
R9161t3208 n9162 n3209 R=1.145e+01 
R9162t3964 n9163 n3965 R=4.165e+00 
R9162t2216 n9163 n2217 R=6.709e+00 
R9162t7042 n9163 n7043 R=2.999e+01 
R9162t6328 n9163 n6329 R=3.819e+00 
R9163t1332 n9164 n1333 R=8.263e+00 
R9163t3274 n9164 n3275 R=4.929e+00 
R9163t1718 n9164 n1719 R=3.252e+01 
R9163t7028 n9164 n7029 R=3.423e+00 
R9164t303 n9165 n304 R=3.473e+00 
R9164t13 n9165 n14 R=6.242e+00 
R9164t9016 n9165 n9017 R=1.120e+01 
R9165t1085 n9166 n1086 R=5.787e+00 
R9165t2079 n9166 n2080 R=4.643e+00 
R9165t8454 n9166 n8455 R=7.721e+01 
R9165t2224 n9166 n2225 R=1.075e+01 
R9165t5413 n9166 n5414 R=6.869e+00 
R9165t7723 n9166 n7724 R=6.825e+00 
R9166t6328 n9167 n6329 R=5.760e+00 
R9166t6767 n9167 n6768 R=2.702e+00 
R9166t9162 n9167 n9163 R=7.695e+00 
R9166t3964 n9167 n3965 R=1.013e+01 
R9166t5232 n9167 n5233 R=1.074e+01 
R9166t5601 n9167 n5602 R=5.952e+00 
R9167t1545 n9168 n1546 R=1.506e+01 
R9167t1739 n9168 n1740 R=1.937e+01 
R9167t947 n9168 n948 R=4.027e+01 
R9167t6325 n9168 n6326 R=5.182e+00 
R9167t6259 n9168 n6260 R=3.753e+00 
R9167t8506 n9168 n8507 R=7.578e+01 
R9167t5098 n9168 n5099 R=2.525e+00 
R9168t1593 n9169 n1594 R=7.724e+01 
R9168t3247 n9169 n3248 R=5.379e+00 
R9168t668 n9169 n669 R=4.268e+00 
R9168t2052 n9169 n2053 R=6.979e+00 
R9169t3298 n9170 n3299 R=1.937e+00 
R9169t5560 n9170 n5561 R=8.353e+00 
R9169t8526 n9170 n8527 R=3.937e+01 
R9169t3222 n9170 n3223 R=4.847e+00 
R9170t806 n9171 n807 R=2.668e+01 
R9170t384 n9171 n385 R=1.898e+01 
R9170t9106 n9171 n9107 R=2.785e+01 
R9170t756 n9171 n757 R=1.002e+01 
R9170t3931 n9171 n3932 R=2.251e+00 
R9171t1718 n9172 n1719 R=4.811e+00 
R9171t3751 n9172 n3752 R=7.259e+00 
R9171t9163 n9172 n9164 R=8.077e+00 
R9171t7028 n9172 n7029 R=1.059e+01 
R9171t7332 n9172 n7333 R=2.773e+00 
R9172t4935 n9173 n4936 R=8.963e+00 
R9172t7290 n9173 n7291 R=3.512e+00 
R9172t1312 n9173 n1313 R=6.080e+01 
R9172t9143 n9173 n9144 R=3.090e+00 
R9172t3680 n9173 n3681 R=7.973e+00 
R9173t541 n9174 n542 R=7.965e+00 
R9173t5075 n9174 n5076 R=2.300e+01 
R9173t1202 n9174 n1203 R=3.322e+00 
R9173t2371 n9174 n2372 R=5.856e+00 
R9173t2011 n9174 n2012 R=4.690e+00 
R9174t4905 n9175 n4906 R=7.738e+00 
R9174t7571 n9175 n7572 R=6.851e+01 
R9174t2717 n9175 n2718 R=1.628e+01 
R9174t564 n9175 n565 R=3.842e+02 
R9174t6 n9175 n7 R=8.562e+00 
R9174t799 n9175 n800 R=7.296e+00 
R9174t4071 n9175 n4072 R=7.236e+00 
R9174t7003 n9175 n7004 R=1.232e+01 
R9175t1692 n9176 n1693 R=2.430e+01 
R9175t7238 n9176 n7239 R=2.826e+00 
R9175t1375 n9176 n1376 R=4.586e+00 
R9175t8600 n9176 n8601 R=4.493e+01 
R9176t7370 n9177 n7371 R=6.206e+00 
R9176t8221 n9177 n8222 R=1.152e+01 
R9176t7866 n9177 n7867 R=5.565e+00 
R9176t6269 n9177 n6270 R=1.170e+01 
R9176t1455 n9177 n1456 R=9.388e+00 
R9176t5349 n9177 n5350 R=5.170e+00 
R9176t4274 n9177 n4275 R=1.813e+02 
R9177t711 n9178 n712 R=5.873e+00 
R9177t7667 n9178 n7668 R=2.970e+01 
R9177t2477 n9178 n2478 R=7.755e+00 
R9177t8927 n9178 n8928 R=1.385e+01 
R9177t2967 n9178 n2968 R=3.441e+00 
R9177t3784 n9178 n3785 R=1.073e+02 
R9178t2623 n9179 n2624 R=5.541e+01 
R9178t4424 n9179 n4425 R=2.244e+00 
R9178t4660 n9179 n4661 R=4.560e+01 
R9178t994 n9179 n995 R=1.465e+02 
R9178t1736 n9179 n1737 R=4.713e+00 
R9178t5629 n9179 n5630 R=6.573e+00 
R9178t6540 n9179 n6541 R=4.577e+01 
R9178t5171 n9179 n5172 R=1.782e+01 
R9179t6444 n9180 n6445 R=3.640e+00 
R9179t7072 n9180 n7073 R=1.319e+01 
R9179t768 n9180 n769 R=8.293e+01 
R9179t8114 n9180 n8115 R=4.844e+00 
R9179t2081 n9180 n2082 R=2.591e+01 
R9179t2373 n9180 n2374 R=3.468e+00 
R9180t6081 n9181 n6082 R=5.144e+01 
R9180t6720 n9181 n6721 R=1.889e+00 
R9180t20 n9181 n21 R=2.477e+01 
R9180t7186 n9181 n7187 R=3.870e+00 
R9180t2737 n9181 n2738 R=7.159e+00 
R9180t5143 n9181 n5144 R=2.327e+01 
R9181t1822 n9182 n1823 R=2.080e+00 
R9181t3738 n9182 n3739 R=3.586e+01 
R9181t7069 n9182 n7070 R=3.084e+01 
R9181t2485 n9182 n2486 R=4.034e+00 
R9181t3130 n9182 n3131 R=2.247e+01 
R9181t1917 n9182 n1918 R=7.254e+00 
R9182t2360 n9183 n2361 R=5.460e+00 
R9182t3090 n9183 n3091 R=2.064e+01 
R9182t2438 n9183 n2439 R=5.575e+00 
R9182t2301 n9183 n2302 R=5.594e+00 
R9183t1098 n9184 n1099 R=1.128e+01 
R9183t3871 n9184 n3872 R=7.461e+00 
R9183t7210 n9184 n7211 R=4.803e+00 
R9183t391 n9184 n392 R=9.187e+00 
R9184t6096 n9185 n6097 R=1.612e+01 
R9184t6740 n9185 n6741 R=1.760e+01 
R9184t4448 n9185 n4449 R=3.187e+00 
R9184t7917 n9185 n7918 R=6.282e+00 
R9185t5700 n9186 n5701 R=5.710e+00 
R9185t7267 n9186 n7268 R=2.294e+01 
R9185t828 n9186 n829 R=6.570e+00 
R9185t7576 n9186 n7577 R=1.132e+01 
R9185t1232 n9186 n1233 R=2.811e+00 
R9185t6841 n9186 n6842 R=4.847e+02 
R9186t1544 n9187 n1545 R=7.360e+00 
R9186t5045 n9187 n5046 R=1.339e+01 
R9186t4321 n9187 n4322 R=2.397e+00 
R9186t3590 n9187 n3591 R=3.932e+01 
R9186t8524 n9187 n8525 R=2.854e+00 
R9187t6447 n9188 n6448 R=9.261e+00 
R9187t6873 n9188 n6874 R=1.447e+01 
R9187t8544 n9188 n8545 R=1.588e+01 
R9187t2087 n9188 n2088 R=4.305e+00 
R9187t1129 n9188 n1130 R=1.929e+01 
R9187t2254 n9188 n2255 R=5.651e+00 
R9188t1680 n9189 n1681 R=2.114e+01 
R9188t7014 n9189 n7015 R=1.050e+01 
R9188t7405 n9189 n7406 R=5.278e+00 
R9188t8104 n9189 n8105 R=6.587e+00 
R9188t5994 n9189 n5995 R=2.133e+01 
R9188t2008 n9189 n2009 R=4.058e+01 
R9188t4701 n9189 n4702 R=4.101e+00 
R9189t8264 n9190 n8265 R=1.128e+02 
R9189t7539 n9190 n7540 R=9.172e+00 
R9189t8704 n9190 n8705 R=2.234e+01 
R9189t1052 n9190 n1053 R=6.323e+00 
R9189t6271 n9190 n6272 R=6.896e+01 
R9189t1698 n9190 n1699 R=1.086e+01 
R9190t2133 n9191 n2134 R=3.742e+00 
R9190t3404 n9191 n3405 R=1.328e+01 
R9190t6676 n9191 n6677 R=3.452e+01 
R9190t7540 n9191 n7541 R=3.585e+00 
R9190t5969 n9191 n5970 R=1.936e+02 
R9191t3260 n9192 n3261 R=2.454e+01 
R9191t4946 n9192 n4947 R=6.056e+00 
R9191t3303 n9192 n3304 R=2.167e+00 
R9191t1082 n9192 n1083 R=4.496e+02 
R9191t7912 n9192 n7913 R=4.477e+00 
R9191t4600 n9192 n4601 R=1.307e+01 
R9192t6268 n9193 n6269 R=6.017e+00 
R9192t8321 n9193 n8322 R=2.751e+01 
R9192t7766 n9193 n7767 R=6.245e+00 
R9192t9083 n9193 n9084 R=2.369e+01 
R9192t8109 n9193 n8110 R=3.634e+00 
R9193t5637 n9194 n5638 R=6.487e+00 
R9193t6727 n9194 n6728 R=1.398e+01 
R9193t189 n9194 n190 R=8.795e+00 
R9193t7325 n9194 n7326 R=4.545e+02 
R9193t8350 n9194 n8351 R=9.155e+00 
R9193t6511 n9194 n6512 R=2.854e+00 
R9194t2914 n9195 n2915 R=5.208e+00 
R9194t5522 n9195 n5523 R=1.868e+01 
R9194t6894 n9195 n6895 R=2.192e+01 
R9194t5692 n9195 n5693 R=1.025e+01 
R9194t5095 n9195 n5096 R=1.011e+01 
R9195t64 n9196 n65 R=4.700e+01 
R9195t3072 n9196 n3073 R=3.781e+00 
R9195t245 n9196 n246 R=3.719e+00 
R9195t460 n9196 n461 R=5.800e+00 
R9196t46 n9197 n47 R=9.248e+00 
R9196t289 n9197 n290 R=3.558e+00 
R9196t4483 n9197 n4484 R=5.461e+00 
R9196t2650 n9197 n2651 R=3.753e+01 
R9196t8611 n9197 n8612 R=9.329e+00 
R9197t1514 n9198 n1515 R=3.033e+01 
R9197t3703 n9198 n3704 R=1.625e+01 
R9197t3199 n9198 n3200 R=5.871e+00 
R9197t6089 n9198 n6090 R=7.742e+00 
R9197t8328 n9198 n8329 R=1.015e+01 
R9197t7123 n9198 n7124 R=6.609e+00 
R9197t5957 n9198 n5958 R=7.233e+00 
R9198t295 n9199 n296 R=5.014e+00 
R9198t4927 n9199 n4928 R=3.191e+00 
R9198t5246 n9199 n5247 R=9.277e+00 
R9198t1350 n9199 n1351 R=7.086e+00 
R9198t872 n9199 n873 R=1.812e+01 
R9199t926 n9200 n927 R=3.315e+00 
R9199t7754 n9200 n7755 R=4.180e+01 
R9199t1594 n9200 n1595 R=4.439e+00 
R9199t6062 n9200 n6063 R=8.005e+00 
R9199t5206 n9200 n5207 R=1.072e+01 
R9200t695 n9201 n696 R=7.158e+00 
R9200t5802 n9201 n5803 R=4.464e+00 
R9200t3129 n9201 n3130 R=9.520e+00 
R9200t5422 n9201 n5423 R=1.255e+01 
R9200t1372 n9201 n1373 R=4.019e+00 
R9201t4924 n9202 n4925 R=6.268e+00 
R9201t5329 n9202 n5330 R=3.246e+00 
R9201t8725 n9202 n8726 R=1.396e+02 
R9201t3510 n9202 n3511 R=5.619e+00 
R9201t1156 n9202 n1157 R=3.691e+00 
R9201t7145 n9202 n7146 R=3.662e+01 
R9202t413 n9203 n414 R=2.567e+01 
R9202t6176 n9203 n6177 R=2.210e+01 
R9202t4485 n9203 n4486 R=4.170e+00 
R9202t7829 n9203 n7830 R=5.939e+00 
R9202t7732 n9203 n7733 R=4.036e+01 
R9202t5769 n9203 n5770 R=6.728e+00 
R9202t8703 n9203 n8704 R=7.044e+00 
R9203t4586 n9204 n4587 R=2.968e+00 
R9203t7307 n9204 n7308 R=5.975e+00 
R9203t7877 n9204 n7878 R=2.183e+01 
R9203t8045 n9204 n8046 R=8.858e+00 
R9203t40 n9204 n41 R=4.212e+00 
R9203t5437 n9204 n5438 R=1.020e+02 
R9204t3085 n9205 n3086 R=5.768e+00 
R9204t6933 n9205 n6934 R=6.134e+00 
R9204t5574 n9205 n5575 R=2.232e+01 
R9204t3384 n9205 n3385 R=1.847e+01 
R9204t2259 n9205 n2260 R=8.011e+00 
R9205t6167 n9206 n6168 R=7.024e+00 
R9205t4012 n9206 n4013 R=8.029e+00 
R9205t5463 n9206 n5464 R=9.948e+01 
R9205t5309 n9206 n5310 R=2.719e+00 
R9205t8697 n9206 n8698 R=1.612e+01 
R9206t1107 n9207 n1108 R=2.384e+01 
R9206t1527 n9207 n1528 R=2.414e+01 
R9206t1329 n9207 n1330 R=2.092e+01 
R9206t4012 n9207 n4013 R=7.232e+00 
R9206t9205 n9207 n9206 R=5.215e+00 
R9206t6167 n9207 n6168 R=1.162e+01 
R9207t8 n9208 n9 R=1.265e+01 
R9207t3026 n9208 n3027 R=9.098e+01 
R9207t6460 n9208 n6461 R=2.708e+00 
R9207t3802 n9208 n3803 R=4.201e+00 
R9208t5658 n9209 n5659 R=4.531e+00 
R9208t7463 n9209 n7464 R=5.733e+00 
R9208t1762 n9209 n1763 R=1.421e+01 
R9208t7909 n9209 n7910 R=2.543e+00 
R9208t7631 n9209 n7632 R=3.171e+01 
R9209t6688 n9210 n6689 R=2.260e+03 
R9209t8065 n9210 n8066 R=4.765e+00 
R9209t8151 n9210 n8152 R=3.594e+01 
R9209t3852 n9210 n3853 R=7.498e+00 
R9209t6062 n9210 n6063 R=7.322e+00 
R9209t469 n9210 n470 R=8.276e+00 
R9209t5689 n9210 n5690 R=6.289e+00 
R9209t4615 n9210 n4616 R=2.064e+02 
R9210t2707 n9211 n2708 R=3.268e+00 
R9210t6130 n9211 n6131 R=1.195e+01 
R9210t2297 n9211 n2298 R=9.068e+00 
R9210t506 n9211 n507 R=3.101e+00 
R9211t171 n9212 n172 R=4.700e+00 
R9211t4509 n9212 n4510 R=7.416e+00 
R9211t2482 n9212 n2483 R=5.293e+01 
R9211t8780 n9212 n8781 R=1.579e+01 
R9211t2715 n9212 n2716 R=2.554e+01 
R9211t7377 n9212 n7378 R=3.043e+00 
R9211t1531 n9212 n1532 R=2.833e+01 
R9211t7078 n9212 n7079 R=1.050e+01 
R9212t7138 n9213 n7139 R=1.639e+01 
R9212t8523 n9213 n8524 R=1.930e+00 
R9212t4362 n9213 n4363 R=4.030e+01 
R9212t1889 n9213 n1 R=6.335e+00 
R9212t42 n9213 n43 R=3.393e+00 
R9213t2714 n9214 n2715 R=2.093e+01 
R9213t4464 n9214 n4465 R=1.034e+01 
R9213t6485 n9214 n6486 R=5.851e+00 
R9213t2099 n9214 n2100 R=3.914e+00 
R9213t952 n9214 n953 R=2.757e+00 
R9214t5821 n9215 n5822 R=1.677e+01 
R9214t8077 n9215 n8078 R=3.650e+00 
R9214t3126 n9215 n3127 R=8.387e+00 
R9214t5111 n9215 n5112 R=3.800e+00 
R9214t8709 n9215 n8710 R=5.365e+01 
R9215t7882 n9216 n7883 R=5.659e+02 
R9215t4510 n9216 n4511 R=8.328e+01 
R9215t4870 n9216 n4871 R=3.515e+00 
R9215t6523 n9216 n6524 R=3.693e+02 
R9215t7718 n9216 n7719 R=3.235e+01 
R9215t9151 n9216 n9152 R=2.960e+00 
R9216t2664 n9217 n2665 R=1.862e+01 
R9216t5266 n9217 n5267 R=1.832e+00 
R9216t96 n9217 n97 R=5.413e+01 
R9216t4256 n9217 n4257 R=8.151e+00 
R9216t1763 n9217 n1764 R=1.969e+00 
R9216t7257 n9217 n7258 R=1.380e+01 
R9217t2715 n9218 n2716 R=1.368e+01 
R9217t6862 n9218 n6863 R=9.752e+00 
R9217t151 n9218 n152 R=3.314e+00 
R9217t6164 n9218 n6165 R=6.314e+01 
R9217t7450 n9218 n7451 R=1.745e+01 
R9217t904 n9218 n905 R=5.461e+00 
R9218t2006 n9219 n2007 R=1.584e+00 
R9218t4651 n9219 n4652 R=3.404e+01 
R9218t8032 n9219 n8033 R=1.161e+01 
R9218t949 n9219 n950 R=1.425e+00 
R9218t4676 n9219 n4677 R=1.829e+02 
R9219t4364 n9220 n4365 R=4.262e+00 
R9219t6289 n9220 n6290 R=1.906e+01 
R9219t6167 n9220 n6168 R=9.624e+00 
R9219t9205 n9220 n9206 R=1.235e+02 
R9219t8697 n9220 n8698 R=9.871e+00 
R9219t6884 n9220 n6885 R=3.506e+01 
R9219t7413 n9220 n7414 R=3.008e+00 
R9220t1205 n9221 n1206 R=2.196e+01 
R9220t4370 n9221 n4371 R=5.079e+01 
R9220t4762 n9221 n4763 R=4.745e+00 
R9220t2311 n9221 n2312 R=3.509e+00 
R9220t7759 n9221 n7760 R=9.572e+00 
R9220t512 n9221 n513 R=3.165e+03 
R9220t1833 n9221 n1834 R=5.579e+00 
R9221t1089 n9222 n1090 R=2.964e+01 
R9221t6551 n9222 n6552 R=3.198e+00 
R9221t6188 n9222 n6189 R=1.164e+02 
R9221t6237 n9222 n6238 R=9.224e+00 
R9221t1286 n9222 n1287 R=1.062e+03 
R9221t90 n9222 n91 R=5.250e+00 
R9221t4757 n9222 n4758 R=6.121e+00 
R9222t1750 n9223 n1751 R=1.018e+01 
R9222t4097 n9223 n4098 R=1.248e+02 
R9222t4605 n9223 n4606 R=3.258e+00 
R9222t6291 n9223 n6292 R=5.600e+00 
R9222t5229 n9223 n5230 R=4.205e+00 
R9223t1086 n9224 n1087 R=5.906e+01 
R9223t9021 n9224 n9022 R=1.414e+01 
R9223t3407 n9224 n3408 R=5.458e+00 
R9223t6373 n9224 n6374 R=5.679e+00 
R9223t2005 n9224 n2006 R=1.719e+01 
R9223t8140 n9224 n8141 R=3.648e+00 
R9224t1831 n9225 n1832 R=3.137e+00 
R9224t4673 n9225 n4674 R=5.227e+00 
R9224t6297 n9225 n6298 R=1.541e+01 
R9224t950 n9225 n951 R=4.061e+00 
R9225t5258 n9226 n5259 R=7.151e+00 
R9225t7812 n9226 n7813 R=1.227e+01 
R9226t491 n9227 n492 R=1.614e+01 
R9226t6173 n9227 n6174 R=2.737e+01 
R9226t7043 n9227 n7044 R=3.649e+01 
R9226t3795 n9227 n3796 R=6.919e+01 
R9226t8019 n9227 n8020 R=5.200e+00 
R9226t526 n9227 n527 R=1.124e+01 
R9227t4802 n9228 n4803 R=3.288e+01 
R9227t6178 n9228 n6179 R=5.900e+01 
R9227t1209 n9228 n1210 R=2.123e+00 
R9227t7419 n9228 n7420 R=1.758e+01 
R9227t4206 n9228 n4207 R=1.884e+01 
R9227t8201 n9228 n8202 R=1.817e+00 
R9228t2327 n9229 n2328 R=2.829e+00 
R9228t7375 n9229 n7376 R=3.634e+00 
R9228t771 n9229 n772 R=4.066e+00 
R9228t5113 n9229 n5114 R=1.290e+01 
R9229t2927 n9230 n2928 R=1.762e+01 
R9229t2967 n9230 n2968 R=9.423e+00 
R9229t510 n9230 n511 R=6.861e+00 
R9229t9004 n9230 n9005 R=1.932e+01 
R9229t2749 n9230 n2750 R=8.848e+00 
R9229t2378 n9230 n2379 R=4.214e+00 
R9230t1447 n9231 n1448 R=8.301e+00 
R9230t9015 n9231 n9016 R=8.659e+00 
R9230t2158 n9231 n2159 R=2.200e+01 
R9230t3873 n9231 n3874 R=2.660e+01 
R9230t121 n9231 n122 R=1.201e+01 
R9230t6723 n9231 n6724 R=1.416e+01 
R9230t7181 n9231 n7182 R=2.538e+00 
R9230t4146 n9231 n4147 R=1.568e+02 
R9231t4245 n9232 n4246 R=1.982e+00 
R9231t4606 n9232 n4607 R=1.571e+01 
R9231t8728 n9232 n8729 R=2.809e+00 
R9231t751 n9232 n752 R=1.101e+01 
R9232t7230 n9233 n7231 R=7.982e+00 
R9232t8442 n9233 n8443 R=1.234e+01 
R9232t6669 n9233 n6670 R=3.762e+00 
R9232t1970 n9233 n1971 R=6.960e+00 
R9232t3216 n9233 n3217 R=3.597e+00 
R9233t16 n9234 n17 R=6.806e+01 
R9233t9121 n9234 n9122 R=4.759e+00 
R9233t6198 n9234 n6199 R=1.556e+01 
R9233t6399 n9234 n6400 R=6.454e+00 
R9233t1855 n9234 n1856 R=8.911e+00 
R9233t5913 n9234 n5914 R=4.283e+00 
R9234t4492 n9235 n4493 R=6.761e+00 
R9234t7263 n9235 n7264 R=1.207e+01 
R9234t8659 n9235 n8660 R=2.871e+00 
R9234t2361 n9235 n2362 R=1.126e+01 
R9235t1805 n9236 n1806 R=1.526e+01 
R9235t8015 n9236 n8016 R=4.498e+00 
R9235t5205 n9236 n5206 R=1.247e+01 
R9235t7031 n9236 n7032 R=1.324e+01 
R9235t8946 n9236 n8947 R=5.533e+00 
R9235t6316 n9236 n6317 R=9.491e+00 
R9236t4717 n9237 n4718 R=1.998e+00 
R9236t4930 n9237 n4931 R=3.837e+00 
R9236t6823 n9237 n6824 R=1.224e+01 
R9236t1846 n9237 n1847 R=1.175e+01 
R9236t4875 n9237 n4876 R=1.303e+01 
R9237t299 n9238 n300 R=3.746e+00 
R9237t8389 n9238 n8390 R=4.620e+01 
R9237t4727 n9238 n4728 R=4.387e+00 
R9237t2908 n9238 n2909 R=3.998e+00 
R9237t3556 n9238 n3557 R=2.705e+01 
R9238t1561 n9239 n1562 R=8.645e+00 
R9238t4872 n9239 n4873 R=1.522e+01 
R9238t1785 n9239 n1786 R=8.087e+00 
R9238t7974 n9239 n7975 R=3.741e+00 
R9239t5518 n9240 n5519 R=1.189e+01 
R9239t7644 n9240 n7645 R=5.923e+00 
R9239t585 n9240 n586 R=1.428e+01 
R9239t3312 n9240 n3313 R=1.948e+00 
R9239t4863 n9240 n4864 R=2.791e+01 
R9239t4544 n9240 n4545 R=7.707e+01 
R9239t5224 n9240 n5225 R=7.207e+00 
R9240t2441 n9241 n2442 R=2.810e+01 
R9240t2478 n9241 n2479 R=6.838e+00 
R9240t2917 n9241 n2918 R=5.841e+00 
R9240t7718 n9241 n7719 R=1.492e+02 
R9240t9215 n9241 n9216 R=1.566e+01 
R9240t6523 n9241 n6524 R=7.381e+00 
R9240t6679 n9241 n6680 R=7.580e+00 
R9241t2384 n9242 n2385 R=2.898e+00 
R9241t5648 n9242 n5649 R=7.222e+00 
R9241t2783 n9242 n2784 R=1.377e+01 
R9241t7643 n9242 n7644 R=6.807e+00 
R9242t3023 n9243 n3024 R=5.173e+00 
R9242t4852 n9243 n4853 R=4.040e+00 
R9242t2335 n9243 n2336 R=1.137e+01 
R9242t8323 n9243 n8324 R=8.440e+00 
R9242t2683 n9243 n2684 R=7.133e+00 
R9243t813 n9244 n814 R=2.000e+01 
R9243t2687 n9244 n2688 R=2.011e+00 
R9243t6694 n9244 n6695 R=8.601e+00 
R9243t6273 n9244 n6274 R=1.065e+01 
R9243t7737 n9244 n7738 R=5.098e+00 
R9244t7083 n9245 n7084 R=1.534e+00 
R9244t7764 n9245 n7765 R=3.357e+01 
R9244t8046 n9245 n8047 R=9.581e+00 
R9244t2905 n9245 n2906 R=5.069e+00 
R9244t1788 n9245 n1789 R=5.163e+00 
R9245t2923 n9246 n2924 R=5.963e+00 
R9245t3411 n9246 n3412 R=2.142e+01 
R9245t5987 n9246 n5988 R=4.380e+00 
R9245t1900 n9246 n1901 R=1.677e+01 
R9245t1608 n9246 n1609 R=6.452e+00 
R9246t2419 n9247 n2420 R=1.284e+01 
R9246t6695 n9247 n6696 R=7.260e+00 
R9246t4440 n9247 n4441 R=7.963e+00 
R9246t4961 n9247 n4962 R=1.542e+01 
R9246t2699 n9247 n2700 R=6.406e+00 
R9246t8524 n9247 n8525 R=7.445e+00 
R9247t908 n9248 n909 R=1.057e+01 
R9247t7732 n9248 n7733 R=1.575e+01 
R9247t5769 n9248 n5770 R=6.248e+01 
R9247t8148 n9248 n8149 R=8.318e+00 
R9247t1885 n9248 n1886 R=1.729e+01 
R9247t388 n9248 n389 R=5.095e+00 
R9247t3616 n9248 n3617 R=1.698e+01 
R9247t8763 n9248 n8764 R=9.159e+00 
R9248t5563 n9249 n5564 R=8.160e+00 
R9248t8219 n9249 n8220 R=2.541e+02 
R9248t3557 n9249 n3558 R=4.549e+00 
R9248t4860 n9249 n4861 R=9.724e+01 
R9248t5577 n9249 n5578 R=3.274e+00 
R9248t2654 n9249 n2655 R=7.658e+00 
R9248t8567 n9249 n8568 R=1.978e+01 
R9249t4696 n9250 n4697 R=3.038e+00 
R9249t5618 n9250 n5619 R=3.829e+00 
R9249t7852 n9250 n7853 R=4.926e+01 
R9249t1656 n9250 n1657 R=5.040e+00 
R9249t9146 n9250 n9147 R=2.584e+01 
R9250t3003 n9251 n3004 R=5.444e+00 
R9250t6980 n9251 n6981 R=1.529e+01 
R9250t1224 n9251 n1225 R=3.985e+00 
R9250t7331 n9251 n7332 R=3.947e+00 
R9251t1426 n9252 n1427 R=5.864e+00 
R9251t6381 n9252 n6382 R=2.838e+00 
R9251t6929 n9252 n6930 R=6.690e+00 
R9251t2191 n9252 n2192 R=9.062e+00 
R9251t8800 n9252 n8801 R=1.546e+01 
R9251t6092 n9252 n6093 R=5.822e+01 
R9252t6614 n9253 n6615 R=3.402e+00 
R9252t3533 n9253 n3534 R=7.104e+00 
R9252t237 n9253 n238 R=7.396e+00 
R9252t7879 n9253 n7880 R=3.217e+00 
R9253t2274 n9254 n2275 R=2.152e+02 
R9253t7970 n9254 n7971 R=3.240e+01 
R9253t3775 n9254 n3776 R=2.430e+00 
R9253t7142 n9254 n7143 R=1.199e+02 
R9253t4406 n9254 n4407 R=3.783e+01 
R9253t1138 n9254 n1139 R=4.904e+00 
R9253t3746 n9254 n3747 R=2.846e+00 
R9254t3621 n9255 n3622 R=1.884e+01 
R9254t8402 n9255 n8403 R=5.121e+00 
R9254t6718 n9255 n6719 R=4.378e+00 
R9254t6643 n9255 n6644 R=4.262e+00 
R9254t8564 n9255 n8565 R=3.976e+02 
R9254t4039 n9255 n4040 R=3.989e+00 
R9255t6182 n9256 n6183 R=6.970e+00 
R9255t8595 n9256 n8596 R=4.404e+00 
R9255t7306 n9256 n7307 R=2.863e+00 
R9255t1594 n9256 n1595 R=2.072e+01 
R9255t9199 n9256 n9200 R=1.380e+01 
R9255t926 n9256 n927 R=1.906e+01 
R9256t3940 n9257 n3941 R=3.328e+00 
R9256t7174 n9257 n7175 R=9.114e+00 
R9256t2345 n9257 n2346 R=4.876e+00 
R9256t7948 n9257 n7949 R=2.362e+01 
R9256t5128 n9257 n5129 R=6.788e+00 
R9256t1875 n9257 n1876 R=2.595e+02 
R9257t7929 n9258 n7930 R=6.375e+00 
R9257t8122 n9258 n8123 R=5.050e+00 
R9257t2400 n9258 n2401 R=1.824e+01 
R9257t1316 n9258 n1317 R=5.356e+00 
R9257t162 n9258 n163 R=7.814e+00 
R9257t2751 n9258 n2752 R=1.455e+01 
R9258t3883 n9259 n3884 R=8.659e+00 
R9258t4185 n9259 n4186 R=6.680e+00 
R9258t4191 n9259 n4192 R=1.552e+02 
R9258t2456 n9259 n2457 R=1.631e+01 
R9258t8408 n9259 n8409 R=8.167e+00 
R9258t466 n9259 n467 R=4.098e+00 
R9259t3921 n9260 n3922 R=3.228e+00 
R9259t5117 n9260 n5118 R=5.028e+00 
R9259t8870 n9260 n8871 R=2.553e+00 
R9260t2758 n9261 n2759 R=1.788e+01 
R9260t7867 n9261 n7868 R=4.910e+00 
R9260t4892 n9261 n4893 R=3.910e+01 
R9260t2819 n9261 n2820 R=5.691e+00 
R9260t4121 n9261 n4122 R=8.753e+00 
R9260t1196 n9261 n1197 R=9.728e+00 
R9261t6004 n9262 n6005 R=5.682e+00 
R9261t6415 n9262 n6416 R=3.582e+00 
R9261t2364 n9262 n2365 R=3.851e+00 
R9261t3018 n9262 n3019 R=9.532e+00 
R9262t1167 n9263 n1168 R=7.553e+01 
R9262t2467 n9263 n2468 R=1.656e+01 
R9262t1854 n9263 n1855 R=6.434e+00 
R9262t6596 n9263 n6597 R=6.601e+00 
R9262t4056 n9263 n4057 R=1.755e+01 
R9262t6547 n9263 n6548 R=1.692e+01 
R9262t5573 n9263 n5574 R=5.145e+00 
R9263t3276 n9264 n3277 R=5.827e+00 
R9263t3374 n9264 n3375 R=5.963e+00 
R9263t1664 n9264 n1665 R=5.610e+00 
R9263t4709 n9264 n4710 R=3.023e+02 
R9263t4516 n9264 n4517 R=2.190e+00 
R9264t5464 n9265 n5465 R=1.442e+01 
R9264t7462 n9265 n7463 R=3.567e+00 
R9264t4113 n9265 n4114 R=1.469e+01 
R9264t4155 n9265 n4156 R=2.205e+00 
R9265t188 n9266 n189 R=1.063e+01 
R9265t428 n9266 n429 R=6.325e+00 
R9265t856 n9266 n857 R=5.567e+00 
R9265t4598 n9266 n4599 R=7.701e+00 
R9265t4640 n9266 n4641 R=4.019e+02 
R9265t6692 n9266 n6693 R=5.334e+00 
R9265t7202 n9266 n7203 R=1.311e+02 
R9266t4543 n9267 n4544 R=2.614e+00 
R9266t6321 n9267 n6322 R=5.943e+01 
R9266t524 n9267 n525 R=2.240e+00 
R9266t2896 n9267 n2897 R=3.897e+01 
R9266t5449 n9267 n5450 R=6.661e+00 
R9267t4706 n9268 n4707 R=1.187e+01 
R9267t8818 n9268 n8819 R=1.883e+01 
R9267t890 n9268 n891 R=5.189e+02 
R9267t5690 n9268 n5691 R=4.031e+00 
R9267t260 n9268 n261 R=3.334e+01 
R9267t3684 n9268 n3685 R=1.039e+01 
R9268t2337 n9269 n2338 R=6.042e+00 
R9268t2774 n9269 n2775 R=1.371e+01 
R9268t1498 n9269 n1499 R=8.640e+00 
R9268t7962 n9269 n7963 R=8.424e+00 
R9268t6836 n9269 n6837 R=1.213e+01 
R9268t5689 n9269 n5690 R=1.593e+01 
R9269t4039 n9270 n4040 R=2.560e+00 
R9269t6443 n9270 n6444 R=2.208e+01 
R9269t3872 n9270 n3873 R=3.038e+00 
R9269t5294 n9270 n5295 R=1.448e+01 
R9270t2886 n9271 n2887 R=2.189e+01 
R9270t7277 n9271 n7278 R=4.901e+00 
R9270t7320 n9271 n7321 R=4.612e+00 
R9270t4611 n9271 n4612 R=1.135e+01 
R9270t8078 n9271 n8079 R=1.342e+01 
R9270t4886 n9271 n4887 R=8.216e+00 
R9271t2390 n9272 n2391 R=1.876e+02 
R9271t8883 n9272 n8884 R=1.735e+01 
R9271t6458 n9272 n6459 R=3.545e+01 
R9271t153 n9272 n154 R=5.059e+00 
R9271t4752 n9272 n4753 R=1.406e+02 
R9271t8606 n9272 n8607 R=3.220e+00 
R9271t556 n9272 n557 R=3.321e+01 
R9271t8325 n9272 n8326 R=4.208e+00 
R9272t1048 n9273 n1049 R=5.861e+02 
R9272t7677 n9273 n7678 R=6.169e+00 
R9272t3778 n9273 n3779 R=7.160e+01 
R9272t6353 n9273 n6354 R=9.157e+00 
R9272t4252 n9273 n4253 R=5.640e+00 
R9272t6197 n9273 n6198 R=2.595e+01 
R9272t6703 n9273 n6704 R=3.455e+00 
R9273t4354 n9274 n4355 R=3.583e+00 
R9273t6896 n9274 n6897 R=8.220e+00 
R9273t3776 n9274 n3777 R=6.346e+01 
R9273t7995 n9274 n7996 R=1.944e+00 
R9273t4637 n9274 n4638 R=2.477e+01 
R9274t4151 n9275 n4152 R=3.127e+01 
R9274t5452 n9275 n5453 R=2.139e+01 
R9274t2585 n9275 n2586 R=6.381e+00 
R9274t5087 n9275 n5088 R=4.708e+00 
R9274t965 n9275 n966 R=1.504e+02 
R9274t1533 n9275 n1534 R=1.252e+01 
R9274t7879 n9275 n7880 R=5.341e+00 
R9274t237 n9275 n238 R=2.405e+01 
R9275t575 n9276 n576 R=2.511e+00 
R9275t6029 n9276 n6030 R=1.365e+01 
R9275t4130 n9276 n4131 R=1.863e+01 
R9275t2532 n9276 n2533 R=3.027e+00 
R9275t7744 n9276 n7745 R=1.551e+01 
R9275t977 n9276 n978 R=1.695e+01 
R9276t973 n9277 n974 R=1.520e+00 
R9276t3733 n9277 n3734 R=1.754e+01 
R9276t5961 n9277 n5962 R=1.368e+01 
R9276t2396 n9277 n2397 R=2.707e+00 
R9277t7025 n9278 n7026 R=2.824e+00 
R9277t7397 n9278 n7398 R=1.727e+01 
R9277t6380 n9278 n6381 R=4.161e+00 
R9278t226 n9279 n227 R=7.945e+01 
R9278t1026 n9279 n1027 R=3.956e+00 
R9278t3065 n9279 n3066 R=5.139e+00 
R9278t1892 n9279 n1893 R=6.752e+00 
R9278t8722 n9279 n8723 R=1.019e+02 
R9279t3968 n9280 n3969 R=2.549e+01 
R9279t4451 n9280 n4452 R=3.463e+00 
R9279t3349 n9280 n3350 R=4.147e+00 
R9280t2 n9281 n3 R=3.166e+00 
R9280t4784 n9281 n4785 R=7.513e+00 
R9280t3086 n9281 n3087 R=7.136e+00 
R9280t7407 n9281 n7408 R=5.459e+00 
R9281t6090 n9282 n6091 R=3.672e+00 
R9281t8791 n9282 n8792 R=1.012e+02 
R9281t6345 n9282 n6346 R=4.344e+01 
R9281t7351 n9282 n7352 R=7.336e+00 
R9281t6445 n9282 n6446 R=4.410e+00 
R9282t211 n9283 n212 R=5.401e+00 
R9282t8490 n9283 n8491 R=1.268e+01 
R9282t808 n9283 n809 R=6.739e+00 
R9282t4064 n9283 n4065 R=3.351e+00 
R9282t7997 n9283 n7998 R=2.021e+01 
R9282t1509 n9283 n1510 R=2.466e+01 
R9283t2616 n9284 n2617 R=7.857e+00 
R9283t7408 n9284 n7409 R=4.694e+01 
R9283t3771 n9284 n3772 R=9.490e+00 
R9283t5703 n9284 n5704 R=7.759e+00 
R9283t4917 n9284 n4918 R=5.801e+00 
R9283t1600 n9284 n1601 R=1.019e+01 
R9283t7619 n9284 n7620 R=1.250e+01 
R9284t2507 n9285 n2508 R=1.087e+01 
R9284t2625 n9285 n2626 R=9.744e+00 
R9284t1947 n9285 n1948 R=5.124e+00 
R9284t2818 n9285 n2819 R=2.228e+02 
R9284t3600 n9285 n3601 R=1.067e+01 
R9284t1570 n9285 n1571 R=8.812e+00 
R9285t8742 n9286 n8743 R=6.001e+01 
R9285t8886 n9286 n8887 R=1.721e+01 
R9285t2039 n9286 n2040 R=1.757e+01 
R9285t3839 n9286 n3840 R=8.254e+00 
R9285t9136 n9286 n9137 R=3.882e+00 
R9285t203 n9286 n204 R=1.094e+01 
R9285t7967 n9286 n7968 R=3.650e+00 
R9286t3583 n9287 n3584 R=3.653e+01 
R9286t5881 n9287 n5882 R=4.879e+01 
R9286t6410 n9287 n6411 R=2.238e+00 
R9286t4937 n9287 n4938 R=8.597e+00 
R9286t7519 n9287 n7520 R=2.232e+02 
R9286t5244 n9287 n5245 R=1.809e+00 
R9287t5850 n9288 n5851 R=3.197e+01 
R9287t6893 n9288 n6894 R=1.609e+02 
R9287t6267 n9288 n6268 R=4.973e+01 
R9287t7449 n9288 n7450 R=2.127e+00 
R9287t3302 n9288 n3303 R=2.319e+02 
R9287t4249 n9288 n4250 R=2.420e+01 
R9287t6685 n9288 n6686 R=4.451e+00 
R9287t5603 n9288 n5604 R=2.663e+01 
R9287t4765 n9288 n4766 R=5.644e+00 
R9287t4823 n9288 n4824 R=5.752e+01 
R9288t871 n9289 n872 R=4.555e+00 
R9288t8844 n9289 n8845 R=1.376e+01 
R9288t69 n9289 n70 R=1.162e+01 
R9288t3791 n9289 n3792 R=5.746e+00 
R9288t194 n9289 n195 R=7.415e+00 
R9288t8478 n9289 n8479 R=8.971e+00 
R9288t5208 n9289 n5209 R=9.612e+01 
R9289t8501 n9290 n8502 R=1.429e+02 
R9289t3149 n9290 n3150 R=5.507e+00 
R9289t7329 n9290 n7330 R=1.251e+01 
R9289t8036 n9290 n8037 R=7.889e+00 
R9289t9101 n9290 n9102 R=1.044e+01 
R9289t1047 n9290 n1048 R=4.328e+00 
R9290t5450 n9291 n5451 R=4.869e+00 
R9290t5542 n9291 n5543 R=4.675e+00 
R9290t6607 n9291 n6608 R=2.661e+00 
R9290t4914 n9291 n4915 R=6.905e+00 
R9291t7263 n9292 n7264 R=1.185e+01 
R9291t9234 n9292 n9235 R=5.480e+00 
R9291t2361 n9292 n2362 R=1.733e+01 
R9291t7859 n9292 n7860 R=1.270e+01 
R9291t7708 n9292 n7709 R=6.611e+00 
R9291t3958 n9292 n3959 R=2.164e+01 
R9291t6817 n9292 n6818 R=1.227e+01 
R9291t5625 n9292 n5626 R=9.310e+00 
R9292t179 n9293 n180 R=5.214e+01 
R9292t6364 n9293 n6365 R=5.586e+00 
R9292t1541 n9293 n1542 R=5.332e+00 
R9292t8729 n9293 n8730 R=3.538e+00 
R9292t5999 n9293 n6000 R=8.723e+01 
R9292t236 n9293 n237 R=9.413e+00 
R9293t4410 n9294 n4411 R=4.353e+00 
R9293t7314 n9294 n7315 R=3.366e+01 
R9293t7154 n9294 n7155 R=7.206e+00 
R9293t7243 n9294 n7244 R=1.702e+01 
R9293t5356 n9294 n5357 R=1.566e+00 
R9293t3998 n9294 n3999 R=7.116e+01 
R9294t8277 n9295 n8278 R=2.831e+01 
R9294t8699 n9295 n8700 R=3.509e+01 
R9294t6411 n9295 n6412 R=2.827e+00 
R9294t7498 n9295 n7499 R=9.066e+00 
R9294t616 n9295 n617 R=1.623e+01 
R9294t2413 n9295 n2414 R=2.231e+00 
R9295t3427 n9296 n3428 R=1.895e+01 
R9295t4431 n9296 n4432 R=4.933e+00 
R9295t945 n9296 n946 R=5.076e+00 
R9295t3038 n9296 n3039 R=8.695e+00 
R9295t703 n9296 n704 R=7.943e+00 
R9295t9140 n9296 n9141 R=9.499e+00 
R9296t1090 n9297 n1091 R=9.338e+00 
R9296t8773 n9297 n8774 R=3.197e+00 
R9297t6511 n9298 n6512 R=2.989e+00 
R9297t8350 n9298 n8351 R=7.434e+00 
R9297t6379 n9298 n6380 R=1.133e+01 
R9297t7620 n9298 n7621 R=4.525e+00 
R9297t550 n9298 n551 R=1.228e+01 
R9297t7305 n9298 n7306 R=1.195e+02 
R9298t5565 n9299 n5566 R=3.849e+00 
R9298t7057 n9299 n7058 R=1.089e+01 
R9298t8404 n9299 n8405 R=1.175e+01 
R9298t1923 n9299 n1924 R=7.290e+00 
R9298t8710 n9299 n8711 R=9.039e+00 
R9298t2012 n9299 n2013 R=1.767e+01 
R9298t3464 n9299 n3465 R=2.100e+01 
R9298t7284 n9299 n7285 R=1.880e+01 
R9299t891 n9300 n892 R=1.134e+01 
R9299t6999 n9300 n7000 R=5.419e+00 
R9299t2435 n9300 n2436 R=1.445e+01 
R9299t7224 n9300 n7225 R=3.760e+00 
R9300t2926 n9301 n2927 R=4.501e+00 
R9300t5364 n9301 n5365 R=6.994e+00 
R9300t6495 n9301 n6496 R=5.193e+00 
R9300t9036 n9301 n9037 R=2.835e+01 
R9301t684 n9302 n685 R=2.663e+00 
R9301t8535 n9302 n8536 R=3.838e+02 
R9301t5985 n9302 n5986 R=3.754e+00 
R9301t553 n9302 n554 R=1.026e+01 
R9301t3481 n9302 n3482 R=5.424e+01 
R9301t8808 n9302 n8809 R=5.358e+00 
R9302t1679 n9303 n1680 R=7.347e+00 
R9302t6976 n9303 n6977 R=3.601e+00 
R9302t6995 n9303 n6996 R=9.770e+00 
R9302t8486 n9303 n8487 R=2.035e+00 
R9302t154 n9303 n155 R=5.800e+01 
R9303t3221 n9304 n3222 R=9.262e+00 
R9303t5500 n9304 n5501 R=2.998e+00 
R9303t7575 n9304 n7576 R=2.656e+01 
R9303t809 n9304 n810 R=8.385e+01 
R9303t5123 n9304 n5124 R=5.934e+00 
R9303t2521 n9304 n2522 R=5.216e+00 
R9304t51 n9305 n52 R=4.100e+01 
R9304t6667 n9305 n6668 R=1.772e+01 
R9304t3409 n9305 n3410 R=1.797e+00 
R9304t1463 n9305 n1464 R=1.839e+01 
R9304t8130 n9305 n8131 R=1.172e+01 
R9304t4825 n9305 n4826 R=3.884e+00 
R9305t3997 n9306 n3998 R=6.641e+00 
R9305t9022 n9306 n9023 R=2.750e+00 
R9305t680 n9306 n681 R=2.732e+01 
R9305t3528 n9306 n3529 R=1.312e+01 
R9305t3275 n9306 n3276 R=2.353e+00 
R9306t2835 n9307 n2836 R=4.192e+02 
R9306t8411 n9307 n8412 R=4.772e+00 
R9306t3903 n9307 n3904 R=4.746e+00 
R9306t4994 n9307 n4995 R=1.019e+01 
R9306t354 n9307 n355 R=5.302e+01 
R9306t8631 n9307 n8632 R=3.206e+00 
R9306t5875 n9307 n5876 R=1.675e+01 
R9307t6402 n9308 n6403 R=3.116e+00 
R9307t6853 n9308 n6854 R=1.174e+01 
R9307t3257 n9308 n3258 R=4.679e+00 
R9307t8286 n9308 n8287 R=1.077e+01 
R9308t197 n9309 n198 R=8.696e+01 
R9308t4154 n9309 n4155 R=1.477e+01 
R9308t8654 n9309 n8655 R=5.006e+00 
R9308t437 n9309 n438 R=2.592e+01 
R9308t6735 n9309 n6736 R=4.261e+01 
R9308t2693 n9309 n2694 R=3.902e+00 
R9308t4815 n9309 n4816 R=6.216e+01 
R9308t6662 n9309 n6663 R=4.214e+00 
R9309t2021 n9310 n2022 R=4.751e+01 
R9309t8974 n9310 n8975 R=1.914e+01 
R9309t5401 n9310 n5402 R=4.827e+00 
R9309t9036 n9310 n9037 R=8.546e+00 
R9309t2303 n9310 n2304 R=1.612e+00 
R9310t8518 n9311 n8519 R=5.330e+00 
R9310t8683 n9311 n8684 R=9.372e+00 
R9310t212 n9311 n213 R=4.202e+00 
R9310t7456 n9311 n7457 R=1.683e+01 
R9310t3259 n9311 n3260 R=7.297e+02 
R9310t4595 n9311 n4596 R=1.694e+01 
R9310t484 n9311 n485 R=5.818e+00 
R9311t4293 n9312 n4294 R=2.753e+01 
R9311t8578 n9312 n8579 R=2.309e+01 
R9311t7580 n9312 n7581 R=5.353e+00 
R9311t7074 n9312 n7075 R=7.226e+00 
R9311t8572 n9312 n8573 R=5.987e+00 
R9312t80 n9313 n81 R=4.677e+00 
R9312t7632 n9313 n7633 R=1.476e+01 
R9312t2294 n9313 n2295 R=1.611e+01 
R9312t2286 n9313 n2287 R=6.266e+00 
R9312t3038 n9313 n3039 R=4.105e+01 
R9312t945 n9313 n946 R=1.583e+02 
R9312t5567 n9313 n5568 R=7.510e+00 
R9312t4745 n9313 n4746 R=6.057e+00 
R9313t3753 n9314 n3754 R=9.780e+00 
R9313t6812 n9314 n6813 R=2.150e+00 
R9313t8098 n9314 n8099 R=4.194e+00 
R9313t6106 n9314 n6107 R=7.241e+00 
R9314t491 n9315 n492 R=4.941e+00 
R9314t6173 n9315 n6174 R=1.896e+02 
R9314t7670 n9315 n7671 R=7.962e+00 
R9314t6629 n9315 n6630 R=1.578e+01 
R9314t3106 n9315 n3107 R=1.548e+01 
R9314t5010 n9315 n5011 R=3.260e+00 
R9314t526 n9315 n527 R=1.546e+01 
R9315t2362 n9316 n2363 R=2.486e+00 
R9315t2436 n9316 n2437 R=9.973e+00 
R9315t8308 n9316 n8309 R=6.546e+00 
R9315t6034 n9316 n6035 R=3.965e+00 
R9315t4577 n9316 n4578 R=1.432e+01 
R9315t2803 n9316 n2804 R=4.862e+01 
R9316t3292 n9317 n3293 R=3.872e+00 
R9316t5942 n9317 n5943 R=2.336e+02 
R9316t4817 n9317 n4818 R=2.127e+01 
R9316t6552 n9317 n6553 R=7.014e+00 
R9316t5032 n9317 n5033 R=1.828e+00 
R9316t2659 n9317 n2660 R=2.569e+01 
R9317t280 n9318 n281 R=2.201e+00 
R9317t1595 n9318 n1596 R=2.648e+01 
R9317t7049 n9318 n7050 R=2.405e+01 
R9317t2094 n9318 n2095 R=1.154e+02 
R9317t5126 n9318 n5127 R=2.321e+00 
R9317t3447 n9318 n3448 R=7.774e+00 
R9318t2019 n9319 n2020 R=1.445e+01 
R9318t3276 n9319 n3277 R=1.139e+01 
R9318t6546 n9319 n6547 R=4.730e+00 
R9318t7075 n9319 n7076 R=1.499e+01 
R9318t5959 n9319 n5960 R=8.959e+00 
R9318t5619 n9319 n5620 R=9.269e+00 
R9318t6389 n9319 n6390 R=3.936e+01 
R9319t4242 n9320 n4243 R=7.559e+01 
R9319t7158 n9320 n7159 R=5.020e+00 
R9319t8768 n9320 n8769 R=5.935e+01 
R9319t7687 n9320 n7688 R=3.538e+00 
R9319t6562 n9320 n6563 R=2.194e+01 
R9319t1432 n9320 n1433 R=6.701e+00 
R9319t4537 n9320 n4538 R=7.007e+01 
R9319t1043 n9320 n1044 R=6.576e+00 
R9320t2488 n9321 n2489 R=3.635e+00 
R9320t8881 n9321 n8882 R=4.098e+00 
R9320t2195 n9321 n2196 R=3.387e+02 
R9320t4596 n9321 n4597 R=5.496e+00 
R9320t3370 n9321 n3371 R=2.766e+01 
R9320t5753 n9321 n5754 R=1.026e+01 
R9321t2760 n9322 n2761 R=8.802e+00 
R9321t3718 n9322 n3719 R=1.578e+01 
R9321t7213 n9322 n7214 R=9.542e+00 
R9321t330 n9322 n331 R=6.601e+00 
R9321t2215 n9322 n2216 R=5.548e+00 
R9321t9082 n9322 n9083 R=6.369e+02 
R9321t1756 n9322 n1757 R=3.308e+01 
R9321t4615 n9322 n4616 R=7.661e+00 
R9322t2394 n9323 n2395 R=1.137e+01 
R9322t5429 n9323 n5430 R=2.290e+00 
R9322t218 n9323 n219 R=9.084e+00 
R9323t1871 n9324 n1872 R=5.946e+00 
R9323t7006 n9324 n7007 R=4.689e+02 
R9323t1309 n9324 n1310 R=5.557e+00 
R9323t2889 n9324 n2890 R=4.647e+00 
R9323t1101 n9324 n1102 R=1.422e+01 
R9323t8414 n9324 n8415 R=8.570e+00 
R9324t6368 n1 n6369 R=2.175e+02 
R9325t5852 n9326 n5853 R=2.039e+02 
R9325t6690 n9326 n6691 R=3.121e+00 
R9325t5312 n9326 n5313 R=4.429e+02 
R9325t3636 n9326 n3637 R=6.027e+00 
R9325t2637 n9326 n2638 R=1.161e+01 
R9325t5837 n9326 n5838 R=2.329e+02 
R9325t2748 n9326 n2749 R=1.025e+01 
R9326t2507 n9327 n2508 R=1.335e+02 
R9326t3768 n9327 n3769 R=5.839e+00 
R9326t5636 n9327 n5637 R=1.167e+01 
R9326t1202 n9327 n1203 R=9.010e+00 
R9326t2371 n9327 n2372 R=3.582e+02 
R9326t267 n9327 n268 R=2.171e+00 
R9326t2993 n9327 n2994 R=2.207e+01 
R9327t4932 n9328 n4933 R=7.093e+00 
R9327t1329 n9328 n1330 R=3.254e+01 
R9327t5572 n9328 n5573 R=9.058e+00 
R9328t1641 n9329 n1642 R=2.984e+00 
R9328t1852 n9329 n1853 R=2.658e+01 
R9328t2394 n9329 n2395 R=1.956e+01 
R9328t8733 n9329 n8734 R=2.817e+01 
R9328t5711 n9329 n5712 R=1.816e+00 
R9328t5768 n9329 n5769 R=2.316e+01 
R9329t1155 n9330 n1156 R=4.063e+02 
R9329t4569 n9330 n4570 R=1.234e+01 
R9329t2232 n9330 n2233 R=4.946e+00 
R9329t4789 n9330 n4790 R=5.871e+00 
R9329t7226 n9330 n7227 R=4.764e+00 
R9330t2858 n9331 n2859 R=2.010e+01 
R9330t3436 n9331 n3437 R=5.083e+00 
R9330t7613 n9331 n7614 R=8.722e+00 
R9330t935 n9331 n936 R=3.991e+00 
R9331t3115 n9332 n3116 R=6.696e+00 
R9331t9088 n9332 n9089 R=1.440e+01 
R9331t5970 n9332 n5971 R=2.668e+00 
R9331t1370 n9332 n1371 R=4.010e+00 
R9331t2183 n9332 n2184 R=1.741e+01 
R9332t6590 n9333 n6591 R=3.290e+00 
R9332t6614 n9333 n6615 R=1.476e+02 
R9332t6969 n9333 n6970 R=4.095e+00 
R9332t2288 n9333 n2289 R=7.592e+00 
R9332t3533 n9333 n3534 R=4.421e+00 
R9332t9252 n9333 n9253 R=2.401e+01 
R9333t809 n9334 n810 R=2.013e+01 
R9333t8738 n9334 n8739 R=3.714e+00 
R9333t3949 n9334 n3950 R=1.295e+03 
R9333t3191 n9334 n3192 R=9.674e+00 
R9333t8280 n9334 n8281 R=8.532e+00 
R9333t7575 n9334 n7576 R=7.627e+00 
R9334t2510 n9335 n2511 R=5.935e+00 
R9334t6339 n9335 n6340 R=9.470e+00 
R9334t56 n9335 n57 R=4.094e+00 
R9334t975 n9335 n976 R=4.148e+00 
R9335t3914 n9336 n3915 R=2.972e+00 
R9335t5215 n9336 n5216 R=6.513e+00 
R9336t5215 n9337 n5216 R=3.277e+01 
R9336t9335 n9337 n9336 R=1.286e+00 
R9336t892 n9337 n893 R=2.894e+01 
R9336t1317 n9337 n1318 R=2.108e+00 
R9336t8116 n9337 n8117 R=2.585e+01 
R9336t6795 n9337 n6796 R=2.372e+01 
R9336t3914 n9337 n3915 R=1.326e+01 
R9337t4689 n9338 n4690 R=1.456e+00 
R9337t7386 n9338 n7387 R=1.039e+02 
R9337t6309 n9338 n6310 R=2.294e+00 
R9337t7835 n9338 n7836 R=8.530e+00 
R9337t7616 n9338 n7617 R=5.340e+01 
R9337t9043 n9338 n9044 R=1.959e+01 
R9338t3307 n9339 n3308 R=9.082e+00 
R9338t8320 n9339 n8321 R=1.309e+01 
R9338t453 n9339 n454 R=4.806e+00 
R9338t4918 n9339 n4919 R=6.711e+00 
R9338t8668 n9339 n8669 R=5.239e+00 
R9338t4682 n9339 n4683 R=2.565e+02 
R9339t6190 n9340 n6191 R=5.270e+00 
R9339t9049 n9340 n9050 R=4.289e+01 
R9339t248 n9340 n249 R=2.197e+01 
R9339t4233 n9340 n4234 R=4.121e+00 
R9339t8826 n9340 n8827 R=3.887e+00 
R9340t64 n9341 n65 R=4.419e+01 
R9340t3072 n9341 n3073 R=3.376e+00 
R9340t9014 n9341 n9015 R=3.923e+00 
R9340t4019 n9341 n4020 R=6.028e+00 
R9340t5375 n9341 n5376 R=8.761e+00 
R9341t504 n9342 n505 R=1.832e+01 
R9341t792 n9342 n793 R=1.005e+01 
R9341t1867 n9342 n1868 R=3.087e+01 
R9341t8725 n9342 n8726 R=3.986e+00 
R9341t591 n9342 n592 R=5.465e+00 
R9341t3510 n9342 n3511 R=2.418e+01 
R9341t3351 n9342 n3352 R=7.328e+00 
R9341t4708 n9342 n4709 R=1.515e+01 
R9342t5117 n9343 n5118 R=5.480e+00 
R9342t8620 n9343 n8621 R=7.795e+00 
R9342t8807 n9343 n8808 R=5.065e+00 
R9342t7548 n9343 n7549 R=4.622e+00 
R9343t3170 n9344 n3171 R=7.303e+00 
R9343t7473 n9344 n7474 R=8.322e+00 
R9343t573 n9344 n574 R=6.866e+00 
R9343t8966 n9344 n8967 R=2.610e+01 
R9343t1818 n9344 n1819 R=2.777e+00 
R9344t2169 n9345 n2170 R=7.324e+00 
R9344t8129 n9345 n8130 R=5.377e+01 
R9344t505 n9345 n506 R=2.797e+01 
R9344t1753 n9345 n1754 R=2.611e+00 
R9344t5739 n9345 n5740 R=9.724e+00 
R9344t191 n9345 n192 R=3.281e+01 
R9344t3646 n9345 n3647 R=1.904e+02 
R9344t4923 n9345 n4924 R=4.137e+02 
R9344t4334 n9345 n4335 R=8.628e+00 
R9344t5199 n9345 n5200 R=3.852e+00 
R9345t2157 n9346 n2158 R=1.002e+01 
R9345t6080 n9346 n6081 R=5.685e+00 
R9345t946 n9346 n947 R=7.735e+00 
R9345t954 n9346 n955 R=2.826e+01 
R9345t3016 n9346 n3017 R=2.012e+02 
R9345t4706 n9346 n4707 R=7.747e+00 
R9345t1137 n9346 n1138 R=5.609e+00 
R9346t4138 n9347 n4139 R=9.229e+00 
R9346t4344 n9347 n4345 R=3.467e+00 
R9346t2523 n9347 n2524 R=8.157e+00 
R9346t8507 n9347 n8508 R=8.179e+00 
R9346t804 n9347 n805 R=8.344e+00 
R9346t228 n9347 n229 R=7.101e+00 
R9347t1971 n9348 n1972 R=2.318e+01 
R9347t9083 n9348 n9084 R=8.509e+00 
R9347t7244 n9348 n7245 R=5.369e+00 
R9348t3792 n9349 n3793 R=4.053e+00 
R9348t6492 n9349 n6493 R=2.552e+01 
R9348t414 n9349 n415 R=1.722e+03 
R9348t6388 n9349 n6389 R=2.810e+00 
R9348t8826 n9349 n8827 R=8.536e+00 
R9348t4539 n9349 n4540 R=2.556e+01 
R9348t6491 n9349 n6492 R=8.414e+00 
R9349t2020 n9350 n2021 R=1.200e+01 
R9349t3005 n9350 n3006 R=1.770e+01 
R9349t8815 n9350 n8816 R=3.459e+00 
R9349t6170 n9350 n6171 R=3.563e+00 
R9349t6747 n9350 n6748 R=6.363e+00 
R9350t2901 n9351 n2902 R=2.301e+01 
R9350t5405 n9351 n5406 R=4.679e+00 
R9350t6649 n9351 n6650 R=4.390e+00 
R9350t1195 n9351 n1196 R=2.543e+00 
R9351t29 n9352 n30 R=7.773e+01 
R9351t3930 n9352 n3931 R=5.829e+00 
R9351t811 n9352 n812 R=9.946e+00 
R9351t3887 n9352 n3888 R=8.965e+00 
R9351t5297 n9352 n5298 R=3.242e+00 
R9352t2579 n9353 n2580 R=2.261e+01 
R9352t7883 n9353 n7884 R=3.637e+00 
R9352t8676 n9353 n8677 R=1.281e+01 
R9352t5904 n9353 n5905 R=7.823e+00 
R9352t7949 n9353 n7950 R=3.004e+00 
R9352t6786 n9353 n6787 R=2.154e+02 
R9352t8882 n9353 n8883 R=4.146e+01 
R9353t5128 n9354 n5129 R=1.986e+01 
R9353t7948 n9354 n7949 R=1.448e+01 
R9353t4283 n9354 n4284 R=1.794e+01 
R9353t4065 n9354 n4066 R=1.477e+01 
R9353t1207 n9354 n1208 R=2.142e+01 
R9353t5339 n9354 n5340 R=6.074e+00 
R9353t4086 n9354 n4087 R=6.292e+00 
R9353t7341 n9354 n7342 R=2.055e+01 
R9354t2907 n9355 n2908 R=1.042e+01 
R9354t9008 n9355 n9009 R=7.874e+00 
R9354t1505 n9355 n1506 R=1.113e+02 
R9354t4283 n9355 n4284 R=5.463e+01 
R9354t5128 n9355 n5129 R=5.615e+00 
R9354t9256 n9355 n9257 R=1.436e+01 
R9354t1875 n9355 n1876 R=4.002e+00 
R9355t8 n9356 n9 R=7.468e+00 
R9355t9207 n9356 n9208 R=4.294e+00 
R9355t7775 n9356 n7776 R=5.220e+00 
R9355t5324 n9356 n5325 R=4.387e+00 
R9355t3026 n9356 n3027 R=1.809e+02 
R9356t3279 n9357 n3280 R=3.016e+00 
R9356t8430 n9357 n8431 R=6.079e+01 
R9356t928 n9357 n929 R=1.027e+01 
R9356t5093 n9357 n5094 R=2.276e+00 
R9357t2754 n9358 n2755 R=5.257e+00 
R9357t7557 n9358 n7558 R=2.083e+00 
R9357t524 n9358 n525 R=6.768e+00 
R9358t364 n9359 n365 R=8.708e+00 
R9358t7011 n9359 n7012 R=5.308e+00 
R9358t4549 n9359 n4550 R=1.669e+01 
R9358t7652 n9359 n7653 R=3.398e+00 
R9358t7065 n9359 n7066 R=3.958e+00 
R9359t7374 n9360 n7375 R=3.896e+00 
R9359t8557 n9360 n8558 R=5.306e+00 
R9359t1126 n9360 n1127 R=2.407e+00 
R9360t7395 n9361 n7396 R=4.365e+01 
R9360t7860 n9361 n7861 R=5.291e+00 
R9360t3229 n9361 n3230 R=4.694e+00 
R9360t218 n9361 n219 R=2.067e+02 
R9360t6458 n9361 n6459 R=2.131e+02 
R9360t8026 n9361 n8027 R=2.127e+01 
R9361t1107 n9362 n1108 R=1.435e+01 
R9361t7746 n9362 n7747 R=2.938e+00 
R9361t1058 n9362 n1059 R=2.959e+00 
R9361t8301 n9362 n8302 R=1.068e+01 
R9361t2590 n9362 n2591 R=1.861e+01 
R9361t7840 n9362 n7841 R=6.026e+01 
R9362t4792 n9363 n4793 R=6.675e+00 
R9362t8299 n9363 n8300 R=5.370e+00 
R9362t1612 n9363 n1613 R=8.881e+00 
R9362t8966 n9363 n8967 R=1.101e+01 
R9362t5619 n9363 n5620 R=1.696e+01 
R9362t6797 n9363 n6798 R=1.030e+01 
R9362t4220 n9363 n4221 R=1.372e+01 
R9363t4212 n9364 n4213 R=1.342e+01 
R9363t5643 n9364 n5644 R=2.211e+01 
R9363t4294 n9364 n4295 R=7.587e+00 
R9363t7089 n9364 n7090 R=8.163e+00 
R9363t8843 n9364 n8844 R=7.742e+00 
R9363t7166 n9364 n7167 R=5.183e+00 
R9364t297 n9365 n298 R=6.173e+00 
R9364t1494 n9365 n1495 R=3.429e+00 
R9364t6246 n9365 n6247 R=1.645e+01 
R9364t6367 n9365 n6368 R=3.064e+01 
R9364t5003 n9365 n5004 R=6.653e+00 
R9364t4915 n9365 n4916 R=8.320e+00 
R9365t5439 n9366 n5440 R=1.463e+01 
R9365t6359 n9366 n6360 R=5.728e+00 
R9365t5860 n9366 n5861 R=3.614e+00 
R9365t4386 n9366 n4387 R=5.074e+00 
R9365t1973 n9366 n1974 R=1.170e+01 
R9366t4528 n9367 n4529 R=4.480e+00 
R9366t8814 n9367 n8815 R=7.802e+00 
R9366t2500 n9367 n2501 R=8.929e+00 
R9366t3209 n9367 n3210 R=4.146e+00 
R9366t460 n9367 n461 R=7.932e+01 
R9367t1870 n9368 n1871 R=3.601e+00 
R9367t4135 n9368 n4136 R=6.669e+00 
R9367t8293 n9368 n8294 R=1.210e+01 
R9367t6228 n9368 n6229 R=4.789e+00 
R9367t5292 n9368 n5293 R=2.679e+01 
R9367t8632 n9368 n8633 R=3.089e+01 
R9368t1602 n9369 n1603 R=1.058e+02 
R9368t2855 n9369 n2856 R=3.842e+00 
R9368t4957 n9369 n4958 R=2.366e+00 
R9368t2101 n9369 n2102 R=1.416e+01 
R9368t4728 n9369 n4729 R=3.626e+00 
R9369t168 n9370 n169 R=5.381e+01 
R9369t1048 n9370 n1049 R=2.371e+01 
R9369t226 n9370 n227 R=6.087e+00 
R9369t9278 n9370 n9279 R=7.207e+00 
R9369t8722 n9370 n8723 R=4.619e+00 
R9369t1218 n9370 n1219 R=1.183e+01 
R9369t746 n9370 n747 R=1.262e+01 
R9370t561 n9371 n562 R=2.342e+02 
R9370t1534 n9371 n1535 R=6.037e+00 
R9370t7495 n9371 n7496 R=7.520e+00 
R9370t3299 n9371 n3300 R=9.063e+00 
R9370t4315 n9371 n4316 R=3.650e+00 
R9371t1411 n9372 n1412 R=2.411e+00 
R9371t4070 n9372 n4071 R=1.152e+01 
R9371t7951 n9372 n7952 R=1.229e+02 
R9371t7684 n9372 n7685 R=3.328e+01 
R9371t1001 n9372 n1002 R=3.545e+00 
R9371t6292 n9372 n6293 R=1.237e+01 
R9372t1217 n9373 n1218 R=2.224e+00 
R9372t7546 n9373 n7547 R=4.180e+01 
R9372t8508 n9373 n8509 R=1.060e+01 
R9372t4300 n9373 n4301 R=5.180e+01 
R9372t956 n9373 n957 R=4.219e+00 
R9372t6772 n9373 n6773 R=3.890e+00 
R9373t4549 n9374 n4550 R=1.240e+02 
R9373t6299 n9374 n6300 R=1.534e+01 
R9373t7135 n9374 n7136 R=5.377e+00 
R9373t797 n9374 n798 R=1.475e+01 
R9373t518 n9374 n519 R=7.161e+00 
R9373t6745 n9374 n6746 R=7.580e+00 
R9373t7011 n9374 n7012 R=2.760e+01 
R9374t115 n9375 n116 R=3.326e+01 
R9374t4190 n9375 n4191 R=1.208e+02 
R9374t2730 n9375 n2731 R=1.157e+01 
R9374t8527 n9375 n8528 R=3.253e+00 
R9374t1566 n9375 n1567 R=7.524e+00 
R9374t7800 n9375 n7801 R=4.309e+00 
R9375t3113 n9376 n3114 R=1.136e+01 
R9375t4793 n9376 n4794 R=4.563e+01 
R9375t5101 n9376 n5102 R=3.301e+00 
R9375t1298 n9376 n1299 R=3.608e+01 
R9375t7087 n9376 n7088 R=1.966e+01 
R9375t249 n9376 n250 R=4.528e+00 
R9376t2465 n9377 n2466 R=5.383e+01 
R9376t6510 n9377 n6511 R=2.408e+00 
R9376t5391 n9377 n5392 R=2.174e+00 
R9376t7107 n9377 n7108 R=9.951e+00 
R9376t8994 n9377 n8995 R=2.543e+01 
R9377t4834 n9378 n4835 R=3.977e+01 
R9377t6898 n9378 n6899 R=5.038e+00 
R9377t685 n9378 n686 R=7.048e+00 
R9377t361 n9378 n362 R=6.762e+00 
R9377t1861 n9378 n1862 R=4.677e+01 
R9377t7685 n9378 n7686 R=1.245e+01 
R9377t9102 n9378 n9103 R=1.049e+02 
R9377t8875 n9378 n8876 R=7.196e+00 
R9378t4450 n9379 n4451 R=5.611e+00 
R9378t9099 n9379 n9100 R=1.008e+01 
R9378t8275 n9379 n8276 R=2.173e+00 
R9378t4143 n9379 n4144 R=1.411e+02 
R9378t5418 n9379 n5419 R=2.477e+01 
R9378t834 n9379 n835 R=4.864e+00 
R9379t4932 n9380 n4933 R=1.501e+01 
R9379t6084 n9380 n6085 R=5.974e+00 
R9379t9327 n9380 n9328 R=3.482e+00 
R9379t1329 n9380 n1330 R=4.519e+01 
R9379t3677 n9380 n3678 R=3.111e+00 
R9379t4088 n9380 n4089 R=2.842e+01 
R9379t7033 n9380 n7034 R=1.863e+01 
R9380t4732 n9381 n4733 R=6.209e+00 
R9380t5965 n9381 n5966 R=2.157e+01 
R9380t3782 n9381 n3783 R=2.881e+01 
R9380t1255 n9381 n1256 R=4.108e+00 
R9380t7096 n9381 n7097 R=1.650e+01 
R9380t8156 n9381 n8157 R=4.942e+00 
R9381t3544 n9382 n3545 R=1.048e+01 
R9381t8142 n9382 n8143 R=3.914e+01 
R9381t7812 n9382 n7813 R=9.771e+00 
R9381t9225 n9382 n9226 R=5.408e+00 
R9381t5258 n9382 n5259 R=3.472e+00 
R9382t3530 n9383 n3531 R=2.095e+01 
R9382t3594 n9383 n3595 R=1.479e+01 
R9382t8923 n9383 n8924 R=6.966e+00 
R9382t8328 n9383 n8329 R=5.254e+00 
R9382t8771 n9383 n8772 R=1.283e+01 
R9382t7941 n9383 n7942 R=2.214e+01 
R9382t1804 n9383 n1805 R=4.759e+00 
R9383t5426 n9384 n5427 R=2.391e+00 
R9383t7182 n9384 n7183 R=3.691e+01 
R9383t5257 n9384 n5258 R=1.602e+00 
R9383t5888 n9384 n5889 R=2.218e+01 
R9383t6487 n9384 n6488 R=1.082e+01 
R9384t663 n9385 n664 R=1.827e+01 
R9384t2940 n9385 n2941 R=1.398e+01 
R9384t3201 n9385 n3202 R=3.293e+00 
R9384t1135 n9385 n1136 R=2.490e+01 
R9384t5439 n9385 n5440 R=3.862e+01 
R9384t5860 n9385 n5861 R=2.553e+00 
R9385t8094 n9386 n8095 R=3.606e+00 
R9385t8449 n9386 n8450 R=5.366e+01 
R9385t7379 n9386 n7380 R=5.173e+01 
R9385t540 n9386 n541 R=1.178e+01 
R9385t2640 n9386 n2641 R=8.645e+00 
R9385t2769 n9386 n2770 R=2.576e+00 
R9386t2140 n9387 n2141 R=2.088e+01 
R9386t2407 n9387 n2408 R=1.300e+02 
R9386t3264 n9387 n3265 R=1.495e+01 
R9386t2075 n9387 n2076 R=4.465e+00 
R9386t210 n9387 n211 R=2.796e+01 
R9386t6345 n9387 n6346 R=1.425e+01 
R9386t9281 n9387 n9282 R=3.547e+00 
R9386t7351 n9387 n7352 R=8.818e+00 
R9387t687 n9388 n688 R=7.686e+00 
R9387t2709 n9388 n2710 R=7.091e+00 
R9387t4646 n9388 n4647 R=1.424e+01 
R9387t6568 n9388 n6569 R=4.173e+00 
R9387t7412 n9388 n7413 R=1.388e+01 
R9387t1380 n9388 n1381 R=7.117e+00 
R9388t4604 n9389 n4605 R=9.757e+00 
R9388t8514 n9389 n8515 R=6.117e+00 
R9388t7717 n9389 n7718 R=2.100e+00 
R9388t4645 n9389 n4646 R=1.561e+01 
R9388t6628 n9389 n6629 R=9.630e+00 
R9388t571 n9389 n572 R=7.556e+00 
R9389t2272 n9390 n2273 R=1.070e+01 
R9389t8965 n9390 n8966 R=4.538e+00 
R9389t1391 n9390 n1392 R=4.020e+00 
R9389t9027 n9390 n9028 R=4.230e+00 
R9390t448 n9391 n449 R=6.688e+00 
R9390t3523 n9391 n3524 R=1.015e+01 
R9390t7268 n9391 n7269 R=1.360e+01 
R9390t1916 n9391 n1917 R=6.326e+00 
R9390t3939 n9391 n3940 R=1.435e+02 
R9390t8021 n9391 n8022 R=2.040e+00 
R9391t2553 n9392 n2554 R=3.273e+00 
R9391t4375 n9392 n4376 R=1.943e+01 
R9391t5993 n9392 n5994 R=1.350e+01 
R9391t1260 n9392 n1261 R=3.554e+00 
R9391t1249 n9392 n1250 R=9.566e+00 
R9392t2671 n9393 n2672 R=2.020e+00 
R9392t8669 n9393 n8670 R=7.778e+00 
R9392t811 n9393 n812 R=2.069e+01 
R9392t9351 n9393 n9352 R=2.293e+02 
R9392t3887 n9393 n3888 R=2.168e+00 
R9392t7362 n9393 n7363 R=6.175e+00 
R9392t3180 n9393 n3181 R=2.154e+02 
R9393t6402 n9394 n6403 R=5.094e+00 
R9393t9307 n9394 n9308 R=1.681e+01 
R9393t44 n9394 n45 R=9.206e+00 
R9393t6673 n9394 n6674 R=1.820e+01 
R9393t8286 n9394 n8287 R=3.733e+00 
R9394t3572 n9395 n3573 R=2.378e+01 
R9394t7942 n9395 n7943 R=1.605e+01 
R9394t5639 n9395 n5640 R=7.525e+00 
R9394t7904 n9395 n7905 R=3.323e+00 
R9394t1571 n9395 n1572 R=2.473e+01 
R9394t7560 n9395 n7561 R=2.384e+00 
R9395t5727 n9396 n5728 R=7.593e+00 
R9395t8419 n9396 n8420 R=7.585e+00 
R9395t5212 n9396 n5213 R=1.028e+01 
R9395t1711 n9396 n1712 R=3.881e+00 
R9396t1315 n9397 n1316 R=1.751e+01 
R9396t7892 n9397 n7893 R=3.794e+02 
R9396t1698 n9397 n1699 R=4.790e+00 
R9396t9189 n9397 n9190 R=4.057e+00 
R9396t8264 n9397 n8265 R=7.716e+00 
R9397t7964 n9398 n7965 R=1.022e+01 
R9397t8600 n9398 n8601 R=3.935e+00 
R9397t9175 n9398 n9176 R=3.817e+00 
R9397t1375 n9398 n1376 R=8.884e+00 
R9398t2269 n9399 n2270 R=1.499e+01 
R9398t3123 n9399 n3124 R=6.815e+00 
R9398t1055 n9399 n1056 R=3.514e+01 
R9398t3360 n9399 n3361 R=2.367e+00 
R9398t8529 n9399 n8530 R=5.282e+03 
R9398t8580 n9399 n8581 R=4.993e+00 
R9399t982 n9400 n983 R=2.123e+01 
R9399t1568 n9400 n1569 R=8.228e+00 
R9399t7435 n9400 n7436 R=1.636e+01 
R9399t8459 n9400 n8460 R=1.120e+01 
R9399t2188 n9400 n2189 R=9.267e+00 
R9399t6663 n9400 n6664 R=1.387e+01 
R9399t5032 n9400 n5033 R=2.380e+02 
R9399t7001 n9400 n7002 R=3.916e+00 
R9400t5172 n9401 n5173 R=6.082e+00 
R9400t6670 n9401 n6671 R=3.494e+00 
R9400t7770 n9401 n7771 R=2.366e+01 
R9400t2678 n9401 n2679 R=2.898e+00 
R9401t1844 n9402 n1845 R=4.283e+00 
R9401t6419 n9402 n6420 R=1.221e+01 
R9401t4755 n9402 n4756 R=3.702e+00 
R9401t3412 n9402 n3413 R=6.421e+00 
R9401t5012 n9402 n5013 R=2.025e+01 
R9402t784 n9403 n785 R=6.485e+00 
R9402t6163 n9403 n6164 R=4.237e+00 
R9402t4728 n9403 n4729 R=6.948e+00 
R9402t2101 n9403 n2102 R=1.022e+01 
R9402t5897 n9403 n5898 R=2.613e+01 
R9403t1823 n9404 n1824 R=6.691e+00 
R9403t120 n9404 n121 R=4.956e+00 
R9403t4314 n9404 n4315 R=1.841e+01 
R9403t3717 n9404 n3718 R=1.086e+01 
R9404t2276 n9405 n2277 R=9.528e+00 
R9404t6029 n9405 n6030 R=1.252e+01 
R9404t4081 n9405 n4082 R=1.073e+01 
R9404t611 n9405 n612 R=4.145e+00 
R9404t2460 n9405 n2461 R=3.537e+01 
R9404t7094 n9405 n7095 R=1.190e+01 
R9404t4130 n9405 n4131 R=8.123e+00 
R9405t468 n9406 n469 R=2.335e+00 
R9405t6946 n9406 n6947 R=1.015e+02 
R9405t3479 n9406 n3480 R=6.115e+00 
R9405t6031 n9406 n6032 R=2.837e+01 
R9405t1132 n9406 n1133 R=4.018e+00 
R9405t4109 n9406 n4110 R=3.448e+01 
R9406t621 n9407 n622 R=9.977e+00 
R9406t7761 n9407 n7762 R=5.789e+00 
R9406t7177 n9407 n7178 R=4.042e+00 
R9406t6478 n9407 n6479 R=1.558e+01 
R9406t6242 n9407 n6243 R=4.855e+00 
R9406t4676 n9407 n4677 R=2.565e+01 
R9406t4651 n9407 n4652 R=8.350e+01 
R9407t1743 n9408 n1744 R=5.274e+00 
R9407t7849 n9408 n7850 R=5.608e+00 
R9407t1335 n9408 n1336 R=1.032e+01 
R9407t1800 n9408 n1801 R=2.819e+01 
R9407t5594 n9408 n5595 R=1.933e+00 
R9408t1804 n9409 n1805 R=5.510e+00 
R9408t7941 n9409 n7942 R=2.516e+01 
R9408t3530 n9409 n3531 R=7.355e+00 
R9408t3945 n9409 n3946 R=7.601e+00 
R9408t3051 n9409 n3052 R=7.491e+00 
R9408t8347 n9409 n8348 R=2.299e+01 
R9408t5376 n9409 n5377 R=1.334e+01 
R9409t5268 n9410 n5269 R=3.978e+00 
R9409t7376 n9410 n7377 R=1.898e+01 
R9409t4780 n9410 n4781 R=3.769e+00 
R9409t7002 n9410 n7003 R=4.393e+01 
R9409t4567 n9410 n4568 R=3.607e+00 
R9410t1696 n9411 n1697 R=1.291e+01 
R9410t7874 n9411 n7875 R=2.263e+00 
R9410t1047 n9411 n1048 R=1.856e+01 
R9410t9289 n9411 n9290 R=2.805e+01 
R9410t8501 n9411 n8502 R=3.348e+00 
R9410t5046 n9411 n5047 R=4.427e+01 
R9411t1328 n9412 n1329 R=1.224e+01 
R9411t7676 n9412 n7677 R=3.130e+00 
R9411t6855 n9412 n6856 R=7.392e+00 
R9411t2328 n9412 n2329 R=1.000e+01 
R9411t2551 n9412 n2552 R=9.299e+00 
R9411t163 n9412 n164 R=1.546e+01 
R9412t4325 n9413 n4326 R=1.167e+01 
R9412t7852 n9413 n7853 R=2.267e+00 
R9412t493 n9413 n494 R=9.490e+00 
R9412t1185 n9413 n1186 R=7.736e+00 
R9412t2563 n9413 n2564 R=4.484e+01 
R9412t1656 n9413 n1657 R=6.127e+00 
R9413t1327 n9414 n1328 R=1.963e+01 
R9413t3863 n9414 n3864 R=1.534e+01 
R9413t2319 n9414 n2320 R=3.725e+00 
R9413t6807 n9414 n6808 R=4.114e+00 
R9413t5724 n9414 n5725 R=1.460e+01 
R9414t2754 n9415 n2755 R=6.392e+00 
R9414t9357 n9415 n9358 R=6.119e+00 
R9414t5574 n9415 n5575 R=2.306e+01 
R9414t7533 n9415 n7534 R=2.965e+00 
R9414t524 n9415 n525 R=9.769e+00 
R9415t1071 n9416 n1072 R=2.376e+00 
R9415t5141 n9416 n5142 R=1.499e+01 
R9415t2700 n9416 n2701 R=6.026e+00 
R9415t3368 n9416 n3369 R=4.923e+01 
R9415t3640 n9416 n3641 R=1.049e+01 
R9415t2477 n9416 n2478 R=2.601e+01 
R9416t4248 n9417 n4249 R=4.493e+01 
R9416t7348 n9417 n7349 R=2.022e+00 
R9416t4041 n9417 n4042 R=4.218e+00 
R9416t1621 n9417 n1622 R=8.535e+00 
R9416t4987 n9417 n4988 R=8.805e+00 
R9416t1166 n9417 n1167 R=2.583e+01 
R9417t4801 n9418 n4802 R=9.275e+00 
R9417t6146 n9418 n6147 R=4.997e+00 
R9417t2581 n9418 n2582 R=2.494e+00 
R9417t1514 n9418 n1515 R=3.651e+01 
R9417t5210 n9418 n5211 R=4.469e+00 
R9417t1140 n9418 n1141 R=1.054e+02 
R9418t2422 n9419 n2423 R=3.923e+00 
R9418t6523 n9419 n6524 R=1.626e+01 
R9418t7471 n9419 n7472 R=1.424e+02 
R9418t1117 n9419 n1118 R=1.341e+02 
R9418t5555 n9419 n5556 R=1.030e+01 
R9418t4960 n9419 n4961 R=1.057e+01 
R9418t3355 n9419 n3356 R=6.783e+00 
R9419t494 n9420 n495 R=2.666e+00 
R9419t1390 n9420 n1391 R=9.148e+01 
R9419t6732 n9420 n6733 R=7.940e+00 
R9419t5133 n9420 n5134 R=5.343e+00 
R9419t4722 n9420 n4723 R=9.896e+01 
R9419t7026 n9420 n7027 R=7.209e+00 
R9420t6173 n9421 n6174 R=1.839e+01 
R9420t9226 n9421 n9227 R=2.318e+00 
R9420t7043 n9421 n7044 R=4.057e+00 
R9420t3702 n9421 n3703 R=7.408e+00 
R9421t2178 n9422 n2179 R=2.973e+00 
R9421t4590 n9422 n4591 R=1.014e+01 
R9421t287 n9422 n288 R=7.775e+00 
R9421t8938 n9422 n8939 R=7.954e+00 
R9421t7167 n9422 n7168 R=2.395e+01 
R9421t4776 n9422 n4777 R=2.619e+01 
R9422t5576 n9423 n5577 R=8.709e+00 
R9422t8990 n9423 n8991 R=7.584e+01 
R9422t4268 n9423 n4269 R=3.021e+00 
R9422t8937 n9423 n8938 R=8.716e+00 
R9423t5544 n9424 n5545 R=2.899e+01 
R9423t3968 n9424 n3969 R=2.247e+00 
R9423t9279 n9424 n9280 R=5.214e+01 
R9423t7460 n9424 n7461 R=2.392e+01 
R9424t8504 n9425 n8505 R=3.024e+00 
R9424t7071 n9425 n7072 R=1.521e+01 
R9424t5664 n9425 n5665 R=1.192e+01 
R9424t574 n9425 n575 R=8.156e+00 
R9424t1257 n9425 n1258 R=4.534e+00 
R9424t7129 n9425 n7130 R=2.764e+02 
R9425t517 n9426 n518 R=2.032e+00 
R9425t1497 n9426 n1498 R=3.917e+00 
R9426t28 n9427 n29 R=6.504e+00 
R9426t6611 n9427 n6612 R=7.567e+00 
R9426t1230 n9427 n1231 R=1.196e+01 
R9426t8232 n9427 n8233 R=2.164e+00 
R9426t3562 n9427 n3563 R=1.857e+02 
R9426t6951 n9427 n6952 R=1.253e+01 
R9427t1692 n9428 n1693 R=8.101e+00 
R9427t3396 n9428 n3397 R=4.778e+00 
R9427t2765 n9428 n2766 R=1.648e+01 
R9427t7238 n9428 n7239 R=5.992e+00 
R9427t9175 n9428 n9176 R=9.667e+00 
R9428t2149 n9429 n2150 R=2.626e+00 
R9428t8234 n9429 n8235 R=3.206e+00 
R9428t3377 n9429 n3378 R=7.908e+01 
R9429t291 n9430 n292 R=8.031e+01 
R9429t3609 n9430 n3610 R=3.677e+00 
R9429t5700 n9430 n5701 R=1.088e+01 
R9429t8631 n9430 n8632 R=1.121e+02 
R9429t2569 n9430 n2570 R=3.173e+00 
R9429t6281 n9430 n6282 R=1.225e+01 
R9430t3260 n9431 n3261 R=1.187e+01 
R9430t6277 n9431 n6278 R=2.915e+00 
R9430t2604 n9431 n2605 R=4.983e+00 
R9430t3854 n9431 n3855 R=1.608e+01 
R9430t1931 n9431 n1932 R=1.834e+01 
R9430t47 n9431 n48 R=5.604e+00 
R9431t630 n9432 n631 R=3.506e+00 
R9431t1007 n9432 n1008 R=6.461e+01 
R9431t3207 n9432 n3208 R=5.229e+00 
R9431t6998 n9432 n6999 R=4.379e+00 
R9431t8552 n9432 n8553 R=3.578e+02 
R9431t4444 n9432 n4445 R=8.694e+00 
R9432t6908 n9433 n6909 R=3.399e+00 
R9432t3468 n9433 n3469 R=4.383e+01 
R9432t7990 n9433 n7991 R=5.197e+00 
R9432t3183 n9433 n3184 R=5.966e+00 
R9433t5574 n9434 n5575 R=5.314e+00 
R9433t9204 n9434 n9205 R=3.044e+00 
R9433t9154 n9434 n9155 R=5.567e+00 
R9433t7728 n9434 n7729 R=5.586e+00 
R9433t3384 n9434 n3385 R=1.261e+02 
R9434t18 n9435 n19 R=6.419e+00 
R9434t1852 n9435 n1853 R=2.709e+01 
R9434t7316 n9435 n7317 R=9.919e+00 
R9434t218 n9435 n219 R=1.257e+01 
R9434t9322 n9435 n9323 R=3.483e+00 
R9434t2394 n9435 n2395 R=1.489e+02 
R9434t1641 n9435 n1642 R=1.143e+02 
R9435t104 n9436 n105 R=4.212e+00 
R9435t2005 n9436 n2006 R=6.035e+00 
R9435t7269 n9436 n7270 R=1.979e+02 
R9435t4847 n9436 n4848 R=2.307e+01 
R9435t2824 n9436 n2825 R=9.837e+00 
R9435t8208 n9436 n8209 R=5.580e+00 
R9435t159 n9436 n160 R=1.240e+01 
R9435t1291 n9436 n1292 R=2.457e+01 
R9436t4273 n9437 n4274 R=3.499e+00 
R9436t5220 n9437 n5221 R=3.921e+00 
R9436t4760 n9437 n4761 R=1.223e+01 
R9436t1348 n9437 n1349 R=4.785e+00 
R9436t4073 n9437 n4074 R=7.453e+01 
R9437t6496 n9438 n6497 R=8.695e+00 
R9437t7962 n9438 n7963 R=1.515e+01 
R9437t1794 n9438 n1795 R=1.108e+01 
R9437t8480 n9438 n8481 R=5.433e+00 
R9438t4358 n9439 n4359 R=6.690e+02 
R9438t7098 n9439 n7099 R=2.851e+00 
R9438t6734 n9439 n6735 R=2.765e+00 
R9438t2211 n9439 n2212 R=1.152e+01 
R9438t2140 n9439 n2141 R=1.455e+02 
R9438t7579 n9439 n7580 R=8.605e+00 
R9439t4690 n9440 n4691 R=4.335e+00 
R9439t6129 n9440 n6130 R=2.463e+01 
R9439t1374 n9440 n1375 R=1.585e+01 
R9439t68 n9440 n69 R=3.384e+00 
R9440t2453 n9441 n2454 R=3.469e+00 
R9440t7842 n9441 n7843 R=8.053e+00 
R9440t8763 n9441 n8764 R=4.516e+01 
R9440t3616 n9441 n3617 R=1.074e+01 
R9440t9103 n9441 n9104 R=1.566e+01 
R9440t7907 n9441 n7908 R=5.222e+00 
R9441t141 n9442 n142 R=7.196e+00 
R9441t8769 n9442 n8770 R=9.671e+00 
R9441t7690 n9442 n7691 R=5.822e+01 
R9441t3649 n9442 n3650 R=2.656e+00 
R9441t8370 n9442 n8371 R=5.604e+00 
R9442t1798 n9443 n1799 R=1.473e+01 
R9442t3575 n9443 n3576 R=5.896e+00 
R9442t5364 n9443 n5365 R=7.385e+00 
R9442t9300 n9443 n9301 R=8.381e+00 
R9442t6495 n9443 n6496 R=5.555e+00 
R9442t6132 n9443 n6133 R=9.264e+00 
R9443t3062 n9444 n3063 R=5.012e+02 
R9443t5607 n9444 n5608 R=2.151e+01 
R9443t5511 n9444 n5512 R=2.785e+00 
R9443t8636 n9444 n8637 R=6.097e+00 
R9443t5299 n9444 n5300 R=2.713e+01 
R9443t4398 n9444 n4399 R=5.833e+00 
R9443t1502 n9444 n1503 R=2.901e+01 
R9443t1746 n9444 n1747 R=1.596e+01 
R9444t5637 n9445 n5638 R=3.002e+00 
R9444t6727 n9445 n6728 R=2.130e+01 
R9444t8089 n9445 n8090 R=1.808e+01 
R9444t375 n9445 n376 R=1.684e+01 
R9444t6803 n9445 n6804 R=3.146e+01 
R9444t5254 n9445 n5255 R=3.510e+01 
R9444t7521 n9445 n7522 R=3.660e+00 
R9444t7305 n9445 n7306 R=2.649e+01 
R9444t9297 n9445 n9298 R=2.171e+01 
R9444t6511 n9445 n6512 R=2.038e+02 
R9444t9193 n9445 n9194 R=1.125e+01 
R9445t3764 n9446 n3765 R=5.748e+00 
R9445t5074 n9446 n5075 R=9.055e+00 
R9445t159 n9446 n160 R=1.133e+01 
R9445t9435 n9446 n9436 R=8.285e+01 
R9445t1291 n9446 n1292 R=2.663e+00 
R9445t5270 n9446 n5271 R=1.299e+01 
R9445t1737 n9446 n1738 R=7.649e+00 
R9446t620 n9447 n621 R=2.375e+00 
R9446t6620 n9447 n6621 R=3.095e+01 
R9446t900 n9447 n901 R=1.472e+01 
R9446t6448 n9447 n6449 R=2.707e+00 
R9446t5260 n9447 n5261 R=1.762e+01 
R9447t2987 n9448 n2988 R=8.719e+00 
R9447t8234 n9448 n8235 R=1.239e+01 
R9447t9428 n9448 n9429 R=1.352e+01 
R9447t769 n9448 n770 R=1.190e+02 
R9447t1683 n9448 n1684 R=3.874e+00 
R9447t3465 n9448 n3466 R=9.619e+00 
R9448t397 n9449 n398 R=7.651e+00 
R9448t4177 n9449 n4178 R=4.023e+01 
R9448t2728 n9449 n2729 R=2.449e+01 
R9448t4148 n9449 n4149 R=5.785e+00 
R9448t3856 n9449 n3857 R=6.446e+00 
R9448t1198 n9449 n1199 R=1.268e+01 
R9448t4711 n9449 n4712 R=1.858e+01 
R9448t4110 n9449 n4111 R=6.486e+00 
R9449t2828 n9450 n2829 R=4.345e+00 
R9449t3094 n9450 n3095 R=1.479e+01 
R9449t907 n9450 n908 R=4.205e+00 
R9449t5264 n9450 n5265 R=1.103e+01 
R9449t1181 n9450 n1182 R=1.284e+01 
R9449t2164 n9450 n2165 R=3.112e+01 
R9450t1269 n9451 n1270 R=5.797e+00 
R9450t7124 n9451 n7125 R=5.088e+00 
R9450t8909 n9451 n8910 R=3.381e+01 
R9450t1556 n9451 n1557 R=1.892e+01 
R9450t8522 n9451 n8523 R=5.496e+00 
R9450t805 n9451 n806 R=2.529e+01 
R9450t4704 n9451 n4705 R=1.022e+02 
R9450t2757 n9451 n2758 R=3.397e+01 
R9450t2636 n9451 n2637 R=1.765e+01 
R9451t3269 n9452 n3270 R=7.188e+00 
R9451t8534 n9452 n8535 R=1.374e+01 
R9451t5958 n9452 n5959 R=8.956e+00 
R9451t1669 n9452 n1670 R=4.128e+00 
R9451t5241 n9452 n5242 R=4.089e+00 
R9451t4212 n9452 n4213 R=2.209e+01 
R9452t1052 n9453 n1053 R=7.398e+00 
R9452t9189 n9453 n9190 R=2.897e+01 
R9452t1378 n9453 n1379 R=1.651e+01 
R9452t3155 n9453 n3156 R=1.496e+01 
R9452t4176 n9453 n4177 R=4.505e+01 
R9452t1262 n9453 n1263 R=4.863e+00 
R9452t8704 n9453 n8705 R=2.771e+00 
R9453t2543 n9454 n2544 R=1.916e+00 
R9453t8794 n9454 n8795 R=5.460e+01 
R9453t8120 n9454 n8121 R=9.187e+00 
R9453t850 n9454 n851 R=5.716e+00 
R9453t4606 n9454 n4607 R=8.513e+00 
R9454t7520 n9455 n7521 R=6.100e+00 
R9454t7982 n9455 n7983 R=2.484e+01 
R9454t2696 n9455 n2697 R=4.263e+00 
R9454t8336 n9455 n8337 R=2.052e+01 
R9454t7372 n9455 n7373 R=1.177e+01 
R9455t6449 n9456 n6450 R=1.519e+01 
R9455t8383 n9456 n8384 R=3.640e+00 
R9455t5121 n9456 n5122 R=4.601e+01 
R9455t2447 n9456 n2448 R=6.250e+00 
R9455t7721 n9456 n7722 R=2.382e+01 
R9455t7578 n9456 n7579 R=4.533e+00 
R9455t1382 n9456 n1383 R=3.752e+01 
R9456t2252 n9457 n2253 R=8.865e+00 
R9456t6744 n9457 n6745 R=2.947e+00 
R9456t3568 n9457 n3569 R=4.810e+00 
R9456t6349 n9457 n6350 R=4.794e+00 
R9457t7054 n9458 n7055 R=1.218e+01 
R9457t7271 n9458 n7272 R=3.619e+00 
R9457t1073 n9458 n1074 R=3.828e+01 
R9457t7957 n9458 n7958 R=1.865e+01 
R9457t5839 n9458 n5840 R=6.168e+00 
R9458t4834 n9459 n4835 R=2.129e+00 
R9458t6898 n9459 n6899 R=2.088e+01 
R9458t8773 n9459 n8774 R=9.093e+00 
R9458t9296 n9459 n9297 R=4.566e+00 
R9458t8875 n9459 n8876 R=1.776e+01 
R9459t867 n9460 n868 R=5.174e+00 
R9459t8718 n9460 n8719 R=4.886e+00 
R9459t54 n9460 n55 R=8.805e+00 
R9459t148 n9460 n149 R=4.427e+00 
R9459t4 n9460 n5 R=3.481e+01 
R9459t4285 n9460 n4286 R=5.998e+01 
R9460t2285 n9461 n2286 R=4.271e+01 
R9460t3816 n9461 n3817 R=7.315e+01 
R9460t3576 n9461 n3577 R=9.219e+00 
R9460t5849 n9461 n5850 R=8.367e+00 
R9460t196 n9461 n197 R=7.511e+00 
R9460t7640 n9461 n7641 R=6.782e+00 
R9461t3437 n9462 n3438 R=6.557e+00 
R9461t6012 n9462 n6013 R=5.403e+00 
R9461t888 n9462 n889 R=2.945e+02 
R9461t5548 n9462 n5549 R=2.466e+00 
R9461t4744 n9462 n4745 R=1.259e+01 
R9462t805 n9463 n806 R=2.576e+00 
R9462t9450 n9463 n9451 R=1.050e+01 
R9462t495 n9463 n496 R=1.328e+01 
R9462t7566 n9463 n7567 R=1.227e+01 
R9462t8522 n9463 n8523 R=2.912e+00 
R9463t1364 n9464 n1365 R=2.186e+01 
R9463t7530 n9464 n7531 R=2.413e+00 
R9463t7293 n9464 n7294 R=1.010e+01 
R9463t1517 n9464 n1518 R=3.397e+00 
R9463t8902 n9464 n8903 R=9.857e+00 
R9463t6006 n9464 n6007 R=3.555e+01 
R9464t2277 n9465 n2278 R=1.877e+01 
R9464t6355 n9465 n6356 R=7.713e+00 
R9464t3817 n9465 n3818 R=8.994e+00 
R9464t4939 n9465 n4940 R=2.928e+00 
R9464t2112 n9465 n2113 R=4.964e+00 
R9465t2848 n9466 n2849 R=3.082e+00 
R9465t7208 n9466 n7209 R=4.560e+01 
R9465t3717 n9466 n3718 R=8.541e+00 
R9465t9403 n9466 n9404 R=4.647e+00 
R9465t1823 n9466 n1824 R=1.078e+01 
R9466t667 n9467 n668 R=3.529e+00 
R9466t5538 n9467 n5539 R=2.834e+01 
R9466t559 n9467 n560 R=3.001e+00 
R9466t8551 n9467 n8552 R=3.200e+00 
R9467t622 n9468 n623 R=2.816e+00 
R9467t7478 n9468 n7479 R=5.010e+01 
R9467t7740 n9468 n7741 R=3.228e+00 
R9467t93 n9468 n94 R=1.015e+01 
R9467t2147 n9468 n2148 R=2.105e+01 
R9467t2349 n9468 n2350 R=4.224e+01 
R9468t7025 n9469 n7026 R=8.374e+00 
R9468t9277 n9469 n9278 R=2.273e+01 
R9468t5983 n9469 n5984 R=1.388e+02 
R9468t4412 n9469 n4413 R=8.456e+01 
R9468t6635 n9469 n6636 R=6.581e+00 
R9468t131 n9469 n132 R=1.508e+01 
R9468t6380 n9469 n6381 R=4.803e+00 
R9469t784 n9470 n785 R=8.504e+00 
R9469t9402 n9470 n9403 R=3.037e+01 
R9469t3078 n9470 n3079 R=2.288e+01 
R9469t1301 n9470 n1302 R=3.646e+00 
R9469t5897 n9470 n5898 R=1.675e+00 
R9470t70 n9471 n71 R=2.888e+00 
R9470t2054 n9471 n2055 R=7.760e+00 
R9470t5269 n9471 n5270 R=6.233e+00 
R9470t4092 n9471 n4093 R=5.139e+00 
R9471t5544 n9472 n5545 R=9.357e+00 
R9471t9423 n9472 n9424 R=4.354e+00 
R9471t7460 n9472 n7461 R=1.218e+01 
R9471t2402 n9472 n2403 R=4.365e+00 
R9471t3033 n9472 n3034 R=5.843e+00 
R9472t1167 n9473 n1168 R=2.758e+01 
R9472t6421 n9473 n6422 R=7.231e+01 
R9472t3996 n9473 n3997 R=5.000e+01 
R9472t8306 n9473 n8307 R=7.829e+00 
R9472t5612 n9473 n5613 R=3.362e+00 
R9472t6393 n9473 n6394 R=1.019e+02 
R9472t3713 n9473 n3714 R=1.608e+01 
R9472t5194 n9473 n5195 R=3.438e+01 
R9472t8610 n9473 n8611 R=4.708e+00 
R9473t1184 n9474 n1185 R=6.680e+00 
R9473t4848 n9474 n4849 R=4.789e+00 
R9473t4951 n9474 n4952 R=5.384e+00 
R9473t4231 n9474 n4232 R=3.674e+02 
R9473t1307 n9474 n1308 R=2.191e+01 
R9473t3824 n9474 n3825 R=1.010e+01 
R9474t1561 n9475 n1562 R=5.930e+01 
R9474t9238 n9475 n9239 R=4.392e+00 
R9474t4872 n9475 n4873 R=2.298e+01 
R9474t3118 n9475 n3119 R=1.006e+01 
R9474t2966 n9475 n2967 R=1.329e+01 
R9474t2931 n9475 n2932 R=4.811e+02 
R9474t6522 n9475 n6523 R=1.478e+01 
R9474t8416 n9475 n8417 R=4.787e+00 
R9475t6289 n9476 n6290 R=4.981e+00 
R9475t8690 n9476 n8691 R=6.679e+00 
R9475t6417 n9476 n6418 R=6.049e+00 
R9475t8998 n9476 n8999 R=5.749e+00 
R9476t157 n9477 n158 R=3.663e+00 
R9476t5816 n9477 n5817 R=7.362e+00 
R9476t5136 n9477 n5137 R=1.106e+02 
R9476t2733 n9477 n2734 R=1.913e+01 
R9476t5165 n9477 n5166 R=4.840e+00 
R9476t451 n9477 n452 R=5.568e+00 
R9476t6767 n9477 n6768 R=8.248e+01 
R9477t81 n9478 n82 R=2.534e+01 
R9477t5200 n9478 n5201 R=3.531e+00 
R9477t4729 n9478 n4730 R=2.559e+00 
R9477t7159 n9478 n7160 R=7.017e+00 
R9478t8448 n9479 n8449 R=5.457e+00 
R9478t8604 n9479 n8605 R=4.781e+01 
R9478t2173 n9479 n2174 R=6.025e+00 
R9478t652 n9479 n653 R=3.319e+01 
R9478t9016 n9479 n9017 R=1.639e+01 
R9478t1109 n9479 n1110 R=2.372e+01 
R9478t4277 n9479 n4278 R=4.265e+00 
R9478t7635 n9479 n7636 R=2.891e+01 
R9479t3632 n9480 n3633 R=7.929e+00 
R9479t8736 n9480 n8737 R=1.613e+01 
R9479t874 n9480 n875 R=2.012e+01 
R9479t4977 n9480 n4978 R=6.117e+00 
R9479t3211 n9480 n3212 R=8.565e+00 
R9479t5594 n9480 n5595 R=5.038e+00 
R9479t9407 n9480 n9408 R=4.556e+01 
R9479t1743 n9480 n1744 R=3.021e+02 
R9479t3022 n9480 n3023 R=1.272e+02 
R9480t1372 n9481 n1373 R=5.835e+00 
R9480t8912 n9481 n8913 R=5.879e+00 
R9480t4067 n9481 n4068 R=1.153e+01 
R9480t4989 n9481 n4990 R=4.038e+00 
R9480t71 n9481 n72 R=6.556e+00 
R9481t605 n9482 n606 R=4.859e+00 
R9481t3286 n9482 n3287 R=6.879e+00 
R9481t4379 n9482 n4380 R=2.364e+00 
R9481t2596 n9482 n2597 R=7.083e+00 
R9482t1849 n9483 n1850 R=5.604e+00 
R9482t7365 n9483 n7366 R=1.832e+01 
R9482t2151 n9483 n2152 R=1.075e+01 
R9482t8801 n9483 n8802 R=3.556e+00 
R9482t1690 n9483 n1691 R=4.956e+00 
R9482t7599 n9483 n7600 R=5.204e+01 
R9482t2973 n9483 n2974 R=3.541e+01 
R9483t620 n9484 n621 R=1.349e+01 
R9483t2042 n9484 n2043 R=3.605e+00 
R9483t6611 n9484 n6612 R=1.978e+01 
R9483t8833 n9484 n8834 R=2.192e+00 
R9483t8653 n9484 n8654 R=2.188e+01 
R9484t4050 n9485 n4051 R=2.214e+01 
R9484t6235 n9485 n6236 R=4.910e+00 
R9484t7818 n9485 n7819 R=1.644e+01 
R9484t6910 n9485 n6911 R=6.451e+00 
R9484t3937 n9485 n3938 R=2.252e+01 
R9484t2146 n9485 n2147 R=2.923e+01 
R9484t8067 n9485 n8068 R=4.224e+00 
R9485t2952 n9486 n2953 R=3.563e+00 
R9485t8622 n9486 n8623 R=2.200e+01 
R9485t8831 n9486 n8832 R=3.258e+00 
R9485t3266 n9486 n3267 R=4.552e+00 
R9486t218 n9487 n219 R=9.818e+00 
R9486t9360 n9487 n9361 R=1.798e+00 
R9486t6458 n9487 n6459 R=2.817e+01 
R9486t5044 n9487 n5045 R=9.228e+00 
R9486t7316 n9487 n7317 R=2.304e+01 
R9486t9434 n9487 n9435 R=4.878e+00 
R9487t4268 n9488 n4269 R=2.411e+02 
R9487t7025 n9488 n7026 R=1.051e+03 
R9487t9422 n9488 n9423 R=3.615e+00 
R9487t8937 n9488 n8938 R=1.716e+02 
R9487t5983 n9488 n5984 R=1.535e+00 
R9487t9468 n9488 n9469 R=5.685e+00 
R9488t5947 n9489 n5948 R=4.776e+00 
R9488t6622 n9489 n6623 R=9.243e+00 
R9488t2842 n9489 n2843 R=6.288e+00 
R9488t6114 n9489 n6115 R=2.556e+01 
R9488t7528 n9489 n7529 R=1.582e+03 
R9488t2038 n9489 n2039 R=4.448e+00 
R9489t971 n9490 n972 R=3.128e+00 
R9489t5368 n9490 n5369 R=2.233e+01 
R9489t4986 n9490 n4987 R=2.554e+02 
R9489t4069 n9490 n4070 R=3.024e+00 
R9489t2423 n9490 n2424 R=2.484e+00 
R9490t1494 n9491 n1495 R=1.979e+00 
R9490t8804 n9491 n8805 R=1.229e+01 
R9490t4546 n9491 n4547 R=1.063e+01 
R9490t7885 n9491 n7886 R=4.243e+01 
R9490t8092 n9491 n8093 R=3.019e+00 
R9490t465 n9491 n466 R=8.910e+01 
R9491t29 n9492 n30 R=4.116e+00 
R9491t9351 n9492 n9352 R=1.048e+01 
R9491t5297 n9492 n5298 R=4.388e+00 
R9491t4800 n9492 n4801 R=6.591e+01 
R9491t1099 n9492 n1100 R=2.778e+00 
R9492t3029 n9493 n3030 R=4.081e+00 
R9492t7620 n9493 n7621 R=4.936e+00 
R9492t373 n9493 n374 R=1.035e+01 
R9492t550 n9493 n551 R=3.460e+00 
R9492t9297 n9493 n9298 R=2.365e+01 
R9493t6792 n9494 n6793 R=1.094e+01 
R9493t7596 n9494 n7597 R=2.024e+01 
R9493t6204 n9494 n6205 R=4.295e+00 
R9493t9041 n9494 n9042 R=8.022e+01 
R9493t6457 n9494 n6458 R=6.550e+00 
R9493t2530 n9494 n2531 R=1.134e+01 
R9494t515 n9495 n516 R=7.333e+00 
R9494t3158 n9495 n3159 R=4.361e+00 
R9494t5477 n9495 n5478 R=9.406e+00 
R9494t3823 n9495 n3824 R=4.976e+00 
R9494t2339 n9495 n2340 R=1.506e+01 
R9494t2520 n9495 n2521 R=1.478e+01 
R9495t836 n9496 n837 R=2.442e+01 
R9495t3908 n9496 n3909 R=9.464e+00 
R9495t8818 n9496 n8819 R=8.375e+00 
R9495t9267 n9496 n9268 R=3.628e+00 
R9495t4706 n9496 n4707 R=1.691e+02 
R9495t8137 n9496 n8138 R=4.197e+00 
R9496t8798 n9497 n8799 R=4.204e+00 
R9496t8951 n9497 n8952 R=1.415e+02 
R9496t6046 n9497 n6047 R=1.598e+01 
R9496t3400 n9497 n3401 R=5.238e+00 
R9496t2359 n9497 n2360 R=2.629e+00 
R9497t2852 n9498 n2853 R=3.091e+01 
R9497t8513 n9498 n8514 R=1.395e+01 
R9497t7134 n9498 n7135 R=8.151e+00 
R9497t419 n9498 n420 R=4.895e+00 
R9497t7054 n9498 n7055 R=4.516e+00 
R9498t2370 n9499 n2371 R=3.364e+00 
R9498t4613 n9499 n4614 R=5.640e+00 
R9498t7379 n9499 n7380 R=2.486e+01 
R9498t1832 n9499 n1833 R=2.107e+00 
R9499t6738 n9500 n6739 R=1.990e+00 
R9499t8238 n9500 n8239 R=4.893e+01 
R9499t27 n9500 n28 R=2.167e+00 
R9499t625 n9500 n626 R=1.359e+01 
R9500t329 n9501 n330 R=2.152e+01 
R9500t3474 n9501 n3475 R=3.776e+00 
R9500t2284 n9501 n2285 R=1.862e+01 
R9500t442 n9501 n443 R=2.963e+01 
R9500t3537 n9501 n3538 R=2.988e+00 
R9500t5377 n9501 n5378 R=2.451e+01 
R9501t134 n9502 n135 R=2.145e+00 
R9501t7215 n9502 n7216 R=6.423e+00 
R9501t8355 n9502 n8356 R=1.595e+00 
R9502t5806 n9503 n5807 R=9.623e+00 
R9502t6302 n9503 n6303 R=1.876e+01 
R9502t8317 n9503 n8318 R=3.253e+00 
R9502t2339 n9503 n2340 R=6.379e+00 
R9502t3823 n9503 n3824 R=8.285e+01 
R9502t8031 n9503 n8032 R=3.386e+00 
R9503t1368 n9504 n1369 R=2.258e+01 
R9503t2652 n9504 n2653 R=8.249e+00 
R9503t1799 n9504 n1800 R=2.926e+00 
R9503t3353 n9504 n3354 R=4.950e+01 
R9503t7063 n9504 n7064 R=1.770e+00 
R9504t4995 n9505 n4996 R=5.664e+00 
R9504t8901 n9505 n8902 R=1.120e+01 
R9504t9004 n9505 n9005 R=4.632e+00 
R9504t510 n9505 n511 R=1.615e+02 
R9504t1767 n9505 n1768 R=2.558e+00 
R9505t7617 n9506 n7618 R=1.181e+01 
R9505t8176 n9506 n8177 R=1.890e+01 
R9505t2944 n9506 n2945 R=5.003e+00 
R9505t3717 n9506 n3718 R=1.118e+01 
R9505t3661 n9506 n3662 R=3.032e+01 
R9505t8401 n9506 n8402 R=5.269e+00 
R9505t6301 n9506 n6302 R=5.548e+00 
R9506t7141 n9507 n7142 R=2.348e+01 
R9506t7914 n9507 n7915 R=3.138e+00 
R9506t847 n9507 n848 R=6.369e+00 
R9506t5100 n9507 n5101 R=9.972e+00 
R9506t6563 n9507 n6564 R=1.114e+01 
R9506t4054 n9507 n4055 R=9.316e+00 
R9507t1655 n9508 n1656 R=2.974e+00 
R9507t8753 n9508 n8754 R=1.224e+01 
R9507t4880 n9508 n4881 R=2.387e+02 
R9507t1118 n9508 n1119 R=1.988e+00 
R9507t2982 n9508 n2983 R=6.989e+00 
R9508t1041 n9509 n1042 R=2.120e+01 
R9508t6721 n9509 n6722 R=5.074e+00 
R9508t2868 n9509 n2869 R=2.486e+00 
R9508t2641 n9509 n2642 R=4.639e+00 
R9509t1439 n9510 n1440 R=2.885e+03 
R9509t2847 n9510 n2848 R=3.584e+00 
R9509t1652 n9510 n1653 R=2.315e+01 
R9509t2570 n9510 n2571 R=7.595e+00 
R9509t5295 n9510 n5296 R=8.292e+00 
R9509t5863 n9510 n5864 R=8.705e+00 
R9509t6952 n9510 n6953 R=2.654e+01 
R9509t9100 n9510 n9101 R=1.262e+01 
R9509t4021 n9510 n4022 R=1.184e+01 
R9510t42 n1 n43 R=2.901e+01 
R9510t4042 n1 n4043 R=8.107e+01 
R9511t1691 n9512 n1692 R=6.215e+00 
R9511t2176 n9512 n2177 R=7.187e+00 
R9511t322 n9512 n323 R=8.609e+00 
R9511t4329 n9512 n4330 R=6.507e+00 
R9511t8403 n9512 n8404 R=5.182e+00 
R9511t8665 n9512 n8666 R=5.499e+01 
R9511t1111 n9512 n1112 R=7.051e+01 
R9512t1841 n9513 n1842 R=3.360e+00 
R9512t2649 n9513 n2650 R=1.557e+01 
R9512t5502 n9513 n5503 R=1.192e+01 
R9512t7353 n9513 n7354 R=4.108e+01 
R9512t1853 n9513 n1854 R=2.847e+00 
R9512t876 n9513 n877 R=1.931e+01 
R9512t7663 n9513 n7664 R=2.491e+01 
R9513t1596 n9514 n1597 R=2.250e+00 
R9513t7054 n9514 n7055 R=9.123e+01 
R9513t9457 n9514 n9458 R=3.649e+00 
R9513t5839 n9514 n5840 R=1.656e+01 
R9513t6180 n9514 n6181 R=2.059e+01 
R9514t6000 n9515 n6001 R=6.279e+01 
R9514t6655 n9515 n6656 R=4.196e+00 
R9514t5933 n9515 n5934 R=4.465e+00 
R9514t951 n9515 n952 R=2.031e+01 
R9514t1350 n9515 n1351 R=1.403e+02 
R9514t8930 n9515 n8931 R=9.366e+00 
R9514t1307 n9515 n1308 R=6.283e+00 
R9514t6111 n9515 n6112 R=1.250e+01 
R9515t2357 n9516 n2358 R=3.583e+01 
R9515t5271 n9516 n5272 R=2.702e+00 
R9515t8224 n9516 n8225 R=8.751e+00 
R9515t1467 n9516 n1468 R=1.382e+01 
R9515t1421 n9516 n1422 R=6.728e+00 
R9515t8230 n9516 n8231 R=1.421e+01 
R9516t4044 n9517 n4045 R=6.947e+00 
R9516t4160 n9517 n4161 R=1.133e+02 
R9516t4545 n9517 n4546 R=3.929e+00 
R9516t7250 n9517 n7251 R=1.018e+01 
R9516t252 n9517 n253 R=1.213e+01 
R9516t4739 n9517 n4740 R=3.071e+00 
R9517t3188 n9518 n3189 R=4.318e+00 
R9517t7200 n9518 n7201 R=1.298e+01 
R9517t2121 n9518 n2122 R=1.497e+01 
R9517t4861 n9518 n4862 R=3.385e+00 
R9517t4404 n9518 n4405 R=4.215e+01 
R9517t4771 n9518 n4772 R=2.625e+02 
R9517t8550 n9518 n8551 R=6.990e+00 
R9518t1992 n9519 n1993 R=8.330e+00 
R9518t7934 n9519 n7935 R=4.827e+00 
R9518t8045 n9519 n8046 R=6.494e+00 
R9518t285 n9519 n286 R=2.289e+00 
R9519t1252 n9520 n1253 R=1.063e+01 
R9519t5883 n9520 n5884 R=2.297e+00 
R9519t4011 n9520 n4012 R=2.362e+00 
R9519t8888 n9520 n8889 R=7.390e+00 
R9520t7569 n9521 n7570 R=1.154e+01 
R9520t8337 n9521 n8338 R=1.560e+01 
R9520t8063 n9521 n8064 R=5.510e+01 
R9520t5275 n9521 n5276 R=4.697e+00 
R9520t7595 n9521 n7596 R=9.356e+00 
R9520t6901 n9521 n6902 R=4.007e+00 
R9520t8168 n9521 n8169 R=2.124e+01 
R9521t2922 n9522 n2923 R=3.775e+02 
R9521t7882 n9522 n7883 R=6.906e+00 
R9521t4134 n9522 n4135 R=4.294e+00 
R9521t4510 n9522 n4511 R=3.159e+00 
R9521t9215 n9522 n9216 R=4.963e+00 
R9522t925 n9523 n926 R=2.544e+01 
R9522t6280 n9523 n6281 R=2.119e+01 
R9522t8672 n9523 n8673 R=1.627e+00 
R9522t8348 n9523 n8349 R=1.153e+01 
R9522t2372 n9523 n2373 R=3.815e+00 
R9522t4129 n9523 n4130 R=1.238e+02 
R9523t2149 n9524 n2150 R=1.352e+01 
R9523t9428 n9524 n9429 R=5.201e+00 
R9523t9447 n9524 n9448 R=6.217e+01 
R9523t769 n9524 n770 R=3.600e+00 
R9523t7214 n9524 n7215 R=2.641e+00 
R9523t1764 n9524 n1765 R=6.728e+02 
R9524t5526 n9525 n5527 R=1.261e+01 
R9524t7445 n9525 n7446 R=1.431e+01 
R9524t6340 n9525 n6341 R=1.084e+02 
R9524t156 n9525 n157 R=3.347e+00 
R9525t3279 n9526 n3280 R=2.032e+01 
R9525t8430 n9526 n8431 R=2.050e+00 
R9525t8056 n9526 n8057 R=3.474e+00 
R9525t7022 n9526 n7023 R=6.726e+01 
R9525t814 n9526 n815 R=6.337e+00 
R9525t2083 n9526 n2084 R=1.677e+02 
R9525t5465 n9526 n5466 R=5.070e+01 
R9526t2285 n9527 n2286 R=1.519e+01 
R9526t9460 n9527 n9461 R=4.389e+00 
R9526t7640 n9527 n7641 R=7.121e+00 
R9526t4911 n9527 n4912 R=1.270e+01 
R9526t6780 n9527 n6781 R=4.125e+00 
R9527t1327 n9528 n1328 R=1.026e+01 
R9527t3863 n9528 n3864 R=7.597e+00 
R9527t2107 n9528 n2108 R=1.303e+01 
R9527t639 n9528 n640 R=7.693e+00 
R9527t6637 n9528 n6638 R=6.541e+01 
R9527t6267 n9528 n6268 R=2.778e+00 
R9527t6893 n9528 n6894 R=2.334e+01 
R9528t3694 n9529 n3695 R=7.851e+00 
R9528t4382 n9529 n4383 R=1.790e+04 
R9528t257 n9529 n258 R=3.242e+00 
R9528t9056 n9529 n9057 R=7.728e+00 
R9528t1949 n9529 n1950 R=7.546e+00 
R9528t7275 n9529 n7276 R=3.018e+01 
R9528t1010 n9529 n1011 R=8.373e+00 
R9529t3559 n9530 n3560 R=1.739e+01 
R9529t7419 n9530 n7420 R=2.298e+00 
R9529t8570 n9530 n8571 R=5.939e+00 
R9529t2779 n9530 n2780 R=3.849e+00 
R9529t1893 n9530 n1894 R=4.492e+01 
R9530t2956 n9531 n2957 R=5.729e+00 
R9530t4101 n9531 n4102 R=7.383e+01 
R9530t5180 n9531 n5181 R=1.761e+02 
R9530t5792 n9531 n5793 R=1.759e+01 
R9530t8824 n9531 n8825 R=3.422e+00 
R9531t5268 n9532 n5269 R=6.605e+00 
R9531t7376 n9532 n7377 R=2.116e+01 
R9531t7516 n9532 n7517 R=5.364e+00 
R9531t6217 n9532 n6218 R=4.084e+01 
R9531t3783 n9532 n3784 R=7.494e+01 
R9531t546 n9532 n547 R=8.122e+00 
R9531t3281 n9532 n3282 R=8.978e+00 
R9531t4222 n9532 n4223 R=8.574e+00 
R9532t1707 n9533 n1708 R=6.026e+00 
R9532t8491 n9533 n8492 R=3.535e+00 
R9532t3913 n9533 n3914 R=1.051e+01 
R9532t4272 n9533 n4273 R=1.062e+01 
R9532t377 n9533 n378 R=3.131e+01 
R9532t6551 n9533 n6552 R=2.880e+01 
R9533t3331 n9534 n3332 R=6.584e+00 
R9533t5848 n9534 n5849 R=2.406e+00 
R9533t4936 n9534 n4937 R=2.723e+01 
R9533t4922 n9534 n4923 R=3.185e+00 
R9533t4430 n9534 n4431 R=1.706e+01 
R9534t3389 n9535 n1 R=7.560e+00 
R9534t8817 n9535 n8818 R=1.380e+01 
R9534t8612 n9535 n8613 R=3.704e+00 
R9534t2247 n9535 n2248 R=1.480e+01 
R9534t5531 n9535 n5532 R=3.626e+01 
R9534t3819 n9535 n3820 R=9.478e+00 
R9534t2964 n9535 n2965 R=8.871e+00 
R9535t7293 n9536 n7294 R=2.109e+00 
R9535t8897 n9536 n8898 R=2.266e+01 
R9535t9128 n9536 n9129 R=5.817e+00 
R9535t2351 n9536 n2352 R=2.654e+00 
R9536t6180 n9537 n6181 R=2.820e+00 
R9536t9513 n9537 n9514 R=9.006e+00 
R9536t5839 n9537 n5840 R=8.007e+00 
R9536t1976 n9537 n1977 R=1.872e+01 
R9536t1400 n9537 n1401 R=6.747e+00 
R9536t6660 n9537 n6661 R=9.842e+01 
R9537t1749 n9538 n1750 R=3.504e+00 
R9537t4471 n9538 n4472 R=2.766e+01 
R9537t3834 n9538 n3835 R=1.080e+01 
R9537t581 n9538 n582 R=1.744e+02 
R9537t2056 n9538 n2057 R=3.446e+00 
R9537t5763 n9538 n5764 R=4.786e+00 
R9538t1841 n9539 n1842 R=4.945e+00 
R9538t2649 n9539 n2650 R=5.719e+00 
R9538t6579 n9539 n6580 R=1.246e+01 
R9538t7695 n9539 n7696 R=6.078e+00 
R9538t8258 n9539 n8259 R=1.484e+01 
R9539t5139 n9540 n5140 R=1.794e+01 
R9539t6556 n9540 n6557 R=7.568e+01 
R9539t2214 n9540 n2215 R=2.627e+00 
R9539t7927 n9540 n7928 R=8.562e+00 
R9539t1581 n9540 n1582 R=9.178e+00 
R9539t7357 n9540 n7358 R=3.625e+00 
R9540t5709 n9541 n5710 R=7.882e+00 
R9540t5735 n9541 n5736 R=1.866e+02 
R9540t1003 n9541 n1004 R=2.273e+00 
R9540t2665 n9541 n2666 R=6.630e+03 
R9540t6298 n9541 n6299 R=1.564e+01 
R9540t7826 n9541 n7827 R=3.095e+00 
R9541t209 n9542 n210 R=1.353e+01 
R9541t8252 n9542 n8253 R=3.370e+02 
R9541t8330 n9542 n8331 R=6.128e+01 
R9541t202 n9542 n203 R=1.077e+01 
R9541t6683 n9542 n6684 R=6.242e+00 
R9541t3586 n9542 n3587 R=4.852e+00 
R9541t873 n9542 n874 R=8.553e+01 
R9541t6885 n9542 n6886 R=2.501e+00 
R9542t993 n9543 n994 R=4.900e+00 
R9542t8553 n9543 n8554 R=3.710e+00 
R9542t1326 n9543 n1327 R=1.967e+01 
R9542t3508 n9543 n3509 R=2.198e+01 
R9542t1830 n9543 n1831 R=3.463e+00 
R9542t3899 n9543 n3900 R=3.655e+01 
R9543t2047 n9544 n2048 R=2.861e+00 
R9543t4162 n9544 n4163 R=4.260e+01 
R9543t1645 n9544 n1646 R=9.988e+01 
R9543t7655 n9544 n7656 R=3.054e+00 
R9543t7259 n9544 n7260 R=4.948e+00 
R9544t9027 n9545 n9028 R=5.850e+00 
R9544t9389 n9545 n9390 R=4.142e+01 
R9544t1442 n9545 n1443 R=1.627e+01 
R9544t7647 n9545 n7648 R=5.711e+00 
R9544t7983 n9545 n7984 R=2.485e+00 
R9544t1391 n9545 n1392 R=1.384e+02 
R9545t2549 n9546 n2550 R=3.508e+01 
R9545t5669 n9546 n5670 R=4.522e+00 
R9545t8968 n9546 n8969 R=3.944e+00 
R9545t3005 n9546 n3006 R=8.153e+00 
R9545t12 n9546 n13 R=6.337e+01 
R9545t8451 n9546 n8452 R=3.857e+00 
R9546t382 n9547 n383 R=3.003e+01 
R9546t4649 n9547 n4650 R=1.246e+01 
R9546t4693 n9547 n4694 R=3.642e+00 
R9546t479 n9547 n480 R=1.440e+01 
R9546t9114 n9547 n9115 R=1.660e+02 
R9546t4742 n9547 n4743 R=3.592e+00 
R9546t5552 n9547 n5553 R=9.028e+00 
R9547t6924 n9548 n6925 R=2.838e+00 
R9547t8295 n9548 n8296 R=1.201e+01 
R9547t8536 n9548 n8537 R=6.882e+00 
R9547t5014 n9548 n5015 R=3.642e+00 
R9547t7782 n9548 n7783 R=1.584e+01 
R9548t5643 n9549 n5644 R=3.262e+00 
R9548t7166 n9549 n7167 R=3.832e+01 
R9548t5800 n9549 n5801 R=8.077e+00 
R9548t2734 n9549 n2735 R=6.649e+00 
R9548t79 n9549 n80 R=8.044e+00 
R9548t4893 n9549 n4894 R=1.652e+01 
R9549t9439 n9550 n9440 R=8.009e+00 
R9549t1374 n9550 n1375 R=4.133e+01 
R9549t1311 n9550 n1312 R=5.609e+00 
R9549t8424 n9550 n8425 R=1.774e+01 
R9549t2161 n9550 n2162 R=2.587e+00 
R9550t808 n9551 n809 R=5.756e+00 
R9550t8431 n9551 n8432 R=1.016e+01 
R9550t3411 n9551 n3412 R=2.447e+01 
R9550t9245 n9551 n9246 R=9.124e+00 
R9550t5987 n9551 n5988 R=1.515e+01 
R9550t3582 n9551 n3583 R=7.733e+00 
R9550t619 n9551 n620 R=3.861e+00 
R9550t1382 n9551 n1383 R=5.130e+02 
R9551t1303 n9552 n1304 R=1.526e+01 
R9551t7559 n9552 n7560 R=9.208e+01 
R9551t4562 n9552 n4563 R=4.576e+00 
R9551t1299 n9552 n1300 R=4.141e+00 
R9551t378 n9552 n379 R=3.408e+00 
R9552t517 n9553 n518 R=1.996e+02 
R9552t7583 n9553 n7584 R=3.245e+00 
R9552t3607 n9553 n3608 R=2.124e+00 
R9552t1914 n9553 n1915 R=8.885e+01 
R9552t1497 n9553 n1498 R=3.089e+01 
R9552t9425 n9553 n9426 R=5.140e+00 
R9553t6947 n9554 n6948 R=6.917e+00 
R9553t6985 n9554 n6986 R=1.094e+01 
R9553t6221 n9554 n6222 R=6.969e+00 
R9553t1733 n9554 n1734 R=6.625e+00 
R9553t276 n9554 n277 R=2.710e+01 
R9553t8949 n9554 n8950 R=3.595e+02 
R9554t2331 n9555 n2332 R=3.813e+00 
R9554t3895 n9555 n3896 R=1.308e+01 
R9554t964 n9555 n965 R=9.557e+00 
R9554t3401 n9555 n3402 R=1.454e+00 
R9555t2567 n9556 n2568 R=1.614e+02 
R9555t6610 n9556 n6611 R=2.439e+00 
R9555t7165 n9556 n7166 R=9.060e+00 
R9555t182 n9556 n183 R=8.172e+00 
R9555t2705 n9556 n2706 R=6.691e+00 
R9556t3810 n9557 n3811 R=9.148e+00 
R9556t8227 n9557 n8228 R=1.431e+01 
R9556t7992 n9557 n7993 R=4.739e+00 
R9556t8751 n9557 n8752 R=1.888e+00 
R9557t3165 n9558 n3166 R=3.950e+00 
R9557t1008 n9558 n1009 R=2.765e+00 
R9557t1895 n9558 n1896 R=2.714e+01 
R9557t4683 n9558 n4684 R=7.656e+02 
R9557t3185 n9558 n3186 R=8.675e+01 
R9558t5115 n9559 n5116 R=1.923e+01 
R9558t7832 n9559 n7833 R=1.206e+01 
R9558t2161 n9559 n2162 R=3.502e+01 
R9558t9549 n9559 n9550 R=7.348e+00 
R9558t9439 n9559 n9440 R=2.565e+01 
R9558t4690 n9559 n4691 R=5.902e+00 
R9558t5668 n9559 n5669 R=6.237e+00 
R9558t8058 n9559 n8059 R=7.636e+00 
R9559t5706 n9560 n5707 R=2.210e+01 
R9559t8933 n9560 n8934 R=1.752e+02 
R9559t618 n9560 n619 R=2.112e+01 
R9559t3372 n9560 n3373 R=4.385e+00 
R9559t2014 n9560 n2015 R=2.284e+01 
R9559t3817 n9560 n3818 R=3.902e+00 
R9559t4292 n9560 n4293 R=3.239e+00 
R9560t6868 n9561 n6869 R=5.056e+00 
R9560t7776 n9561 n7777 R=8.926e+00 
R9560t3019 n9561 n3020 R=5.428e+01 
R9560t766 n9561 n767 R=2.216e+01 
R9560t1579 n9561 n1580 R=2.574e+00 
R9560t4529 n9561 n4530 R=2.209e+01 
R9561t724 n9562 n725 R=2.642e+01 
R9561t8646 n9562 n8647 R=1.654e+00 
R9561t1433 n9562 n1434 R=2.445e+01 
R9561t7207 n9562 n7208 R=6.399e+00 
R9561t4741 n9562 n4742 R=6.876e+00 
R9561t833 n9562 n834 R=1.118e+01 
R9562t2417 n9563 n2418 R=3.010e+02 
R9562t5149 n9563 n5150 R=1.478e+01 
R9562t4996 n9563 n1 R=2.690e+00 
R9562t8679 n9563 n1 R=5.067e+00 
R9562t8281 n9563 n8282 R=6.116e+00 
R9562t7715 n9563 n7716 R=9.934e+00 
R9563t2466 n9564 n2467 R=2.221e+01 
R9563t3467 n9564 n3468 R=3.205e+00 
R9563t3889 n9564 n3890 R=5.185e+00 
R9563t4599 n9564 n4600 R=1.017e+01 
R9564t5023 n9565 n5024 R=1.827e+01 
R9564t5355 n9565 n5356 R=6.694e+00 
R9564t6791 n9565 n6792 R=1.174e+01 
R9564t751 n9565 n752 R=2.388e+00 
R9564t4993 n9565 n4994 R=6.506e+00 
R9565t4533 n9566 n4534 R=7.415e+00 
R9565t7493 n9566 n7494 R=9.899e+00 
R9565t6805 n9566 n6806 R=1.479e+01 
R9565t963 n9566 n964 R=2.348e+01 
R9565t6081 n9566 n6082 R=1.343e+01 
R9565t7573 n9566 n7574 R=6.582e+00 
R9565t7621 n9566 n7622 R=1.715e+02 
R9565t984 n9566 n985 R=5.436e+00 
R9565t5540 n9566 n5541 R=3.071e+01 
R9566t8009 n9567 n8010 R=7.882e+00 
R9566t8353 n9567 n8354 R=5.983e+00 
R9566t4062 n9567 n4063 R=5.598e+01 
R9566t2853 n9567 n2854 R=3.732e+00 
R9567t1705 n9568 n1706 R=1.293e+01 
R9567t8749 n9568 n8750 R=4.019e+00 
R9567t6172 n9568 n6173 R=6.595e+00 
R9567t5610 n9568 n5611 R=8.317e+01 
R9567t8936 n9568 n8937 R=5.940e+00 
R9567t1523 n9568 n1524 R=1.758e+01 
R9567t3729 n9568 n3730 R=1.018e+01 
R9567t4865 n9568 n4866 R=1.283e+01 
R9568t5256 n9569 n5257 R=2.326e+01 
R9568t8476 n9569 n8477 R=7.024e+00 
R9568t5899 n9569 n5900 R=1.936e+00 
R9568t5626 n9569 n5627 R=8.813e+00 
R9568t8515 n9569 n8516 R=3.504e+00 
R9569t7613 n9570 n7614 R=6.928e+00 
R9569t9330 n9570 n9331 R=5.683e+00 
R9569t4619 n9570 n4620 R=5.927e+00 
R9569t4445 n9570 n4446 R=4.238e+00 
R9569t2858 n9570 n2859 R=7.930e+00 
R9570t242 n9571 n243 R=1.553e+02 
R9570t6626 n9571 n6627 R=1.772e+01 
R9570t2711 n9571 n2712 R=3.654e+00 
R9570t8279 n9571 n8280 R=2.809e+00 
R9570t1162 n9571 n1163 R=3.633e+00 
R9571t3128 n9572 n3129 R=2.516e+01 
R9571t8038 n9572 n8039 R=2.944e+00 
R9571t1051 n9572 n1052 R=3.234e+02 
R9571t6883 n9572 n6884 R=2.217e+00 
R9571t8356 n9572 n8357 R=5.974e+00 
R9572t4027 n9573 n4028 R=1.832e+01 
R9572t6320 n9573 n6321 R=7.443e+00 
R9572t4163 n9573 n4164 R=9.792e+00 
R9572t103 n9573 n104 R=2.371e+01 
R9572t7625 n9573 n7626 R=3.467e+00 
R9572t7458 n9573 n7459 R=7.912e+00 
R9572t7911 n9573 n7912 R=2.637e+01 
R9573t5323 n9574 n5324 R=6.555e+00 
R9573t6210 n9574 n6211 R=6.728e+01 
R9573t7741 n9574 n7742 R=3.624e+02 
R9573t6465 n9574 n6466 R=7.558e+00 
R9573t8044 n9574 n8045 R=7.103e+00 
R9573t2117 n9574 n2118 R=4.494e+00 
R9574t4695 n9575 n4696 R=1.977e+01 
R9574t7781 n9575 n7782 R=1.496e+01 
R9574t1978 n9575 n1979 R=1.742e+00 
R9574t3099 n9575 n3100 R=1.545e+00 
R9575t5859 n9576 n5860 R=1.144e+01 
R9575t8180 n9576 n8181 R=4.061e+00 
R9575t2886 n9576 n2887 R=2.144e+00 
R9575t1654 n9576 n1655 R=1.284e+01 
R9575t4512 n9576 n4513 R=7.892e+00 
R9576t1592 n9577 n1593 R=1.073e+02 
R9576t6598 n9577 n6599 R=2.577e+00 
R9576t2638 n9577 n2639 R=8.477e+01 
R9576t2480 n9577 n2481 R=1.356e+01 
R9576t1288 n9577 n1289 R=3.918e+00 
R9576t8235 n9577 n8236 R=7.630e+00 
R9577t235 n9578 n236 R=2.619e+01 
R9577t5652 n9578 n5653 R=7.318e+02 
R9577t6207 n9578 n6208 R=5.666e+00 
R9577t2748 n9578 n2749 R=2.169e+01 
R9577t8642 n9578 n8643 R=5.503e+00 
R9577t5988 n9578 n5989 R=6.593e+00 
R9577t5153 n9578 n5154 R=5.226e+01 
R9577t2673 n9578 n2674 R=5.436e+00 
R9578t3628 n9579 n3629 R=9.662e+00 
R9578t8070 n9579 n8071 R=1.095e+01 
R9578t1555 n9579 n1556 R=6.124e+00 
R9578t3874 n9579 n3875 R=5.238e+00 
R9578t1776 n9579 n1777 R=2.110e+02 
R9578t2206 n9579 n2207 R=8.572e+00 
R9578t3359 n9579 n3360 R=1.126e+01 
R9579t2686 n9580 n2687 R=4.546e+01 
R9579t6483 n9580 n6484 R=2.162e+00 
R9579t3843 n9580 n3844 R=3.480e+01 
R9579t4008 n9580 n4009 R=6.507e+00 
R9579t9025 n9580 n9026 R=3.404e+00 
R9579t1601 n9580 n1602 R=1.704e+01 
R9579t873 n9580 n874 R=4.128e+01 
R9580t2526 n9581 n2527 R=1.845e+00 
R9580t5920 n9581 n5921 R=3.695e+01 
R9580t6719 n9581 n6720 R=6.877e+01 
R9580t4125 n9581 n4126 R=4.480e+00 
R9580t8057 n9581 n8058 R=1.432e+02 
R9580t2736 n9581 n2737 R=5.869e+00 
R9580t7621 n9581 n7622 R=1.018e+01 
R9581t8219 n9582 n8220 R=2.814e+00 
R9581t8670 n9582 n8671 R=9.127e+00 
R9581t4261 n9582 n4262 R=6.446e+01 
R9581t2268 n9582 n2269 R=8.471e+00 
R9581t2430 n9582 n2431 R=4.076e+00 
R9582t598 n9583 n599 R=2.031e+01 
R9582t790 n9583 n791 R=3.047e+01 
R9582t8851 n9583 n8852 R=4.320e+00 
R9582t4328 n9583 n4329 R=9.282e+01 
R9582t7158 n9583 n7159 R=8.741e+00 
R9582t4242 n9583 n4243 R=3.791e+00 
R9582t4933 n9583 n4934 R=4.482e+00 
R9583t5180 n9584 n5181 R=5.266e+00 
R9583t9530 n9584 n9531 R=5.238e+00 
R9583t6346 n9584 n6347 R=3.263e+01 
R9583t8521 n9584 n8522 R=3.936e+00 
R9583t2341 n9584 n2342 R=1.494e+01 
R9583t2956 n9584 n2957 R=1.546e+01 
R9584t515 n9585 n516 R=3.574e+00 
R9584t3158 n9585 n3159 R=1.545e+01 
R9584t5477 n9585 n5478 R=1.066e+01 
R9584t8193 n9585 n8194 R=2.265e+00 
R9584t3180 n9585 n3181 R=3.152e+01 
R9584t624 n9585 n625 R=9.877e+00 
R9585t344 n9586 n345 R=1.112e+01 
R9585t6935 n9586 n6936 R=2.427e+01 
R9585t1110 n9586 n1111 R=3.667e+01 
R9585t5472 n9586 n5473 R=6.869e+00 
R9585t89 n9586 n90 R=9.366e+00 
R9585t4124 n9586 n4125 R=1.986e+01 
R9585t176 n9586 n177 R=4.597e+00 
R9585t4003 n9586 n4004 R=2.011e+01 
R9586t6947 n9587 n6948 R=6.769e+00 
R9586t9553 n9587 n9554 R=7.888e+00 
R9586t4300 n9587 n4301 R=4.290e+00 
R9586t8949 n9587 n8950 R=3.376e+00 
R9587t557 n9588 n558 R=1.337e+01 
R9587t8910 n9588 n8911 R=7.928e+00 
R9587t7071 n9588 n7072 R=3.173e+00 
R9587t9424 n9588 n9425 R=4.331e+02 
R9587t8504 n9588 n8505 R=7.118e+00 
R9587t4552 n9588 n4553 R=8.375e+00 
R9587t3512 n9588 n3513 R=2.803e+01 
R9588t8775 n9589 n8776 R=4.525e+00 
R9588t8827 n9589 n8828 R=7.360e+00 
R9588t2376 n9589 n2377 R=4.015e+02 
R9588t5219 n9589 n5220 R=2.743e+02 
R9588t6206 n9589 n6207 R=4.562e+00 
R9588t8855 n9589 n8856 R=7.988e+00 
R9588t5460 n9589 n5461 R=1.940e+01 
R9589t351 n9590 n352 R=5.491e+00 
R9589t7273 n9590 n7274 R=5.823e+00 
R9589t4833 n9590 n4834 R=6.860e+00 
R9589t3232 n9590 n3233 R=7.449e+01 
R9589t4772 n9590 n4773 R=1.012e+01 
R9589t6609 n9590 n6610 R=4.975e+00 
R9589t3478 n9590 n3479 R=2.362e+01 
R9589t477 n9590 n478 R=5.975e+01 
R9590t1900 n9591 n1901 R=1.562e+01 
R9590t2265 n9591 n2266 R=3.760e+00 
R9590t2801 n9591 n2802 R=4.205e+01 
R9590t1688 n9591 n1689 R=5.883e+00 
R9590t4673 n9591 n4674 R=3.473e+02 
R9590t1831 n9591 n1832 R=7.874e+00 
R9590t5948 n9591 n5949 R=1.092e+01 
R9590t4712 n9591 n4713 R=3.363e+01 
R9590t1608 n9591 n1609 R=1.744e+01 
R9591t5417 n9592 n5418 R=2.942e+01 
R9591t6128 n9592 n6129 R=3.269e+00 
R9591t3080 n9592 n3081 R=5.180e+00 
R9591t6652 n9592 n6653 R=9.161e+01 
R9591t5335 n9592 n5336 R=1.250e+02 
R9591t3615 n9592 n3616 R=5.124e+00 
R9591t2721 n9592 n2722 R=1.844e+01 
R9592t1790 n9593 n1791 R=1.093e+01 
R9592t8801 n9593 n8802 R=2.789e+00 
R9592t2800 n9593 n2801 R=2.229e+01 
R9592t7966 n9593 n7967 R=3.311e+00 
R9592t3725 n9593 n3726 R=8.298e+00 
R9593t6363 n9594 n6364 R=2.506e+00 
R9593t6370 n9594 n6371 R=3.690e+00 
R9593t4495 n9594 n4496 R=2.935e+02 
R9593t1206 n9594 n1207 R=3.183e+02 
R9593t2668 n9594 n2669 R=2.936e+00 
R9594t2987 n9595 n2988 R=9.117e+00 
R9594t9447 n9595 n9448 R=1.201e+01 
R9594t3465 n9595 n3466 R=4.583e+00 
R9594t8156 n9595 n8157 R=5.613e+00 
R9594t9380 n9595 n9381 R=8.533e+01 
R9594t7096 n9595 n7097 R=5.293e+00 
R9595t4727 n9596 n4728 R=2.156e+00 
R9595t8389 n9596 n8390 R=9.861e+00 
R9595t1193 n9596 n1194 R=9.802e+01 
R9595t8182 n9596 n8183 R=4.807e+00 
R9595t6516 n9596 n6517 R=6.267e+00 
R9595t7857 n9596 n7858 R=5.358e+01 
R9596t110 n9597 n111 R=2.743e+00 
R9596t5616 n9597 n5617 R=7.052e+00 
R9596t7052 n9597 n7053 R=1.112e+01 
R9596t4860 n9597 n4861 R=1.337e+01 
R9596t3104 n9597 n3105 R=1.153e+01 
R9597t3027 n9598 n3028 R=2.985e+01 
R9597t5895 n9598 n5896 R=2.026e+01 
R9597t4691 n9598 n4692 R=4.916e+00 
R9597t4049 n9598 n4050 R=5.317e+00 
R9597t5214 n9598 n5215 R=1.159e+02 
R9597t7374 n9598 n7375 R=1.128e+01 
R9597t9359 n9598 n9360 R=2.056e+01 
R9597t1126 n9598 n1127 R=6.712e+00 
R9598t1413 n9599 n1414 R=5.519e+01 
R9598t7833 n9599 n7834 R=2.940e+00 
R9598t48 n9599 n49 R=6.708e+00 
R9598t2892 n9599 n2893 R=1.990e+01 
R9598t8464 n9599 n8465 R=3.337e+01 
R9598t2464 n9599 n2465 R=6.865e+00 
R9598t2660 n9599 n2661 R=1.334e+01 
R9599t273 n9600 n274 R=4.657e+00 
R9599t8053 n9600 n8054 R=2.218e+02 
R9599t3 n9600 n4 R=1.704e+01 
R9599t6028 n9600 n6029 R=1.116e+01 
R9599t4172 n9600 n4173 R=1.249e+01 
R9599t6047 n9600 n6048 R=5.208e+00 
R9599t1655 n9600 n1656 R=1.000e+01 
R9600t1602 n9601 n1603 R=4.854e+00 
R9600t2855 n9601 n2856 R=4.440e+00 
R9600t9028 n9601 n9029 R=7.335e+00 
R9600t6519 n9601 n6520 R=9.015e+01 
R9600t3008 n9601 n3009 R=3.019e+00 
R9601t6597 n9602 n6598 R=1.175e+01 
R9601t8215 n9602 n8216 R=4.180e+00 
R9601t7612 n9602 n7613 R=1.036e+01 
R9601t6141 n9602 n6142 R=5.888e+00 
R9602t6384 n9603 n6385 R=5.923e+00 
R9602t9074 n9603 n9075 R=4.777e+00 
R9602t4769 n9603 n4770 R=3.115e+01 
R9602t6188 n9603 n6189 R=3.732e+00 
R9602t4262 n9603 n4263 R=7.172e+00 
R9603t6908 n9604 n6909 R=4.903e+00 
R9603t9432 n9604 n9433 R=2.195e+01 
R9603t8969 n9604 n8970 R=3.387e+01 
R9603t1723 n9604 n1724 R=3.832e+00 
R9603t3028 n9604 n3029 R=1.439e+02 
R9604t806 n9605 n807 R=1.149e+02 
R9604t9170 n9605 n9171 R=2.988e+00 
R9604t384 n9605 n385 R=6.730e+00 
R9604t9078 n9605 n9079 R=6.465e+00 
R9604t8629 n9605 n8630 R=4.389e+01 
R9604t3315 n9605 n3316 R=1.572e+01 
R9604t3003 n9605 n3004 R=1.168e+01 
R9605t7460 n9606 n7461 R=2.774e+00 
R9605t9423 n9606 n9424 R=7.684e+00 
R9605t9279 n9606 n9280 R=4.364e+00 
R9605t3349 n9606 n3350 R=1.866e+01 
R9605t2667 n9606 n2668 R=6.683e+00 
R9606t1388 n9607 n1389 R=5.902e+00 
R9606t6514 n9607 n6515 R=1.636e+01 
R9606t2424 n9607 n2425 R=5.784e+00 
R9606t6624 n9607 n6625 R=2.992e+02 
R9606t7771 n9607 n7772 R=1.118e+01 
R9606t1881 n9607 n1882 R=1.457e+01 
R9606t1572 n9607 n1573 R=4.242e+00 
R9607t5699 n9608 n5700 R=2.611e+01 
R9607t6742 n9608 n6743 R=4.635e+00 
R9607t4114 n9608 n4115 R=8.739e+00 
R9607t6229 n9608 n6230 R=4.998e+00 
R9607t1610 n9608 n1611 R=8.658e+00 
R9607t4967 n9608 n4968 R=9.539e+00 
R9608t527 n9609 n528 R=1.149e+02 
R9608t6848 n9609 n6849 R=6.471e+00 
R9608t4686 n9609 n4687 R=9.250e+00 
R9608t7871 n9609 n7872 R=2.592e+01 
R9608t4026 n9609 n4027 R=9.576e+00 
R9608t6964 n9609 n6965 R=2.943e+00 
R9608t4062 n9609 n4063 R=1.995e+01 
R9609t8548 n9610 n8549 R=1.032e+01 
R9609t9043 n9610 n9044 R=7.119e+00 
R9609t4689 n9610 n4690 R=2.192e+00 
R9609t8165 n9610 n8166 R=4.053e+00 
R9610t3800 n9611 n3801 R=5.508e+00 
R9610t6443 n9611 n6444 R=3.268e+00 
R9610t7058 n9611 n7059 R=8.784e+00 
R9610t5475 n9611 n5476 R=4.196e+01 
R9610t3872 n9611 n3873 R=2.046e+01 
R9610t9269 n9611 n9270 R=8.195e+00 
R9611t3792 n9612 n3793 R=1.290e+01 
R9611t7173 n9612 n7174 R=1.153e+01 
R9611t7950 n9612 n7951 R=2.452e+00 
R9611t8433 n9612 n8434 R=3.856e+02 
R9611t54 n9612 n55 R=2.185e+01 
R9611t161 n9612 n162 R=2.186e+01 
R9611t7163 n9612 n7164 R=4.838e+00 
R9612t3113 n9613 n3114 R=1.015e+01 
R9612t5785 n9613 n5786 R=6.522e+00 
R9612t3391 n9613 n3392 R=1.361e+01 
R9612t9116 n9613 n9117 R=2.029e+00 
R9612t4374 n9613 n4375 R=3.191e+02 
R9612t4793 n9613 n4794 R=6.560e+00 
R9613t72 n9614 n73 R=1.981e+00 
R9613t7034 n9614 n7035 R=9.497e+00 
R9613t1019 n9614 n1020 R=1.437e+01 
R9613t7745 n9614 n7746 R=1.237e+01 
R9613t6575 n9614 n6576 R=4.082e+00 
R9614t5741 n9615 n5742 R=2.758e+00 
R9614t8084 n9615 n8085 R=4.288e+00 
R9614t8580 n9615 n8581 R=5.951e+00 
R9614t1402 n9615 n1403 R=1.118e+01 
R9614t3358 n9615 n3359 R=1.655e+01 
R9615t2843 n9616 n2844 R=2.553e+00 
R9615t8132 n9616 n8133 R=3.197e+00 
R9615t7752 n9616 n7753 R=7.647e+00 
R9615t7224 n9616 n7225 R=2.685e+01 
R9616t886 n9617 n887 R=1.527e+01 
R9616t2820 n9617 n2821 R=2.673e+00 
R9616t4710 n9617 n4711 R=1.912e+01 
R9616t4047 n9617 n4048 R=5.123e+00 
R9616t4907 n9617 n4908 R=2.592e+01 
R9616t6588 n9617 n6589 R=7.760e+00 
R9617t928 n9618 n929 R=5.513e+00 
R9617t5973 n9618 n5974 R=2.243e+01 
R9617t9356 n9618 n9357 R=1.897e+01 
R9617t5093 n9618 n5094 R=6.828e+00 
R9617t2399 n9618 n2400 R=1.625e+01 
R9617t6644 n9618 n6645 R=4.549e+00 
R9618t5833 n9619 n5834 R=8.422e+00 
R9618t8785 n9619 n8786 R=1.488e+01 
R9618t8706 n9619 n8707 R=1.083e+01 
R9618t3132 n9619 n3133 R=1.146e+01 
R9618t2912 n9619 n2913 R=5.028e+00 
R9618t1594 n9619 n1595 R=2.034e+01 
R9618t7306 n9619 n7307 R=7.810e+00 
R9619t2507 n9620 n2508 R=6.108e+00 
R9619t9284 n9620 n9285 R=7.912e+00 
R9619t1947 n9620 n1948 R=1.901e+01 
R9619t7454 n9620 n7455 R=1.611e+01 
R9619t8074 n9620 n8075 R=1.550e+01 
R9619t8386 n9620 n8387 R=2.418e+01 
R9619t3768 n9620 n3769 R=6.967e+00 
R9619t9326 n9620 n9327 R=1.392e+01 
R9620t4062 n9621 n4063 R=1.562e+01 
R9620t4196 n9621 n4197 R=4.480e+00 
R9620t9566 n9621 n9567 R=4.170e+00 
R9620t2853 n9621 n2854 R=1.577e+01 
R9620t796 n9621 n797 R=7.882e+00 
R9620t8977 n9621 n8978 R=3.170e+01 
R9620t527 n9621 n528 R=2.626e+01 
R9621t2651 n9622 n2652 R=8.975e+00 
R9621t6948 n9622 n6949 R=1.375e+01 
R9621t843 n9622 n844 R=2.900e+00 
R9621t8252 n9622 n8253 R=9.932e+00 
R9621t2986 n9622 n2987 R=1.486e+01 
R9621t6979 n9622 n6980 R=6.922e+00 
R9622t2260 n9623 n2261 R=4.904e+00 
R9622t8707 n9623 n8708 R=7.355e+00 
R9622t3650 n9623 n3651 R=4.444e+00 
R9622t739 n9623 n740 R=3.067e+00 
R9623t3196 n9624 n3197 R=4.582e+00 
R9623t3203 n9624 n3204 R=1.318e+01 
R9623t2369 n9624 n2370 R=1.185e+01 
R9623t8724 n9624 n8725 R=2.979e+00 
R9623t112 n9624 n113 R=7.352e+00 
R9623t7862 n9624 n7863 R=1.694e+01 
R9624t2665 n9625 n2666 R=1.740e+01 
R9624t5667 n9625 n5668 R=2.385e+01 
R9624t2189 n9625 n2190 R=3.096e+00 
R9624t934 n9625 n935 R=3.569e+00 
R9625t1493 n9626 n1494 R=6.459e+00 
R9625t2152 n9626 n2153 R=1.034e+01 
R9625t3522 n9626 n3523 R=5.093e+00 
R9625t5276 n9626 n5277 R=4.015e+01 
R9625t4100 n9626 n4101 R=1.054e+01 
R9625t4804 n9626 n4805 R=5.890e+00 
R9625t5544 n9626 n5545 R=6.398e+01 
R9626t2906 n9627 n2907 R=2.280e+01 
R9626t4576 n9627 n4577 R=2.307e+00 
R9626t5015 n9627 n5016 R=2.762e+00 
R9626t7572 n9627 n7573 R=6.917e+00 
R9627t428 n9628 n429 R=5.447e+01 
R9627t2938 n9628 n2939 R=2.059e+00 
R9627t4096 n9628 n4097 R=1.205e+01 
R9627t1929 n9628 n1930 R=3.365e+01 
R9627t856 n9628 n857 R=3.150e+00 
R9627t9265 n9628 n9266 R=2.376e+01 
R9628t711 n9629 n712 R=6.640e+00 
R9628t3034 n9629 n3035 R=6.103e+00 
R9628t9177 n9629 n9178 R=5.888e+00 
R9628t2477 n9629 n2478 R=7.177e+00 
R9629t5009 n9630 n5010 R=9.027e+00 
R9629t6065 n9630 n6066 R=4.392e+01 
R9629t3089 n9630 n3090 R=6.013e+00 
R9629t7709 n9630 n7710 R=7.599e+00 
R9629t1399 n9630 n1400 R=1.627e+01 
R9629t8613 n9630 n8614 R=1.181e+01 
R9629t1730 n9630 n1731 R=3.401e+01 
R9629t3378 n9630 n3379 R=4.717e+00 
R9630t4013 n9631 n4014 R=1.458e+01 
R9630t5408 n9631 n5409 R=1.447e+03 
R9630t8688 n9631 n8689 R=6.025e+00 
R9630t2410 n9631 n2411 R=4.703e+00 
R9630t7288 n9631 n7289 R=4.471e+00 
R9630t6591 n9631 n6592 R=7.319e+00 
R9631t6454 n9632 n6455 R=7.002e+00 
R9631t6994 n9632 n6995 R=1.694e+01 
R9631t3227 n9632 n3228 R=8.719e+00 
R9631t8890 n9632 n8891 R=4.020e+00 
R9631t3569 n9632 n3570 R=1.883e+02 
R9631t6079 n9632 n6080 R=1.214e+01 
R9631t6608 n9632 n6609 R=2.474e+01 
R9632t7868 n9633 n7869 R=1.363e+01 
R9632t8394 n9633 n8395 R=4.893e+01 
R9632t572 n9633 n573 R=8.106e+00 
R9632t749 n9633 n750 R=4.346e+00 
R9632t2723 n9633 n2724 R=6.283e+00 
R9632t6709 n9633 n6710 R=6.954e+01 
R9632t2355 n9633 n2356 R=4.803e+00 
R9633t1699 n9634 n1700 R=3.703e+00 
R9633t4467 n9634 n4468 R=8.419e+00 
R9633t6116 n9634 n6117 R=1.043e+02 
R9633t6653 n9634 n6654 R=2.761e+00 
R9633t5856 n9634 n5857 R=2.116e+01 
R9634t573 n9635 n574 R=9.702e+00 
R9634t9343 n9635 n9344 R=1.617e+01 
R9634t3239 n9635 n3240 R=5.697e+00 
R9634t5887 n9635 n5888 R=6.608e+00 
R9634t5757 n9635 n5758 R=5.107e+00 
R9634t3170 n9635 n3171 R=1.427e+01 
R9635t1329 n9636 n1330 R=5.602e+00 
R9635t9327 n9636 n9328 R=9.746e+00 
R9635t9206 n9636 n9207 R=5.042e+00 
R9635t4012 n9636 n4013 R=8.892e+00 
R9635t7712 n9636 n7713 R=2.945e+01 
R9635t5572 n9636 n5573 R=4.281e+00 
R9636t5332 n9637 n5333 R=1.220e+01 
R9636t7905 n9637 n7906 R=1.526e+01 
R9636t5809 n9637 n5810 R=2.265e+00 
R9636t7296 n9637 n7297 R=1.600e+02 
R9636t8856 n9637 n8857 R=1.659e+02 
R9636t8285 n9637 n8286 R=3.465e+00 
R9637t3702 n9638 n3703 R=3.640e+00 
R9637t7043 n9638 n7044 R=1.620e+01 
R9637t7603 n9638 n7604 R=4.153e+00 
R9637t4009 n9638 n4010 R=2.828e+01 
R9637t268 n9638 n269 R=7.786e+00 
R9638t6214 n9639 n6215 R=4.560e+00 
R9638t7915 n9639 n7916 R=9.734e+00 
R9638t6915 n9639 n6916 R=1.428e+01 
R9638t4255 n9639 n4256 R=1.337e+01 
R9638t1793 n9639 n1794 R=5.284e+00 
R9639t7983 n9640 n7984 R=6.028e+00 
R9639t9544 n9640 n9545 R=4.889e+01 
R9639t7647 n9640 n7648 R=9.234e+00 
R9639t1448 n9640 n1449 R=3.154e+00 
R9639t7890 n9640 n7891 R=1.160e+01 
R9639t8364 n9640 n8365 R=1.380e+01 
R9640t551 n9641 n552 R=4.671e+00 
R9640t683 n9641 n684 R=8.799e+00 
R9640t480 n9641 n481 R=8.478e+01 
R9640t82 n9641 n83 R=9.168e+00 
R9640t8177 n9641 n8178 R=8.736e+00 
R9640t1840 n9641 n1841 R=5.136e+00 
R9640t6018 n9641 n6019 R=7.838e+01 
R9641t387 n9642 n388 R=1.507e+01 
R9641t1942 n9642 n1943 R=3.922e+00 
R9641t1456 n9642 n1457 R=3.236e+01 
R9641t3108 n9642 n3109 R=4.961e+00 
R9641t7496 n9642 n7497 R=8.075e+00 
R9641t3263 n9642 n3264 R=6.131e+00 
R9642t2872 n9643 n2873 R=1.110e+01 
R9642t3869 n9643 n3870 R=2.458e+00 
R9642t2568 n9643 n2569 R=2.156e+01 
R9642t6914 n9643 n6915 R=2.581e+00 
R9643t830 n9644 n831 R=4.548e+00 
R9643t6521 n9644 n6522 R=5.857e+00 
R9643t7500 n9644 n7501 R=1.756e+02 
R9643t7812 n9644 n7813 R=6.194e+00 
R9643t9225 n9644 n9226 R=2.930e+00 
R9643t5258 n9644 n5259 R=3.158e+01 
R9644t3476 n9645 n3477 R=4.798e+00 
R9644t7138 n9645 n7139 R=1.316e+02 
R9644t4042 n9645 n4043 R=5.740e+00 
R9644t9510 n9645 n1 R=6.528e+00 
R9644t42 n9645 n43 R=6.790e+00 
R9644t9212 n9645 n9213 R=7.381e+01 
R9645t1176 n9646 n1177 R=7.135e+00 
R9645t2176 n9646 n2177 R=8.837e+00 
R9645t6102 n9646 n6103 R=3.632e+00 
R9645t7251 n9646 n7252 R=1.516e+01 
R9645t1691 n9646 n1692 R=7.267e+00 
R9646t4635 n9647 n4636 R=1.642e+00 
R9646t6256 n9647 n6257 R=2.723e+00 
R9646t1165 n9647 n1166 R=5.947e+00 
R9647t5254 n9648 n5255 R=3.906e+00 
R9647t6774 n9648 n6775 R=4.496e+00 
R9647t7922 n9648 n7923 R=4.569e+01 
R9647t5646 n9648 n5647 R=4.393e+00 
R9648t3638 n9649 n3639 R=3.469e+00 
R9648t8427 n9649 n8428 R=6.590e+00 
R9648t2738 n9649 n2739 R=5.414e+01 
R9648t3356 n9649 n3357 R=3.779e+00 
R9648t1727 n9649 n1 R=9.791e+01 
R9648t2063 n9649 n1 R=5.215e+00 
R9649t2282 n9650 n2283 R=3.178e+01 
R9649t4959 n9650 n4960 R=1.628e+01 
R9649t1972 n9650 n1973 R=6.911e+00 
R9649t8793 n9650 n8794 R=2.230e+00 
R9649t5181 n9650 n5182 R=3.376e+01 
R9649t3818 n9650 n3819 R=9.069e+00 
R9649t1139 n9650 n1140 R=1.720e+01 
R9650t9432 n9651 n9433 R=1.053e+01 
R9650t9603 n9651 n9604 R=5.127e+00 
R9650t3028 n9651 n3029 R=6.563e+00 
R9650t6752 n9651 n6753 R=9.884e+00 
R9650t2317 n9651 n2318 R=1.612e+01 
R9650t3183 n9651 n3184 R=3.800e+00 
R9651t2463 n9652 n2464 R=1.851e+01 
R9651t7701 n9652 n7702 R=6.335e+00 
R9651t9007 n9652 n9008 R=5.644e+00 
R9651t1220 n9652 n1221 R=2.015e+01 
R9651t4633 n9652 n4634 R=2.181e+00 
R9651t5512 n9652 n5513 R=5.422e+01 
R9652t3061 n9653 n3062 R=1.140e+01 
R9652t7897 n9653 n7898 R=1.471e+01 
R9652t764 n9653 n765 R=2.283e+00 
R9652t8895 n9653 n8896 R=1.230e+01 
R9652t914 n9653 n915 R=7.303e+01 
R9652t7698 n9653 n7699 R=4.251e+00 
R9653t1729 n9654 n1730 R=6.366e+00 
R9653t8596 n9654 n8597 R=2.534e+00 
R9653t4181 n9654 n4182 R=3.123e+00 
R9654t7747 n9655 n7748 R=2.016e+03 
R9654t8957 n9655 n8958 R=4.746e+00 
R9654t5086 n9655 n5087 R=4.880e+00 
R9654t3833 n9655 n3834 R=4.118e+01 
R9654t2342 n9655 n2343 R=1.043e+01 
R9654t8581 n9655 n8582 R=4.605e+00 
R9654t5741 n9655 n5742 R=4.376e+01 
R9655t665 n9656 n666 R=1.068e+02 
R9655t8643 n9656 n8644 R=6.923e+00 
R9655t325 n9656 n326 R=5.894e+00 
R9655t6259 n9656 n6260 R=5.922e+00 
R9655t5961 n9656 n5962 R=4.073e+00 
R9655t6357 n9656 n6358 R=2.656e+01 
R9656t2131 n9657 n2132 R=3.405e+00 
R9656t4950 n9657 n4951 R=3.431e+00 
R9656t5447 n9657 n5448 R=3.190e+01 
R9656t7217 n9657 n7218 R=2.413e+00 
R9656t5373 n9657 n5374 R=3.436e+01 
R9657t982 n9658 n983 R=4.531e+00 
R9657t7208 n9658 n7209 R=3.843e+00 
R9657t1568 n9658 n1569 R=3.108e+00 
R9658t3565 n9659 n3566 R=2.499e+00 
R9658t4598 n9659 n4599 R=5.681e+00 
R9658t5363 n9659 n5364 R=8.208e+00 
R9658t1979 n9659 n1980 R=6.602e+00 
R9659t3472 n9660 n3473 R=5.860e+00 
R9659t4493 n9660 n4494 R=2.547e+01 
R9659t7105 n9660 n7106 R=1.204e+01 
R9659t8921 n9660 n8922 R=9.456e+00 
R9659t4827 n9660 n4828 R=8.102e+00 
R9659t4427 n9660 n4428 R=6.902e+00 
R9659t2066 n9660 n2067 R=4.124e+01 
R9660t2143 n9661 n2144 R=3.566e+00 
R9660t7278 n9661 n7279 R=6.296e+00 
R9660t423 n9661 n424 R=1.228e+01 
R9660t6291 n9661 n6292 R=3.510e+01 
R9660t2404 n9661 n2405 R=3.344e+00 
R9660t6708 n9661 n6709 R=1.688e+01 
R9660t8125 n9661 n8126 R=2.538e+01 
R9661t1109 n9662 n1110 R=2.212e+00 
R9661t5710 n9662 n5711 R=1.062e+02 
R9661t9016 n9662 n9017 R=5.444e+00 
R9661t9164 n9662 n9165 R=3.316e+00 
R9661t303 n9662 n304 R=1.753e+01 
R9662t653 n9663 n654 R=1.718e+01 
R9662t6101 n9663 n6102 R=1.625e+00 
R9662t4285 n9663 n4286 R=2.234e+02 
R9662t9459 n9663 n9460 R=9.486e+01 
R9662t867 n9663 n868 R=1.258e+01 
R9662t8617 n9663 n8618 R=3.924e+00 
R9663t2786 n9664 n2787 R=6.763e+00 
R9663t6463 n9664 n6464 R=1.535e+01 
R9663t172 n9664 n173 R=3.065e+00 
R9663t4744 n9664 n4745 R=1.098e+01 
R9663t9461 n9664 n9462 R=9.384e+00 
R9663t5548 n9664 n5549 R=2.596e+01 
R9663t7431 n9664 n7432 R=9.232e+01 
R9664t2558 n9665 n2559 R=1.268e+01 
R9664t4305 n9665 n4306 R=3.664e+00 
R9664t2653 n9665 n2654 R=8.250e+00 
R9664t6044 n9665 n6045 R=8.160e+00 
R9664t2392 n9665 n2393 R=2.740e+01 
R9664t1927 n9665 n1928 R=5.526e+00 
R9665t5082 n9666 n5083 R=4.104e+00 
R9665t9102 n9666 n9103 R=1.743e+01 
R9665t8875 n9666 n8876 R=2.564e+01 
R9665t9458 n9666 n9459 R=9.127e+00 
R9665t9296 n9666 n9297 R=6.813e+00 
R9665t1090 n9666 n1091 R=2.049e+01 
R9665t1967 n9666 n1968 R=8.619e+00 
R9665t7304 n9666 n7305 R=1.130e+01 
R9666t1436 n9667 n1437 R=2.964e+00 
R9666t7540 n9667 n7541 R=1.070e+02 
R9667t1026 n9668 n1027 R=1.315e+01 
R9667t3165 n9668 n3166 R=2.581e+01 
R9667t3730 n9668 n3731 R=8.453e+00 
R9667t3185 n9668 n3186 R=3.158e+00 
R9667t9557 n9668 n9558 R=3.106e+00 
R9668t331 n9669 n332 R=5.846e+00 
R9668t582 n9669 n583 R=7.195e+01 
R9668t1016 n9669 n1017 R=2.381e+01 
R9668t8447 n9669 n8448 R=2.331e+00 
R9668t6299 n9669 n6300 R=2.122e+02 
R9668t4610 n9669 n4611 R=2.504e+01 
R9668t7758 n9669 n7759 R=3.938e+00 
R9669t565 n9670 n566 R=1.984e+02 
R9669t6961 n9670 n6962 R=1.486e+01 
R9669t8118 n9670 n8119 R=4.105e+00 
R9669t6525 n9670 n6526 R=1.075e+01 
R9669t5058 n9670 n5059 R=1.164e+01 
R9669t5288 n9670 n5289 R=1.208e+01 
R9669t4098 n9670 n4099 R=2.608e+01 
R9669t425 n9670 n426 R=5.984e+00 
R9670t2141 n9671 n2142 R=7.040e+00 
R9670t3169 n9671 n3170 R=1.386e+01 
R9670t7542 n9671 n7543 R=7.132e+00 
R9670t7471 n9671 n7472 R=2.981e+00 
R9670t9418 n9671 n9419 R=6.063e+00 
R9670t2422 n9671 n2423 R=5.590e+01 
R9671t4871 n9672 n4872 R=3.796e+00 
R9671t6938 n9672 n6939 R=8.644e+00 
R9671t4466 n9672 n4467 R=1.955e+00 
R9671t2611 n9672 n2612 R=1.455e+01 
R9672t8734 n9673 n8735 R=3.156e+00 
R9672t8745 n9673 n8746 R=1.013e+01 
R9672t3680 n9673 n3681 R=1.797e+01 
R9672t6475 n9673 n6476 R=2.876e+00 
R9672t7871 n9673 n7872 R=9.446e+00 
R9673t3613 n9674 n3614 R=6.274e+00 
R9673t3625 n9674 n3626 R=1.591e+01 
R9673t827 n9674 n828 R=1.876e+01 
R9673t6897 n9674 n6898 R=2.658e+01 
R9673t1521 n9674 n1522 R=8.656e+00 
R9673t6365 n9674 n6366 R=2.712e+01 
R9673t4122 n9674 n4123 R=1.485e+01 
R9673t7487 n9674 n7488 R=1.138e+01 
R9673t6127 n9674 n6128 R=9.729e+00 
R9674t669 n9675 n670 R=4.601e+00 
R9674t7184 n9675 n7185 R=1.077e+01 
R9674t1141 n9675 n1142 R=5.008e+00 
R9674t1820 n9675 n1821 R=1.946e+01 
R9674t1905 n9675 n1906 R=1.244e+01 
R9674t3400 n9675 n3401 R=3.980e+01 
R9675t6309 n9676 n6310 R=7.914e+00 
R9675t8128 n9676 n8129 R=1.728e+01 
R9675t4974 n9676 n4975 R=5.198e+00 
R9675t1935 n9676 n1936 R=8.609e+00 
R9675t8864 n9676 n8865 R=7.613e+00 
R9675t6741 n9676 n6742 R=1.005e+02 
R9675t6362 n9676 n6363 R=6.921e+00 
R9676t784 n9677 n785 R=2.749e+01 
R9676t5028 n9677 n5029 R=4.056e+00 
R9676t8315 n9677 n8316 R=2.630e+00 
R9676t3762 n9677 n3763 R=1.778e+01 
R9676t3175 n9677 n3176 R=9.307e+00 
R9676t3980 n9677 n3981 R=6.302e+00 
R9677t2457 n9678 n2458 R=6.018e+01 
R9677t4031 n9678 n4032 R=2.170e+00 
R9677t5515 n9678 n5516 R=4.884e+01 
R9677t2255 n9678 n2256 R=3.283e+00 
R9677t4435 n9678 n4436 R=1.102e+01 
R9677t4901 n9678 n4902 R=1.411e+01 
R9678t4779 n9679 n4780 R=6.076e+00 
R9678t7150 n9679 n7151 R=5.635e+01 
R9678t8356 n9679 n8357 R=4.574e+01 
R9678t3669 n9679 n3670 R=8.613e+00 
R9678t3365 n9679 n3366 R=6.059e+00 
R9678t7679 n9679 n7680 R=1.027e+01 
R9678t2745 n9679 n2746 R=4.161e+00 
R9679t3874 n9680 n3875 R=7.690e+01 
R9679t4170 n9680 n4171 R=2.303e+01 
R9679t9578 n9680 n9579 R=8.225e+01 
R9679t1555 n9680 n1556 R=3.671e+00 
R9679t5237 n9680 n5238 R=2.231e+01 
R9679t670 n9680 n671 R=4.937e+00 
R9679t2125 n9680 n2126 R=8.598e+00 
R9679t5721 n9680 n5722 R=8.208e+00 
R9680t2154 n9681 n2155 R=6.840e+01 
R9680t3947 n9681 n3948 R=2.125e+00 
R9680t7625 n9681 n7626 R=8.132e+01 
R9680t9572 n9681 n9573 R=2.730e+01 
R9680t7458 n9681 n7459 R=2.981e+00 
R9680t1620 n9681 n1621 R=4.708e+00 
R9681t5116 n9682 n5117 R=4.814e+00 
R9681t6434 n9682 n6435 R=3.531e+00 
R9681t6835 n9682 n6836 R=1.895e+01 
R9681t8293 n9682 n8294 R=7.582e+00 
R9681t9367 n9682 n9368 R=5.783e+00 
R9681t1870 n9682 n1871 R=5.187e+01 
R9681t4169 n9682 n4170 R=7.717e+01 
R9682t3385 n9683 n3386 R=9.580e+00 
R9682t7905 n9683 n7906 R=1.842e+00 
R9682t5332 n9683 n5333 R=4.808e+01 
R9682t2854 n9683 n2855 R=2.752e+02 
R9682t8183 n9683 n8184 R=1.452e+01 
R9682t7519 n9683 n7520 R=4.367e+00 
R9682t4937 n9683 n4938 R=1.120e+01 
R9683t6532 n9684 n6533 R=1.312e+01 
R9683t8463 n9684 n8464 R=3.883e+00 
R9683t37 n9684 n38 R=1.725e+01 
R9683t9034 n9684 n9035 R=3.217e+01 
R9683t6911 n9684 n6912 R=1.421e+01 
R9683t6617 n9684 n6618 R=2.308e+00 
R9683t4405 n9684 n4406 R=1.709e+01 
R9683t8836 n9684 n8837 R=4.418e+01 
R9684t5300 n9685 n5301 R=2.003e+01 
R9684t5493 n9685 n5494 R=6.917e+00 
R9684t1609 n9685 n1610 R=2.004e+01 
R9684t8062 n9685 n8063 R=1.241e+01 
R9684t4866 n9685 n4867 R=1.116e+01 
R9684t1138 n9685 n1139 R=3.119e+00 
R9685t3521 n9686 n3522 R=4.131e+00 
R9685t6381 n9686 n6382 R=5.439e+00 
R9685t8578 n9686 n8579 R=3.537e+00 
R9685t9311 n9686 n9312 R=3.370e+01 
R9685t4293 n9686 n4294 R=6.160e+00 
R9685t2602 n9686 n2603 R=1.881e+01 
R9686t286 n9687 n287 R=1.938e+00 
R9686t6219 n9687 n6220 R=7.790e+01 
R9686t1553 n9687 n1554 R=3.227e+01 
R9686t3549 n9687 n3550 R=5.788e+01 
R9686t8165 n9687 n8166 R=2.516e+00 
R9686t8548 n9687 n8549 R=2.368e+01 
R9686t2574 n9687 n2575 R=2.561e+01 
R9687t4522 n9688 n4523 R=1.479e+01 
R9687t4888 n9688 n4889 R=5.155e+00 
R9687t5787 n9688 n5788 R=7.304e+00 
R9687t5396 n9688 n5397 R=2.884e+00 
R9687t210 n9688 n211 R=1.361e+01 
R9688t5638 n9689 n5639 R=3.868e+01 
R9688t6517 n9689 n6518 R=6.601e+00 
R9688t496 n9689 n497 R=7.990e+00 
R9688t1922 n9689 n1923 R=4.362e+01 
R9688t3912 n9689 n3913 R=4.305e+00 
R9688t4590 n9689 n4591 R=6.061e+00 
R9688t4776 n9689 n4777 R=9.510e+00 
R9689t2480 n9690 n2481 R=2.540e+00 
R9689t8889 n9690 n8890 R=3.081e+01 
R9689t1288 n9690 n1289 R=1.238e+01 
R9689t83 n9690 n84 R=2.256e+00 
R9689t1451 n9690 n1452 R=7.439e+00 
R9690t4163 n9691 n4164 R=2.702e+00 
R9690t6346 n9691 n6347 R=3.265e+01 
R9690t3589 n9691 n3590 R=1.225e+01 
R9690t2534 n9691 n2535 R=4.514e+00 
R9690t8243 n9691 n8244 R=2.480e+03 
R9690t103 n9691 n104 R=9.267e+00 
R9691t7987 n9692 n7988 R=3.917e+00 
R9691t8043 n9692 n8044 R=4.362e+01 
R9691t8117 n9692 n8118 R=1.248e+01 
R9691t3326 n9692 n3327 R=5.049e+00 
R9691t1425 n9692 n1426 R=6.250e+00 
R9692t1183 n9693 n1184 R=6.998e+00 
R9692t5073 n9693 n5074 R=6.244e+01 
R9692t1703 n9693 n1704 R=6.321e+00 
R9692t5758 n9693 n5759 R=9.343e+01 
R9692t851 n9693 n852 R=5.321e+00 
R9692t7032 n9693 n7033 R=1.111e+01 
R9692t3395 n9693 n3396 R=2.765e+01 
R9692t6076 n9693 n6077 R=8.516e+00 
R9693t1229 n9694 n1230 R=3.013e+00 
R9693t6280 n9694 n6281 R=1.375e+01 
R9693t5929 n9694 n5930 R=7.085e+00 
R9693t6391 n9694 n6392 R=2.833e+00 

*** contact connections

*** simulation 
*.op 
*.dc Vdd 0 1 0.02 
.dc Vdd 0 0 0.02 

*** options 

.print DC v(n1) i(Vdd) V(n1) V(n2) V(n3) V(n4) V(n5) V(n6) V(n7) V(n8) V(n9) V(n10) V(n11) V(n12) V(n13) V(n14) V(n15) V(n16) V(n17) V(n18) V(n19) V(n20) V(n21) V(n22) V(n23) V(n24) V(n25) V(n26) V(n27) V(n28) V(n29) V(n30) V(n31) V(n32) V(n33) V(n34) V(n35) V(n36) V(n37) V(n38) V(n39) V(n40) V(n41) V(n42) V(n43) V(n44) V(n45) V(n46) V(n47) V(n48) V(n49) V(n50) V(n51) V(n52) V(n53) V(n54) V(n55) V(n56) V(n57) V(n58) V(n59) V(n60) V(n61) V(n62) V(n63) V(n64) V(n65) V(n66) V(n67) V(n68) V(n69) V(n70) V(n71) V(n72) V(n73) V(n74) V(n75) V(n76) V(n77) V(n78) V(n79) V(n80) V(n81) V(n82) V(n83) V(n84) V(n85) V(n86) V(n87) V(n88) V(n89) V(n90) V(n91) V(n92) V(n93) V(n94) V(n95) V(n96) V(n97) V(n98) V(n99) V(n100) V(n101) V(n102) V(n103) V(n104) V(n105) V(n106) V(n107) V(n108) V(n109) V(n110) V(n111) V(n112) V(n113) V(n114) V(n115) V(n116) V(n117) V(n118) V(n119) V(n120) V(n121) V(n122) V(n123) V(n124) V(n125) V(n126) V(n127) V(n128) V(n129) V(n130) V(n131) V(n132) V(n133) V(n134) V(n135) V(n136) V(n137) V(n138) V(n139) V(n140) V(n141) V(n142) V(n143) V(n144) V(n145) V(n146) V(n147) V(n148) V(n149) V(n150) V(n151) V(n152) V(n153) V(n154) V(n155) V(n156) V(n157) V(n158) V(n159) V(n160) V(n161) V(n162) V(n163) V(n164) V(n165) V(n166) V(n167) V(n168) V(n169) V(n170) V(n171) V(n172) V(n173) V(n174) V(n1) V(n176) V(n177) V(n178) V(n179) V(n180) V(n181) V(n182) V(n183) V(n184) V(n185) V(n186) V(n187) V(n188) V(n189) V(n190) V(n191) V(n192) V(n193) V(n194) V(n195) V(n196) V(n197) V(n198) V(n199) V(n200) V(n201) V(n202) V(n203) V(n204) V(n205) V(n206) V(n207) V(n208) V(n209) V(n210) V(n211) V(n212) V(n213) V(n214) V(n215) V(n216) V(n217) V(n218) V(n219) V(n220) V(n221) V(n222) V(n223) V(n224) V(n225) V(n226) V(n227) V(n228) V(n229) V(n230) V(n231) V(n1) V(n233) V(n234) V(n235) V(n236) V(n237) V(n238) V(n239) V(n240) V(n241) V(n242) V(n243) V(n244) V(n245) V(n246) V(n247) V(n248) V(n249) V(n250) V(n251) V(n252) V(n253) V(n254) V(n255) V(n256) V(n257) V(n258) V(n259) V(n260) V(n261) V(n262) V(n263) V(n264) V(n265) V(n266) V(n267) V(n268) V(n269) V(n270) V(n271) V(n272) V(n273) V(n274) V(n275) V(n276) V(n277) V(n278) V(n1) V(n280) V(n281) V(n282) V(n283) V(n284) V(n285) V(n286) V(n287) V(n288) V(n289) V(n290) V(n291) V(n292) V(n293) V(n294) V(n295) V(n296) V(n297) V(n298) V(n299) V(n300) V(n301) V(n302) V(n303) V(n304) V(n305) V(n306) V(n307) V(n308) V(n309) V(n310) V(n311) V(n312) V(n313) V(n314) V(n315) V(n1) V(n317) V(n318) V(n319) V(n320) V(n321) V(n322) V(n323) V(n324) V(n325) V(n326) V(n327) V(n328) V(n329) V(n330) V(n331) V(n332) V(n333) V(n334) V(n335) V(n336) V(n337) V(n338) V(n339) V(n340) V(n341) V(n342) V(n343) V(n344) V(n345) V(n346) V(n347) V(n348) V(n349) V(n350) V(n351) V(n352) V(n353) V(n354) V(n355) V(n356) V(n357) V(n358) V(n359) V(n360) V(n361) V(n362) V(n363) V(n364) V(n365) V(n366) V(n367) V(n368) V(n369) V(n370) V(n371) V(n372) V(n373) V(n374) V(n375) V(n376) V(n377) V(n378) V(n379) V(n380) V(n381) V(n382) V(n383) V(n384) V(n385) V(n386) V(n387) V(n388) V(n389) V(n390) V(n391) V(n392) V(n393) V(n394) V(n395) V(n396) V(n397) V(n398) V(n1) V(n400) V(n401) V(n402) V(n403) V(n404) V(n405) V(n406) V(n407) V(n408) V(n409) V(n410) V(n411) V(n412) V(n413) V(n414) V(n415) V(n416) V(n417) V(n418) V(n419) V(n420) V(n421) V(n422) V(n423) V(n424) V(n425) V(n426) V(n427) V(n428) V(n429) V(n430) V(n431) V(n432) V(n433) V(n434) V(n435) V(n436) V(n437) V(n438) V(n439) V(n440) V(n441) V(n442) V(n443) V(n444) V(n445) V(n446) V(n447) V(n448) V(n449) V(n450) V(n451) V(n452) V(n453) V(n454) V(n455) V(n456) V(n457) V(n458) V(n459) V(n460) V(n461) V(n462) V(n463) V(n464) V(n465) V(n466) V(n467) V(n468) V(n469) V(n470) V(n471) V(n472) V(n473) V(n474) V(n475) V(n476) V(n477) V(n478) V(n479) V(n480) V(n481) V(n482) V(n483) V(n1) V(n485) V(n486) V(n487) V(n488) V(n489) V(n490) V(n491) V(n492) V(n493) V(n494) V(n495) V(n496) V(n497) V(n498) V(n499) V(n500) V(n501) V(n502) V(n503) V(n504) V(n505) V(n506) V(n507) V(n508) V(n509) V(n510) V(n511) V(n512) V(n513) V(n514) V(n515) V(n516) V(n517) V(n518) V(n519) V(n520) V(n521) V(n522) V(n523) V(n524) V(n525) V(n526) V(n527) V(n528) V(n529) V(n530) V(n531) V(n532) V(n533) V(n534) V(n535) V(n536) V(n537) V(n538) V(n539) V(n540) V(n541) V(n542) V(n543) V(n544) V(n545) V(n546) V(n547) V(n548) V(n549) V(n550) V(n551) V(n552) V(n553) V(n554) V(n555) V(n556) V(n557) V(n558) V(n559) V(n560) V(n561) V(n562) V(n563) V(n564) V(n565) V(n566) V(n567) V(n568) V(n569) V(n570) V(n571) V(n572) V(n573) V(n574) V(n575) V(n576) V(n577) V(n578) V(n579) V(n580) V(n581) V(n582) V(n583) V(n584) V(n585) V(n586) V(n587) V(n588) V(n589) V(n590) V(n591) V(n592) V(n593) V(n594) V(n595) V(n596) V(n597) V(n598) V(n599) V(n600) V(n601) V(n602) V(n603) V(n604) V(n605) V(n606) V(n607) V(n608) V(n609) V(n610) V(n611) V(n612) V(n613) V(n614) V(n615) V(n616) V(n617) V(n618) V(n619) V(n620) V(n621) V(n622) V(n623) V(n624) V(n625) V(n626) V(n627) V(n628) V(n629) V(n630) V(n631) V(n632) V(n633) V(n634) V(n635) V(n636) V(n637) V(n638) V(n639) V(n640) V(n641) V(n642) V(n643) V(n644) V(n645) V(n646) V(n647) V(n648) V(n649) V(n650) V(n651) V(n652) V(n653) V(n654) V(n655) V(n656) V(n657) V(n658) V(n659) V(n660) V(n661) V(n662) V(n663) V(n664) V(n665) V(n666) V(n667) V(n668) V(n669) V(n670) V(n671) V(n672) V(n673) V(n674) V(n675) V(n676) V(n677) V(n678) V(n679) V(n680) V(n681) V(n682) V(n683) V(n684) V(n685) V(n686) V(n687) V(n688) V(n689) V(n690) V(n691) V(n692) V(n1) V(n694) V(n695) V(n696) V(n697) V(n698) V(n699) V(n700) V(n701) V(n702) V(n703) V(n704) V(n705) V(n706) V(n707) V(n708) V(n709) V(n710) V(n711) V(n712) V(n713) V(n714) V(n715) V(n716) V(n717) V(n718) V(n719) V(n720) V(n721) V(n722) V(n723) V(n724) V(n725) V(n726) V(n727) V(n728) V(n729) V(n730) V(n731) V(n732) V(n733) V(n734) V(n735) V(n736) V(n737) V(n738) V(n739) V(n740) V(n741) V(n742) V(n743) V(n744) V(n745) V(n746) V(n747) V(n748) V(n749) V(n750) V(n751) V(n752) V(n753) V(n754) V(n755) V(n756) V(n757) V(n758) V(n759) V(n760) V(n761) V(n762) V(n763) V(n764) V(n765) V(n766) V(n767) V(n768) V(n769) V(n770) V(n771) V(n772) V(n773) V(n774) V(n775) V(n776) V(n777) V(n778) V(n779) V(n780) V(n781) V(n782) V(n783) V(n784) V(n785) V(n786) V(n787) V(n788) V(n789) V(n790) V(n791) V(n792) V(n793) V(n794) V(n795) V(n796) V(n797) V(n798) V(n799) V(n800) V(n801) V(n802) V(n803) V(n804) V(n805) V(n806) V(n807) V(n808) V(n809) V(n810) V(n811) V(n812) V(n813) V(n814) V(n815) V(n816) V(n817) V(n818) V(n819) V(n820) V(n821) V(n822) V(n823) V(n824) V(n825) V(n826) V(n827) V(n828) V(n829) V(n830) V(n831) V(n832) V(n833) V(n834) V(n835) V(n836) V(n837) V(n838) V(n839) V(n840) V(n841) V(n842) V(n843) V(n844) V(n845) V(n846) V(n847) V(n848) V(n849) V(n850) V(n851) V(n852) V(n853) V(n854) V(n855) V(n856) V(n857) V(n858) V(n859) V(n860) V(n861) V(n862) V(n863) V(n864) V(n865) V(n866) V(n867) V(n868) V(n869) V(n870) V(n871) V(n872) V(n873) V(n874) V(n875) V(n876) V(n877) V(n878) V(n879) V(n880) V(n881) V(n882) V(n883) V(n884) V(n885) V(n886) V(n887) V(n888) V(n889) V(n890) V(n891) V(n892) V(n893) V(n894) V(n895) V(n896) V(n897) V(n1) V(n899) V(n900) V(n901) V(n902) V(n903) V(n904) V(n905) V(n906) V(n907) V(n908) V(n909) V(n910) V(n911) V(n912) V(n913) V(n914) V(n915) V(n916) V(n917) V(n918) V(n919) V(n920) V(n921) V(n922) V(n923) V(n924) V(n925) V(n926) V(n927) V(n928) V(n929) V(n930) V(n931) V(n932) V(n933) V(n934) V(n935) V(n936) V(n937) V(n938) V(n939) V(n940) V(n941) V(n942) V(n943) V(n944) V(n945) V(n946) V(n947) V(n948) V(n949) V(n950) V(n951) V(n952) V(n953) V(n954) V(n955) V(n956) V(n957) V(n958) V(n959) V(n960) V(n961) V(n962) V(n963) V(n964) V(n965) V(n966) V(n967) V(n968) V(n969) V(n970) V(n971) V(n972) V(n973) V(n974) V(n975) V(n976) V(n977) V(n978) V(n979) V(n980) V(n981) V(n982) V(n983) V(n984) V(n985) V(n986) V(n987) V(n988) V(n989) V(n990) V(n991) V(n992) V(n993) V(n994) V(n995) V(n996) V(n997) V(n998) V(n999) V(n1000) V(n1001) V(n1002) V(n1003) V(n1004) V(n1005) V(n1006) V(n1007) V(n1008) V(n1009) V(n1010) V(n1011) V(n1012) V(n1013) V(n1014) V(n1015) V(n1016) V(n1017) V(n1018) V(n1019) V(n1020) V(n1021) V(n1022) V(n1023) V(n1024) V(n1025) V(n1026) V(n1027) V(n1028) V(n1029) V(n1030) V(n1031) V(n1032) V(n1033) V(n1034) V(n1035) V(n1036) V(n1037) V(n1038) V(n1039) V(n1040) V(n1041) V(n1042) V(n1043) V(n1044) V(n1045) V(n1046) V(n1047) V(n1048) V(n1049) V(n1050) V(n1051) V(n1052) V(n1053) V(n1054) V(n1055) V(n1056) V(n1057) V(n1058) V(n1059) V(n1060) V(n1061) V(n1062) V(n1063) V(n1064) V(n1065) V(n1066) V(n1067) V(n1068) V(n1069) V(n1070) V(n1071) V(n1072) V(n1073) V(n1074) V(n1075) V(n1076) V(n1077) V(n1078) V(n1079) V(n1080) V(n1081) V(n1082) V(n1083) V(n1084) V(n1085) V(n1086) V(n1087) V(n1088) V(n1089) V(n1090) V(n1091) V(n1092) V(n1093) V(n1094) V(n1095) V(n1096) V(n1097) V(n1098) V(n1099) V(n1100) V(n1101) V(n1102) V(n1103) V(n1104) V(n1105) V(n1106) V(n1107) V(n1108) V(n1109) V(n1110) V(n1111) V(n1112) V(n1113) V(n1114) V(n1115) V(n1116) V(n1117) V(n1118) V(n1119) V(n1120) V(n1121) V(n1122) V(n1123) V(n1124) V(n1125) V(n1126) V(n1127) V(n1128) V(n1129) V(n1130) V(n1131) V(n1132) V(n1133) V(n1134) V(n1135) V(n1136) V(n1137) V(n1138) V(n1139) V(n1140) V(n1141) V(n1142) V(n1143) V(n1144) V(n1145) V(n1146) V(n1147) V(n1148) V(n1149) V(n1150) V(n1151) V(n1152) V(n1153) V(n1154) V(n1) V(n1156) V(n1157) V(n1158) V(n1159) V(n1160) V(n1161) V(n1162) V(n1163) V(n1164) V(n1165) V(n1166) V(n1167) V(n1168) V(n1169) V(n1170) V(n1171) V(n1172) V(n1173) V(n1174) V(n1175) V(n1176) V(n1177) V(n1178) V(n1179) V(n1) V(n1181) V(n1182) V(n1183) V(n1184) V(n1185) V(n1186) V(n1187) V(n1188) V(n1189) V(n1190) V(n1191) V(n1192) V(n1193) V(n1194) V(n1195) V(n1196) V(n1197) V(n1198) V(n1199) V(n1200) V(n1201) V(n1) V(n1203) V(n1204) V(n1205) V(n1206) V(n1207) V(n1208) V(n1209) V(n1210) V(n1211) V(n1212) V(n1213) V(n1214) V(n1215) V(n1216) V(n1217) V(n1218) V(n1219) V(n1220) V(n1221) V(n1222) V(n1223) V(n1224) V(n1225) V(n1226) V(n1227) V(n1228) V(n1229) V(n1230) V(n1231) V(n1232) V(n1233) V(n1234) V(n1235) V(n1236) V(n1237) V(n1238) V(n1239) V(n1240) V(n1241) V(n1242) V(n1243) V(n1244) V(n1245) V(n1246) V(n1247) V(n1248) V(n1249) V(n1250) V(n1251) V(n1252) V(n1253) V(n1254) V(n1255) V(n1256) V(n1257) V(n1258) V(n1259) V(n1260) V(n1261) V(n1262) V(n1263) V(n1264) V(n1265) V(n1266) V(n1267) V(n1268) V(n1269) V(n1270) V(n1271) V(n1) V(n1273) V(n1) V(n1275) V(n1276) V(n1277) V(n1278) V(n1279) V(n1280) V(n1281) V(n1282) V(n1283) V(n1284) V(n1285) V(n1286) V(n1287) V(n1288) V(n1289) V(n1290) V(n1291) V(n1292) V(n1293) V(n1294) V(n1295) V(n1296) V(n1297) V(n1298) V(n1299) V(n1300) V(n1301) V(n1302) V(n1303) V(n1304) V(n1305) V(n1306) V(n1307) V(n1308) V(n1309) V(n1310) V(n1311) V(n1312) V(n1313) V(n1314) V(n1315) V(n1316) V(n1317) V(n1318) V(n1319) V(n1320) V(n1321) V(n1322) V(n1) V(n1324) V(n1325) V(n1326) V(n1327) V(n1328) V(n1329) V(n1330) V(n1331) V(n1332) V(n1333) V(n1334) V(n1335) V(n1336) V(n1337) V(n1338) V(n1339) V(n1340) V(n1341) V(n1342) V(n1343) V(n1344) V(n1345) V(n1346) V(n1347) V(n1348) V(n1349) V(n1350) V(n1351) V(n1352) V(n1353) V(n1354) V(n1355) V(n1356) V(n1357) V(n1358) V(n1359) V(n1360) V(n1361) V(n1362) V(n1363) V(n1364) V(n1365) V(n1366) V(n1367) V(n1368) V(n1369) V(n1370) V(n1371) V(n1372) V(n1373) V(n1374) V(n1375) V(n1376) V(n1377) V(n1378) V(n1379) V(n1380) V(n1381) V(n1382) V(n1383) V(n1384) V(n1385) V(n1386) V(n1387) V(n1388) V(n1389) V(n1390) V(n1391) V(n1392) V(n1393) V(n1394) V(n1395) V(n1396) V(n1397) V(n1398) V(n1399) V(n1400) V(n1401) V(n1402) V(n1403) V(n1404) V(n1405) V(n1406) V(n1407) V(n1408) V(n1409) V(n1410) V(n1411) V(n1412) V(n1413) V(n1414) V(n1415) V(n1416) V(n1417) V(n1418) V(n1419) V(n1420) V(n1421) V(n1422) V(n1423) V(n1424) V(n1425) V(n1426) V(n1427) V(n1428) V(n1429) V(n1430) V(n1431) V(n1432) V(n1433) V(n1434) V(n1435) V(n1436) V(n1437) V(n1438) V(n1439) V(n1440) V(n1441) V(n1442) V(n1443) V(n1444) V(n1445) V(n1446) V(n1447) V(n1448) V(n1449) V(n1450) V(n1451) V(n1452) V(n1453) V(n1454) V(n1455) V(n1456) V(n1457) V(n1458) V(n1459) V(n1460) V(n1461) V(n1462) V(n1463) V(n1464) V(n1465) V(n1466) V(n1467) V(n1468) V(n1469) V(n1470) V(n1471) V(n1472) V(n1473) V(n1474) V(n1475) V(n1476) V(n1477) V(n1478) V(n1479) V(n1480) V(n1481) V(n1482) V(n1483) V(n1484) V(n1) V(n1486) V(n1487) V(n1488) V(n1489) V(n1490) V(n1491) V(n1492) V(n1493) V(n1494) V(n1495) V(n1496) V(n1497) V(n1498) V(n1499) V(n1500) V(n1501) V(n1502) V(n1503) V(n1504) V(n1505) V(n1506) V(n1507) V(n1508) V(n1509) V(n1510) V(n1511) V(n1512) V(n1513) V(n1514) V(n1515) V(n1516) V(n1517) V(n1518) V(n1519) V(n1520) V(n1521) V(n1522) V(n1523) V(n1524) V(n1525) V(n1526) V(n1527) V(n1528) V(n1529) V(n1530) V(n1531) V(n1532) V(n1533) V(n1534) V(n1535) V(n1536) V(n1537) V(n1538) V(n1539) V(n1540) V(n1541) V(n1542) V(n1543) V(n1544) V(n1545) V(n1546) V(n1547) V(n1548) V(n1549) V(n1550) V(n1551) V(n1552) V(n1553) V(n1554) V(n1555) V(n1556) V(n1557) V(n1558) V(n1559) V(n1560) V(n1561) V(n1562) V(n1563) V(n1564) V(n1565) V(n1566) V(n1567) V(n1568) V(n1569) V(n1570) V(n1571) V(n1572) V(n1573) V(n1574) V(n1575) V(n1576) V(n1577) V(n1578) V(n1579) V(n1580) V(n1581) V(n1582) V(n1583) V(n1584) V(n1585) V(n1586) V(n1587) V(n1588) V(n1589) V(n1590) V(n1591) V(n1592) V(n1593) V(n1594) V(n1595) V(n1596) V(n1597) V(n1598) V(n1599) V(n1600) V(n1601) V(n1602) V(n1603) V(n1604) V(n1605) V(n1606) V(n1607) V(n1608) V(n1609) V(n1610) V(n1611) V(n1612) V(n1613) V(n1614) V(n1615) V(n1616) V(n1617) V(n1618) V(n1619) V(n1620) V(n1621) V(n1622) V(n1623) V(n1624) V(n1625) V(n1626) V(n1627) V(n1628) V(n1629) V(n1630) V(n1631) V(n1632) V(n1633) V(n1634) V(n1635) V(n1636) V(n1637) V(n1638) V(n1639) V(n1640) V(n1641) V(n1642) V(n1643) V(n1644) V(n1645) V(n1646) V(n1647) V(n1648) V(n1649) V(n1650) V(n1651) V(n1652) V(n1653) V(n1654) V(n1655) V(n1656) V(n1657) V(n1658) V(n1659) V(n1660) V(n1661) V(n1662) V(n1663) V(n1664) V(n1665) V(n1666) V(n1667) V(n1668) V(n1669) V(n1670) V(n1671) V(n1672) V(n1673) V(n1674) V(n1675) V(n1676) V(n1677) V(n1678) V(n1679) V(n1680) V(n1681) V(n1682) V(n1683) V(n1684) V(n1685) V(n1686) V(n1687) V(n1688) V(n1689) V(n1690) V(n1691) V(n1692) V(n1693) V(n1694) V(n1695) V(n1696) V(n1697) V(n1698) V(n1699) V(n1700) V(n1701) V(n1702) V(n1703) V(n1704) V(n1705) V(n1706) V(n1707) V(n1708) V(n1) V(n1710) V(n1711) V(n1712) V(n1713) V(n1714) V(n1715) V(n1716) V(n1717) V(n1718) V(n1719) V(n1720) V(n1721) V(n1722) V(n1723) V(n1724) V(n1725) V(n1726) V(n1727) V(n1) V(n1729) V(n1730) V(n1731) V(n1732) V(n1733) V(n1734) V(n1735) V(n1736) V(n1737) V(n1738) V(n1739) V(n1740) V(n1741) V(n1742) V(n1743) V(n1744) V(n1745) V(n1746) V(n1747) V(n1748) V(n1749) V(n1750) V(n1751) V(n1752) V(n1753) V(n1754) V(n1755) V(n1756) V(n1757) V(n1758) V(n1759) V(n1760) V(n1761) V(n1762) V(n1763) V(n1764) V(n1765) V(n1766) V(n1767) V(n1768) V(n1769) V(n1770) V(n1771) V(n1772) V(n1773) V(n1774) V(n1775) V(n1776) V(n1777) V(n1778) V(n1779) V(n1) V(n1781) V(n1782) V(n1783) V(n1784) V(n1785) V(n1786) V(n1787) V(n1788) V(n1789) V(n1790) V(n1791) V(n1792) V(n1793) V(n1794) V(n1795) V(n1796) V(n1797) V(n1798) V(n1799) V(n1800) V(n1801) V(n1802) V(n1803) V(n1804) V(n1805) V(n1806) V(n1807) V(n1808) V(n1809) V(n1810) V(n1811) V(n1812) V(n1813) V(n1814) V(n1815) V(n1816) V(n1817) V(n1818) V(n1819) V(n1820) V(n1821) V(n1822) V(n1823) V(n1824) V(n1825) V(n1826) V(n1827) V(n1828) V(n1829) V(n1830) V(n1831) V(n1832) V(n1833) V(n1834) V(n1835) V(n1836) V(n1837) V(n1838) V(n1839) V(n1) V(n1841) V(n1842) V(n1843) V(n1844) V(n1845) V(n1846) V(n1847) V(n1848) V(n1849) V(n1850) V(n1851) V(n1852) V(n1853) V(n1854) V(n1855) V(n1856) V(n1857) V(n1858) V(n1859) V(n1860) V(n1861) V(n1862) V(n1863) V(n1864) V(n1865) V(n1866) V(n1867) V(n1868) V(n1869) V(n1870) V(n1871) V(n1872) V(n1873) V(n1874) V(n1875) V(n1876) V(n1877) V(n1878) V(n1879) V(n1880) V(n1881) V(n1882) V(n1883) V(n1884) V(n1885) V(n1886) V(n1887) V(n1888) V(n1889) V(n1) V(n1891) V(n1892) V(n1893) V(n1894) V(n1895) V(n1896) V(n1897) V(n1898) V(n1899) V(n1900) V(n1901) V(n1902) V(n1903) V(n1904) V(n1905) V(n1906) V(n1907) V(n1908) V(n1909) V(n1910) V(n1911) V(n1912) V(n1913) V(n1914) V(n1915) V(n1916) V(n1917) V(n1918) V(n1919) V(n1920) V(n1921) V(n1922) V(n1923) V(n1924) V(n1925) V(n1926) V(n1927) V(n1928) V(n1929) V(n1930) V(n1931) V(n1932) V(n1933) V(n1934) V(n1935) V(n1936) V(n1937) V(n1938) V(n1939) V(n1940) V(n1941) V(n1942) V(n1943) V(n1944) V(n1945) V(n1946) V(n1947) V(n1948) V(n1949) V(n1950) V(n1951) V(n1952) V(n1953) V(n1954) V(n1955) V(n1956) V(n1957) V(n1958) V(n1959) V(n1960) V(n1961) V(n1962) V(n1963) V(n1964) V(n1965) V(n1966) V(n1967) V(n1968) V(n1969) V(n1970) V(n1971) V(n1972) V(n1973) V(n1974) V(n1975) V(n1976) V(n1977) V(n1978) V(n1979) V(n1980) V(n1981) V(n1982) V(n1983) V(n1984) V(n1985) V(n1986) V(n1987) V(n1988) V(n1989) V(n1990) V(n1991) V(n1992) V(n1993) V(n1994) V(n1995) V(n1996) V(n1) V(n1998) V(n1999) V(n2000) V(n2001) V(n2002) V(n2003) V(n2004) V(n2005) V(n2006) V(n2007) V(n2008) V(n2009) V(n2010) V(n2011) V(n2012) V(n2013) V(n2014) V(n2015) V(n2016) V(n2017) V(n2018) V(n2019) V(n2020) V(n2021) V(n2022) V(n2023) V(n2024) V(n2025) V(n2026) V(n2027) V(n2028) V(n2029) V(n2030) V(n2031) V(n2032) V(n2033) V(n2034) V(n2035) V(n2036) V(n2037) V(n2038) V(n2039) V(n2040) V(n2041) V(n2042) V(n2043) V(n2044) V(n2045) V(n2046) V(n1) V(n2048) V(n2049) V(n2050) V(n2051) V(n2052) V(n2053) V(n2054) V(n2055) V(n2056) V(n2057) V(n2058) V(n2059) V(n2060) V(n2061) V(n2062) V(n2063) V(n1) V(n2065) V(n2066) V(n2067) V(n2068) V(n2069) V(n2070) V(n2071) V(n2072) V(n2073) V(n2074) V(n2075) V(n2076) V(n2077) V(n2078) V(n2079) V(n2080) V(n2081) V(n2082) V(n2083) V(n2084) V(n2085) V(n2086) V(n2087) V(n2088) V(n2089) V(n2090) V(n2091) V(n1) V(n2093) V(n2094) V(n2095) V(n2096) V(n2097) V(n2098) V(n2099) V(n2100) V(n2101) V(n2102) V(n2103) V(n2104) V(n2105) V(n2106) V(n2107) V(n2108) V(n2109) V(n2110) V(n2111) V(n2112) V(n2113) V(n2114) V(n2115) V(n2116) V(n2117) V(n2118) V(n2119) V(n2120) V(n2121) V(n2122) V(n2123) V(n2124) V(n2125) V(n2126) V(n2127) V(n2128) V(n2129) V(n2130) V(n2131) V(n2132) V(n2133) V(n2134) V(n2135) V(n2136) V(n2137) V(n2138) V(n2139) V(n2140) V(n2141) V(n2142) V(n2143) V(n2144) V(n2145) V(n2146) V(n2147) V(n2148) V(n2149) V(n2150) V(n2151) V(n2152) V(n2153) V(n2154) V(n2155) V(n2156) V(n2157) V(n2158) V(n2159) V(n2160) V(n2161) V(n2162) V(n2163) V(n2164) V(n2165) V(n2166) V(n2167) V(n2168) V(n2169) V(n2170) V(n2171) V(n2172) V(n2173) V(n2174) V(n2175) V(n2176) V(n2177) V(n2178) V(n2179) V(n2180) V(n2181) V(n2182) V(n2183) V(n2184) V(n2185) V(n2186) V(n2187) V(n2188) V(n2189) V(n2190) V(n2191) V(n2192) V(n2193) V(n2194) V(n2195) V(n2196) V(n2197) V(n2198) V(n1) V(n2200) V(n2201) V(n2202) V(n2203) V(n2204) V(n2205) V(n2206) V(n2207) V(n2208) V(n2209) V(n2210) V(n2211) V(n2212) V(n2213) V(n2214) V(n2215) V(n2216) V(n2217) V(n2218) V(n2219) V(n2220) V(n2221) V(n2222) V(n2223) V(n2224) V(n2225) V(n2226) V(n2227) V(n2228) V(n2229) V(n2230) V(n2231) V(n2232) V(n2233) V(n2234) V(n2235) V(n2236) V(n2237) V(n2238) V(n2239) V(n2240) V(n2241) V(n2242) V(n2243) V(n2244) V(n2245) V(n2246) V(n2247) V(n2248) V(n2249) V(n2250) V(n2251) V(n2252) V(n2253) V(n2254) V(n2255) V(n2256) V(n2257) V(n2258) V(n2259) V(n2260) V(n2261) V(n2262) V(n2263) V(n2264) V(n2265) V(n2266) V(n2267) V(n2268) V(n2269) V(n2270) V(n2271) V(n2272) V(n2273) V(n2274) V(n2275) V(n2276) V(n2277) V(n2278) V(n2279) V(n2280) V(n2281) V(n2282) V(n2283) V(n2284) V(n2285) V(n2286) V(n2287) V(n2288) V(n2289) V(n2290) V(n2291) V(n2292) V(n2293) V(n2294) V(n2295) V(n2296) V(n2297) V(n2298) V(n2299) V(n2300) V(n2301) V(n2302) V(n2303) V(n2304) V(n2305) V(n2306) V(n2307) V(n2308) V(n2309) V(n2310) V(n2311) V(n2312) V(n2313) V(n2314) V(n2315) V(n2316) V(n2317) V(n2318) V(n2319) V(n2320) V(n2321) V(n2322) V(n2323) V(n2324) V(n2325) V(n2326) V(n2327) V(n2328) V(n2329) V(n2330) V(n2331) V(n2332) V(n2333) V(n2334) V(n2335) V(n2336) V(n2337) V(n2338) V(n2339) V(n2340) V(n2341) V(n2342) V(n2343) V(n2344) V(n2345) V(n2346) V(n2347) V(n2348) V(n2349) V(n2350) V(n2351) V(n2352) V(n2353) V(n2354) V(n2355) V(n2356) V(n2357) V(n2358) V(n2359) V(n2360) V(n2361) V(n2362) V(n2363) V(n2364) V(n2365) V(n2366) V(n2367) V(n2368) V(n2369) V(n2370) V(n2371) V(n2372) V(n2373) V(n2374) V(n2375) V(n2376) V(n2377) V(n2378) V(n2379) V(n2380) V(n2381) V(n2382) V(n2383) V(n2384) V(n2385) V(n2386) V(n2387) V(n2388) V(n2389) V(n2390) V(n2391) V(n2392) V(n2393) V(n2394) V(n2395) V(n1) V(n2397) V(n2398) V(n2399) V(n2400) V(n2401) V(n2402) V(n2403) V(n2404) V(n2405) V(n2406) V(n2407) V(n2408) V(n2409) V(n2410) V(n2411) V(n2412) V(n2413) V(n2414) V(n2415) V(n2416) V(n2417) V(n2418) V(n2419) V(n2420) V(n2421) V(n2422) V(n2423) V(n2424) V(n2425) V(n2426) V(n2427) V(n2428) V(n2429) V(n2430) V(n2431) V(n2432) V(n2433) V(n2434) V(n2435) V(n2436) V(n2437) V(n2438) V(n2439) V(n1) V(n2441) V(n2442) V(n2443) V(n2444) V(n2445) V(n2446) V(n1) V(n2448) V(n2449) V(n2450) V(n2451) V(n2452) V(n2453) V(n2454) V(n2455) V(n2456) V(n2457) V(n2458) V(n2459) V(n2460) V(n2461) V(n2462) V(n2463) V(n2464) V(n2465) V(n2466) V(n2467) V(n2468) V(n2469) V(n2470) V(n2471) V(n2472) V(n2473) V(n2474) V(n2475) V(n2476) V(n2477) V(n2478) V(n2479) V(n2480) V(n2481) V(n2482) V(n2483) V(n2484) V(n2485) V(n2486) V(n2487) V(n2488) V(n2489) V(n2490) V(n2491) V(n2492) V(n2493) V(n2494) V(n2495) V(n2496) V(n2497) V(n2498) V(n2499) V(n2500) V(n2501) V(n2502) V(n2503) V(n2504) V(n2505) V(n2506) V(n2507) V(n2508) V(n2509) V(n2510) V(n2511) V(n2512) V(n2513) V(n2514) V(n2515) V(n2516) V(n2517) V(n2518) V(n2519) V(n2520) V(n2521) V(n2522) V(n2523) V(n2524) V(n2525) V(n2526) V(n2527) V(n2528) V(n2529) V(n2530) V(n2531) V(n2532) V(n2533) V(n2534) V(n2535) V(n2536) V(n2537) V(n2538) V(n2539) V(n2540) V(n2541) V(n2542) V(n2543) V(n2544) V(n2545) V(n2546) V(n2547) V(n2548) V(n2549) V(n2550) V(n2551) V(n2552) V(n2553) V(n2554) V(n2555) V(n2556) V(n2557) V(n2558) V(n2559) V(n2560) V(n2561) V(n2562) V(n2563) V(n2564) V(n2565) V(n2566) V(n2567) V(n2568) V(n2569) V(n2570) V(n2571) V(n1) V(n2573) V(n2574) V(n2575) V(n2576) V(n2577) V(n2578) V(n2579) V(n2580) V(n2581) V(n2582) V(n2583) V(n2584) V(n2585) V(n2586) V(n2587) V(n2588) V(n2589) V(n2590) V(n2591) V(n2592) V(n2593) V(n2594) V(n2595) V(n2596) V(n2597) V(n2598) V(n2599) V(n2600) V(n2601) V(n2602) V(n2603) V(n2604) V(n2605) V(n2606) V(n2607) V(n2608) V(n2609) V(n2610) V(n1) V(n2612) V(n2613) V(n2614) V(n2615) V(n2616) V(n2617) V(n2618) V(n2619) V(n2620) V(n2621) V(n2622) V(n2623) V(n2624) V(n2625) V(n2626) V(n2627) V(n2628) V(n2629) V(n2630) V(n2631) V(n2632) V(n2633) V(n2634) V(n2635) V(n2636) V(n2637) V(n2638) V(n2639) V(n2640) V(n2641) V(n2642) V(n2643) V(n2644) V(n2645) V(n2646) V(n2647) V(n2648) V(n2649) V(n2650) V(n2651) V(n2652) V(n2653) V(n2654) V(n2655) V(n2656) V(n2657) V(n2658) V(n2659) V(n2660) V(n2661) V(n2662) V(n2663) V(n2664) V(n2665) V(n2666) V(n2667) V(n2668) V(n2669) V(n2670) V(n2671) V(n2672) V(n2673) V(n2674) V(n2675) V(n2676) V(n2677) V(n2678) V(n2679) V(n2680) V(n2681) V(n2682) V(n2683) V(n2684) V(n2685) V(n2686) V(n2687) V(n2688) V(n2689) V(n2690) V(n2691) V(n2692) V(n2693) V(n2694) V(n2695) V(n2696) V(n2697) V(n2698) V(n2699) V(n2700) V(n2701) V(n2702) V(n2703) V(n2704) V(n2705) V(n2706) V(n2707) V(n2708) V(n2709) V(n2710) V(n2711) V(n2712) V(n2713) V(n2714) V(n2715) V(n2716) V(n2717) V(n2718) V(n2719) V(n2720) V(n2721) V(n2722) V(n2723) V(n2724) V(n2725) V(n2726) V(n2727) V(n2728) V(n2729) V(n2730) V(n2731) V(n2732) V(n2733) V(n2734) V(n2735) V(n2736) V(n2737) V(n2738) V(n2739) V(n2740) V(n2741) V(n2742) V(n2743) V(n2744) V(n2745) V(n2746) V(n2747) V(n1) V(n2749) V(n2750) V(n2751) V(n2752) V(n2753) V(n2754) V(n2755) V(n2756) V(n2757) V(n2758) V(n2759) V(n2760) V(n2761) V(n2762) V(n2763) V(n2764) V(n2765) V(n2766) V(n2767) V(n2768) V(n2769) V(n2770) V(n2771) V(n2772) V(n2773) V(n2774) V(n2775) V(n2776) V(n2777) V(n2778) V(n2779) V(n2780) V(n2781) V(n2782) V(n2783) V(n2784) V(n2785) V(n2786) V(n2787) V(n2788) V(n2789) V(n2790) V(n2791) V(n2792) V(n2793) V(n2794) V(n2795) V(n2796) V(n2797) V(n2798) V(n2799) V(n2800) V(n2801) V(n2802) V(n2803) V(n2804) V(n2805) V(n2806) V(n2807) V(n2808) V(n2809) V(n2810) V(n2811) V(n2812) V(n2813) V(n2814) V(n2815) V(n2816) V(n2817) V(n2818) V(n2819) V(n2820) V(n2821) V(n2822) V(n2823) V(n2824) V(n2825) V(n2826) V(n2827) V(n2828) V(n2829) V(n2830) V(n2831) V(n2832) V(n2833) V(n2834) V(n2835) V(n2836) V(n2837) V(n2838) V(n2839) V(n2840) V(n2841) V(n2842) V(n2843) V(n2844) V(n2845) V(n2846) V(n2847) V(n2848) V(n2849) V(n2850) V(n1) V(n2852) V(n2853) V(n2854) V(n2855) V(n2856) V(n2857) V(n2858) V(n2859) V(n2860) V(n2861) V(n2862) V(n2863) V(n2864) V(n2865) V(n2866) V(n2867) V(n2868) V(n2869) V(n1) V(n2871) V(n2872) V(n2873) V(n2874) V(n2875) V(n2876) V(n2877) V(n2878) V(n2879) V(n2880) V(n2881) V(n2882) V(n2883) V(n2884) V(n2885) V(n2886) V(n2887) V(n2888) V(n2889) V(n2890) V(n2891) V(n2892) V(n2893) V(n2894) V(n2895) V(n2896) V(n2897) V(n2898) V(n2899) V(n2900) V(n1) V(n2902) V(n2903) V(n2904) V(n2905) V(n2906) V(n2907) V(n2908) V(n2909) V(n2910) V(n2911) V(n2912) V(n2913) V(n2914) V(n2915) V(n2916) V(n2917) V(n2918) V(n2919) V(n2920) V(n2921) V(n2922) V(n2923) V(n2924) V(n2925) V(n2926) V(n2927) V(n2928) V(n2929) V(n2930) V(n2931) V(n2932) V(n2933) V(n2934) V(n2935) V(n2936) V(n2937) V(n2938) V(n2939) V(n2940) V(n2941) V(n2942) V(n2943) V(n1) V(n2945) V(n2946) V(n2947) V(n2948) V(n2949) V(n2950) V(n2951) V(n2952) V(n2953) V(n2954) V(n2955) V(n2956) V(n2957) V(n2958) V(n2959) V(n2960) V(n2961) V(n2962) V(n2963) V(n2964) V(n2965) V(n2966) V(n2967) V(n2968) V(n2969) V(n2970) V(n2971) V(n2972) V(n2973) V(n2974) V(n2975) V(n2976) V(n2977) V(n2978) V(n2979) V(n2980) V(n2981) V(n2982) V(n2983) V(n2984) V(n2985) V(n2986) V(n2987) V(n2988) V(n2989) V(n2990) V(n2991) V(n2992) V(n2993) V(n2994) V(n2995) V(n2996) V(n2997) V(n2998) V(n2999) V(n3000) V(n3001) V(n3002) V(n3003) V(n3004) V(n3005) V(n3006) V(n3007) V(n3008) V(n3009) V(n3010) V(n3011) V(n3012) V(n3013) V(n3014) V(n3015) V(n3016) V(n3017) V(n3018) V(n3019) V(n3020) V(n3021) V(n3022) V(n3023) V(n3024) V(n3025) V(n3026) V(n3027) V(n3028) V(n3029) V(n3030) V(n3031) V(n3032) V(n3033) V(n3034) V(n3035) V(n3036) V(n3037) V(n3038) V(n3039) V(n1) V(n3041) V(n3042) V(n3043) V(n3044) V(n3045) V(n3046) V(n3047) V(n3048) V(n3049) V(n3050) V(n3051) V(n3052) V(n3053) V(n3054) V(n3055) V(n3056) V(n3057) V(n3058) V(n3059) V(n3060) V(n3061) V(n3062) V(n3063) V(n3064) V(n3065) V(n3066) V(n3067) V(n3068) V(n3069) V(n3070) V(n3071) V(n3072) V(n3073) V(n3074) V(n3075) V(n3076) V(n3077) V(n3078) V(n3079) V(n3080) V(n3081) V(n3082) V(n3083) V(n3084) V(n3085) V(n3086) V(n3087) V(n3088) V(n3089) V(n3090) V(n3091) V(n3092) V(n3093) V(n3094) V(n3095) V(n3096) V(n3097) V(n1) V(n3099) V(n3100) V(n3101) V(n3102) V(n3103) V(n3104) V(n3105) V(n3106) V(n3107) V(n3108) V(n3109) V(n3110) V(n3111) V(n1) V(n3113) V(n3114) V(n3115) V(n3116) V(n3117) V(n3118) V(n3119) V(n3120) V(n3121) V(n3122) V(n3123) V(n3124) V(n3125) V(n3126) V(n3127) V(n3128) V(n3129) V(n3130) V(n3131) V(n3132) V(n3133) V(n3134) V(n3135) V(n3136) V(n3137) V(n3138) V(n3139) V(n3140) V(n3141) V(n3142) V(n3143) V(n3144) V(n3145) V(n3146) V(n3147) V(n3148) V(n3149) V(n3150) V(n3151) V(n3152) V(n3153) V(n3154) V(n3155) V(n3156) V(n3157) V(n3158) V(n3159) V(n3160) V(n3161) V(n3162) V(n3163) V(n3164) V(n3165) V(n3166) V(n3167) V(n3168) V(n1) V(n3170) V(n3171) V(n3172) V(n3173) V(n3174) V(n3175) V(n3176) V(n3177) V(n3178) V(n3179) V(n3180) V(n3181) V(n3182) V(n3183) V(n3184) V(n3185) V(n3186) V(n3187) V(n3188) V(n3189) V(n3190) V(n3191) V(n3192) V(n3193) V(n3194) V(n3195) V(n3196) V(n3197) V(n3198) V(n3199) V(n3200) V(n3201) V(n3202) V(n3203) V(n3204) V(n3205) V(n3206) V(n3207) V(n3208) V(n3209) V(n3210) V(n3211) V(n3212) V(n3213) V(n3214) V(n3215) V(n3216) V(n3217) V(n3218) V(n3219) V(n3220) V(n3221) V(n3222) V(n3223) V(n1) V(n3225) V(n3226) V(n3227) V(n3228) V(n3229) V(n3230) V(n3231) V(n3232) V(n3233) V(n3234) V(n3235) V(n3236) V(n3237) V(n3238) V(n3239) V(n3240) V(n3241) V(n3242) V(n3243) V(n3244) V(n3245) V(n3246) V(n3247) V(n3248) V(n3249) V(n3250) V(n3251) V(n3252) V(n3253) V(n3254) V(n3255) V(n3256) V(n3257) V(n3258) V(n3259) V(n3260) V(n3261) V(n3262) V(n3263) V(n3264) V(n3265) V(n3266) V(n3267) V(n3268) V(n3269) V(n3270) V(n3271) V(n3272) V(n3273) V(n3274) V(n3275) V(n3276) V(n3277) V(n3278) V(n3279) V(n3280) V(n3281) V(n3282) V(n3283) V(n3284) V(n3285) V(n3286) V(n3287) V(n3288) V(n3289) V(n3290) V(n3291) V(n3292) V(n3293) V(n3294) V(n3295) V(n3296) V(n3297) V(n3298) V(n3299) V(n3300) V(n3301) V(n3302) V(n3303) V(n3304) V(n3305) V(n3306) V(n3307) V(n3308) V(n1) V(n3310) V(n3311) V(n3312) V(n3313) V(n3314) V(n3315) V(n3316) V(n3317) V(n3318) V(n3319) V(n3320) V(n3321) V(n3322) V(n3323) V(n3324) V(n3325) V(n3326) V(n3327) V(n3328) V(n3329) V(n3330) V(n3331) V(n3332) V(n3333) V(n3334) V(n3335) V(n3336) V(n3337) V(n3338) V(n3339) V(n3340) V(n3341) V(n3342) V(n3343) V(n3344) V(n3345) V(n3346) V(n3347) V(n3348) V(n3349) V(n3350) V(n3351) V(n3352) V(n3353) V(n3354) V(n3355) V(n3356) V(n3357) V(n3358) V(n3359) V(n3360) V(n3361) V(n3362) V(n3363) V(n3364) V(n3365) V(n3366) V(n3367) V(n3368) V(n3369) V(n3370) V(n3371) V(n3372) V(n3373) V(n3374) V(n3375) V(n3376) V(n3377) V(n3378) V(n3379) V(n3380) V(n3381) V(n3382) V(n3383) V(n3384) V(n3385) V(n3386) V(n3387) V(n3388) V(n3389) V(n1) V(n3391) V(n3392) V(n3393) V(n3394) V(n3395) V(n3396) V(n3397) V(n3398) V(n3399) V(n3400) V(n3401) V(n3402) V(n3403) V(n3404) V(n3405) V(n3406) V(n3407) V(n3408) V(n3409) V(n3410) V(n3411) V(n3412) V(n3413) V(n3414) V(n3415) V(n3416) V(n3417) V(n3418) V(n3419) V(n3420) V(n3421) V(n3422) V(n3423) V(n3424) V(n3425) V(n3426) V(n3427) V(n3428) V(n3429) V(n3430) V(n3431) V(n3432) V(n3433) V(n3434) V(n3435) V(n3436) V(n3437) V(n3438) V(n3439) V(n3440) V(n3441) V(n3442) V(n3443) V(n3444) V(n3445) V(n3446) V(n3447) V(n3448) V(n3449) V(n3450) V(n3451) V(n3452) V(n3453) V(n3454) V(n3455) V(n3456) V(n3457) V(n3458) V(n3459) V(n3460) V(n3461) V(n3462) V(n3463) V(n3464) V(n3465) V(n3466) V(n3467) V(n3468) V(n3469) V(n3470) V(n3471) V(n3472) V(n3473) V(n3474) V(n3475) V(n3476) V(n3477) V(n3478) V(n3479) V(n3480) V(n3481) V(n3482) V(n3483) V(n3484) V(n3485) V(n3486) V(n3487) V(n3488) V(n3489) V(n3490) V(n3491) V(n3492) V(n1) V(n3494) V(n3495) V(n3496) V(n3497) V(n3498) V(n3499) V(n3500) V(n3501) V(n3502) V(n3503) V(n3504) V(n3505) V(n3506) V(n3507) V(n3508) V(n3509) V(n3510) V(n3511) V(n3512) V(n3513) V(n3514) V(n3515) V(n3516) V(n3517) V(n3518) V(n3519) V(n3520) V(n3521) V(n3522) V(n3523) V(n3524) V(n3525) V(n3526) V(n3527) V(n3528) V(n3529) V(n3530) V(n3531) V(n3532) V(n3533) V(n3534) V(n3535) V(n3536) V(n3537) V(n3538) V(n3539) V(n3540) V(n3541) V(n3542) V(n3543) V(n3544) V(n3545) V(n3546) V(n3547) V(n3548) V(n3549) V(n3550) V(n3551) V(n3552) V(n3553) V(n3554) V(n3555) V(n3556) V(n3557) V(n3558) V(n3559) V(n3560) V(n3561) V(n3562) V(n3563) V(n3564) V(n3565) V(n3566) V(n3567) V(n3568) V(n3569) V(n3570) V(n3571) V(n3572) V(n3573) V(n3574) V(n3575) V(n3576) V(n3577) V(n3578) V(n3579) V(n3580) V(n3581) V(n3582) V(n3583) V(n3584) V(n3585) V(n3586) V(n3587) V(n3588) V(n3589) V(n3590) V(n3591) V(n3592) V(n3593) V(n3594) V(n3595) V(n3596) V(n3597) V(n3598) V(n3599) V(n3600) V(n3601) V(n3602) V(n3603) V(n3604) V(n3605) V(n3606) V(n3607) V(n3608) V(n3609) V(n3610) V(n3611) V(n3612) V(n3613) V(n3614) V(n3615) V(n3616) V(n3617) V(n3618) V(n3619) V(n3620) V(n3621) V(n3622) V(n3623) V(n3624) V(n3625) V(n3626) V(n3627) V(n3628) V(n3629) V(n3630) V(n3631) V(n3632) V(n3633) V(n3634) V(n3635) V(n3636) V(n3637) V(n3638) V(n3639) V(n3640) V(n3641) V(n3642) V(n3643) V(n3644) V(n3645) V(n3646) V(n3647) V(n3648) V(n3649) V(n3650) V(n3651) V(n3652) V(n3653) V(n3654) V(n3655) V(n3656) V(n3657) V(n3658) V(n3659) V(n3660) V(n3661) V(n3662) V(n3663) V(n3664) V(n3665) V(n3666) V(n3667) V(n3668) V(n3669) V(n3670) V(n3671) V(n3672) V(n3673) V(n3674) V(n3675) V(n3676) V(n3677) V(n3678) V(n3679) V(n3680) V(n3681) V(n3682) V(n3683) V(n3684) V(n3685) V(n3686) V(n3687) V(n3688) V(n3689) V(n3690) V(n3691) V(n3692) V(n3693) V(n3694) V(n3695) V(n3696) V(n3697) V(n3698) V(n3699) V(n3700) V(n3701) V(n3702) V(n3703) V(n3704) V(n3705) V(n3706) V(n3707) V(n3708) V(n3709) V(n3710) V(n3711) V(n3712) V(n3713) V(n3714) V(n3715) V(n3716) V(n3717) V(n3718) V(n3719) V(n3720) V(n3721) V(n3722) V(n3723) V(n3724) V(n3725) V(n3726) V(n3727) V(n3728) V(n3729) V(n3730) V(n3731) V(n3732) V(n3733) V(n3734) V(n3735) V(n3736) V(n3737) V(n3738) V(n3739) V(n3740) V(n3741) V(n3742) V(n3743) V(n3744) V(n3745) V(n3746) V(n3747) V(n3748) V(n3749) V(n3750) V(n3751) V(n3752) V(n3753) V(n3754) V(n3755) V(n3756) V(n3757) V(n3758) V(n3759) V(n3760) V(n3761) V(n3762) V(n3763) V(n3764) V(n3765) V(n3766) V(n3767) V(n3768) V(n3769) V(n3770) V(n3771) V(n3772) V(n3773) V(n3774) V(n3775) V(n3776) V(n3777) V(n3778) V(n3779) V(n3780) V(n3781) V(n3782) V(n3783) V(n3784) V(n3785) V(n3786) V(n3787) V(n3788) V(n3789) V(n3790) V(n3791) V(n3792) V(n3793) V(n3794) V(n3795) V(n3796) V(n3797) V(n3798) V(n3799) V(n3800) V(n3801) V(n3802) V(n3803) V(n3804) V(n3805) V(n3806) V(n3807) V(n3808) V(n3809) V(n3810) V(n3811) V(n3812) V(n3813) V(n3814) V(n3815) V(n3816) V(n3817) V(n3818) V(n3819) V(n3820) V(n3821) V(n3822) V(n3823) V(n3824) V(n3825) V(n3826) V(n3827) V(n3828) V(n3829) V(n3830) V(n3831) V(n3832) V(n3833) V(n3834) V(n3835) V(n3836) V(n3837) V(n3838) V(n3839) V(n3840) V(n3841) V(n3842) V(n3843) V(n3844) V(n3845) V(n3846) V(n3847) V(n3848) V(n3849) V(n3850) V(n3851) V(n3852) V(n3853) V(n3854) V(n3855) V(n3856) V(n3857) V(n3858) V(n3859) V(n3860) V(n3861) V(n3862) V(n3863) V(n3864) V(n3865) V(n3866) V(n3867) V(n3868) V(n3869) V(n3870) V(n3871) V(n3872) V(n3873) V(n3874) V(n3875) V(n3876) V(n3877) V(n3878) V(n3879) V(n3880) V(n3881) V(n3882) V(n3883) V(n3884) V(n3885) V(n3886) V(n3887) V(n3888) V(n3889) V(n3890) V(n3891) V(n3892) V(n3893) V(n3894) V(n3895) V(n3896) V(n3897) V(n3898) V(n3899) V(n3900) V(n3901) V(n3902) V(n3903) V(n3904) V(n3905) V(n3906) V(n3907) V(n3908) V(n3909) V(n3910) V(n3911) V(n3912) V(n3913) V(n3914) V(n3915) V(n3916) V(n3917) V(n3918) V(n3919) V(n3920) V(n3921) V(n3922) V(n3923) V(n3924) V(n3925) V(n3926) V(n3927) V(n3928) V(n3929) V(n3930) V(n3931) V(n3932) V(n3933) V(n3934) V(n3935) V(n3936) V(n3937) V(n3938) V(n3939) V(n3940) V(n3941) V(n3942) V(n3943) V(n3944) V(n3945) V(n3946) V(n3947) V(n3948) V(n3949) V(n3950) V(n3951) V(n1) V(n3953) V(n3954) V(n3955) V(n3956) V(n3957) V(n3958) V(n3959) V(n3960) V(n3961) V(n3962) V(n3963) V(n3964) V(n3965) V(n3966) V(n3967) V(n3968) V(n3969) V(n3970) V(n3971) V(n3972) V(n3973) V(n3974) V(n3975) V(n3976) V(n3977) V(n3978) V(n3979) V(n3980) V(n3981) V(n3982) V(n3983) V(n3984) V(n3985) V(n3986) V(n3987) V(n3988) V(n3989) V(n3990) V(n3991) V(n3992) V(n3993) V(n3994) V(n3995) V(n3996) V(n3997) V(n3998) V(n3999) V(n4000) V(n4001) V(n4002) V(n4003) V(n4004) V(n4005) V(n4006) V(n4007) V(n4008) V(n4009) V(n4010) V(n4011) V(n4012) V(n4013) V(n4014) V(n4015) V(n4016) V(n4017) V(n4018) V(n4019) V(n4020) V(n4021) V(n4022) V(n4023) V(n4024) V(n4025) V(n4026) V(n4027) V(n4028) V(n4029) V(n4030) V(n4031) V(n4032) V(n4033) V(n4034) V(n4035) V(n4036) V(n4037) V(n4038) V(n4039) V(n4040) V(n4041) V(n4042) V(n4043) V(n4044) V(n4045) V(n4046) V(n4047) V(n4048) V(n4049) V(n4050) V(n4051) V(n4052) V(n4053) V(n4054) V(n4055) V(n4056) V(n4057) V(n4058) V(n4059) V(n4060) V(n4061) V(n4062) V(n4063) V(n4064) V(n4065) V(n4066) V(n4067) V(n4068) V(n4069) V(n4070) V(n4071) V(n4072) V(n4073) V(n4074) V(n4075) V(n4076) V(n4077) V(n4078) V(n4079) V(n4080) V(n4081) V(n4082) V(n4083) V(n4084) V(n4085) V(n4086) V(n4087) V(n4088) V(n4089) V(n4090) V(n4091) V(n4092) V(n4093) V(n4094) V(n4095) V(n4096) V(n4097) V(n4098) V(n4099) V(n4100) V(n4101) V(n4102) V(n4103) V(n4104) V(n4105) V(n4106) V(n4107) V(n4108) V(n4109) V(n4110) V(n4111) V(n4112) V(n4113) V(n4114) V(n4115) V(n4116) V(n4117) V(n4118) V(n4119) V(n4120) V(n4121) V(n4122) V(n4123) V(n4124) V(n4125) V(n4126) V(n4127) V(n4128) V(n4129) V(n4130) V(n4131) V(n4132) V(n4133) V(n4134) V(n4135) V(n4136) V(n4137) V(n4138) V(n4139) V(n4140) V(n4141) V(n4142) V(n4143) V(n4144) V(n4145) V(n4146) V(n4147) V(n4148) V(n4149) V(n4150) V(n4151) V(n4152) V(n4153) V(n4154) V(n4155) V(n4156) V(n4157) V(n4158) V(n4159) V(n4160) V(n4161) V(n4162) V(n4163) V(n4164) V(n4165) V(n4166) V(n4167) V(n4168) V(n4169) V(n4170) V(n4171) V(n4172) V(n4173) V(n4174) V(n4175) V(n4176) V(n4177) V(n4178) V(n4179) V(n4180) V(n4181) V(n4182) V(n4183) V(n4184) V(n4185) V(n4186) V(n4187) V(n4188) V(n4189) V(n1) V(n4191) V(n4192) V(n4193) V(n4194) V(n4195) V(n4196) V(n4197) V(n4198) V(n4199) V(n4200) V(n4201) V(n4202) V(n4203) V(n4204) V(n4205) V(n4206) V(n4207) V(n4208) V(n4209) V(n4210) V(n4211) V(n4212) V(n4213) V(n4214) V(n4215) V(n4216) V(n4217) V(n4218) V(n4219) V(n4220) V(n4221) V(n4222) V(n4223) V(n4224) V(n4225) V(n4226) V(n4227) V(n4228) V(n4229) V(n4230) V(n4231) V(n4232) V(n4233) V(n4234) V(n4235) V(n4236) V(n4237) V(n4238) V(n4239) V(n4240) V(n4241) V(n4242) V(n4243) V(n4244) V(n4245) V(n4246) V(n4247) V(n4248) V(n4249) V(n4250) V(n4251) V(n4252) V(n4253) V(n4254) V(n4255) V(n4256) V(n4257) V(n4258) V(n4259) V(n4260) V(n4261) V(n4262) V(n4263) V(n4264) V(n4265) V(n4266) V(n4267) V(n4268) V(n4269) V(n4270) V(n4271) V(n4272) V(n4273) V(n4274) V(n4275) V(n4276) V(n4277) V(n4278) V(n4279) V(n4280) V(n4281) V(n4282) V(n4283) V(n4284) V(n4285) V(n4286) V(n4287) V(n4288) V(n4289) V(n4290) V(n4291) V(n4292) V(n4293) V(n4294) V(n4295) V(n4296) V(n4297) V(n4298) V(n4299) V(n4300) V(n4301) V(n4302) V(n4303) V(n4304) V(n4305) V(n4306) V(n4307) V(n4308) V(n4309) V(n4310) V(n4311) V(n4312) V(n4313) V(n4314) V(n4315) V(n4316) V(n4317) V(n4318) V(n4319) V(n4320) V(n4321) V(n4322) V(n4323) V(n4324) V(n4325) V(n4326) V(n4327) V(n4328) V(n4329) V(n4330) V(n1) V(n1) V(n4333) V(n4334) V(n4335) V(n4336) V(n4337) V(n4338) V(n1) V(n4340) V(n4341) V(n4342) V(n4343) V(n4344) V(n4345) V(n4346) V(n4347) V(n4348) V(n4349) V(n4350) V(n4351) V(n4352) V(n4353) V(n4354) V(n4355) V(n4356) V(n4357) V(n4358) V(n4359) V(n4360) V(n4361) V(n4362) V(n4363) V(n4364) V(n4365) V(n4366) V(n4367) V(n4368) V(n4369) V(n4370) V(n4371) V(n4372) V(n4373) V(n4374) V(n4375) V(n4376) V(n4377) V(n4378) V(n4379) V(n4380) V(n4381) V(n4382) V(n4383) V(n4384) V(n4385) V(n1) V(n4387) V(n4388) V(n4389) V(n4390) V(n4391) V(n4392) V(n4393) V(n4394) V(n4395) V(n4396) V(n4397) V(n4398) V(n4399) V(n4400) V(n4401) V(n4402) V(n4403) V(n4404) V(n4405) V(n4406) V(n4407) V(n4408) V(n4409) V(n4410) V(n4411) V(n4412) V(n4413) V(n4414) V(n4415) V(n4416) V(n4417) V(n4418) V(n4419) V(n4420) V(n4421) V(n4422) V(n4423) V(n4424) V(n4425) V(n4426) V(n4427) V(n4428) V(n4429) V(n4430) V(n4431) V(n4432) V(n4433) V(n4434) V(n4435) V(n4436) V(n4437) V(n4438) V(n4439) V(n4440) V(n4441) V(n4442) V(n4443) V(n4444) V(n4445) V(n4446) V(n4447) V(n4448) V(n4449) V(n4450) V(n4451) V(n4452) V(n4453) V(n4454) V(n4455) V(n4456) V(n4457) V(n4458) V(n4459) V(n4460) V(n4461) V(n4462) V(n4463) V(n4464) V(n4465) V(n4466) V(n4467) V(n4468) V(n4469) V(n4470) V(n4471) V(n4472) V(n4473) V(n4474) V(n4475) V(n4476) V(n4477) V(n4478) V(n4479) V(n4480) V(n4481) V(n4482) V(n4483) V(n4484) V(n4485) V(n4486) V(n4487) V(n4488) V(n4489) V(n4490) V(n4491) V(n4492) V(n4493) V(n4494) V(n4495) V(n4496) V(n4497) V(n4498) V(n4499) V(n4500) V(n4501) V(n4502) V(n4503) V(n4504) V(n4505) V(n4506) V(n4507) V(n4508) V(n4509) V(n4510) V(n4511) V(n4512) V(n4513) V(n4514) V(n4515) V(n4516) V(n4517) V(n4518) V(n4519) V(n4520) V(n4521) V(n4522) V(n4523) V(n4524) V(n4525) V(n4526) V(n4527) V(n4528) V(n4529) V(n4530) V(n1) V(n4532) V(n4533) V(n4534) V(n4535) V(n4536) V(n4537) V(n4538) V(n4539) V(n4540) V(n4541) V(n4542) V(n4543) V(n4544) V(n4545) V(n4546) V(n4547) V(n4548) V(n4549) V(n4550) V(n4551) V(n4552) V(n4553) V(n4554) V(n4555) V(n4556) V(n4557) V(n4558) V(n4559) V(n4560) V(n4561) V(n4562) V(n4563) V(n4564) V(n4565) V(n4566) V(n4567) V(n4568) V(n4569) V(n4570) V(n4571) V(n4572) V(n4573) V(n4574) V(n4575) V(n4576) V(n4577) V(n4578) V(n4579) V(n4580) V(n4581) V(n4582) V(n4583) V(n4584) V(n4585) V(n4586) V(n4587) V(n4588) V(n4589) V(n4590) V(n4591) V(n4592) V(n4593) V(n4594) V(n4595) V(n4596) V(n4597) V(n4598) V(n4599) V(n4600) V(n4601) V(n4602) V(n4603) V(n4604) V(n4605) V(n4606) V(n4607) V(n4608) V(n4609) V(n1) V(n4611) V(n4612) V(n4613) V(n4614) V(n4615) V(n4616) V(n4617) V(n4618) V(n4619) V(n4620) V(n4621) V(n4622) V(n4623) V(n4624) V(n4625) V(n4626) V(n4627) V(n4628) V(n4629) V(n4630) V(n4631) V(n4632) V(n4633) V(n4634) V(n4635) V(n4636) V(n4637) V(n4638) V(n4639) V(n4640) V(n4641) V(n4642) V(n4643) V(n4644) V(n4645) V(n4646) V(n4647) V(n4648) V(n4649) V(n4650) V(n4651) V(n4652) V(n4653) V(n4654) V(n4655) V(n4656) V(n4657) V(n4658) V(n4659) V(n4660) V(n4661) V(n4662) V(n4663) V(n4664) V(n4665) V(n4666) V(n1) V(n4668) V(n4669) V(n4670) V(n4671) V(n4672) V(n4673) V(n4674) V(n4675) V(n4676) V(n4677) V(n4678) V(n4679) V(n4680) V(n4681) V(n4682) V(n4683) V(n4684) V(n4685) V(n4686) V(n4687) V(n4688) V(n4689) V(n4690) V(n4691) V(n4692) V(n4693) V(n4694) V(n4695) V(n4696) V(n4697) V(n4698) V(n4699) V(n4700) V(n4701) V(n4702) V(n4703) V(n4704) V(n4705) V(n4706) V(n4707) V(n4708) V(n4709) V(n4710) V(n4711) V(n4712) V(n4713) V(n4714) V(n4715) V(n4716) V(n4717) V(n4718) V(n4719) V(n4720) V(n4721) V(n4722) V(n4723) V(n4724) V(n4725) V(n4726) V(n4727) V(n4728) V(n4729) V(n4730) V(n4731) V(n4732) V(n4733) V(n4734) V(n4735) V(n4736) V(n4737) V(n4738) V(n4739) V(n4740) V(n4741) V(n4742) V(n4743) V(n4744) V(n4745) V(n4746) V(n4747) V(n4748) V(n4749) V(n4750) V(n4751) V(n4752) V(n4753) V(n4754) V(n4755) V(n4756) V(n4757) V(n4758) V(n4759) V(n4760) V(n4761) V(n4762) V(n4763) V(n4764) V(n4765) V(n4766) V(n4767) V(n4768) V(n4769) V(n4770) V(n4771) V(n4772) V(n4773) V(n4774) V(n4775) V(n4776) V(n4777) V(n4778) V(n1) V(n4780) V(n4781) V(n4782) V(n4783) V(n4784) V(n4785) V(n4786) V(n4787) V(n4788) V(n4789) V(n4790) V(n4791) V(n4792) V(n4793) V(n4794) V(n4795) V(n4796) V(n4797) V(n4798) V(n4799) V(n4800) V(n4801) V(n4802) V(n4803) V(n4804) V(n4805) V(n4806) V(n4807) V(n1) V(n4809) V(n4810) V(n4811) V(n4812) V(n4813) V(n4814) V(n4815) V(n4816) V(n4817) V(n4818) V(n4819) V(n4820) V(n4821) V(n4822) V(n4823) V(n4824) V(n4825) V(n4826) V(n4827) V(n4828) V(n4829) V(n4830) V(n4831) V(n4832) V(n4833) V(n4834) V(n4835) V(n4836) V(n4837) V(n4838) V(n4839) V(n4840) V(n4841) V(n4842) V(n4843) V(n4844) V(n4845) V(n4846) V(n4847) V(n4848) V(n4849) V(n4850) V(n4851) V(n4852) V(n4853) V(n4854) V(n4855) V(n4856) V(n4857) V(n4858) V(n4859) V(n4860) V(n4861) V(n4862) V(n4863) V(n4864) V(n4865) V(n4866) V(n4867) V(n4868) V(n4869) V(n4870) V(n4871) V(n4872) V(n4873) V(n4874) V(n4875) V(n4876) V(n4877) V(n4878) V(n4879) V(n4880) V(n4881) V(n4882) V(n4883) V(n4884) V(n4885) V(n4886) V(n4887) V(n4888) V(n4889) V(n4890) V(n4891) V(n4892) V(n4893) V(n4894) V(n4895) V(n4896) V(n4897) V(n4898) V(n4899) V(n4900) V(n4901) V(n4902) V(n4903) V(n4904) V(n4905) V(n4906) V(n4907) V(n4908) V(n4909) V(n4910) V(n4911) V(n4912) V(n4913) V(n4914) V(n4915) V(n4916) V(n4917) V(n4918) V(n4919) V(n1) V(n4921) V(n4922) V(n4923) V(n4924) V(n4925) V(n4926) V(n4927) V(n4928) V(n4929) V(n4930) V(n4931) V(n4932) V(n4933) V(n4934) V(n4935) V(n4936) V(n4937) V(n4938) V(n4939) V(n4940) V(n4941) V(n4942) V(n4943) V(n4944) V(n4945) V(n4946) V(n4947) V(n4948) V(n4949) V(n4950) V(n4951) V(n4952) V(n4953) V(n4954) V(n4955) V(n4956) V(n4957) V(n4958) V(n4959) V(n4960) V(n4961) V(n4962) V(n4963) V(n4964) V(n4965) V(n4966) V(n4967) V(n4968) V(n4969) V(n4970) V(n4971) V(n4972) V(n4973) V(n4974) V(n4975) V(n4976) V(n4977) V(n4978) V(n4979) V(n4980) V(n4981) V(n4982) V(n4983) V(n4984) V(n4985) V(n4986) V(n4987) V(n4988) V(n4989) V(n4990) V(n4991) V(n4992) V(n4993) V(n4994) V(n4995) V(n4996) V(n1) V(n4998) V(n4999) V(n5000) V(n5001) V(n5002) V(n5003) V(n5004) V(n5005) V(n5006) V(n5007) V(n5008) V(n5009) V(n5010) V(n5011) V(n5012) V(n5013) V(n5014) V(n5015) V(n5016) V(n5017) V(n5018) V(n5019) V(n5020) V(n5021) V(n5022) V(n5023) V(n5024) V(n5025) V(n5026) V(n5027) V(n5028) V(n5029) V(n5030) V(n5031) V(n5032) V(n5033) V(n5034) V(n5035) V(n5036) V(n5037) V(n5038) V(n5039) V(n5040) V(n5041) V(n5042) V(n5043) V(n5044) V(n5045) V(n5046) V(n5047) V(n5048) V(n5049) V(n5050) V(n5051) V(n5052) V(n5053) V(n5054) V(n5055) V(n5056) V(n5057) V(n5058) V(n5059) V(n5060) V(n5061) V(n5062) V(n5063) V(n5064) V(n5065) V(n5066) V(n5067) V(n5068) V(n5069) V(n5070) V(n5071) V(n5072) V(n5073) V(n5074) V(n5075) V(n5076) V(n5077) V(n5078) V(n5079) V(n5080) V(n5081) V(n5082) V(n5083) V(n5084) V(n5085) V(n5086) V(n5087) V(n5088) V(n5089) V(n5090) V(n5091) V(n5092) V(n5093) V(n5094) V(n1) V(n5096) V(n5097) V(n5098) V(n5099) V(n5100) V(n5101) V(n5102) V(n5103) V(n5104) V(n5105) V(n5106) V(n5107) V(n5108) V(n5109) V(n5110) V(n5111) V(n5112) V(n5113) V(n5114) V(n5115) V(n5116) V(n5117) V(n5118) V(n5119) V(n5120) V(n5121) V(n5122) V(n5123) V(n5124) V(n5125) V(n5126) V(n5127) V(n5128) V(n5129) V(n5130) V(n5131) V(n5132) V(n5133) V(n5134) V(n5135) V(n5136) V(n5137) V(n5138) V(n5139) V(n5140) V(n5141) V(n5142) V(n5143) V(n5144) V(n5145) V(n5146) V(n5147) V(n5148) V(n5149) V(n5150) V(n5151) V(n5152) V(n5153) V(n5154) V(n5155) V(n5156) V(n5157) V(n5158) V(n5159) V(n5160) V(n5161) V(n5162) V(n5163) V(n5164) V(n5165) V(n5166) V(n5167) V(n5168) V(n5169) V(n5170) V(n5171) V(n5172) V(n5173) V(n5174) V(n5175) V(n5176) V(n5177) V(n5178) V(n5179) V(n5180) V(n5181) V(n5182) V(n5183) V(n5184) V(n5185) V(n5186) V(n5187) V(n5188) V(n5189) V(n5190) V(n5191) V(n5192) V(n5193) V(n5194) V(n5195) V(n5196) V(n5197) V(n5198) V(n5199) V(n5200) V(n5201) V(n5202) V(n5203) V(n5204) V(n5205) V(n5206) V(n5207) V(n5208) V(n5209) V(n1) V(n5211) V(n5212) V(n5213) V(n5214) V(n5215) V(n5216) V(n5217) V(n5218) V(n5219) V(n5220) V(n5221) V(n5222) V(n5223) V(n5224) V(n5225) V(n5226) V(n5227) V(n5228) V(n5229) V(n5230) V(n5231) V(n5232) V(n5233) V(n5234) V(n5235) V(n5236) V(n5237) V(n5238) V(n5239) V(n5240) V(n5241) V(n5242) V(n5243) V(n1) V(n5245) V(n5246) V(n5247) V(n5248) V(n5249) V(n5250) V(n5251) V(n5252) V(n5253) V(n5254) V(n5255) V(n5256) V(n5257) V(n5258) V(n5259) V(n5260) V(n5261) V(n5262) V(n5263) V(n5264) V(n5265) V(n5266) V(n5267) V(n5268) V(n5269) V(n5270) V(n5271) V(n5272) V(n5273) V(n5274) V(n5275) V(n5276) V(n5277) V(n5278) V(n5279) V(n5280) V(n5281) V(n5282) V(n5283) V(n5284) V(n5285) V(n5286) V(n5287) V(n5288) V(n5289) V(n5290) V(n5291) V(n5292) V(n5293) V(n5294) V(n5295) V(n5296) V(n5297) V(n5298) V(n5299) V(n5300) V(n5301) V(n5302) V(n5303) V(n5304) V(n5305) V(n5306) V(n5307) V(n5308) V(n5309) V(n5310) V(n5311) V(n5312) V(n5313) V(n5314) V(n5315) V(n5316) V(n5317) V(n5318) V(n5319) V(n5320) V(n5321) V(n5322) V(n5323) V(n5324) V(n5325) V(n5326) V(n5327) V(n5328) V(n5329) V(n5330) V(n5331) V(n5332) V(n5333) V(n5334) V(n5335) V(n5336) V(n5337) V(n5338) V(n5339) V(n5340) V(n5341) V(n5342) V(n5343) V(n5344) V(n5345) V(n5346) V(n5347) V(n5348) V(n5349) V(n5350) V(n5351) V(n5352) V(n5353) V(n5354) V(n5355) V(n5356) V(n5357) V(n5358) V(n5359) V(n5360) V(n5361) V(n5362) V(n5363) V(n5364) V(n5365) V(n5366) V(n5367) V(n5368) V(n5369) V(n5370) V(n5371) V(n5372) V(n5373) V(n5374) V(n5375) V(n5376) V(n5377) V(n5378) V(n5379) V(n5380) V(n5381) V(n5382) V(n5383) V(n5384) V(n5385) V(n5386) V(n5387) V(n5388) V(n5389) V(n5390) V(n5391) V(n5392) V(n5393) V(n5394) V(n5395) V(n5396) V(n5397) V(n5398) V(n5399) V(n5400) V(n5401) V(n5402) V(n5403) V(n5404) V(n5405) V(n5406) V(n5407) V(n5408) V(n5409) V(n5410) V(n5411) V(n5412) V(n5413) V(n5414) V(n5415) V(n5416) V(n5417) V(n5418) V(n5419) V(n5420) V(n5421) V(n5422) V(n5423) V(n5424) V(n5425) V(n5426) V(n5427) V(n5428) V(n5429) V(n5430) V(n5431) V(n5432) V(n5433) V(n5434) V(n5435) V(n5436) V(n5437) V(n5438) V(n5439) V(n5440) V(n5441) V(n5442) V(n5443) V(n5444) V(n5445) V(n5446) V(n5447) V(n5448) V(n5449) V(n5450) V(n5451) V(n5452) V(n5453) V(n5454) V(n5455) V(n5456) V(n5457) V(n5458) V(n5459) V(n5460) V(n5461) V(n5462) V(n1) V(n5464) V(n5465) V(n5466) V(n5467) V(n5468) V(n5469) V(n5470) V(n5471) V(n5472) V(n5473) V(n5474) V(n5475) V(n5476) V(n5477) V(n5478) V(n5479) V(n5480) V(n5481) V(n5482) V(n5483) V(n5484) V(n5485) V(n5486) V(n5487) V(n5488) V(n5489) V(n5490) V(n5491) V(n5492) V(n5493) V(n5494) V(n5495) V(n5496) V(n5497) V(n5498) V(n5499) V(n5500) V(n5501) V(n5502) V(n5503) V(n1) V(n5505) V(n5506) V(n5507) V(n5508) V(n5509) V(n5510) V(n5511) V(n5512) V(n5513) V(n5514) V(n5515) V(n5516) V(n5517) V(n5518) V(n5519) V(n5520) V(n5521) V(n5522) V(n5523) V(n1) V(n5525) V(n5526) V(n5527) V(n5528) V(n5529) V(n5530) V(n5531) V(n5532) V(n5533) V(n5534) V(n5535) V(n5536) V(n5537) V(n5538) V(n5539) V(n5540) V(n5541) V(n5542) V(n5543) V(n5544) V(n5545) V(n5546) V(n5547) V(n5548) V(n5549) V(n5550) V(n5551) V(n5552) V(n5553) V(n5554) V(n5555) V(n5556) V(n5557) V(n5558) V(n5559) V(n5560) V(n5561) V(n5562) V(n5563) V(n5564) V(n5565) V(n5566) V(n5567) V(n5568) V(n5569) V(n5570) V(n1) V(n5572) V(n5573) V(n5574) V(n5575) V(n5576) V(n5577) V(n5578) V(n5579) V(n5580) V(n5581) V(n5582) V(n5583) V(n5584) V(n5585) V(n5586) V(n5587) V(n5588) V(n5589) V(n5590) V(n5591) V(n5592) V(n5593) V(n5594) V(n5595) V(n5596) V(n5597) V(n5598) V(n5599) V(n5600) V(n5601) V(n5602) V(n1) V(n5604) V(n5605) V(n5606) V(n5607) V(n5608) V(n5609) V(n5610) V(n5611) V(n5612) V(n5613) V(n5614) V(n5615) V(n5616) V(n5617) V(n5618) V(n5619) V(n5620) V(n5621) V(n5622) V(n5623) V(n5624) V(n5625) V(n5626) V(n5627) V(n5628) V(n5629) V(n5630) V(n5631) V(n5632) V(n5633) V(n5634) V(n5635) V(n5636) V(n5637) V(n5638) V(n5639) V(n5640) V(n5641) V(n5642) V(n5643) V(n5644) V(n5645) V(n5646) V(n5647) V(n5648) V(n5649) V(n5650) V(n5651) V(n5652) V(n5653) V(n5654) V(n5655) V(n5656) V(n5657) V(n5658) V(n5659) V(n5660) V(n5661) V(n5662) V(n5663) V(n5664) V(n5665) V(n5666) V(n5667) V(n5668) V(n5669) V(n5670) V(n5671) V(n5672) V(n5673) V(n5674) V(n5675) V(n5676) V(n5677) V(n5678) V(n5679) V(n5680) V(n5681) V(n5682) V(n5683) V(n5684) V(n5685) V(n5686) V(n5687) V(n5688) V(n5689) V(n5690) V(n5691) V(n5692) V(n5693) V(n5694) V(n5695) V(n5696) V(n5697) V(n5698) V(n5699) V(n5700) V(n5701) V(n5702) V(n5703) V(n5704) V(n5705) V(n5706) V(n5707) V(n1) V(n5709) V(n5710) V(n5711) V(n5712) V(n5713) V(n5714) V(n5715) V(n5716) V(n5717) V(n5718) V(n5719) V(n5720) V(n5721) V(n5722) V(n5723) V(n5724) V(n5725) V(n5726) V(n5727) V(n5728) V(n5729) V(n5730) V(n5731) V(n5732) V(n5733) V(n5734) V(n5735) V(n5736) V(n5737) V(n5738) V(n5739) V(n5740) V(n5741) V(n5742) V(n5743) V(n5744) V(n5745) V(n5746) V(n5747) V(n5748) V(n5749) V(n5750) V(n5751) V(n5752) V(n5753) V(n5754) V(n5755) V(n5756) V(n5757) V(n5758) V(n5759) V(n5760) V(n5761) V(n5762) V(n5763) V(n5764) V(n5765) V(n5766) V(n5767) V(n5768) V(n5769) V(n5770) V(n5771) V(n5772) V(n5773) V(n5774) V(n5775) V(n5776) V(n5777) V(n5778) V(n5779) V(n5780) V(n5781) V(n5782) V(n5783) V(n5784) V(n5785) V(n5786) V(n5787) V(n5788) V(n5789) V(n5790) V(n5791) V(n5792) V(n5793) V(n5794) V(n5795) V(n5796) V(n5797) V(n5798) V(n5799) V(n5800) V(n5801) V(n5802) V(n5803) V(n5804) V(n5805) V(n5806) V(n5807) V(n5808) V(n5809) V(n5810) V(n5811) V(n5812) V(n5813) V(n5814) V(n5815) V(n5816) V(n5817) V(n5818) V(n5819) V(n5820) V(n5821) V(n5822) V(n5823) V(n5824) V(n5825) V(n5826) V(n5827) V(n5828) V(n5829) V(n5830) V(n5831) V(n5832) V(n5833) V(n5834) V(n5835) V(n5836) V(n5837) V(n5838) V(n5839) V(n5840) V(n5841) V(n5842) V(n5843) V(n5844) V(n5845) V(n5846) V(n5847) V(n5848) V(n5849) V(n5850) V(n5851) V(n5852) V(n5853) V(n5854) V(n5855) V(n5856) V(n5857) V(n5858) V(n5859) V(n5860) V(n5861) V(n5862) V(n5863) V(n5864) V(n5865) V(n5866) V(n5867) V(n5868) V(n5869) V(n5870) V(n5871) V(n5872) V(n5873) V(n5874) V(n5875) V(n5876) V(n5877) V(n5878) V(n5879) V(n5880) V(n5881) V(n5882) V(n5883) V(n5884) V(n5885) V(n5886) V(n5887) V(n5888) V(n5889) V(n5890) V(n5891) V(n5892) V(n5893) V(n5894) V(n5895) V(n5896) V(n5897) V(n5898) V(n5899) V(n5900) V(n5901) V(n5902) V(n5903) V(n5904) V(n5905) V(n5906) V(n5907) V(n5908) V(n5909) V(n1) V(n5911) V(n5912) V(n5913) V(n5914) V(n5915) V(n5916) V(n5917) V(n5918) V(n5919) V(n5920) V(n5921) V(n5922) V(n5923) V(n5924) V(n5925) V(n5926) V(n5927) V(n5928) V(n5929) V(n5930) V(n5931) V(n5932) V(n1) V(n5934) V(n5935) V(n5936) V(n5937) V(n5938) V(n5939) V(n5940) V(n5941) V(n5942) V(n5943) V(n5944) V(n5945) V(n5946) V(n5947) V(n5948) V(n5949) V(n5950) V(n5951) V(n5952) V(n5953) V(n5954) V(n5955) V(n5956) V(n5957) V(n5958) V(n5959) V(n5960) V(n5961) V(n5962) V(n5963) V(n5964) V(n5965) V(n5966) V(n5967) V(n5968) V(n5969) V(n5970) V(n5971) V(n5972) V(n5973) V(n5974) V(n5975) V(n5976) V(n5977) V(n5978) V(n5979) V(n5980) V(n5981) V(n5982) V(n5983) V(n5984) V(n5985) V(n5986) V(n5987) V(n5988) V(n5989) V(n5990) V(n5991) V(n5992) V(n5993) V(n5994) V(n5995) V(n5996) V(n5997) V(n5998) V(n5999) V(n6000) V(n6001) V(n6002) V(n6003) V(n6004) V(n6005) V(n6006) V(n6007) V(n6008) V(n6009) V(n6010) V(n6011) V(n6012) V(n6013) V(n6014) V(n6015) V(n6016) V(n6017) V(n6018) V(n6019) V(n6020) V(n6021) V(n6022) V(n6023) V(n6024) V(n6025) V(n6026) V(n6027) V(n6028) V(n6029) V(n6030) V(n6031) V(n6032) V(n6033) V(n6034) V(n6035) V(n6036) V(n6037) V(n6038) V(n6039) V(n6040) V(n6041) V(n1) V(n6043) V(n6044) V(n6045) V(n6046) V(n6047) V(n6048) V(n6049) V(n6050) V(n6051) V(n6052) V(n6053) V(n6054) V(n6055) V(n6056) V(n6057) V(n6058) V(n6059) V(n6060) V(n6061) V(n6062) V(n6063) V(n6064) V(n6065) V(n6066) V(n6067) V(n6068) V(n6069) V(n6070) V(n6071) V(n6072) V(n6073) V(n6074) V(n6075) V(n6076) V(n6077) V(n6078) V(n6079) V(n6080) V(n6081) V(n6082) V(n6083) V(n6084) V(n6085) V(n6086) V(n6087) V(n6088) V(n6089) V(n6090) V(n6091) V(n6092) V(n6093) V(n6094) V(n6095) V(n6096) V(n6097) V(n6098) V(n6099) V(n6100) V(n6101) V(n6102) V(n6103) V(n6104) V(n6105) V(n6106) V(n6107) V(n6108) V(n6109) V(n6110) V(n6111) V(n6112) V(n6113) V(n6114) V(n6115) V(n6116) V(n6117) V(n6118) V(n6119) V(n1) V(n6121) V(n6122) V(n6123) V(n6124) V(n6125) V(n6126) V(n6127) V(n6128) V(n6129) V(n6130) V(n6131) V(n6132) V(n6133) V(n6134) V(n6135) V(n6136) V(n6137) V(n6138) V(n6139) V(n6140) V(n6141) V(n6142) V(n6143) V(n6144) V(n6145) V(n6146) V(n6147) V(n6148) V(n6149) V(n6150) V(n6151) V(n6152) V(n6153) V(n6154) V(n6155) V(n6156) V(n6157) V(n6158) V(n6159) V(n6160) V(n6161) V(n6162) V(n6163) V(n6164) V(n6165) V(n6166) V(n6167) V(n6168) V(n6169) V(n6170) V(n6171) V(n6172) V(n6173) V(n6174) V(n1) V(n6176) V(n6177) V(n6178) V(n6179) V(n6180) V(n6181) V(n6182) V(n6183) V(n6184) V(n6185) V(n6186) V(n6187) V(n6188) V(n6189) V(n6190) V(n6191) V(n6192) V(n6193) V(n6194) V(n6195) V(n6196) V(n6197) V(n6198) V(n6199) V(n6200) V(n6201) V(n6202) V(n6203) V(n6204) V(n6205) V(n6206) V(n6207) V(n6208) V(n6209) V(n6210) V(n6211) V(n6212) V(n6213) V(n6214) V(n6215) V(n6216) V(n6217) V(n6218) V(n6219) V(n6220) V(n6221) V(n6222) V(n6223) V(n6224) V(n6225) V(n6226) V(n6227) V(n6228) V(n6229) V(n6230) V(n6231) V(n6232) V(n6233) V(n6234) V(n6235) V(n6236) V(n6237) V(n6238) V(n6239) V(n6240) V(n6241) V(n6242) V(n6243) V(n6244) V(n6245) V(n6246) V(n6247) V(n6248) V(n6249) V(n6250) V(n6251) V(n6252) V(n6253) V(n6254) V(n6255) V(n6256) V(n6257) V(n6258) V(n6259) V(n6260) V(n6261) V(n6262) V(n6263) V(n6264) V(n6265) V(n6266) V(n6267) V(n6268) V(n6269) V(n6270) V(n6271) V(n6272) V(n6273) V(n6274) V(n6275) V(n6276) V(n6277) V(n6278) V(n6279) V(n6280) V(n6281) V(n6282) V(n6283) V(n6284) V(n6285) V(n6286) V(n6287) V(n6288) V(n6289) V(n6290) V(n6291) V(n6292) V(n6293) V(n6294) V(n6295) V(n6296) V(n6297) V(n6298) V(n6299) V(n6300) V(n6301) V(n6302) V(n6303) V(n6304) V(n6305) V(n6306) V(n6307) V(n6308) V(n6309) V(n6310) V(n6311) V(n6312) V(n6313) V(n6314) V(n6315) V(n6316) V(n6317) V(n6318) V(n6319) V(n6320) V(n6321) V(n6322) V(n6323) V(n6324) V(n6325) V(n6326) V(n6327) V(n6328) V(n6329) V(n6330) V(n6331) V(n6332) V(n6333) V(n6334) V(n6335) V(n6336) V(n6337) V(n6338) V(n6339) V(n6340) V(n6341) V(n6342) V(n1) V(n6344) V(n6345) V(n6346) V(n6347) V(n6348) V(n6349) V(n6350) V(n6351) V(n6352) V(n6353) V(n6354) V(n6355) V(n6356) V(n6357) V(n6358) V(n6359) V(n6360) V(n6361) V(n6362) V(n6363) V(n6364) V(n6365) V(n6366) V(n6367) V(n6368) V(n6369) V(n6370) V(n6371) V(n6372) V(n6373) V(n6374) V(n6375) V(n6376) V(n6377) V(n6378) V(n6379) V(n6380) V(n6381) V(n6382) V(n6383) V(n6384) V(n6385) V(n6386) V(n6387) V(n6388) V(n6389) V(n6390) V(n6391) V(n6392) V(n6393) V(n6394) V(n6395) V(n6396) V(n6397) V(n6398) V(n6399) V(n6400) V(n6401) V(n6402) V(n6403) V(n6404) V(n6405) V(n6406) V(n6407) V(n6408) V(n6409) V(n6410) V(n6411) V(n6412) V(n6413) V(n6414) V(n6415) V(n6416) V(n6417) V(n6418) V(n6419) V(n6420) V(n6421) V(n6422) V(n6423) V(n6424) V(n6425) V(n6426) V(n6427) V(n6428) V(n6429) V(n6430) V(n6431) V(n6432) V(n6433) V(n6434) V(n6435) V(n6436) V(n6437) V(n6438) V(n6439) V(n6440) V(n6441) V(n6442) V(n6443) V(n6444) V(n6445) V(n6446) V(n6447) V(n6448) V(n6449) V(n6450) V(n6451) V(n6452) V(n6453) V(n6454) V(n6455) V(n6456) V(n6457) V(n6458) V(n6459) V(n6460) V(n6461) V(n6462) V(n6463) V(n6464) V(n6465) V(n6466) V(n6467) V(n6468) V(n6469) V(n1) V(n6471) V(n6472) V(n6473) V(n6474) V(n6475) V(n6476) V(n6477) V(n6478) V(n6479) V(n6480) V(n6481) V(n6482) V(n6483) V(n6484) V(n6485) V(n6486) V(n6487) V(n6488) V(n6489) V(n6490) V(n6491) V(n6492) V(n6493) V(n6494) V(n6495) V(n6496) V(n6497) V(n6498) V(n6499) V(n6500) V(n6501) V(n6502) V(n6503) V(n6504) V(n6505) V(n6506) V(n6507) V(n6508) V(n6509) V(n6510) V(n6511) V(n6512) V(n6513) V(n6514) V(n6515) V(n6516) V(n6517) V(n6518) V(n6519) V(n6520) V(n6521) V(n6522) V(n6523) V(n6524) V(n6525) V(n6526) V(n6527) V(n6528) V(n6529) V(n6530) V(n6531) V(n6532) V(n6533) V(n6534) V(n6535) V(n6536) V(n6537) V(n6538) V(n6539) V(n6540) V(n6541) V(n6542) V(n6543) V(n6544) V(n6545) V(n6546) V(n6547) V(n6548) V(n6549) V(n6550) V(n6551) V(n6552) V(n6553) V(n6554) V(n6555) V(n6556) V(n6557) V(n6558) V(n6559) V(n6560) V(n6561) V(n6562) V(n6563) V(n6564) V(n6565) V(n6566) V(n6567) V(n6568) V(n6569) V(n6570) V(n6571) V(n6572) V(n6573) V(n6574) V(n6575) V(n6576) V(n6577) V(n6578) V(n6579) V(n6580) V(n6581) V(n6582) V(n6583) V(n6584) V(n6585) V(n6586) V(n6587) V(n6588) V(n6589) V(n6590) V(n6591) V(n6592) V(n6593) V(n6594) V(n6595) V(n6596) V(n6597) V(n6598) V(n6599) V(n6600) V(n6601) V(n6602) V(n6603) V(n6604) V(n6605) V(n6606) V(n6607) V(n6608) V(n6609) V(n6610) V(n6611) V(n6612) V(n6613) V(n6614) V(n6615) V(n6616) V(n6617) V(n6618) V(n6619) V(n6620) V(n6621) V(n6622) V(n6623) V(n6624) V(n6625) V(n6626) V(n6627) V(n6628) V(n6629) V(n6630) V(n6631) V(n6632) V(n6633) V(n6634) V(n6635) V(n6636) V(n6637) V(n6638) V(n6639) V(n6640) V(n6641) V(n6642) V(n6643) V(n6644) V(n6645) V(n6646) V(n1) V(n6648) V(n6649) V(n6650) V(n6651) V(n6652) V(n6653) V(n6654) V(n6655) V(n6656) V(n6657) V(n6658) V(n6659) V(n6660) V(n6661) V(n6662) V(n6663) V(n6664) V(n6665) V(n6666) V(n6667) V(n6668) V(n6669) V(n6670) V(n6671) V(n6672) V(n6673) V(n6674) V(n6675) V(n6676) V(n6677) V(n6678) V(n6679) V(n6680) V(n6681) V(n6682) V(n6683) V(n6684) V(n6685) V(n6686) V(n6687) V(n6688) V(n6689) V(n6690) V(n6691) V(n6692) V(n6693) V(n6694) V(n6695) V(n6696) V(n6697) V(n6698) V(n6699) V(n6700) V(n6701) V(n6702) V(n6703) V(n6704) V(n6705) V(n6706) V(n6707) V(n6708) V(n6709) V(n6710) V(n6711) V(n6712) V(n6713) V(n6714) V(n6715) V(n6716) V(n6717) V(n6718) V(n6719) V(n6720) V(n6721) V(n6722) V(n6723) V(n6724) V(n6725) V(n6726) V(n6727) V(n6728) V(n6729) V(n6730) V(n6731) V(n6732) V(n6733) V(n6734) V(n6735) V(n6736) V(n6737) V(n6738) V(n6739) V(n6740) V(n6741) V(n6742) V(n6743) V(n6744) V(n6745) V(n6746) V(n6747) V(n6748) V(n6749) V(n6750) V(n6751) V(n6752) V(n6753) V(n6754) V(n6755) V(n6756) V(n6757) V(n6758) V(n6759) V(n6760) V(n6761) V(n6762) V(n6763) V(n6764) V(n6765) V(n6766) V(n6767) V(n6768) V(n6769) V(n6770) V(n6771) V(n6772) V(n6773) V(n6774) V(n6775) V(n6776) V(n6777) V(n6778) V(n6779) V(n6780) V(n6781) V(n6782) V(n6783) V(n6784) V(n6785) V(n6786) V(n6787) V(n6788) V(n6789) V(n6790) V(n6791) V(n6792) V(n6793) V(n6794) V(n6795) V(n6796) V(n6797) V(n6798) V(n6799) V(n6800) V(n6801) V(n6802) V(n6803) V(n6804) V(n6805) V(n6806) V(n6807) V(n6808) V(n6809) V(n6810) V(n6811) V(n6812) V(n6813) V(n6814) V(n6815) V(n6816) V(n6817) V(n6818) V(n6819) V(n6820) V(n6821) V(n6822) V(n6823) V(n6824) V(n6825) V(n6826) V(n6827) V(n6828) V(n6829) V(n6830) V(n6831) V(n6832) V(n6833) V(n6834) V(n6835) V(n6836) V(n6837) V(n6838) V(n6839) V(n6840) V(n6841) V(n6842) V(n6843) V(n6844) V(n6845) V(n6846) V(n6847) V(n6848) V(n6849) V(n6850) V(n6851) V(n6852) V(n6853) V(n6854) V(n6855) V(n6856) V(n6857) V(n6858) V(n6859) V(n6860) V(n6861) V(n6862) V(n6863) V(n6864) V(n6865) V(n6866) V(n6867) V(n6868) V(n6869) V(n6870) V(n6871) V(n6872) V(n6873) V(n6874) V(n6875) V(n6876) V(n6877) V(n6878) V(n6879) V(n6880) V(n6881) V(n6882) V(n6883) V(n6884) V(n6885) V(n6886) V(n6887) V(n6888) V(n6889) V(n6890) V(n6891) V(n6892) V(n6893) V(n6894) V(n6895) V(n6896) V(n6897) V(n6898) V(n6899) V(n6900) V(n6901) V(n6902) V(n6903) V(n6904) V(n6905) V(n6906) V(n6907) V(n6908) V(n6909) V(n6910) V(n6911) V(n6912) V(n6913) V(n6914) V(n6915) V(n6916) V(n6917) V(n6918) V(n6919) V(n6920) V(n6921) V(n6922) V(n6923) V(n6924) V(n6925) V(n6926) V(n6927) V(n6928) V(n6929) V(n6930) V(n6931) V(n6932) V(n6933) V(n6934) V(n6935) V(n6936) V(n6937) V(n6938) V(n6939) V(n6940) V(n6941) V(n6942) V(n6943) V(n6944) V(n6945) V(n6946) V(n6947) V(n6948) V(n6949) V(n6950) V(n6951) V(n6952) V(n6953) V(n6954) V(n6955) V(n6956) V(n6957) V(n6958) V(n6959) V(n6960) V(n6961) V(n6962) V(n6963) V(n6964) V(n6965) V(n6966) V(n1) V(n6968) V(n6969) V(n6970) V(n6971) V(n6972) V(n6973) V(n6974) V(n6975) V(n6976) V(n6977) V(n6978) V(n6979) V(n6980) V(n6981) V(n6982) V(n6983) V(n6984) V(n6985) V(n6986) V(n6987) V(n6988) V(n6989) V(n6990) V(n6991) V(n6992) V(n6993) V(n6994) V(n6995) V(n6996) V(n6997) V(n6998) V(n6999) V(n7000) V(n7001) V(n7002) V(n7003) V(n7004) V(n7005) V(n7006) V(n7007) V(n7008) V(n7009) V(n7010) V(n7011) V(n7012) V(n7013) V(n7014) V(n7015) V(n7016) V(n7017) V(n7018) V(n7019) V(n7020) V(n7021) V(n7022) V(n7023) V(n7024) V(n7025) V(n7026) V(n7027) V(n7028) V(n7029) V(n7030) V(n7031) V(n7032) V(n7033) V(n7034) V(n7035) V(n7036) V(n7037) V(n7038) V(n7039) V(n7040) V(n7041) V(n7042) V(n7043) V(n7044) V(n7045) V(n7046) V(n7047) V(n7048) V(n7049) V(n7050) V(n7051) V(n7052) V(n7053) V(n7054) V(n7055) V(n7056) V(n7057) V(n7058) V(n7059) V(n7060) V(n7061) V(n7062) V(n7063) V(n7064) V(n7065) V(n7066) V(n7067) V(n7068) V(n7069) V(n7070) V(n7071) V(n7072) V(n7073) V(n7074) V(n7075) V(n7076) V(n7077) V(n7078) V(n7079) V(n7080) V(n7081) V(n7082) V(n7083) V(n7084) V(n7085) V(n7086) V(n7087) V(n7088) V(n7089) V(n7090) V(n7091) V(n7092) V(n7093) V(n7094) V(n7095) V(n7096) V(n7097) V(n7098) V(n7099) V(n7100) V(n7101) V(n7102) V(n7103) V(n7104) V(n7105) V(n7106) V(n7107) V(n7108) V(n7109) V(n7110) V(n7111) V(n7112) V(n7113) V(n7114) V(n7115) V(n7116) V(n7117) V(n7118) V(n7119) V(n7120) V(n7121) V(n7122) V(n7123) V(n7124) V(n7125) V(n7126) V(n7127) V(n7128) V(n7129) V(n7130) V(n7131) V(n7132) V(n7133) V(n7134) V(n7135) V(n7136) V(n7137) V(n7138) V(n7139) V(n7140) V(n7141) V(n7142) V(n7143) V(n7144) V(n7145) V(n7146) V(n7147) V(n7148) V(n7149) V(n7150) V(n7151) V(n7152) V(n7153) V(n7154) V(n7155) V(n7156) V(n7157) V(n7158) V(n7159) V(n7160) V(n7161) V(n7162) V(n7163) V(n7164) V(n7165) V(n7166) V(n7167) V(n7168) V(n1) V(n7170) V(n7171) V(n7172) V(n7173) V(n7174) V(n7175) V(n7176) V(n7177) V(n7178) V(n7179) V(n7180) V(n7181) V(n7182) V(n7183) V(n7184) V(n7185) V(n7186) V(n7187) V(n7188) V(n7189) V(n7190) V(n7191) V(n7192) V(n7193) V(n7194) V(n7195) V(n7196) V(n7197) V(n7198) V(n7199) V(n7200) V(n7201) V(n7202) V(n7203) V(n7204) V(n7205) V(n7206) V(n7207) V(n7208) V(n7209) V(n7210) V(n7211) V(n7212) V(n7213) V(n7214) V(n7215) V(n7216) V(n7217) V(n7218) V(n7219) V(n7220) V(n7221) V(n7222) V(n7223) V(n7224) V(n7225) V(n7226) V(n7227) V(n7228) V(n7229) V(n7230) V(n7231) V(n7232) V(n7233) V(n7234) V(n7235) V(n7236) V(n7237) V(n7238) V(n7239) V(n7240) V(n7241) V(n7242) V(n7243) V(n7244) V(n7245) V(n7246) V(n7247) V(n7248) V(n7249) V(n7250) V(n7251) V(n7252) V(n7253) V(n7254) V(n7255) V(n7256) V(n7257) V(n7258) V(n7259) V(n7260) V(n7261) V(n7262) V(n7263) V(n7264) V(n7265) V(n7266) V(n7267) V(n7268) V(n7269) V(n7270) V(n7271) V(n7272) V(n7273) V(n7274) V(n7275) V(n7276) V(n7277) V(n7278) V(n7279) V(n7280) V(n7281) V(n7282) V(n7283) V(n7284) V(n7285) V(n7286) V(n7287) V(n7288) V(n7289) V(n7290) V(n7291) V(n7292) V(n7293) V(n7294) V(n7295) V(n7296) V(n7297) V(n7298) V(n7299) V(n7300) V(n7301) V(n7302) V(n1) V(n7304) V(n7305) V(n7306) V(n7307) V(n7308) V(n7309) V(n7310) V(n7311) V(n7312) V(n7313) V(n7314) V(n7315) V(n7316) V(n7317) V(n7318) V(n7319) V(n7320) V(n7321) V(n7322) V(n7323) V(n7324) V(n7325) V(n7326) V(n7327) V(n7328) V(n7329) V(n7330) V(n7331) V(n7332) V(n7333) V(n7334) V(n7335) V(n7336) V(n7337) V(n7338) V(n7339) V(n7340) V(n7341) V(n7342) V(n7343) V(n7344) V(n7345) V(n7346) V(n7347) V(n7348) V(n7349) V(n7350) V(n7351) V(n7352) V(n7353) V(n7354) V(n7355) V(n7356) V(n7357) V(n7358) V(n1) V(n7360) V(n7361) V(n7362) V(n7363) V(n7364) V(n7365) V(n7366) V(n7367) V(n7368) V(n7369) V(n7370) V(n7371) V(n7372) V(n7373) V(n7374) V(n7375) V(n7376) V(n7377) V(n7378) V(n7379) V(n7380) V(n7381) V(n7382) V(n7383) V(n7384) V(n7385) V(n7386) V(n7387) V(n7388) V(n7389) V(n7390) V(n7391) V(n7392) V(n7393) V(n7394) V(n7395) V(n7396) V(n7397) V(n7398) V(n7399) V(n7400) V(n7401) V(n7402) V(n7403) V(n7404) V(n7405) V(n7406) V(n7407) V(n7408) V(n7409) V(n7410) V(n7411) V(n7412) V(n7413) V(n7414) V(n7415) V(n7416) V(n7417) V(n7418) V(n7419) V(n7420) V(n7421) V(n7422) V(n7423) V(n7424) V(n7425) V(n7426) V(n7427) V(n7428) V(n7429) V(n7430) V(n7431) V(n7432) V(n7433) V(n7434) V(n7435) V(n7436) V(n7437) V(n7438) V(n7439) V(n7440) V(n7441) V(n7442) V(n7443) V(n7444) V(n7445) V(n7446) V(n7447) V(n7448) V(n7449) V(n7450) V(n7451) V(n7452) V(n7453) V(n7454) V(n7455) V(n7456) V(n7457) V(n7458) V(n7459) V(n7460) V(n7461) V(n7462) V(n7463) V(n7464) V(n7465) V(n7466) V(n7467) V(n7468) V(n7469) V(n7470) V(n7471) V(n7472) V(n7473) V(n7474) V(n7475) V(n7476) V(n7477) V(n7478) V(n7479) V(n7480) V(n7481) V(n7482) V(n7483) V(n7484) V(n7485) V(n7486) V(n7487) V(n7488) V(n7489) V(n7490) V(n7491) V(n7492) V(n7493) V(n7494) V(n7495) V(n7496) V(n7497) V(n7498) V(n7499) V(n7500) V(n7501) V(n7502) V(n7503) V(n7504) V(n7505) V(n7506) V(n7507) V(n7508) V(n7509) V(n7510) V(n7511) V(n7512) V(n7513) V(n7514) V(n1) V(n7516) V(n7517) V(n7518) V(n7519) V(n7520) V(n7521) V(n7522) V(n7523) V(n7524) V(n7525) V(n7526) V(n7527) V(n7528) V(n7529) V(n7530) V(n7531) V(n7532) V(n7533) V(n7534) V(n7535) V(n7536) V(n7537) V(n7538) V(n7539) V(n7540) V(n7541) V(n7542) V(n7543) V(n7544) V(n7545) V(n7546) V(n7547) V(n7548) V(n7549) V(n7550) V(n7551) V(n7552) V(n7553) V(n7554) V(n7555) V(n7556) V(n7557) V(n7558) V(n7559) V(n7560) V(n7561) V(n7562) V(n7563) V(n7564) V(n7565) V(n7566) V(n7567) V(n7568) V(n7569) V(n7570) V(n7571) V(n7572) V(n7573) V(n7574) V(n7575) V(n7576) V(n7577) V(n7578) V(n7579) V(n7580) V(n7581) V(n7582) V(n7583) V(n7584) V(n7585) V(n7586) V(n7587) V(n7588) V(n7589) V(n7590) V(n7591) V(n7592) V(n7593) V(n7594) V(n7595) V(n7596) V(n7597) V(n7598) V(n7599) V(n7600) V(n7601) V(n7602) V(n7603) V(n7604) V(n7605) V(n7606) V(n7607) V(n7608) V(n7609) V(n7610) V(n7611) V(n7612) V(n7613) V(n7614) V(n7615) V(n7616) V(n7617) V(n7618) V(n7619) V(n7620) V(n7621) V(n7622) V(n7623) V(n7624) V(n7625) V(n7626) V(n7627) V(n7628) V(n7629) V(n7630) V(n7631) V(n7632) V(n7633) V(n7634) V(n7635) V(n7636) V(n7637) V(n7638) V(n7639) V(n7640) V(n7641) V(n7642) V(n7643) V(n7644) V(n7645) V(n7646) V(n7647) V(n7648) V(n7649) V(n7650) V(n7651) V(n7652) V(n7653) V(n7654) V(n7655) V(n7656) V(n1) V(n7658) V(n7659) V(n7660) V(n7661) V(n7662) V(n1) V(n7664) V(n7665) V(n1) V(n7667) V(n7668) V(n7669) V(n7670) V(n7671) V(n1) V(n7673) V(n7674) V(n7675) V(n7676) V(n7677) V(n7678) V(n7679) V(n7680) V(n7681) V(n7682) V(n7683) V(n7684) V(n7685) V(n7686) V(n7687) V(n7688) V(n7689) V(n7690) V(n7691) V(n7692) V(n7693) V(n7694) V(n7695) V(n7696) V(n7697) V(n7698) V(n7699) V(n7700) V(n7701) V(n7702) V(n7703) V(n7704) V(n7705) V(n7706) V(n7707) V(n7708) V(n7709) V(n7710) V(n7711) V(n7712) V(n7713) V(n7714) V(n7715) V(n7716) V(n7717) V(n7718) V(n7719) V(n7720) V(n7721) V(n7722) V(n7723) V(n7724) V(n7725) V(n7726) V(n7727) V(n7728) V(n7729) V(n7730) V(n7731) V(n7732) V(n7733) V(n7734) V(n7735) V(n7736) V(n7737) V(n7738) V(n7739) V(n7740) V(n7741) V(n7742) V(n7743) V(n7744) V(n7745) V(n7746) V(n7747) V(n7748) V(n7749) V(n7750) V(n7751) V(n7752) V(n7753) V(n7754) V(n7755) V(n7756) V(n7757) V(n7758) V(n7759) V(n7760) V(n7761) V(n7762) V(n7763) V(n7764) V(n7765) V(n7766) V(n7767) V(n7768) V(n7769) V(n7770) V(n7771) V(n7772) V(n7773) V(n7774) V(n7775) V(n7776) V(n7777) V(n7778) V(n7779) V(n7780) V(n7781) V(n7782) V(n7783) V(n7784) V(n7785) V(n7786) V(n7787) V(n7788) V(n7789) V(n7790) V(n7791) V(n7792) V(n7793) V(n7794) V(n7795) V(n7796) V(n7797) V(n7798) V(n7799) V(n7800) V(n7801) V(n7802) V(n7803) V(n7804) V(n7805) V(n7806) V(n1) V(n7808) V(n7809) V(n7810) V(n7811) V(n7812) V(n7813) V(n7814) V(n7815) V(n7816) V(n7817) V(n7818) V(n7819) V(n7820) V(n7821) V(n7822) V(n7823) V(n7824) V(n7825) V(n1) V(n7827) V(n7828) V(n7829) V(n7830) V(n7831) V(n7832) V(n7833) V(n7834) V(n7835) V(n7836) V(n7837) V(n7838) V(n7839) V(n7840) V(n7841) V(n7842) V(n7843) V(n7844) V(n7845) V(n7846) V(n7847) V(n7848) V(n7849) V(n7850) V(n7851) V(n7852) V(n7853) V(n7854) V(n7855) V(n7856) V(n7857) V(n7858) V(n7859) V(n7860) V(n7861) V(n7862) V(n7863) V(n7864) V(n7865) V(n7866) V(n7867) V(n7868) V(n7869) V(n7870) V(n7871) V(n7872) V(n7873) V(n7874) V(n7875) V(n7876) V(n7877) V(n7878) V(n7879) V(n7880) V(n7881) V(n7882) V(n7883) V(n7884) V(n7885) V(n7886) V(n7887) V(n7888) V(n7889) V(n7890) V(n7891) V(n7892) V(n7893) V(n7894) V(n7895) V(n7896) V(n7897) V(n7898) V(n7899) V(n7900) V(n7901) V(n7902) V(n7903) V(n7904) V(n7905) V(n7906) V(n7907) V(n7908) V(n7909) V(n7910) V(n7911) V(n7912) V(n7913) V(n7914) V(n7915) V(n7916) V(n7917) V(n7918) V(n7919) V(n7920) V(n7921) V(n7922) V(n7923) V(n7924) V(n7925) V(n7926) V(n7927) V(n7928) V(n7929) V(n7930) V(n7931) V(n7932) V(n7933) V(n7934) V(n7935) V(n7936) V(n7937) V(n7938) V(n1) V(n7940) V(n7941) V(n7942) V(n7943) V(n7944) V(n7945) V(n7946) V(n7947) V(n7948) V(n7949) V(n7950) V(n7951) V(n7952) V(n7953) V(n7954) V(n7955) V(n7956) V(n7957) V(n7958) V(n7959) V(n7960) V(n7961) V(n7962) V(n7963) V(n7964) V(n7965) V(n7966) V(n7967) V(n7968) V(n7969) V(n7970) V(n7971) V(n7972) V(n7973) V(n7974) V(n7975) V(n7976) V(n7977) V(n7978) V(n7979) V(n7980) V(n7981) V(n7982) V(n7983) V(n7984) V(n7985) V(n7986) V(n7987) V(n7988) V(n7989) V(n7990) V(n7991) V(n7992) V(n7993) V(n7994) V(n7995) V(n7996) V(n7997) V(n7998) V(n7999) V(n8000) V(n8001) V(n8002) V(n8003) V(n8004) V(n8005) V(n8006) V(n8007) V(n8008) V(n8009) V(n8010) V(n8011) V(n8012) V(n8013) V(n8014) V(n8015) V(n8016) V(n8017) V(n8018) V(n8019) V(n8020) V(n8021) V(n8022) V(n8023) V(n8024) V(n8025) V(n8026) V(n8027) V(n8028) V(n8029) V(n8030) V(n8031) V(n8032) V(n8033) V(n8034) V(n8035) V(n8036) V(n8037) V(n8038) V(n8039) V(n8040) V(n8041) V(n8042) V(n8043) V(n8044) V(n8045) V(n8046) V(n8047) V(n8048) V(n8049) V(n8050) V(n8051) V(n8052) V(n8053) V(n8054) V(n8055) V(n8056) V(n8057) V(n8058) V(n8059) V(n8060) V(n8061) V(n8062) V(n8063) V(n8064) V(n8065) V(n8066) V(n8067) V(n8068) V(n8069) V(n8070) V(n8071) V(n8072) V(n8073) V(n8074) V(n8075) V(n8076) V(n8077) V(n8078) V(n8079) V(n8080) V(n8081) V(n8082) V(n8083) V(n8084) V(n8085) V(n8086) V(n8087) V(n8088) V(n8089) V(n8090) V(n8091) V(n8092) V(n8093) V(n8094) V(n8095) V(n8096) V(n8097) V(n8098) V(n8099) V(n8100) V(n8101) V(n8102) V(n8103) V(n8104) V(n8105) V(n8106) V(n8107) V(n8108) V(n8109) V(n8110) V(n8111) V(n8112) V(n8113) V(n8114) V(n8115) V(n8116) V(n8117) V(n8118) V(n8119) V(n8120) V(n8121) V(n8122) V(n8123) V(n8124) V(n8125) V(n8126) V(n8127) V(n8128) V(n8129) V(n8130) V(n8131) V(n8132) V(n8133) V(n8134) V(n8135) V(n8136) V(n8137) V(n8138) V(n8139) V(n8140) V(n8141) V(n8142) V(n8143) V(n8144) V(n8145) V(n8146) V(n8147) V(n8148) V(n8149) V(n8150) V(n8151) V(n8152) V(n8153) V(n8154) V(n8155) V(n8156) V(n8157) V(n8158) V(n8159) V(n8160) V(n8161) V(n8162) V(n8163) V(n8164) V(n8165) V(n8166) V(n8167) V(n8168) V(n8169) V(n8170) V(n8171) V(n8172) V(n8173) V(n8174) V(n8175) V(n8176) V(n8177) V(n8178) V(n8179) V(n8180) V(n8181) V(n8182) V(n8183) V(n8184) V(n8185) V(n8186) V(n8187) V(n8188) V(n8189) V(n8190) V(n8191) V(n8192) V(n8193) V(n8194) V(n8195) V(n8196) V(n8197) V(n8198) V(n8199) V(n8200) V(n8201) V(n8202) V(n8203) V(n8204) V(n8205) V(n8206) V(n8207) V(n8208) V(n8209) V(n8210) V(n8211) V(n8212) V(n8213) V(n8214) V(n8215) V(n8216) V(n8217) V(n8218) V(n8219) V(n8220) V(n8221) V(n8222) V(n8223) V(n8224) V(n8225) V(n8226) V(n8227) V(n8228) V(n8229) V(n8230) V(n8231) V(n8232) V(n8233) V(n8234) V(n8235) V(n8236) V(n8237) V(n8238) V(n8239) V(n8240) V(n8241) V(n8242) V(n8243) V(n8244) V(n8245) V(n8246) V(n8247) V(n8248) V(n8249) V(n8250) V(n8251) V(n8252) V(n8253) V(n8254) V(n8255) V(n8256) V(n8257) V(n8258) V(n8259) V(n8260) V(n8261) V(n8262) V(n8263) V(n8264) V(n8265) V(n8266) V(n8267) V(n8268) V(n8269) V(n8270) V(n8271) V(n8272) V(n8273) V(n8274) V(n8275) V(n8276) V(n8277) V(n8278) V(n8279) V(n8280) V(n8281) V(n8282) V(n8283) V(n8284) V(n8285) V(n8286) V(n8287) V(n8288) V(n8289) V(n8290) V(n8291) V(n8292) V(n8293) V(n8294) V(n8295) V(n8296) V(n8297) V(n8298) V(n8299) V(n8300) V(n8301) V(n8302) V(n8303) V(n8304) V(n8305) V(n8306) V(n8307) V(n8308) V(n8309) V(n8310) V(n8311) V(n8312) V(n8313) V(n8314) V(n8315) V(n8316) V(n8317) V(n8318) V(n8319) V(n8320) V(n8321) V(n8322) V(n8323) V(n8324) V(n8325) V(n8326) V(n8327) V(n8328) V(n8329) V(n8330) V(n8331) V(n8332) V(n8333) V(n8334) V(n8335) V(n1) V(n8337) V(n8338) V(n8339) V(n8340) V(n8341) V(n8342) V(n8343) V(n8344) V(n8345) V(n8346) V(n8347) V(n8348) V(n8349) V(n8350) V(n8351) V(n8352) V(n8353) V(n8354) V(n8355) V(n8356) V(n8357) V(n8358) V(n8359) V(n8360) V(n8361) V(n8362) V(n8363) V(n8364) V(n8365) V(n8366) V(n8367) V(n8368) V(n8369) V(n8370) V(n8371) V(n8372) V(n8373) V(n8374) V(n8375) V(n8376) V(n8377) V(n8378) V(n8379) V(n8380) V(n8381) V(n8382) V(n8383) V(n8384) V(n8385) V(n8386) V(n8387) V(n8388) V(n8389) V(n8390) V(n8391) V(n8392) V(n8393) V(n8394) V(n8395) V(n8396) V(n8397) V(n8398) V(n8399) V(n8400) V(n8401) V(n8402) V(n8403) V(n8404) V(n8405) V(n8406) V(n8407) V(n8408) V(n8409) V(n8410) V(n8411) V(n8412) V(n8413) V(n8414) V(n8415) V(n8416) V(n8417) V(n8418) V(n8419) V(n8420) V(n8421) V(n8422) V(n8423) V(n8424) V(n8425) V(n8426) V(n8427) V(n8428) V(n8429) V(n8430) V(n8431) V(n8432) V(n8433) V(n8434) V(n8435) V(n8436) V(n8437) V(n8438) V(n8439) V(n8440) V(n8441) V(n8442) V(n8443) V(n8444) V(n8445) V(n8446) V(n8447) V(n8448) V(n8449) V(n8450) V(n8451) V(n8452) V(n8453) V(n8454) V(n8455) V(n8456) V(n8457) V(n8458) V(n8459) V(n8460) V(n8461) V(n8462) V(n8463) V(n8464) V(n8465) V(n8466) V(n8467) V(n8468) V(n8469) V(n8470) V(n8471) V(n8472) V(n8473) V(n8474) V(n8475) V(n8476) V(n8477) V(n8478) V(n8479) V(n8480) V(n8481) V(n8482) V(n8483) V(n8484) V(n8485) V(n8486) V(n8487) V(n8488) V(n8489) V(n8490) V(n8491) V(n8492) V(n8493) V(n8494) V(n8495) V(n8496) V(n8497) V(n8498) V(n8499) V(n1) V(n8501) V(n8502) V(n8503) V(n8504) V(n8505) V(n8506) V(n8507) V(n8508) V(n8509) V(n8510) V(n8511) V(n8512) V(n8513) V(n8514) V(n8515) V(n8516) V(n8517) V(n8518) V(n8519) V(n8520) V(n8521) V(n8522) V(n8523) V(n8524) V(n8525) V(n8526) V(n8527) V(n8528) V(n8529) V(n8530) V(n8531) V(n8532) V(n8533) V(n8534) V(n8535) V(n8536) V(n8537) V(n8538) V(n8539) V(n8540) V(n8541) V(n8542) V(n8543) V(n8544) V(n8545) V(n8546) V(n8547) V(n8548) V(n8549) V(n8550) V(n8551) V(n8552) V(n8553) V(n8554) V(n1) V(n8556) V(n8557) V(n8558) V(n8559) V(n8560) V(n8561) V(n8562) V(n8563) V(n8564) V(n8565) V(n8566) V(n8567) V(n8568) V(n8569) V(n8570) V(n8571) V(n8572) V(n8573) V(n8574) V(n8575) V(n8576) V(n8577) V(n8578) V(n8579) V(n8580) V(n8581) V(n8582) V(n8583) V(n8584) V(n8585) V(n8586) V(n8587) V(n8588) V(n8589) V(n8590) V(n8591) V(n8592) V(n8593) V(n8594) V(n8595) V(n8596) V(n8597) V(n8598) V(n8599) V(n8600) V(n8601) V(n8602) V(n1) V(n8604) V(n8605) V(n8606) V(n8607) V(n8608) V(n8609) V(n8610) V(n8611) V(n8612) V(n8613) V(n8614) V(n8615) V(n8616) V(n8617) V(n8618) V(n8619) V(n8620) V(n8621) V(n8622) V(n8623) V(n8624) V(n8625) V(n8626) V(n8627) V(n8628) V(n8629) V(n8630) V(n8631) V(n8632) V(n8633) V(n8634) V(n8635) V(n8636) V(n8637) V(n8638) V(n8639) V(n8640) V(n8641) V(n8642) V(n8643) V(n8644) V(n8645) V(n8646) V(n8647) V(n8648) V(n8649) V(n8650) V(n8651) V(n8652) V(n8653) V(n8654) V(n8655) V(n8656) V(n8657) V(n8658) V(n8659) V(n8660) V(n8661) V(n8662) V(n8663) V(n8664) V(n8665) V(n8666) V(n8667) V(n8668) V(n8669) V(n8670) V(n8671) V(n8672) V(n8673) V(n8674) V(n8675) V(n8676) V(n8677) V(n8678) V(n8679) V(n1) V(n8681) V(n8682) V(n8683) V(n8684) V(n8685) V(n8686) V(n8687) V(n8688) V(n8689) V(n8690) V(n8691) V(n8692) V(n8693) V(n8694) V(n8695) V(n8696) V(n8697) V(n8698) V(n8699) V(n8700) V(n8701) V(n8702) V(n8703) V(n8704) V(n8705) V(n8706) V(n8707) V(n8708) V(n8709) V(n8710) V(n8711) V(n8712) V(n8713) V(n8714) V(n8715) V(n8716) V(n8717) V(n8718) V(n8719) V(n8720) V(n8721) V(n8722) V(n8723) V(n8724) V(n8725) V(n8726) V(n8727) V(n8728) V(n8729) V(n8730) V(n8731) V(n8732) V(n8733) V(n8734) V(n8735) V(n8736) V(n8737) V(n8738) V(n8739) V(n8740) V(n8741) V(n8742) V(n8743) V(n8744) V(n8745) V(n8746) V(n8747) V(n8748) V(n8749) V(n8750) V(n8751) V(n8752) V(n8753) V(n8754) V(n8755) V(n8756) V(n8757) V(n8758) V(n8759) V(n8760) V(n8761) V(n8762) V(n8763) V(n8764) V(n8765) V(n8766) V(n8767) V(n8768) V(n8769) V(n8770) V(n8771) V(n8772) V(n8773) V(n8774) V(n8775) V(n8776) V(n8777) V(n8778) V(n8779) V(n8780) V(n8781) V(n8782) V(n8783) V(n8784) V(n8785) V(n8786) V(n8787) V(n8788) V(n8789) V(n8790) V(n8791) V(n8792) V(n8793) V(n8794) V(n8795) V(n8796) V(n8797) V(n8798) V(n8799) V(n8800) V(n8801) V(n8802) V(n8803) V(n8804) V(n8805) V(n8806) V(n8807) V(n8808) V(n8809) V(n8810) V(n8811) V(n8812) V(n8813) V(n8814) V(n8815) V(n8816) V(n8817) V(n8818) V(n8819) V(n8820) V(n8821) V(n8822) V(n8823) V(n8824) V(n8825) V(n8826) V(n8827) V(n8828) V(n8829) V(n8830) V(n8831) V(n8832) V(n8833) V(n8834) V(n8835) V(n8836) V(n8837) V(n8838) V(n8839) V(n8840) V(n8841) V(n8842) V(n1) V(n8844) V(n8845) V(n8846) V(n8847) V(n8848) V(n8849) V(n8850) V(n8851) V(n8852) V(n8853) V(n8854) V(n8855) V(n8856) V(n8857) V(n8858) V(n8859) V(n8860) V(n8861) V(n8862) V(n8863) V(n8864) V(n8865) V(n8866) V(n8867) V(n8868) V(n8869) V(n8870) V(n8871) V(n8872) V(n8873) V(n8874) V(n8875) V(n8876) V(n8877) V(n8878) V(n8879) V(n8880) V(n8881) V(n8882) V(n8883) V(n8884) V(n8885) V(n8886) V(n8887) V(n8888) V(n8889) V(n8890) V(n8891) V(n8892) V(n8893) V(n8894) V(n8895) V(n8896) V(n8897) V(n8898) V(n8899) V(n8900) V(n8901) V(n8902) V(n8903) V(n8904) V(n8905) V(n8906) V(n8907) V(n8908) V(n8909) V(n8910) V(n8911) V(n8912) V(n8913) V(n8914) V(n8915) V(n8916) V(n8917) V(n8918) V(n8919) V(n8920) V(n8921) V(n8922) V(n8923) V(n8924) V(n8925) V(n1) V(n8927) V(n8928) V(n8929) V(n8930) V(n8931) V(n8932) V(n8933) V(n8934) V(n8935) V(n8936) V(n8937) V(n8938) V(n8939) V(n8940) V(n8941) V(n8942) V(n8943) V(n8944) V(n8945) V(n8946) V(n8947) V(n8948) V(n8949) V(n8950) V(n8951) V(n8952) V(n8953) V(n8954) V(n8955) V(n8956) V(n8957) V(n8958) V(n8959) V(n8960) V(n8961) V(n8962) V(n8963) V(n8964) V(n8965) V(n8966) V(n8967) V(n8968) V(n8969) V(n8970) V(n8971) V(n8972) V(n8973) V(n8974) V(n8975) V(n8976) V(n8977) V(n8978) V(n8979) V(n8980) V(n8981) V(n8982) V(n8983) V(n8984) V(n8985) V(n8986) V(n8987) V(n8988) V(n8989) V(n8990) V(n8991) V(n8992) V(n8993) V(n8994) V(n8995) V(n8996) V(n8997) V(n8998) V(n8999) V(n9000) V(n9001) V(n9002) V(n9003) V(n9004) V(n9005) V(n9006) V(n9007) V(n9008) V(n9009) V(n9010) V(n9011) V(n9012) V(n9013) V(n9014) V(n9015) V(n9016) V(n9017) V(n9018) V(n9019) V(n9020) V(n9021) V(n9022) V(n9023) V(n9024) V(n9025) V(n9026) V(n9027) V(n9028) V(n9029) V(n9030) V(n9031) V(n9032) V(n9033) V(n9034) V(n9035) V(n9036) V(n9037) V(n9038) V(n9039) V(n9040) V(n9041) V(n9042) V(n9043) V(n9044) V(n9045) V(n9046) V(n9047) V(n9048) V(n9049) V(n9050) V(n9051) V(n9052) V(n9053) V(n9054) V(n9055) V(n9056) V(n9057) V(n9058) V(n9059) V(n9060) V(n9061) V(n9062) V(n9063) V(n9064) V(n9065) V(n9066) V(n9067) V(n9068) V(n9069) V(n9070) V(n9071) V(n9072) V(n9073) V(n9074) V(n9075) V(n9076) V(n9077) V(n9078) V(n9079) V(n9080) V(n9081) V(n1) V(n9083) V(n9084) V(n9085) V(n9086) V(n9087) V(n9088) V(n9089) V(n9090) V(n9091) V(n9092) V(n9093) V(n9094) V(n9095) V(n9096) V(n9097) V(n9098) V(n9099) V(n9100) V(n9101) V(n9102) V(n9103) V(n9104) V(n9105) V(n9106) V(n9107) V(n9108) V(n9109) V(n9110) V(n9111) V(n9112) V(n9113) V(n9114) V(n9115) V(n9116) V(n9117) V(n9118) V(n9119) V(n9120) V(n9121) V(n9122) V(n9123) V(n9124) V(n9125) V(n9126) V(n9127) V(n9128) V(n9129) V(n9130) V(n9131) V(n9132) V(n9133) V(n9134) V(n9135) V(n9136) V(n9137) V(n1) V(n9139) V(n9140) V(n9141) V(n9142) V(n9143) V(n9144) V(n9145) V(n9146) V(n9147) V(n9148) V(n9149) V(n9150) V(n9151) V(n9152) V(n9153) V(n9154) V(n9155) V(n9156) V(n9157) V(n9158) V(n9159) V(n9160) V(n9161) V(n9162) V(n9163) V(n9164) V(n9165) V(n9166) V(n9167) V(n9168) V(n9169) V(n9170) V(n9171) V(n9172) V(n9173) V(n9174) V(n9175) V(n9176) V(n9177) V(n9178) V(n9179) V(n9180) V(n9181) V(n9182) V(n9183) V(n9184) V(n9185) V(n9186) V(n9187) V(n9188) V(n9189) V(n9190) V(n9191) V(n9192) V(n9193) V(n9194) V(n9195) V(n9196) V(n9197) V(n9198) V(n9199) V(n9200) V(n9201) V(n9202) V(n9203) V(n9204) V(n9205) V(n9206) V(n9207) V(n9208) V(n9209) V(n9210) V(n9211) V(n9212) V(n9213) V(n9214) V(n9215) V(n9216) V(n9217) V(n9218) V(n9219) V(n9220) V(n9221) V(n9222) V(n9223) V(n9224) V(n9225) V(n9226) V(n9227) V(n9228) V(n9229) V(n9230) V(n9231) V(n9232) V(n9233) V(n9234) V(n9235) V(n9236) V(n9237) V(n9238) V(n9239) V(n9240) V(n9241) V(n9242) V(n9243) V(n9244) V(n9245) V(n9246) V(n9247) V(n9248) V(n9249) V(n9250) V(n9251) V(n9252) V(n9253) V(n9254) V(n9255) V(n9256) V(n9257) V(n9258) V(n9259) V(n9260) V(n9261) V(n9262) V(n9263) V(n9264) V(n9265) V(n9266) V(n9267) V(n9268) V(n9269) V(n9270) V(n9271) V(n9272) V(n9273) V(n9274) V(n9275) V(n9276) V(n9277) V(n9278) V(n9279) V(n9280) V(n9281) V(n9282) V(n9283) V(n9284) V(n9285) V(n9286) V(n9287) V(n9288) V(n9289) V(n9290) V(n9291) V(n9292) V(n9293) V(n9294) V(n9295) V(n9296) V(n9297) V(n9298) V(n9299) V(n9300) V(n9301) V(n9302) V(n9303) V(n9304) V(n9305) V(n9306) V(n9307) V(n9308) V(n9309) V(n9310) V(n9311) V(n9312) V(n9313) V(n9314) V(n9315) V(n9316) V(n9317) V(n9318) V(n9319) V(n9320) V(n9321) V(n9322) V(n9323) V(n9324) V(n1) V(n9326) V(n9327) V(n9328) V(n9329) V(n9330) V(n9331) V(n9332) V(n9333) V(n9334) V(n9335) V(n9336) V(n9337) V(n9338) V(n9339) V(n9340) V(n9341) V(n9342) V(n9343) V(n9344) V(n9345) V(n9346) V(n9347) V(n9348) V(n9349) V(n9350) V(n9351) V(n9352) V(n9353) V(n9354) V(n9355) V(n9356) V(n9357) V(n9358) V(n9359) V(n9360) V(n9361) V(n9362) V(n9363) V(n9364) V(n9365) V(n9366) V(n9367) V(n9368) V(n9369) V(n9370) V(n9371) V(n9372) V(n9373) V(n9374) V(n9375) V(n9376) V(n9377) V(n9378) V(n9379) V(n9380) V(n9381) V(n9382) V(n9383) V(n9384) V(n9385) V(n9386) V(n9387) V(n9388) V(n9389) V(n9390) V(n9391) V(n9392) V(n9393) V(n9394) V(n9395) V(n9396) V(n9397) V(n9398) V(n9399) V(n9400) V(n9401) V(n9402) V(n9403) V(n9404) V(n9405) V(n9406) V(n9407) V(n9408) V(n9409) V(n9410) V(n9411) V(n9412) V(n9413) V(n9414) V(n9415) V(n9416) V(n9417) V(n9418) V(n9419) V(n9420) V(n9421) V(n9422) V(n9423) V(n9424) V(n9425) V(n9426) V(n9427) V(n9428) V(n9429) V(n9430) V(n9431) V(n9432) V(n9433) V(n9434) V(n9435) V(n9436) V(n9437) V(n9438) V(n9439) V(n9440) V(n9441) V(n9442) V(n9443) V(n9444) V(n9445) V(n9446) V(n9447) V(n9448) V(n9449) V(n9450) V(n9451) V(n9452) V(n9453) V(n9454) V(n9455) V(n9456) V(n9457) V(n9458) V(n9459) V(n9460) V(n9461) V(n9462) V(n9463) V(n9464) V(n9465) V(n9466) V(n9467) V(n9468) V(n9469) V(n9470) V(n9471) V(n9472) V(n9473) V(n9474) V(n9475) V(n9476) V(n9477) V(n9478) V(n9479) V(n9480) V(n9481) V(n9482) V(n9483) V(n9484) V(n9485) V(n9486) V(n9487) V(n9488) V(n9489) V(n9490) V(n9491) V(n9492) V(n9493) V(n9494) V(n9495) V(n9496) V(n9497) V(n9498) V(n9499) V(n9500) V(n9501) V(n9502) V(n9503) V(n9504) V(n9505) V(n9506) V(n9507) V(n9508) V(n9509) V(n9510) V(n1) V(n9512) V(n9513) V(n9514) V(n9515) V(n9516) V(n9517) V(n9518) V(n9519) V(n9520) V(n9521) V(n9522) V(n9523) V(n9524) V(n9525) V(n9526) V(n9527) V(n9528) V(n9529) V(n9530) V(n9531) V(n9532) V(n9533) V(n9534) V(n9535) V(n9536) V(n9537) V(n9538) V(n9539) V(n9540) V(n9541) V(n9542) V(n9543) V(n9544) V(n9545) V(n9546) V(n9547) V(n9548) V(n9549) V(n9550) V(n9551) V(n9552) V(n9553) V(n9554) V(n9555) V(n9556) V(n9557) V(n9558) V(n9559) V(n9560) V(n9561) V(n9562) V(n9563) V(n9564) V(n9565) V(n9566) V(n9567) V(n9568) V(n9569) V(n9570) V(n9571) V(n9572) V(n9573) V(n9574) V(n9575) V(n9576) V(n9577) V(n9578) V(n9579) V(n9580) V(n9581) V(n9582) V(n9583) V(n9584) V(n9585) V(n9586) V(n9587) V(n9588) V(n9589) V(n9590) V(n9591) V(n9592) V(n9593) V(n9594) V(n9595) V(n9596) V(n9597) V(n9598) V(n9599) V(n9600) V(n9601) V(n9602) V(n9603) V(n9604) V(n9605) V(n9606) V(n9607) V(n9608) V(n9609) V(n9610) V(n9611) V(n9612) V(n9613) V(n9614) V(n9615) V(n9616) V(n9617) V(n9618) V(n9619) V(n9620) V(n9621) V(n9622) V(n9623) V(n9624) V(n9625) V(n9626) V(n9627) V(n9628) V(n9629) V(n9630) V(n9631) V(n9632) V(n9633) V(n9634) V(n9635) V(n9636) V(n9637) V(n9638) V(n9639) V(n9640) V(n9641) V(n9642) V(n9643) V(n9644) V(n9645) V(n9646) V(n9647) V(n9648) V(n9649) V(n9650) V(n9651) V(n9652) V(n9653) V(n9654) V(n9655) V(n9656) V(n9657) V(n9658) V(n9659) V(n9660) V(n9661) V(n9662) V(n9663) V(n9664) V(n9665) V(n9666) V(n9667) V(n9668) V(n9669) V(n9670) V(n9671) V(n9672) V(n9673) V(n9674) V(n9675) V(n9676) V(n9677) V(n9678) V(n9679) V(n9680) V(n9681) V(n9682) V(n9683) V(n9684) V(n9685) V(n9686) V(n9687) V(n9688) V(n9689) V(n9690) V(n9691) V(n9692) V(n9693) V(n9694) I(R91t61) I(R114t47) I(R148t4) I(R148t54) I(R154t89) I(R161t54) I(R193t184) I(R208t124) I(R226t168) I(R236t158) I(R236t179) I(R254t243) I(R266t28) I(R271t119) I(R275t48) I(R289t46) I(R292t173) I(R297t255) I(R303t13) I(R306t20) I(R308t290) I(R320t144) I(R321t186) I(R321t319) I(R346t114) I(R360t185) I(R365t334) I(R367t51) I(R370t279) I(R373t199) I(R376t39) I(R377t270) I(R378t272) I(R380t240) I(R385t194) I(R389t347) I(R393t57) I(R409t274) I(R411t87) I(R418t390) I(R423t65) I(R428t188) I(R434t430) I(R435t147) I(R443t49) I(R445t133) I(R445t35) I(R454t133) I(R457t58) I(R460t64) I(R460t245) I(R465t129) I(R467t312) I(R473t406) I(R475t362) I(R477t281) I(R480t82) I(R485t332) I(R489t10) I(R492t314) I(R495t442) I(R503t396) I(R507t468) I(R521t466) I(R526t491) I(R528t70) I(R529t242) I(R531t101) I(R533t239) I(R534t185) I(R539t505) I(R543t418) I(R549t438) I(R550t373) I(R551t480) I(R558t383) I(R560t429) I(R564t6) I(R565t425) I(R566t520) I(R566t411) I(R580t271) I(R582t331) I(R582t75) I(R584t77) I(R584t272) I(R587t100) I(R589t31) I(R589t580) I(R592t318) I(R592t55) I(R595t393) I(R595t57) I(R596t587) I(R596t100) I(R599t458) I(R600t15) I(R601t496) I(R601t159) I(R606t382) I(R609t238) I(R610t141) I(R613t55) I(R619t581) I(R625t27) I(R627t292) I(R637t264) I(R641t412) I(R647t197) I(R649t17) I(R652t33) I(R656t188) I(R656t428) I(R658t454) I(R660t241) I(R662t284) I(R665t325) I(R666t311) I(R667t559) I(R671t358) I(R673t13) I(R677t213) I(R679t127) I(R680t528) I(R681t5) I(R683t551) I(R685t361) I(R685t488) I(R690t542) I(R693t659) I(R694t525) I(R697t545) I(R699t95) I(R707t623) I(R714t675) I(R714t41) I(R716t145) I(R718t172) I(R721t650) I(R721t203) I(R724t595) I(R724t393) I(R726t130) I(R729t359) I(R729t252) I(R730t271) I(R731t714) I(R731t412) I(R736t162) I(R738t183) I(R738t169) I(R740t633) I(R743t198) I(R745t686) I(R745t548) I(R747t576) I(R749t572) I(R751t175) I(R752t328) I(R754t641) I(R755t36) I(R758t52) I(R758t673) I(R758t13) I(R759t535) I(R762t436) I(R763t659) I(R764t671) I(R764t358) I(R767t45) I(R767t457) I(R772t194) I(R772t385) I(R773t53) I(R775t509) I(R779t444) I(R781t402) I(R782t512) I(R783t244) I(R785t541) I(R786t172) I(R790t598) I(R792t504) I(R792t713) I(R797t518) I(R798t500) I(R798t661) I(R799t6) I(R801t22) I(R803t26) I(R804t228) I(R805t495) I(R807t753) I(R813t688) I(R816t763) I(R816t659) I(R817t88) I(R817t14) I(R819t26) I(R821t609) I(R822t17) I(R823t460) I(R823t245) I(R829t332) I(R829t485) I(R833t724) I(R835t135) I(R838t372) I(R839t118) I(R839t266) I(R840t714) I(R840t731) I(R842t206) I(R843t209) I(R844t781) I(R844t402) I(R845t807) I(R845t753) I(R849t138) I(R850t666) I(R852t580) I(R852t589) I(R853t825) I(R857t583) I(R858t26) I(R858t803) I(R859t785) I(R860t386) I(R860t66) I(R861t435) I(R861t537) I(R862t411) I(R863t164) I(R863t487) I(R864t284) I(R868t441) I(R868t129) I(R868t465) I(R869t366) I(R869t247) I(R871t69) I(R872t295) I(R875t200) I(R878t117) I(R878t736) I(R879t390) I(R883t370) I(R883t392) I(R884t184) I(R884t193) I(R887t400) I(R890t155) I(R892t274) I(R892t409) I(R894t877) I(R897t42) I(R900t757) I(R901t750) I(R904t116) I(R904t292) I(R906t569) I(R909t441) I(R909t868) I(R910t485) I(R911t880) I(R912t695) I(R913t648) I(R915t599) I(R917t789) I(R922t392) I(R929t138) I(R931t135) I(R931t835) I(R934t49) I(R937t562) I(R938t596) I(R939t900) I(R941t531) I(R942t299) I(R942t221) I(R947t521) I(R947t466) I(R948t437) I(R950t559) I(R954t946) I(R955t809) I(R955t462) I(R957t351) I(R960t855) I(R961t440) I(R961t732) I(R967t707) I(R967t623) I(R968t608) I(R968t444) I(R969t737) I(R969t771) I(R970t4) I(R971t953) I(R972t139) I(R972t820) I(R973t324) I(R974t576) I(R975t889) I(R975t56) I(R976t76) I(R977t575) I(R977t393) I(R977t709) I(R979t860) I(R981t586) I(R984t248) I(R985t251) I(R987t399) I(R988t472) I(R990t943) I(R993t980) I(R995t461) I(R998t76) I(R998t456) I(R999t688) I(R999t470) I(R999t813) I(R1005t388) I(R1005t319) I(R1006t972) I(R1006t820) I(R1007t630) I(R1011t395) I(R1015t11) I(R1016t389) I(R1016t582) I(R1017t602) I(R1018t992) I(R1019t629) I(R1019t72) I(R1020t638) I(R1022t206) I(R1023t965) I(R1026t226) I(R1029t803) I(R1036t1024) I(R1039t674) I(R1040t490) I(R1042t177) I(R1044t403) I(R1045t21) I(R1046t408) I(R1048t746) I(R1048t168) I(R1050t282) I(R1051t501) I(R1060t244) I(R1060t783) I(R1062t986) I(R1066t333) I(R1067t396) I(R1067t503) I(R1070t837) I(R1070t537) I(R1072t16) I(R1074t980) I(R1074t747) I(R1075t333) I(R1075t1066) I(R1077t547) I(R1079t696) I(R1081t542) I(R1085t700) I(R1086t1024) I(R1089t270) I(R1090t488) I(R1091t698) I(R1091t497) I(R1094t698) I(R1095t605) I(R1097t78) I(R1097t1021) I(R1098t391) I(R1099t29) I(R1101t238) I(R1102t895) I(R1105t379) I(R1107t1058) I(R1119t614) I(R1123t925) I(R1128t390) I(R1128t879) I(R1129t644) I(R1130t164) I(R1134t116) I(R1136t399) I(R1136t987) I(R1137t587) I(R1137t596) I(R1140t678) I(R1143t538) I(R1144t136) I(R1149t845) I(R1149t807) I(R1150t1115) I(R1153t234) I(R1153t170) I(R1154t1037) I(R1155t1064) I(R1158t12) I(R1160t332) I(R1161t692) I(R1161t706) I(R1163t770) I(R1164t290) I(R1165t184) I(R1165t193) I(R1166t334) I(R1168t1112) I(R1169t499) I(R1170t269) I(R1171t884) I(R1172t335) I(R1173t921) I(R1174t1124) I(R1175t417) I(R1176t881) I(R1178t438) I(R1178t549) I(R1180t117) I(R1181t1020) I(R1181t638) I(R1185t493) I(R1186t530) I(R1188t1187) I(R1191t820) I(R1192t1021) I(R1192t1097) I(R1194t309) I(R1195t1084) I(R1197t1190) I(R1199t107) I(R1200t281) I(R1202t541) I(R1204t1122) I(R1208t614) I(R1208t1119) I(R1209t338) I(R1210t791) I(R1212t704) I(R1212t363) I(R1213t21) I(R1213t1045) I(R1214t98) I(R1215t1039) I(R1218t1056) I(R1218t746) I(R1220t559) I(R1220t667) I(R1222t989) I(R1223t478) I(R1223t719) I(R1224t433) I(R1224t806) I(R1225t953) I(R1225t971) I(R1226t705) I(R1226t149) I(R1227t1145) I(R1230t939) I(R1231t857) I(R1236t160) I(R1238t290) I(R1239t580) I(R1240t1034) I(R1241t511) I(R1241t557) I(R1244t634) I(R1248t718) I(R1251t335) I(R1253t804) I(R1253t199) I(R1253t373) I(R1254t599) I(R1254t915) I(R1257t574) I(R1258t124) I(R1260t1249) I(R1261t225) I(R1264t514) I(R1265t522) I(R1267t1242) I(R1267t76) I(R1270t268) I(R1272t1215) I(R1272t674) I(R1272t1039) I(R1273t327) I(R1275t376) I(R1275t39) I(R1277t781) I(R1277t844) I(R1278t792) I(R1278t1264) I(R1278t713) I(R1279t614) I(R1279t791) I(R1281t738) I(R1282t793) I(R1283t916) I(R1286t90) I(R1287t892) I(R1287t409) I(R1288t345) I(R1288t83) I(R1291t104) I(R1293t472) I(R1294t855) I(R1294t1221) I(R1295t786) I(R1295t1031) I(R1296t330) I(R1298t788) I(R1299t378) I(R1300t1210) I(R1301t352) I(R1306t1004) I(R1308t731) I(R1311t730) I(R1312t220) I(R1313t236) I(R1313t158) I(R1314t959) I(R1316t162) I(R1316t736) I(R1316t878) I(R1317t892) I(R1320t178) I(R1324t800) I(R1326t665) I(R1326t482) I(R1326t993) I(R1328t735) I(R1329t1058) I(R1329t1107) I(R1330t1300) I(R1330t1279) I(R1330t791) I(R1330t1210) I(R1331t1092) I(R1331t136) I(R1331t1144) I(R1334t755) I(R1335t988) I(R1337t1277) I(R1338t23) I(R1338t471) I(R1340t675) I(R1340t1164) I(R1344t740) I(R1346t784) I(R1347t1319) I(R1348t839) I(R1348t266) I(R1349t258) I(R1350t872) I(R1350t951) I(R1352t454) I(R1352t133) I(R1353t60) I(R1353t920) I(R1354t1000) I(R1355t113) I(R1355t585) I(R1356t690) I(R1356t259) I(R1360t423) I(R1365t392) I(R1366t741) I(R1367t1237) I(R1370t1035) I(R1372t695) I(R1372t71) I(R1374t68) I(R1374t1311) I(R1374t271) I(R1374t119) I(R1378t1052) I(R1380t71) I(R1382t619) I(R1384t654) I(R1386t730) I(R1387t22) I(R1388t1178) I(R1388t1145) I(R1389t1104) I(R1390t494) I(R1392t976) I(R1393t547) I(R1393t1077) I(R1395t1298) I(R1396t796) I(R1396t636) I(R1402t224) I(R1405t275) I(R1405t59) I(R1406t1206) I(R1409t1088) I(R1410t253) I(R1412t960) I(R1413t48) I(R1413t600) I(R1413t15) I(R1414t696) I(R1415t230) I(R1418t545) I(R1418t697) I(R1418t633) I(R1420t1244) I(R1420t634) I(R1421t1415) I(R1424t584) I(R1424t77) I(R1426t866) I(R1429t463) I(R1430t938) I(R1431t357) I(R1432t1064) I(R1433t1265) I(R1433t1030) I(R1434t790) I(R1434t1113) I(R1438t1142) I(R1439t402) I(R1439t844) I(R1439t1277) I(R1439t1337) I(R1441t1427) I(R1442t933) I(R1443t1409) I(R1443t1210) I(R1443t791) I(R1444t653) I(R1445t725) I(R1446t763) I(R1446t693) I(R1447t795) I(R1448t430) I(R1448t434) I(R1449t264) I(R1449t637) I(R1451t83) I(R1451t241) I(R1451t5) I(R1452t196) I(R1453t935) I(R1453t340) I(R1454t293) I(R1457t429) I(R1457t800) I(R1457t1324) I(R1458t1437) I(R1460t208) I(R1461t1278) I(R1461t713) I(R1464t376) I(R1464t701) I(R1464t39) I(R1465t486) I(R1466t102) I(R1467t1002) I(R1467t547) I(R1467t1415) I(R1467t1421) I(R1468t1116) I(R1469t1128) I(R1470t169) I(R1471t1175) I(R1471t417) I(R1475t73) I(R1476t352) I(R1478t420) I(R1480t1360) I(R1481t1033) I(R1481t207) I(R1482t56) I(R1482t400) I(R1483t461) I(R1484t1383) I(R1485t280) I(R1486t1391) I(R1488t1159) I(R1489t1430) I(R1494t465) I(R1494t297) I(R1497t517) I(R1497t261) I(R1499t642) I(R1501t803) I(R1501t1029) I(R1504t197) I(R1504t647) I(R1506t124) I(R1508t516) I(R1509t777) I(R1509t1417) I(R1509t211) I(R1510t572) I(R1515t1250) I(R1516t316) I(R1518t855) I(R1518t960) I(R1518t1465) I(R1519t1416) I(R1519t877) I(R1519t631) I(R1525t716) I(R1525t1194) I(R1525t145) I(R1527t1107) I(R1528t145) I(R1529t959) I(R1529t1314) I(R1530t787) I(R1530t1069) I(R1533t1023) I(R1533t965) I(R1534t561) I(R1535t261) I(R1536t802) I(R1541t470) I(R1542t1495) I(R1543t1348) I(R1544t53) I(R1545t466) I(R1545t947) I(R1546t430) I(R1546t147) I(R1549t1536) I(R1549t720) I(R1549t802) I(R1550t941) I(R1550t101) I(R1551t367) I(R1552t1201) I(R1552t398) I(R1553t286) I(R1556t214) I(R1557t435) I(R1557t919) I(R1557t861) I(R1558t265) I(R1560t245) I(R1562t810) I(R1563t1493) I(R1563t728) I(R1564t180) I(R1565t753) I(R1565t1361) I(R1566t1123) I(R1567t241) I(R1567t660) I(R1567t1451) I(R1567t1056) I(R1568t982) I(R1569t837) I(R1572t1388) I(R1573t369) I(R1573t190) I(R1574t835) I(R1574t931) I(R1576t695) I(R1576t912) I(R1578t312) I(R1578t166) I(R1579t766) I(R1580t232) I(R1583t1400) I(R1584t74) I(R1586t1584) I(R1586t832) I(R1587t742) I(R1590t586) I(R1591t1392) I(R1592t972) I(R1592t820) I(R1592t1191) I(R1592t681) I(R1593t1490) I(R1594t469) I(R1595t280) I(R1595t1485) I(R1595t698) I(R1597t69) I(R1598t207) I(R1601t873) I(R1601t824) I(R1603t234) I(R1605t334) I(R1606t1244) I(R1609t1531) I(R1610t1591) I(R1612t573) I(R1615t1472) I(R1616t1360) I(R1622t1607) I(R1623t1187) I(R1623t1188) I(R1626t1419) I(R1627t1240) I(R1628t1094) I(R1629t167) I(R1629t361) I(R1630t629) I(R1631t98) I(R1631t1214) I(R1631t302) I(R1634t865) I(R1634t537) I(R1634t861) I(R1635t644) I(R1635t1617) I(R1635t439) I(R1636t340) I(R1636t1453) I(R1636t935) I(R1637t1200) I(R1639t483) I(R1640t1191) I(R1640t681) I(R1640t1592) I(R1642t328) I(R1643t126) I(R1643t1061) I(R1644t317) I(R1645t678) I(R1646t986) I(R1646t1062) I(R1648t1110) I(R1648t1096) I(R1649t788) I(R1650t1) I(R1651t440) I(R1655t273) I(R1658t1239) I(R1658t927) I(R1661t1597) I(R1662t353) I(R1666t1019) I(R1667t717) I(R1667t1106) I(R1669t1618) I(R1673t1627) I(R1673t114) I(R1675t655) I(R1676t1657) I(R1677t1211) I(R1677t317) I(R1677t1548) I(R1680t1604) I(R1680t362) I(R1681t1289) I(R1682t1147) I(R1682t484) I(R1683t509) I(R1683t769) I(R1684t1558) I(R1685t1575) I(R1687t866) I(R1688t40) I(R1689t77) I(R1691t373) I(R1691t322) I(R1694t522) I(R1694t1265) I(R1694t1433) I(R1694t57) I(R1695t283) I(R1697t1220) I(R1698t1315) I(R1699t41) I(R1702t499) I(R1702t1169) I(R1703t1183) I(R1706t1290) I(R1707t587) I(R1708t1626) I(R1709t85) I(R1709t1456) I(R1710t326) I(R1710t486) I(R1713t1401) I(R1714t1437) I(R1717t487) I(R1718t1332) I(R1721t1679) I(R1722t1503) I(R1724t466) I(R1724t521) I(R1724t947) I(R1725t737) I(R1725t1700) I(R1725t404) I(R1727t106) I(R1728t692) I(R1728t1161) I(R1730t794) I(R1731t966) I(R1732t985) I(R1733t276) I(R1733t1054) I(R1734t310) I(R1735t543) I(R1736t994) I(R1738t1108) I(R1739t1545) I(R1739t339) I(R1740t105) I(R1742t1224) I(R1744t79) I(R1746t1502) I(R1748t39) I(R1748t1454) I(R1751t249) I(R1753t505) I(R1754t1522) I(R1756t1027) I(R1758t1603) I(R1758t1153) I(R1758t1414) I(R1758t696) I(R1759t1172) I(R1760t1146) I(R1760t1502) I(R1760t1746) I(R1762t518) I(R1762t797) I(R1762t227) I(R1766t1638) I(R1766t1127) I(R1767t510) I(R1767t123) I(R1768t275) I(R1768t48) I(R1768t1413) I(R1768t600) I(R1769t848) I(R1770t1471) I(R1771t1194) I(R1771t1525) I(R1771t145) I(R1771t309) I(R1772t90) I(R1772t1286) I(R1772t162) I(R1773t1438) I(R1773t1237) I(R1773t1142) I(R1774t1637) I(R1775t201) I(R1777t176) I(R1780t215) I(R1784t794) I(R1785t1005) I(R1790t1690) I(R1791t779) I(R1791t1083) I(R1791t1343) I(R1792t779) I(R1792t1343) I(R1792t1791) I(R1793t126) I(R1793t1643) I(R1795t1173) I(R1796t30) I(R1797t1416) I(R1797t1519) I(R1799t1615) I(R1800t1335) I(R1802t203) I(R1803t1065) I(R1805t653) I(R1806t1551) I(R1807t432) I(R1808t765) I(R1812t1645) I(R1814t1713) I(R1817t918) I(R1817t1535) I(R1820t1141) I(R1821t1795) I(R1823t120) I(R1825t362) I(R1828t1234) I(R1828t1617) I(R1829t500) I(R1829t798) I(R1829t1583) I(R1832t313) I(R1833t512) I(R1833t782) I(R1834t455) I(R1836t964) I(R1836t998) I(R1837t955) I(R1837t809) I(R1839t1084) I(R1840t1700) I(R1844t222) I(R1845t1496) I(R1845t1066) I(R1847t1628) I(R1848t768) I(R1850t1478) I(R1850t246) I(R1850t420) I(R1851t910) I(R1852t18) I(R1852t1641) I(R1853t876) I(R1856t1647) I(R1858t125) I(R1859t1522) I(R1860t1585) I(R1861t361) I(R1861t1629) I(R1862t1263) I(R1862t338) I(R1863t1624) I(R1863t223) I(R1863t347) I(R1864t1714) I(R1864t1437) I(R1864t1458) I(R1865t234) I(R1865t1153) I(R1866t1385) I(R1867t752) I(R1867t504) I(R1868t1341) I(R1868t366) I(R1869t1472) I(R1874t834) I(R1876t1038) I(R1877t238) I(R1877t609) I(R1877t821) I(R1879t578) I(R1879t870) I(R1880t506) I(R1880t1284) I(R1881t1572) I(R1882t936) I(R1883t91) I(R1883t901) I(R1883t750) I(R1884t422) I(R1885t1005) I(R1885t388) I(R1887t1489) I(R1887t1430) I(R1887t938) I(R1888t455) I(R1889t42) I(R1893t338) I(R1893t1209) I(R1894t1605) I(R1895t437) I(R1895t1008) I(R1897t416) I(R1900t1608) I(R1901t263) I(R1902t813) I(R1902t617) I(R1903t1876) I(R1905t294) I(R1905t1820) I(R1906t648) I(R1906t913) I(R1907t399) I(R1908t453) I(R1908t415) I(R1909t275) I(R1909t48) I(R1910t535) I(R1911t37) I(R1912t1104) I(R1914t1497) I(R1914t1738) I(R1917t216) I(R1917t356) I(R1918t503) I(R1919t1744) I(R1920t701) I(R1921t252) I(R1921t729) I(R1922t601) I(R1922t496) I(R1924t989) I(R1924t1222) I(R1925t1776) I(R1926t328) I(R1926t752) I(R1926t1867) I(R1926t651) I(R1927t458) I(R1928t288) I(R1929t856) I(R1930t1631) I(R1930t302) I(R1931t47) I(R1931t114) I(R1932t203) I(R1932t1802) I(R1933t1834) I(R1933t1739) I(R1934t167) I(R1934t1629) I(R1934t361) I(R1934t685) I(R1935t1381) I(R1937t193) I(R1937t1165) I(R1938t1100) I(R1938t914) I(R1940t1025) I(R1941t1390) I(R1942t387) I(R1942t1456) I(R1944t1744) I(R1944t1919) I(R1948t638) I(R1950t1303) I(R1952t1710) I(R1952t326) I(R1954t1093) I(R1955t1049) I(R1956t221) I(R1957t1539) I(R1957t962) I(R1960t983) I(R1961t728) I(R1962t1746) I(R1962t1760) I(R1963t948) I(R1964t474) I(R1967t1090) I(R1968t1401) I(R1969t1681) I(R1970t456) I(R1973t50) I(R1974t1131) I(R1975t459) I(R1976t1400) I(R1976t661) I(R1977t1033) I(R1977t1481) I(R1977t481) I(R1979t856) I(R1979t1929) I(R1980t1607) I(R1980t1622) I(R1980t1716) I(R1981t742) I(R1981t1587) I(R1982t1335) I(R1982t1800) I(R1982t988) I(R1983t1229) I(R1985t972) I(R1985t1006) I(R1985t139) I(R1986t929) I(R1986t697) I(R1987t936) I(R1988t1685) I(R1988t1032) I(R1989t577) I(R1989t873) I(R1991t1598) I(R1992t40) I(R1993t1369) I(R1995t990) I(R1995t943) I(R1995t131) I(R1999t1214) I(R2000t350) I(R2001t1463) I(R2002t345) I(R2004t463) I(R2004t1429) I(R2005t104) I(R2006t1984) I(R2007t733) I(R2009t810) I(R2009t1562) I(R2009t439) I(R2010t347) I(R2010t1863) I(R2011t1503) I(R2011t1722) I(R2012t885) I(R2015t1577) I(R2016t733) I(R2016t1589) I(R2017t1428) I(R2018t477) I(R2019t1664) I(R2022t735) I(R2022t1328) I(R2024t946) I(R2024t954) I(R2025t723) I(R2026t306) I(R2027t536) I(R2028t855) I(R2028t1518) I(R2028t1294) I(R2030t594) I(R2031t1754) I(R2033t196) I(R2035t1937) I(R2036t459) I(R2036t793) I(R2042t620) I(R2043t1757) I(R2044t309) I(R2045t350) I(R2047t1812) I(R2047t1645) I(R2049t1190) I(R2050t1285) I(R2050t1226) I(R2050t149) I(R2051t529) I(R2052t1593) I(R2053t898) I(R2053t656) I(R2054t1293) I(R2054t1740) I(R2054t105) I(R2054t70) I(R2055t250) I(R2056t581) I(R2059t945) I(R2060t122) I(R2061t1034) I(R2062t1676) I(R2064t1014) I(R2065t766) I(R2066t1459) I(R2068t1950) I(R2068t1303) I(R2071t643) I(R2073t1886) I(R2074t1178) I(R2074t1388) I(R2074t1227) I(R2074t1145) I(R2075t210) I(R2076t657) I(R2077t136) I(R2078t224) I(R2078t1325) I(R2078t1915) I(R2078t1055) I(R2079t1085) I(R2080t1248) I(R2080t327) I(R2081t1967) I(R2082t642) I(R2082t1088) I(R2083t814) I(R2084t99) I(R2085t1384) I(R2086t1893) I(R2087t1828) I(R2087t1617) I(R2087t1635) I(R2087t644) I(R2087t1129) I(R2088t1740) I(R2088t105) I(R2089t401) I(R2092t1858) I(R2094t1373) I(R2097t223) I(R2097t1863) I(R2098t730) I(R2098t271) I(R2099t952) I(R2099t768) I(R2099t1848) I(R2100t154) I(R2100t1777) I(R2101t817) I(R2101t14) I(R2103t474) I(R2103t400) I(R2103t1482) I(R2104t235) I(R2104t1720) I(R2105t1141) I(R2105t669) I(R2105t1903) I(R2106t2105) I(R2106t669) I(R2107t1327) I(R2107t639) I(R2108t1742) I(R2108t1224) I(R2110t1246) I(R2111t1148) I(R2111t720) I(R2111t1549) I(R2112t712) I(R2112t403) I(R2114t362) I(R2114t475) I(R2114t1680) I(R2116t1287) I(R2116t113) I(R2116t1355) I(R2117t1246) I(R2117t2110) I(R2118t1462) I(R2118t732) I(R2118t961) I(R2118t440) I(R2120t1741) I(R2122t1259) I(R2123t399) I(R2123t987) I(R2124t1487) I(R2125t670) I(R2126t637) I(R2126t1449) I(R2127t336) I(R2127t1817) I(R2127t918) I(R2128t1286) I(R2128t2119) I(R2129t654) I(R2130t1570) I(R2132t1611) I(R2133t234) I(R2133t1865) I(R2134t1020) I(R2134t638) I(R2135t1510) I(R2136t1972) I(R2138t983) I(R2138t1960) I(R2138t994) I(R2139t1943) I(R2142t1760) I(R2143t423) I(R2143t65) I(R2144t471) I(R2145t709) I(R2147t25) I(R2147t93) I(R2148t1443) I(R2149t1764) I(R2150t594) I(R2151t207) I(R2151t1481) I(R2152t1493) I(R2153t830) I(R2153t516) I(R2153t1508) I(R2154t1620) I(R2155t233) I(R2156t1168) I(R2156t282) I(R2157t938) I(R2157t596) I(R2157t1137) I(R2158t1447) I(R2159t451) I(R2160t95) I(R2162t2109) I(R2163t32) I(R2164t1181) I(R2166t1820) I(R2166t1905) I(R2167t1765) I(R2167t1806) I(R2168t1775) I(R2168t201) I(R2168t967) I(R2169t523) I(R2170t377) I(R2170t155) I(R2171t1751) I(R2173t652) I(R2174t1494) I(R2174t255) I(R2174t297) I(R2175t215) I(R2175t1780) I(R2176t1176) I(R2176t1691) I(R2176t1111) I(R2177t1176) I(R2177t63) I(R2178t287) I(R2179t1674) I(R2180t311) I(R2181t411) I(R2181t566) I(R2183t1801) I(R2183t1370) I(R2184t1520) I(R2186t1817) I(R2186t1535) I(R2187t2185) I(R2188t1305) I(R2191t1929) I(R2191t1687) I(R2192t191) I(R2192t1753) I(R2192t505) I(R2194t744) I(R2195t126) I(R2195t1643) I(R2195t1061) I(R2199t19) I(R2199t1036) I(R2201t1899) I(R2201t1663) I(R2202t504) I(R2202t792) I(R2202t713) I(R2203t1636) I(R2203t340) I(R2204t1417) I(R2206t1776) I(R2207t487) I(R2207t1347) I(R2207t1717) I(R2208t2136) I(R2209t1243) I(R2210t1158) I(R2211t2140) I(R2212t1696) I(R2213t2017) I(R2213t1053) I(R2215t330) I(R2216t705) I(R2218t2146) I(R2219t316) I(R2219t1516) I(R2219t1299) I(R2220t570) I(R2221t1274) I(R2221t1049) I(R2222t869) I(R2223t380) I(R2224t2065) I(R2226t1808) I(R2227t33) I(R2227t170) I(R2229t1864) I(R2229t1714) I(R2229t705) I(R2230t1289) I(R2231t1395) I(R2231t1298) I(R2231t788) I(R2231t1975) I(R2231t343) I(R2234t366) I(R2234t2130) I(R2235t2182) I(R2236t2150) I(R2236t2030) I(R2236t594) I(R2237t970) I(R2237t484) I(R2238t1729) I(R2239t878) I(R2240t2105) I(R2241t22) I(R2241t1387) I(R2243t280) I(R2243t1485) I(R2244t1983) I(R2244t1943) I(R2245t645) I(R2246t1203) I(R2247t1670) I(R2248t1163) I(R2249t1672) I(R2250t1121) I(R2251t284) I(R2253t22) I(R2253t2241) I(R2253t801) I(R2254t1129) I(R2256t2023) I(R2256t1884) I(R2256t342) I(R2257t2217) I(R2258t60) I(R2258t1318) I(R2259t1175) I(R2260t1397) I(R2261t1146) I(R2261t1502) I(R2261t1760) I(R2262t216) I(R2262t1917) I(R2262t356) I(R2263t217) I(R2263t1634) I(R2264t600) I(R2264t15) I(R2264t1309) I(R2265t1900) I(R2267t316) I(R2267t1516) I(R2268t2048) I(R2269t224) I(R2269t2078) I(R2269t1055) I(R2270t1946) I(R2270t519) I(R2274t2230) I(R2274t499) I(R2275t76) I(R2275t976) I(R2275t1392) I(R2275t456) I(R2275t998) I(R2276t1694) I(R2276t522) I(R2278t1170) I(R2278t269) I(R2279t429) I(R2279t560) I(R2280t472) I(R2280t1293) I(R2280t2109) I(R2281t257) I(R2282t2208) I(R2282t1139) I(R2283t470) I(R2283t999) I(R2284t329) I(R2284t442) I(R2285t449) I(R2287t848) I(R2288t171) I(R2289t2052) I(R2290t906) I(R2291t383) I(R2291t558) I(R2291t476) I(R2292t106) I(R2293t1983) I(R2293t2244) I(R2294t2286) I(R2295t21) I(R2295t1045) I(R2295t1479) I(R2296t823) I(R2296t245) I(R2297t506) I(R2297t605) I(R2297t1880) I(R2298t2093) I(R2299t2030) I(R2299t2236) I(R2300t318) I(R2301t1930) I(R2302t1182) I(R2303t2021) I(R2304t727) I(R2305t397) I(R2305t722) I(R2306t770) I(R2306t1163) I(R2307t2013) I(R2307t1385) I(R2308t960) I(R2308t1518) I(R2308t1412) I(R2308t1465) I(R2311t664) I(R2313t19) I(R2314t1898) I(R2315t1824) I(R2315t2094) I(R2316t1125) I(R2318t1245) I(R2319t1327) I(R2319t2107) I(R2320t523) I(R2320t916) I(R2322t822) I(R2324t1160) I(R2325t368) I(R2326t337) I(R2327t1611) I(R2327t771) I(R2328t1149) I(R2331t108) I(R2332t812) I(R2332t349) I(R2332t1693) I(R2334t1968) I(R2335t1163) I(R2336t2332) I(R2336t349) I(R2338t164) I(R2338t1130) I(R2338t863) I(R2339t1208) I(R2339t1119) I(R2340t1323) I(R2342t1342) I(R2343t1173) I(R2343t1795) I(R2344t2126) I(R2344t1449) I(R2344t1850) I(R2344t246) I(R2345t78) I(R2345t1097) I(R2345t1021) I(R2346t117) I(R2347t2200) I(R2347t2242) I(R2348t513) I(R2348t387) I(R2349t622) I(R2349t2147) I(R2350t1632) I(R2350t7) I(R2351t1887) I(R2351t938) I(R2352t563) I(R2352t1984) I(R2354t370) I(R2354t279) I(R2355t670) I(R2355t391) I(R2356t231) I(R2359t294) I(R2359t1130) I(R2359t164) I(R2360t1990) I(R2360t2301) I(R2363t263) I(R2363t702) I(R2364t1741) I(R2364t2120) I(R2365t409) I(R2366t2239) I(R2366t878) I(R2366t1461) I(R2368t841) I(R2370t635) I(R2370t540) I(R2371t267) I(R2371t1202) I(R2371t2011) I(R2372t1359) I(R2373t2081) I(R2375t1759) I(R2375t1172) I(R2379t1189) I(R2379t395) I(R2380t1945) I(R2380t240) I(R2381t607) I(R2381t1529) I(R2382t2267) I(R2382t316) I(R2382t2219) I(R2383t470) I(R2383t2283) I(R2383t999) I(R2384t509) I(R2384t1683) I(R2385t880) I(R2385t767) I(R2385t457) I(R2386t434) I(R2386t430) I(R2387t2018) I(R2387t2356) I(R2387t706) I(R2388t1968) I(R2388t2334) I(R2389t318) I(R2389t2300) I(R2389t613) I(R2391t1723) I(R2391t841) I(R2391t1978) I(R2392t1936) I(R2392t1927) I(R2392t2005) I(R2392t104) I(R2393t680) I(R2394t1641) I(R2396t1512) I(R2397t5) I(R2397t1451) I(R2397t241) I(R2397t681) I(R2398t502) I(R2398t1158) I(R2398t12) I(R2400t1316) I(R2401t1348) I(R2401t1543) I(R2401t266) I(R2402t181) I(R2404t1073) I(R2405t1302) I(R2406t773) I(R2406t53) I(R2407t1835) I(R2407t2140) I(R2408t2148) I(R2408t1443) I(R2408t791) I(R2409t858) I(R2409t26) I(R2410t253) I(R2411t1731) I(R2411t966) I(R2412t256) I(R2413t616) I(R2414t1936) I(R2415t1961) I(R2415t728) I(R2416t1514) I(R2418t102) I(R2418t1390) I(R2419t1940) I(R2419t1025) I(R2420t1532) I(R2422t2141) I(R2422t365) I(R2423t971) I(R2423t1225) I(R2423t546) I(R2423t109) I(R2426t554) I(R2427t207) I(R2428t1880) I(R2428t1284) I(R2429t2324) I(R2429t296) I(R2430t2268) I(R2432t2194) I(R2432t744) I(R2433t243) I(R2433t254) I(R2433t860) I(R2434t1168) I(R2434t2156) I(R2434t282) I(R2434t1050) I(R2435t1040) I(R2436t2362) I(R2436t449) I(R2437t606) I(R2437t1826) I(R2438t2301) I(R2438t1930) I(R2438t1631) I(R2441t365) I(R2441t334) I(R2442t1500) I(R2443t1403) I(R2444t2321) I(R2445t940) I(R2445t1987) I(R2445t936) I(R2446t1625) I(R2447t969) I(R2448t1189) I(R2449t1934) I(R2449t305) I(R2449t685) I(R2450t1551) I(R2450t1806) I(R2450t824) I(R2450t2167) I(R2454t508) I(R2454t1444) I(R2455t212) I(R2456t1393) I(R2457t2150) I(R2457t2236) I(R2457t2299) I(R2458t1112) I(R2458t1437) I(R2459t172) I(R2459t786) I(R2459t718) I(R2459t1031) I(R2459t1295) I(R2460t611) I(R2460t1474) I(R2461t628) I(R2461t1446) I(R2461t195) I(R2462t1297) I(R2462t679) I(R2462t127) I(R2463t301) I(R2465t442) I(R2465t805) I(R2465t495) I(R2466t2249) I(R2467t1854) I(R2467t1167) I(R2468t2173) I(R2468t652) I(R2468t33) I(R2468t2227) I(R2469t1206) I(R2469t353) I(R2469t1662) I(R2470t1754) I(R2470t2031) I(R2470t1124) I(R2471t787) I(R2472t305) I(R2472t2449) I(R2472t685) I(R2472t488) I(R2473t891) I(R2473t548) I(R2474t1969) I(R2474t2187) I(R2476t987) I(R2476t1136) I(R2477t1071) I(R2478t2441) I(R2479t531) I(R2479t941) I(R2479t101) I(R2479t1550) I(R2480t1288) I(R2483t1147) I(R2483t1682) I(R2483t484) I(R2484t1578) I(R2485t1506) I(R2487t1315) I(R2487t1698) I(R2487t671) I(R2488t126) I(R2488t2195) I(R2489t102) I(R2489t2488) I(R2490t588) I(R2490t374) I(R2491t181) I(R2491t2402) I(R2491t2076) I(R2493t140) I(R2493t1778) I(R2494t1669) I(R2494t1618) I(R2495t2327) I(R2496t2122) I(R2496t924) I(R2497t627) I(R2499t1049) I(R2499t348) I(R2500t614) I(R2500t1279) I(R2500t1119) I(R2501t1324) I(R2502t1552) I(R2502t1201) I(R2503t1884) I(R2503t2256) I(R2503t2023) I(R2504t854) I(R2505t1080) I(R2506t1084) I(R2506t1839) I(R2506t1670) I(R2507t983) I(R2508t826) I(R2509t832) I(R2510t975) I(R2510t1060) I(R2510t783) I(R2511t224) I(R2511t2078) I(R2511t1325) I(R2512t1752) I(R2513t1661) I(R2514t1277) I(R2514t1337) I(R2514t2019) I(R2515t1699) I(R2516t169) I(R2516t738) I(R2516t183) I(R2517t2162) I(R2517t1740) I(R2519t1228) I(R2520t2339) I(R2520t624) I(R2521t390) I(R2521t1357) I(R2522t2121) I(R2523t199) I(R2524t489) I(R2525t83) I(R2525t1892) I(R2528t1938) I(R2529t62) I(R2531t1399) I(R2531t1730) I(R2531t130) I(R2532t383) I(R2532t2291) I(R2533t1354) I(R2533t1000) I(R2533t81) I(R2535t364) I(R2537t177) I(R2537t1042) I(R2538t371) I(R2539t1912) I(R2540t2509) I(R2541t2513) I(R2541t1597) I(R2541t1661) I(R2542t195) I(R2544t1334) I(R2547t1646) I(R2548t53) I(R2549t2527) I(R2550t2510) I(R2550t783) I(R2551t2328) I(R2551t163) I(R2552t971) I(R2552t916) I(R2553t1249) I(R2554t68) I(R2554t119) I(R2554t1374) I(R2556t1068) I(R2557t1891) I(R2557t2535) I(R2559t1838) I(R2560t1577) I(R2561t2122) I(R2561t2496) I(R2561t1259) I(R2563t1656) I(R2563t1185) I(R2564t601) I(R2565t1116) I(R2565t1468) I(R2566t2212) I(R2567t444) I(R2567t968) I(R2568t1912) I(R2568t2539) I(R2568t1104) I(R2570t1652) I(R2571t1084) I(R2572t586) I(R2572t1590) I(R2572t2542) I(R2573t785) I(R2573t859) I(R2573t541) I(R2574t2230) I(R2575t1076) I(R2576t2333) I(R2576t719) I(R2577t1662) I(R2577t1473) I(R2577t1751) I(R2577t2171) I(R2578t1243) I(R2578t2209) I(R2578t94) I(R2579t2048) I(R2579t526) I(R2580t345) I(R2581t1514) I(R2581t243) I(R2582t341) I(R2583t2115) I(R2583t1508) I(R2583t516) I(R2584t2182) I(R2584t399) I(R2584t2123) I(R2586t14) I(R2587t2263) I(R2587t1634) I(R2588t1859) I(R2588t1754) I(R2588t2470) I(R2588t1124) I(R2589t1112) I(R2589t1168) I(R2589t2458) I(R2589t1050) I(R2589t2434) I(R2590t187) I(R2591t394) I(R2592t1283) I(R2592t953) I(R2592t971) I(R2593t1280) I(R2596t551) I(R2596t2102) I(R2598t1787) I(R2599t1385) I(R2601t1276) I(R2602t2262) I(R2602t216) I(R2603t403) I(R2603t1044) I(R2603t712) I(R2603t2112) I(R2605t1575) I(R2605t1856) I(R2608t255) I(R2610t2502) I(R2611t1878) I(R2612t1365) I(R2612t1993) I(R2613t31) I(R2614t2214) I(R2614t1) I(R2614t1625) I(R2615t743) I(R2615t385) I(R2616t2045) I(R2616t2000) I(R2616t350) I(R2617t393) I(R2617t724) I(R2617t977) I(R2619t1681) I(R2619t1969) I(R2620t1719) I(R2622t2208) I(R2622t2282) I(R2622t1139) I(R2625t2507) I(R2625t983) I(R2625t1570) I(R2627t2090) I(R2627t107) I(R2628t433) I(R2629t2442) I(R2630t1904) I(R2631t2432) I(R2631t744) I(R2632t1614) I(R2633t631) I(R2633t1513) I(R2634t1874) I(R2635t359) I(R2635t1782) I(R2638t1592) I(R2638t2480) I(R2639t1794) I(R2640t540) I(R2641t2365) I(R2642t2350) I(R2642t7) I(R2643t1186) I(R2644t2612) I(R2645t2037) I(R2647t2192) I(R2647t191) I(R2647t202) I(R2648t1491) I(R2649t1841) I(R2650t138) I(R2650t929) I(R2651t565) I(R2651t425) I(R2651t843) I(R2652t1368) I(R2652t1799) I(R2654t1636) I(R2654t2203) I(R2655t812) I(R2655t498) I(R2655t349) I(R2655t2332) I(R2656t2040) I(R2657t2626) I(R2657t219) I(R2658t2458) I(R2658t2589) I(R2658t1437) I(R2658t1714) I(R2658t1050) I(R2659t1674) I(R2660t2464) I(R2660t15) I(R2660t1413) I(R2662t304) I(R2663t1306) I(R2663t1004) I(R2665t1003) I(R2665t2189) I(R2666t511) I(R2666t1902) I(R2667t1762) I(R2667t181) I(R2667t2402) I(R2667t645) I(R2668t1206) I(R2668t405) I(R2670t2211) I(R2671t811) I(R2672t1851) I(R2672t910) I(R2672t485) I(R2674t189) I(R2675t509) I(R2675t775) I(R2676t2193) I(R2676t2223) I(R2676t380) I(R2676t240) I(R2677t1575) I(R2677t2605) I(R2677t1856) I(R2678t2093) I(R2678t2163) I(R2679t1286) I(R2679t1772) I(R2679t2128) I(R2680t672) I(R2681t62) I(R2681t2529) I(R2682t2657) I(R2682t2626) I(R2683t166) I(R2685t2240) I(R2685t2545) I(R2685t1903) I(R2685t2105) I(R2686t2192) I(R2686t2647) I(R2686t873) I(R2687t511) I(R2687t1241) I(R2687t813) I(R2687t1902) I(R2687t2666) I(R2688t2092) I(R2689t1843) I(R2689t691) I(R2690t2177) I(R2690t63) I(R2691t854) I(R2692t841) I(R2692t2391) I(R2693t948) I(R2694t138) I(R2694t849) I(R2695t2317) I(R2695t1427) I(R2696t450) I(R2697t1438) I(R2697t1773) I(R2697t2420) I(R2698t2669) I(R2699t2295) I(R2701t459) I(R2701t1649) I(R2701t2036) I(R2702t727) I(R2702t2032) I(R2702t1458) I(R2703t2486) I(R2704t458) I(R2704t599) I(R2704t915) I(R2705t2567) I(R2705t182) I(R2706t1569) I(R2707t944) I(R2707t506) I(R2707t131) I(R2708t1200) I(R2708t281) I(R2709t71) I(R2709t687) I(R2709t1380) I(R2710t1822) I(R2710t1384) I(R2711t242) I(R2712t1213) I(R2714t952) I(R2715t2362) I(R2715t2436) I(R2715t151) I(R2716t1012) I(R2716t1250) I(R2717t2536) I(R2717t564) I(R2718t556) I(R2719t2233) I(R2720t593) I(R2722t1182) I(R2722t2302) I(R2723t749) I(R2724t536) I(R2724t2027) I(R2725t1016) I(R2725t389) I(R2726t1621) I(R2727t1779) I(R2729t826) I(R2729t875) I(R2730t115) I(R2730t1359) I(R2731t832) I(R2731t1586) I(R2732t1553) I(R2733t38) I(R2734t323) I(R2734t79) I(R2734t1744) I(R2734t1919) I(R2735t2636) I(R2735t2233) I(R2735t2719) I(R2737t1807) I(R2738t262) I(R2739t701) I(R2739t293) I(R2742t1490) I(R2742t2630) I(R2742t1904) I(R2743t2437) I(R2744t141) I(R2744t610) I(R2744t2604) I(R2745t1302) I(R2746t966) I(R2746t729) I(R2746t359) I(R2746t2411) I(R2747t1118) I(R2749t2378) I(R2750t896) I(R2751t2679) I(R2751t162) I(R2752t794) I(R2752t585) I(R2753t167) I(R2753t1934) I(R2755t115) I(R2755t1819) I(R2755t1359) I(R2755t2730) I(R2756t2149) I(R2756t1764) I(R2757t2233) I(R2757t2636) I(R2758t931) I(R2758t1574) I(R2759t1333) I(R2759t1856) I(R2759t2605) I(R2761t220) I(R2762t820) I(R2762t2599) I(R2763t1614) I(R2763t2632) I(R2763t552) I(R2764t2358) I(R2765t1775) I(R2765t2168) I(R2767t2095) I(R2768t1631) I(R2768t302) I(R2768t1801) I(R2769t2640) I(R2770t801) I(R2770t22) I(R2770t1387) I(R2771t2458) I(R2771t1196) I(R2771t1458) I(R2771t1437) I(R2773t1460) I(R2773t1520) I(R2774t2337) I(R2774t1498) I(R2775t1488) I(R2776t1312) I(R2777t687) I(R2777t2709) I(R2778t1742) I(R2778t1235) I(R2778t1224) I(R2779t2086) I(R2779t1893) I(R2780t776) I(R2781t2544) I(R2781t1626) I(R2784t121) I(R2785t1957) I(R2785t2251) I(R2785t284) I(R2785t662) I(R2785t1539) I(R2786t786) I(R2786t859) I(R2786t172) I(R2788t815) I(R2788t1807) I(R2788t432) I(R2789t34) I(R2791t820) I(R2791t2762) I(R2792t1763) I(R2792t1599) I(R2793t442) I(R2794t1362) I(R2794t2382) I(R2794t1269) I(R2795t2212) I(R2795t1696) I(R2795t348) I(R2795t2499) I(R2796t96) I(R2796t155) I(R2797t2218) I(R2798t774) I(R2798t2029) I(R2798t1282) I(R2799t1651) I(R2800t2427) I(R2800t207) I(R2800t2151) I(R2801t2265) I(R2801t1688) I(R2801t40) I(R2801t1992) I(R2802t907) I(R2802t251) I(R2803t2362) I(R2803t2715) I(R2803t173) I(R2804t1877) I(R2806t2193) I(R2807t1510) I(R2808t1242) I(R2808t1267) I(R2809t1588) I(R2810t1175) I(R2810t2259) I(R2810t417) I(R2811t631) I(R2811t2633) I(R2811t1513) I(R2812t2312) I(R2812t1199) I(R2813t476) I(R2813t2260) I(R2813t1397) I(R2814t2316) I(R2815t2580) I(R2815t139) I(R2816t542) I(R2818t2234) I(R2818t366) I(R2818t211) I(R2818t1947) I(R2820t886) I(R2820t2688) I(R2821t1034) I(R2821t1240) I(R2821t2061) I(R2822t554) I(R2822t142) I(R2823t1545) I(R2823t466) I(R2824t2313) I(R2825t726) I(R2826t814) I(R2826t2083) I(R2827t2497) I(R2827t1087) I(R2828t2164) I(R2830t2636) I(R2830t2757) I(R2830t2735) I(R2830t2233) I(R2831t2382) I(R2831t2790) I(R2831t2326) I(R2832t2775) I(R2833t1380) I(R2833t930) I(R2834t1344) I(R2834t1843) I(R2836t1131) I(R2836t1302) I(R2837t1280) I(R2837t1358) I(R2838t1484) I(R2839t1990) I(R2839t1339) I(R2840t761) I(R2840t1421) I(R2841t23) I(R2841t1338) I(R2841t471) I(R2841t2144) I(R2842t2585) I(R2843t2034) I(R2844t2780) I(R2845t1615) I(R2845t1799) I(R2845t2652) I(R2846t2528) I(R2846t1938) I(R2846t1100) I(R2846t872) I(R2846t295) I(R2847t1439) I(R2847t1652) I(R2849t1385) I(R2850t1087) I(R2851t1638) I(R2851t2100) I(R2851t1777) I(R2852t420) I(R2853t452) I(R2853t796) I(R2855t1602) I(R2856t1971) I(R2856t708) I(R2857t101) I(R2858t2284) I(R2858t442) I(R2858t2793) I(R2859t1376) I(R2860t2525) I(R2860t1288) I(R2860t345) I(R2860t2002) I(R2861t2632) I(R2861t1614) I(R2863t2192) I(R2863t2686) I(R2863t505) I(R2863t539) I(R2864t2222) I(R2864t1341) I(R2864t1231) I(R2865t968) I(R2865t608) I(R2866t1385) I(R2866t2307) I(R2866t2599) I(R2866t2762) I(R2868t2641) I(R2868t1041) I(R2869t2417) I(R2870t1212) I(R2870t363) I(R2870t2033) I(R2870t2142) I(R2871t2538) I(R2871t2247) I(R2872t1883) I(R2873t1939) I(R2873t127) I(R2873t2656) I(R2873t2040) I(R2873t2358) I(R2874t1806) I(R2875t629) I(R2876t2442) I(R2876t2629) I(R2877t177) I(R2877t2537) I(R2878t1636) I(R2879t1258) I(R2879t1716) I(R2879t1980) I(R2879t1622) I(R2880t359) I(R2880t2635) I(R2882t2606) I(R2882t1623) I(R2882t1188) I(R2883t2566) I(R2884t2588) I(R2884t1559) I(R2884t1174) I(R2884t1124) I(R2886t1654) I(R2887t2527) I(R2887t2549) I(R2888t45) I(R2888t544) I(R2889t1101) I(R2889t2264) I(R2889t1309) I(R2890t1206) I(R2890t2469) I(R2890t2426) I(R2890t353) I(R2891t715) I(R2892t1909) I(R2892t48) I(R2894t2544) I(R2895t229) I(R2896t1215) I(R2896t524) I(R2897t1744) I(R2897t1944) I(R2897t2894) I(R2898t342) I(R2899t833) I(R2901t1195) I(R2902t979) I(R2902t860) I(R2902t2433) I(R2902t243) I(R2903t2200) I(R2903t1260) I(R2904t341) I(R2904t2582) I(R2905t1788) I(R2906t2126) I(R2906t637) I(R2906t264) I(R2906t1416) I(R2906t1519) I(R2906t877) I(R2907t1505) I(R2907t2767) I(R2909t1735) I(R2909t543) I(R2910t1257) I(R2912t759) I(R2912t1594) I(R2913t1674) I(R2914t606) I(R2915t2333) I(R2915t1364) I(R2916t735) I(R2916t2721) I(R2916t163) I(R2917t2478) I(R2918t461) I(R2918t2114) I(R2918t995) I(R2919t561) I(R2920t736) I(R2920t878) I(R2920t2239) I(R2922t1346) I(R2922t784) I(R2923t1890) I(R2923t1608) I(R2924t407) I(R2924t1795) I(R2925t727) I(R2925t2304) I(R2926t2298) I(R2926t2093) I(R2927t510) I(R2928t2194) I(R2929t1480) I(R2929t65) I(R2930t908) I(R2931t2881) I(R2932t769) I(R2932t2783) I(R2933t1990) I(R2933t2360) I(R2933t2301) I(R2934t2325) I(R2934t134) I(R2935t2442) I(R2935t2293) I(R2935t2629) I(R2936t1873) I(R2937t1343) I(R2937t1792) I(R2938t428) I(R2938t1477) I(R2940t663) I(R2942t2777) I(R2942t687) I(R2944t2848) I(R2945t2939) I(R2946t2829) I(R2947t2840) I(R2947t761) I(R2948t339) I(R2948t1739) I(R2948t1545) I(R2949t1466) I(R2950t186) I(R2950t321) I(R2950t1785) I(R2950t2071) I(R2951t58) I(R2951t457) I(R2951t767) I(R2951t45) I(R2952t1867) I(R2953t2667) I(R2953t645) I(R2953t2245) I(R2954t2709) I(R2955t1373) I(R2956t2341) I(R2957t1549) I(R2957t567) I(R2958t2673) I(R2959t854) I(R2959t2504) I(R2960t161) I(R2960t1682) I(R2960t2736) I(R2961t2002) I(R2961t345) I(R2961t2580) I(R2963t535) I(R2963t1910) I(R2963t759) I(R2963t2912) I(R2965t676) I(R2966t643) I(R2966t2931) I(R2966t2881) I(R2967t2378) I(R2967t2927) I(R2969t1304) I(R2971t1389) I(R2972t34) I(R2972t2789) I(R2973t1849) I(R2974t1028) I(R2975t76) I(R2975t1267) I(R2975t1242) I(R2976t1378) I(R2978t1127) I(R2979t1807) I(R2979t815) I(R2979t2788) I(R2980t1500) I(R2980t2091) I(R2980t1154) I(R2980t1037) I(R2981t1404) I(R2981t177) I(R2982t1118) I(R2982t2747) I(R2982t1655) I(R2982t704) I(R2983t1194) I(R2983t994) I(R2983t1736) I(R2984t2483) I(R2985t1024) I(R2985t1086) I(R2986t314) I(R2989t1701) I(R2990t726) I(R2991t2443) I(R2991t2400) I(R2993t2507) I(R2993t267) I(R2994t2787) I(R2995t2690) I(R2995t2597) I(R2996t46) I(R2996t1115) I(R2997t2194) I(R2997t2928) I(R2999t1068) I(R3000t219) I(R3000t1142) I(R3000t831) I(R3001t956) I(R3001t2662) I(R3002t1626) I(R3002t2781) I(R3003t806) I(R3003t1224) I(R3004t493) I(R3005t2020) I(R3005t12) I(R3006t2357) I(R3006t1949) I(R3007t1080) I(R3007t2505) I(R3008t1602) I(R3008t1537) I(R3010t1446) I(R3010t659) I(R3010t693) I(R3011t1475) I(R3011t471) I(R3012t1491) I(R3013t1636) I(R3013t2654) I(R3013t2312) I(R3013t2812) I(R3014t1521) I(R3014t827) I(R3015t431) I(R3016t954) I(R3017t2325) I(R3017t1099) I(R3018t956) I(R3018t2364) I(R3019t2065) I(R3019t766) I(R3019t1668) I(R3020t2501) I(R3020t800) I(R3020t1324) I(R3021t1131) I(R3021t1974) I(R3021t2836) I(R3022t1743) I(R3022t394) I(R3023t2335) I(R3025t2209) I(R3025t1766) I(R3025t1638) I(R3025t2851) I(R3025t2100) I(R3026t1435) I(R3027t1126) I(R3027t1593) I(R3027t2052) I(R3027t2289) I(R3028t1723) I(R3028t1978) I(R3028t2391) I(R3029t881) I(R3029t373) I(R3030t1501) I(R3030t1029) I(R3031t1079) I(R3032t2421) I(R3033t1233) I(R3033t2076) I(R3033t2491) I(R3033t2402) I(R3034t711) I(R3034t2477) I(R3034t634) I(R3035t2732) I(R3036t2210) I(R3036t1158) I(R3037t1290) I(R3037t1872) I(R3038t945) I(R3038t2286) I(R3038t530) I(R3038t703) I(R3039t1625) I(R3041t577) I(R3041t991) I(R3041t2997) I(R3042t1662) I(R3042t353) I(R3043t123) I(R3043t1767) I(R3044t710) I(R3045t2650) I(R3045t929) I(R3047t2390) I(R3048t1783) I(R3049t738) I(R3049t169) I(R3049t1470) I(R3050t2135) I(R3050t1510) I(R3051t2639) I(R3052t2455) I(R3052t212) I(R3053t1125) I(R3053t2031) I(R3054t1587) I(R3055t919) I(R3055t2968) I(R3056t725) I(R3056t1445) I(R3057t2113) I(R3057t1729) I(R3057t2238) I(R3058t324) I(R3058t2898) I(R3058t342) I(R3058t2256) I(R3058t1884) I(R3058t422) I(R3059t962) I(R3060t319) I(R3060t1005) I(R3060t568) I(R3060t388) I(R3062t1452) I(R3062t196) I(R3062t2033) I(R3063t448) I(R3064t1183) I(R3064t2867) I(R3064t1703) I(R3065t1892) I(R3065t1026) I(R3066t1651) I(R3066t2799) I(R3066t1045) I(R3066t1213) I(R3066t2712) I(R3067t427) I(R3067t778) I(R3068t712) I(R3068t2603) I(R3068t2877) I(R3069t801) I(R3069t2770) I(R3070t494) I(R3070t1390) I(R3071t1993) I(R3071t1369) I(R3072t1560) I(R3072t64) I(R3072t245) I(R3073t1062) I(R3073t1646) I(R3073t2547) I(R3073t1234) I(R3074t1039) I(R3074t2678) I(R3074t2163) I(R3075t2872) I(R3076t2392) I(R3076t104) I(R3077t2228) I(R3078t1301) I(R3078t1346) I(R3078t784) I(R3079t1025) I(R3079t2419) I(R3080t2762) I(R3081t2086) I(R3082t881) I(R3082t2314) I(R3083t602) I(R3083t1017) I(R3083t2808) I(R3084t2381) I(R3084t607) I(R3084t2073) I(R3085t2498) I(R3085t2259) I(R3087t921) I(R3089t1495) I(R3090t2360) I(R3090t2438) I(R3090t1631) I(R3090t98) I(R3090t2546) I(R3092t608) I(R3093t2163) I(R3093t2678) I(R3094t907) I(R3094t2828) I(R3095t1078) I(R3095t1685) I(R3095t1575) I(R3096t885) I(R3097t42) I(R3098t2970) I(R3098t537) I(R3098t3055) I(R3099t1978) I(R3100t2353) I(R3101t1030) I(R3102t1047) I(R3102t348) I(R3102t2795) I(R3103t1074) I(R3103t747) I(R3105t866) I(R3105t845) I(R3106t3009) I(R3107t1174) I(R3107t1559) I(R3107t2884) I(R3108t1456) I(R3108t1709) I(R3108t1308) I(R3108t412) I(R3109t2955) I(R3110t2534) I(R3111t3091) I(R3112t2652) I(R3112t2424) I(R3113t1751) I(R3113t249) I(R3115t2183) I(R3117t2808) I(R3117t3083) I(R3117t1267) I(R3117t76) I(R3117t976) I(R3117t1392) I(R3118t643) I(R3118t2966) I(R3119t485) I(R3119t2672) I(R3119t269) I(R3120t879) I(R3120t2909) I(R3120t543) I(R3120t418) I(R3120t390) I(R3122t3035) I(R3123t224) I(R3123t2269) I(R3123t1402) I(R3124t66) I(R3124t860) I(R3124t386) I(R3124t2724) I(R3124t2027) I(R3125t2324) I(R3125t2429) I(R3125t296) I(R3126t2431) I(R3127t2630) I(R3128t2172) I(R3128t1051) I(R3129t2609) I(R3130t356) I(R3130t1917) I(R3130t2485) I(R3131t2405) I(R3131t194) I(R3132t2963) I(R3132t2912) I(R3133t2561) I(R3133t1259) I(R3134t283) I(R3134t1695) I(R3134t2990) I(R3135t1797) I(R3136t604) I(R3137t1911) I(R3137t37) I(R3138t2435) I(R3138t1040) I(R3139t3061) I(R3140t2313) I(R3140t1888) I(R3140t455) I(R3141t929) I(R3141t1986) I(R3142t2204) I(R3143t2017) I(R3143t1428) I(R3145t3128) I(R3145t2172) I(R3146t1041) I(R3146t2868) I(R3147t1054) I(R3148t333) I(R3148t1066) I(R3149t1113) I(R3150t480) I(R3150t82) I(R3151t2752) I(R3152t274) I(R3152t371) I(R3152t2740) I(R3153t230) I(R3153t204) I(R3155t2976) I(R3155t1378) I(R3156t231) I(R3156t2356) I(R3157t3142) I(R3158t515) I(R3158t2520) I(R3158t624) I(R3160t1157) I(R3160t672) I(R3161t1032) I(R3162t471) I(R3162t2144) I(R3163t1672) I(R3163t2271) I(R3164t3088) I(R3164t2681) I(R3164t360) I(R3164t85) I(R3165t1026) I(R3165t226) I(R3165t1008) I(R3167t1356) I(R3167t690) I(R3169t365) I(R3169t2141) I(R3170t2115) I(R3170t2583) I(R3170t1508) I(R3171t2614) I(R3171t1) I(R3172t1507) I(R3174t2023) I(R3174t2256) I(R3174t342) I(R3175t1537) I(R3175t3008) I(R3175t1602) I(R3176t2504) I(R3177t85) I(R3177t3164) I(R3177t534) I(R3177t185) I(R3177t360) I(R3178t754) I(R3179t2572) I(R3179t586) I(R3179t2749) I(R3180t624) I(R3180t2520) I(R3181t484) I(R3181t1682) I(R3181t2237) I(R3181t161) I(R3181t2960) I(R3182t248) I(R3182t2736) I(R3183t2317) I(R3184t447) I(R3184t1121) I(R3185t2243) I(R3186t2058) I(R3186t2166) I(R3187t941) I(R3187t1550) I(R3187t1940) I(R3187t1025) I(R3189t300) I(R3189t1435) I(R3190t2898) I(R3191t2780) I(R3192t992) I(R3193t1422) I(R3194t1162) I(R3197t2049) I(R3198t87) I(R3199t1514) I(R3200t3104) I(R3200t2312) I(R3200t3013) I(R3201t663) I(R3201t1135) I(R3203t3196) I(R3203t2369) I(R3204t227) I(R3204t649) I(R3204t2067) I(R3205t1534) I(R3205t561) I(R3206t1994) I(R3206t1175) I(R3207t1588) I(R3207t1007) I(R3208t1098) I(R3208t3030) I(R3208t819) I(R3208t1332) I(R3209t460) I(R3209t2500) I(R3210t2220) I(R3211t1800) I(R3212t336) I(R3213t2807) I(R3214t1412) I(R3214t855) I(R3214t1294) I(R3214t1221) I(R3215t1789) I(R3216t1836) I(R3216t998) I(R3216t456) I(R3216t1970) I(R3217t2330) I(R3218t1323) I(R3218t2340) I(R3218t1479) I(R3218t2295) I(R3219t54) I(R3219t161) I(R3219t3181) I(R3219t2237) I(R3220t737) I(R3220t1725) I(R3220t404) I(R3221t1128) I(R3221t390) I(R3221t2521) I(R3222t1435) I(R3222t3026) I(R3224t1092) I(R3224t1331) I(R3224t1144) I(R3225t1924) I(R3226t56) I(R3226t1964) I(R3229t1951) I(R3229t218) I(R3229t2084) I(R3231t3144) I(R3232t2598) I(R3232t1787) I(R3233t1750) I(R3233t1441) I(R3233t1427) I(R3233t2695) I(R3235t1366) I(R3235t1181) I(R3235t1020) I(R3235t741) I(R3236t106) I(R3236t1727) I(R3237t3212) I(R3237t336) I(R3237t702) I(R3238t1553) I(R3238t286) I(R3239t573) I(R3240t1258) I(R3240t1716) I(R3240t2879) I(R3241t3063) I(R3242t2155) I(R3243t431) I(R3243t3015) I(R3244t1093) I(R3244t1954) I(R3244t1484) I(R3245t1665) I(R3245t3037) I(R3245t1872) I(R3247t668) I(R3247t1593) I(R3247t1490) I(R3248t1363) I(R3249t2503) I(R3249t2195) I(R3249t1061) I(R3250t1073) I(R3250t2404) I(R3251t1972) I(R3251t2766) I(R3252t290) I(R3252t1164) I(R3252t1340) I(R3254t3251) I(R3254t901) I(R3254t750) I(R3254t2568) I(R3254t2539) I(R3255t1122) I(R3255t2977) I(R3255t1204) I(R3256t392) I(R3256t883) I(R3256t1815) I(R3257t1152) I(R3258t2505) I(R3259t86) I(R3259t2984) I(R3260t2604) I(R3260t1627) I(R3260t1673) I(R3261t1512) I(R3262t3040) I(R3262t2586) I(R3263t387) I(R3263t2348) I(R3263t2611) I(R3263t1878) I(R3264t2075) I(R3264t2140) I(R3264t2211) I(R3265t3078) I(R3265t2917) I(R3266t2952) I(R3266t1867) I(R3267t1416) I(R3267t1797) I(R3267t3135) I(R3269t2051) I(R3270t1624) I(R3270t1863) I(R3270t347) I(R3271t614) I(R3271t1279) I(R3271t791) I(R3271t2408) I(R3272t1009) I(R3272t3050) I(R3274t1332) I(R3275t2160) I(R3275t2088) I(R3275t105) I(R3276t2019) I(R3276t1664) I(R3277t2892) I(R3279t928) I(R3280t3121) I(R3281t3231) I(R3281t3144) I(R3281t546) I(R3282t1778) I(R3282t2493) I(R3282t2968) I(R3282t937) I(R3283t2846) I(R3284t1974) I(R3284t3021) I(R3284t2172) I(R3285t1862) I(R3285t689) I(R3286t605) I(R3286t2596) I(R3286t2102) I(R3286t2453) I(R3287t2651) I(R3287t1665) I(R3287t3245) I(R3288t1611) I(R3288t2327) I(R3288t2495) I(R3290t966) I(R3291t61) I(R3293t1236) I(R3293t3288) I(R3293t2495) I(R3294t2044) I(R3294t309) I(R3294t1771) I(R3295t2716) I(R3295t1860) I(R3295t1585) I(R3296t1734) I(R3297t2844) I(R3299t931) I(R3299t2758) I(R3299t2819) I(R3300t357) I(R3300t1431) I(R3300t1353) I(R3301t660) I(R3301t1567) I(R3301t1056) I(R3303t3260) I(R3303t1082) I(R3304t545) I(R3304t138) I(R3304t2694) I(R3305t530) I(R3306t2100) I(R3306t154) I(R3307t863) I(R3307t1130) I(R3309t2336) I(R3310t2512) I(R3310t94) I(R3310t2578) I(R3310t1243) I(R3311t1788) I(R3312t585) I(R3313t2309) I(R3313t1554) I(R3314t1438) I(R3314t1142) I(R3315t3003) I(R3316t3205) I(R3317t675) I(R3317t112) I(R3317t41) I(R3317t714) I(R3318t2504) I(R3318t519) I(R3319t1362) I(R3319t2794) I(R3320t1755) I(R3321t859) I(R3321t1722) I(R3321t1503) I(R3322t1077) I(R3322t547) I(R3322t1467) I(R3322t1002) I(R3323t1565) I(R3324t112) I(R3325t1552) I(R3325t398) I(R3325t987) I(R3326t2565) I(R3326t1425) I(R3327t1939) I(R3327t1547) I(R3328t887) I(R3329t1835) I(R3330t3143) I(R3330t268) I(R3331t1171) I(R3332t1258) I(R3332t2879) I(R3332t1622) I(R3332t124) I(R3333t729) I(R3333t2746) I(R3333t252) I(R3334t1565) I(R3334t3323) I(R3335t2376) I(R3336t1360) I(R3336t1480) I(R3336t2929) I(R3337t1177) I(R3337t67) I(R3338t2428) I(R3338t1880) I(R3339t1696) I(R3339t2212) I(R3340t2814) I(R3340t2316) I(R3341t426) I(R3341t1047) I(R3342t323) I(R3343t350) I(R3343t2045) I(R3344t1146) I(R3344t1875) I(R3344t2261) I(R3345t1825) I(R3345t461) I(R3346t1297) I(R3346t2462) I(R3346t679) I(R3347t2441) I(R3347t2478) I(R3347t334) I(R3347t1166) I(R3348t2321) I(R3348t2444) I(R3349t2245) I(R3349t645) I(R3349t2667) I(R3350t1191) I(R3351t1264) I(R3353t1881) I(R3353t1615) I(R3353t1799) I(R3353t1368) I(R3354t513) I(R3354t2137) I(R3355t1347) I(R3355t2207) I(R3356t106) I(R3356t2738) I(R3356t1727) I(R3357t1832) I(R3357t313) I(R3358t3137) I(R3358t37) I(R3358t1402) I(R3359t2206) I(R3359t1014) I(R3360t1055) I(R3361t2548) I(R3361t53) I(R3361t1544) I(R3361t2712) I(R3362t2249) I(R3362t2466) I(R3363t1936) I(R3364t3087) I(R3364t982) I(R3364t921) I(R3365t2172) I(R3365t3284) I(R3366t1275) I(R3366t1827) I(R3367t1824) I(R3367t2315) I(R3367t2094) I(R3368t634) I(R3368t2700) I(R3369t825) I(R3369t853) I(R3370t422) I(R3370t1884) I(R3370t2503) I(R3371t1470) I(R3371t3278) I(R3371t16) I(R3372t618) I(R3372t2014) I(R3373t2210) I(R3373t3036) I(R3373t2680) I(R3374t3276) I(R3374t2779) I(R3375t86) I(R3375t3259) I(R3376t2945) I(R3376t1256) I(R3377t1913) I(R3377t2149) I(R3378t1730) I(R3378t794) I(R3379t190) I(R3382t187) I(R3382t2590) I(R3383t2852) I(R3383t420) I(R3383t1850) I(R3384t1175) I(R3384t2259) I(R3384t3206) I(R3385t1923) I(R3386t204) I(R3386t3153) I(R3386t478) I(R3388t1956) I(R3388t221) I(R3389t1639) I(R3390t3251) I(R3391t1406) I(R3391t1473) I(R3392t1686) I(R3392t1566) I(R3394t1379) I(R3394t2576) I(R3396t1692) I(R3396t2765) I(R3396t1775) I(R3397t2617) I(R3397t977) I(R3398t886) I(R3399t2542) I(R3399t2572) I(R3399t3179) I(R3399t195) I(R3400t669) I(R3400t2359) I(R3400t294) I(R3400t1905) I(R3401t2331) I(R3401t964) I(R3402t406) I(R3402t91) I(R3402t1883) I(R3403t1921) I(R3404t234) I(R3404t1603) I(R3404t2133) I(R3405t1782) I(R3405t3054) I(R3406t1440) I(R3406t2583) I(R3407t599) I(R3407t1254) I(R3408t1844) I(R3408t222) I(R3409t1463) I(R3410t3064) I(R3410t2867) I(R3411t1890) I(R3411t2923) I(R3411t808) I(R3412t1378) I(R3413t2049) I(R3413t1190) I(R3413t1197) I(R3413t3197) I(R3414t939) I(R3414t1230) I(R3415t1407) I(R3415t1081) I(R3416t89) I(R3416t1648) I(R3416t1096) I(R3417t3190) I(R3417t2403) I(R3418t628) I(R3418t2412) I(R3418t2461) I(R3419t469) I(R3419t1594) I(R3420t1190) I(R3420t1197) I(R3421t2600) I(R3421t1541) I(R3422t1280) I(R3422t2593) I(R3422t2837) I(R3423t592) I(R3423t2930) I(R3423t908) I(R3423t838) I(R3424t658) I(R3425t1959) I(R3425t1001) I(R3426t3305) I(R3426t2294) I(R3427t1857) I(R3427t945) I(R3428t695) I(R3428t912) I(R3429t891) I(R3429t2882) I(R3430t284) I(R3430t864) I(R3431t2587) I(R3432t3260) I(R3432t3303) I(R3433t1601) I(R3434t318) I(R3434t2300) I(R3434t2623) I(R3435t2387) I(R3435t2356) I(R3435t3156) I(R3436t2284) I(R3436t340) I(R3436t1453) I(R3436t935) I(R3436t2858) I(R3437t888) I(R3438t2731) I(R3438t2342) I(R3438t1342) I(R3439t2340) I(R3439t2374) I(R3439t341) I(R3440t1036) I(R3440t789) I(R3440t1024) I(R3441t2630) I(R3441t3127) I(R3443t995) I(R3443t29) I(R3443t3166) I(R3444t1336) I(R3444t1589) I(R3444t2303) I(R3444t2021) I(R3445t3178) I(R3445t2805) I(R3447t1595) I(R3447t1091) I(R3448t2648) I(R3448t1851) I(R3451t2249) I(R3451t3362) I(R3452t932) I(R3454t2287) I(R3455t3366) I(R3455t1708) I(R3455t1827) I(R3456t1872) I(R3457t536) I(R3457t2951) I(R3458t564) I(R3458t2717) I(R3459t1540) I(R3460t3116) I(R3461t2788) I(R3461t432) I(R3461t2440) I(R3462t93) I(R3463t175) I(R3464t2012) I(R3465t509) I(R3465t2713) I(R3465t1683) I(R3466t3346) I(R3466t127) I(R3466t679) I(R3467t2466) I(R3468t1911) I(R3469t222) I(R3470t1618) I(R3470t2494) I(R3470t1105) I(R3471t2312) I(R3471t34) I(R3472t3454) I(R3473t348) I(R3474t214) I(R3474t329) I(R3475t924) I(R3475t2496) I(R3476t2734) I(R3477t2728) I(R3477t312) I(R3478t477) I(R3478t2018) I(R3479t2628) I(R3479t1096) I(R3480t1765) I(R3480t2167) I(R3480t1806) I(R3480t2874) I(R3481t553) I(R3481t3277) I(R3482t2836) I(R3482t1661) I(R3482t1597) I(R3483t2741) I(R3483t1898) I(R3483t2314) I(R3484t1400) I(R3484t661) I(R3484t1976) I(R3487t63) I(R3487t758) I(R3488t980) I(R3488t1074) I(R3488t616) I(R3488t2413) I(R3489t2725) I(R3489t389) I(R3489t347) I(R3490t7) I(R3490t501) I(R3490t3050) I(R3491t603) I(R3492t2838) I(R3493t2267) I(R3493t1516) I(R3494t1715) I(R3495t1331) I(R3495t2077) I(R3496t1294) I(R3496t1221) I(R3497t981) I(R3497t2378) I(R3497t2749) I(R3498t138) I(R3498t545) I(R3498t3304) I(R3499t1693) I(R3500t222) I(R3500t2273) I(R3500t2867) I(R3501t846) I(R3501t2732) I(R3501t533) I(R3502t3050) I(R3502t1510) I(R3503t1584) I(R3503t1586) I(R3504t2714) I(R3504t1901) I(R3506t1283) I(R3506t523) I(R3506t2320) I(R3506t916) I(R3507t1533) I(R3507t1023) I(R3508t1326) I(R3508t1830) I(R3509t3494) I(R3509t1715) I(R3510t591) I(R3510t1156) I(R3510t3351) I(R3512t3359) I(R3513t3448) I(R3513t1851) I(R3514t944) I(R3515t320) I(R3515t144) I(R3516t3282) I(R3516t2493) I(R3517t621) I(R3517t1984) I(R3517t2006) I(R3518t3515) I(R3519t1415) I(R3519t204) I(R3520t1595) I(R3520t3447) I(R3520t1091) I(R3520t698) I(R3521t216) I(R3521t2602) I(R3522t1493) I(R3523t250) I(R3523t448) I(R3523t1523) I(R3524t3383) I(R3524t1850) I(R3524t246) I(R3525t3163) I(R3525t2271) I(R3526t3246) I(R3527t2664) I(R3527t96) I(R3527t2796) I(R3527t155) I(R3528t680) I(R3528t528) I(R3528t70) I(R3528t2054) I(R3528t105) I(R3528t3275) I(R3529t1266) I(R3529t3215) I(R3529t597) I(R3530t1804) I(R3531t2220) I(R3531t570) I(R3532t1966) I(R3533t2288) I(R3533t237) I(R3534t818) I(R3534t1339) I(R3535t370) I(R3535t883) I(R3535t2354) I(R3536t2154) I(R3536t560) I(R3537t442) I(R3537t495) I(R3538t2346) I(R3538t651) I(R3538t1926) I(R3538t636) I(R3538t436) I(R3539t677) I(R3540t1224) I(R3540t2108) I(R3540t433) I(R3540t507) I(R3541t1398) I(R3541t2893) I(R3542t2123) I(R3542t987) I(R3543t86) I(R3544t1263) I(R3545t17) I(R3545t649) I(R3545t884) I(R3545t1171) I(R3546t416) I(R3547t1613) I(R3547t604) I(R3549t3122) I(R3549t3035) I(R3549t2732) I(R3549t1553) I(R3550t912) I(R3551t1234) I(R3551t3073) I(R3552t3) I(R3552t3244) I(R3552t1484) I(R3552t1383) I(R3553t279) I(R3553t2354) I(R3554t1466) I(R3554t3015) I(R3555t358) I(R3555t2911) I(R3556t299) I(R3556t2908) I(R3556t1956) I(R3556t221) I(R3556t942) I(R3558t170) I(R3558t1153) I(R3558t1758) I(R3558t1414) I(R3559t3541) I(R3559t2893) I(R3560t219) I(R3560t3526) I(R3560t3000) I(R3561t1538) I(R3561t2421) I(R3562t118) I(R3563t757) I(R3563t900) I(R3563t939) I(R3564t3087) I(R3565t1628) I(R3566t1206) I(R3566t2469) I(R3566t1662) I(R3566t2577) I(R3566t1473) I(R3567t296) I(R3568t2252) I(R3569t2385) I(R3569t457) I(R3570t565) I(R3570t192) I(R3571t1215) I(R3571t2896) I(R3573t592) I(R3573t3423) I(R3573t55) I(R3574t3335) I(R3574t1684) I(R3574t2376) I(R3575t1798) I(R3576t2482) I(R3577t811) I(R3578t1961) I(R3578t1233) I(R3578t3033) I(R3579t392) I(R3579t1815) I(R3579t3256) I(R3580t1650) I(R3580t1) I(R3580t3171) I(R3580t1252) I(R3581t3071) I(R3581t597) I(R3582t619) I(R3582t581) I(R3583t1891) I(R3583t17) I(R3584t1216) I(R3584t543) I(R3584t354) I(R3585t2600) I(R3585t569) I(R3586t2647) I(R3586t2686) I(R3586t873) I(R3587t1506) I(R3587t2485) I(R3587t3130) I(R3588t2223) I(R3588t380) I(R3589t263) I(R3589t2534) I(R3589t1901) I(R3590t2419) I(R3590t1367) I(R3590t3079) I(R3591t1114) I(R3591t1108) I(R3592t529) I(R3592t2711) I(R3592t242) I(R3593t542) I(R3593t2816) I(R3593t690) I(R3594t3530) I(R3594t544) I(R3595t3093) I(R3595t2298) I(R3596t2508) I(R3596t1170) I(R3597t2988) I(R3597t300) I(R3598t203) I(R3598t1932) I(R3598t721) I(R3599t2272) I(R3600t2818) I(R3600t2234) I(R3600t2130) I(R3600t1570) I(R3601t1606) I(R3601t1244) I(R3601t1000) I(R3602t1853) I(R3602t793) I(R3602t459) I(R3602t876) I(R3603t654) I(R3603t2129) I(R3603t1571) I(R3604t2033) I(R3605t2316) I(R3605t3340) I(R3605t1123) I(R3605t1566) I(R3606t3557) I(R3606t3009) I(R3607t1914) I(R3608t3095) I(R3608t1078) I(R3609t291) I(R3609t828) I(R3610t2212) I(R3610t2566) I(R3611t399) I(R3611t1136) I(R3611t1907) I(R3612t894) I(R3613t827) I(R3614t643) I(R3614t1812) I(R3614t2881) I(R3614t2966) I(R3615t2721) I(R3615t1747) I(R3616t388) I(R3616t3060) I(R3617t3475) I(R3617t924) I(R3618t3608) I(R3619t630) I(R3619t1007) I(R3620t2547) I(R3620t1646) I(R3621t697) I(R3622t1755) I(R3622t3320) I(R3622t2363) I(R3622t702) I(R3624t2624) I(R3625t3613) I(R3625t827) I(R3626t443) I(R3626t3174) I(R3627t735) I(R3627t2022) I(R3628t3512) I(R3628t3359) I(R3629t1452) I(R3629t3062) I(R3631t2366) I(R3632t874) I(R3633t2945) I(R3634t2321) I(R3634t1812) I(R3634t3348) I(R3635t2970) I(R3635t1569) I(R3635t837) I(R3636t2637) I(R3637t3100) I(R3637t229) I(R3637t2895) I(R3638t262) I(R3638t2738) I(R3639t2981) I(R3639t3068) I(R3640t634) I(R3640t3034) I(R3640t3368) I(R3640t2477) I(R3641t1687) I(R3641t3105) I(R3641t866) I(R3642t2664) I(R3642t260) I(R3642t890) I(R3642t155) I(R3642t3527) I(R3643t429) I(R3643t1457) I(R3643t800) I(R3644t274) I(R3644t409) I(R3644t2365) I(R3645t291) I(R3645t259) I(R3645t1356) I(R3646t191) I(R3647t3119) I(R3647t332) I(R3647t485) I(R3648t2073) I(R3648t1886) I(R3649t2015) I(R3650t2260) I(R3650t1851) I(R3650t3513) I(R3650t739) I(R3651t3234) I(R3652t2188) I(R3653t2659) I(R3653t2706) I(R3654t870) I(R3654t3327) I(R3655t1272) I(R3655t2754) I(R3655t2163) I(R3655t674) I(R3658t458) I(R3658t1927) I(R3658t2558) I(R3659t2290) I(R3660t3468) I(R3661t370) I(R3662t2746) I(R3662t359) I(R3663t1549) I(R3663t2957) I(R3663t567) I(R3663t640) I(R3664t602) I(R3664t3117) I(R3664t1392) I(R3664t1591) I(R3664t1610) I(R3665t96) I(R3665t2796) I(R3666t3496) I(R3666t1294) I(R3666t2028) I(R3667t1182) I(R3668t2946) I(R3669t3128) I(R3669t3365) I(R3670t3516) I(R3670t680) I(R3670t2393) I(R3670t2968) I(R3670t3282) I(R3671t945) I(R3671t3427) I(R3672t108) I(R3673t917) I(R3673t789) I(R3674t1652) I(R3674t2847) I(R3674t1439) I(R3674t1337) I(R3675t109) I(R3676t3228) I(R3676t1198) I(R3677t2241) I(R3677t1329) I(R3677t2253) I(R3678t271) I(R3678t730) I(R3678t1374) I(R3678t1311) I(R3679t2113) I(R3680t1463) I(R3681t1110) I(R3681t756) I(R3682t2296) I(R3683t2563) I(R3683t1185) I(R3684t3016) I(R3684t260) I(R3685t2037) I(R3685t3042) I(R3686t3007) I(R3686t1251) I(R3686t3063) I(R3687t2197) I(R3687t3577) I(R3688t1809) I(R3688t2465) I(R3688t2519) I(R3689t770) I(R3689t1419) I(R3689t1626) I(R3690t142) I(R3691t413) I(R3691t1573) I(R3692t1981) I(R3692t3136) I(R3692t604) I(R3692t3547) I(R3692t1613) I(R3693t107) I(R3693t2627) I(R3693t1870) I(R3694t1010) I(R3695t494) I(R3695t3070) I(R3695t778) I(R3695t126) I(R3696t1952) I(R3696t3387) I(R3697t2442) I(R3697t2876) I(R3698t2992) I(R3699t804) I(R3699t1253) I(R3700t2027) I(R3701t3077) I(R3703t1032) I(R3703t1514) I(R3703t2416) I(R3704t721) I(R3704t3598) I(R3705t546) I(R3705t2423) I(R3705t1225) I(R3706t3304) I(R3706t633) I(R3707t3575) I(R3707t1423) I(R3708t2977) I(R3708t2308) I(R3708t1465) I(R3708t682) I(R3709t2991) I(R3709t2443) I(R3710t3054) I(R3711t980) I(R3711t993) I(R3711t2413) I(R3711t3488) I(R3712t1949) I(R3713t2599) I(R3714t3212) I(R3714t336) I(R3714t2127) I(R3714t1817) I(R3714t2186) I(R3715t1407) I(R3715t3607) I(R3715t2383) I(R3715t1313) I(R3716t275) I(R3716t1405) I(R3716t600) I(R3716t1768) I(R3717t3661) I(R3717t2944) I(R3717t2848) I(R3718t2760) I(R3719t2513) I(R3719t3648) I(R3720t1824) I(R3720t2315) I(R3721t2317) I(R3721t2695) I(R3722t924) I(R3722t3617) I(R3722t3186) I(R3723t1408) I(R3723t3668) I(R3723t2946) I(R3724t1265) I(R3724t801) I(R3725t658) I(R3725t1790) I(R3726t3718) I(R3726t1796) I(R3726t2337) I(R3727t1384) I(R3727t2085) I(R3728t3166) I(R3728t3443) I(R3728t995) I(R3728t461) I(R3729t250) I(R3729t3523) I(R3729t1523) I(R3730t2243) I(R3730t3185) I(R3730t1026) I(R3730t3065) I(R3732t752) I(R3733t1512) I(R3733t2396) I(R3733t973) I(R3733t324) I(R3733t3058) I(R3733t422) I(R3733t1012) I(R3734t114) I(R3734t346) I(R3734t261) I(R3734t1535) I(R3734t1817) I(R3734t918) I(R3735t2067) I(R3735t771) I(R3736t1157) I(R3736t3160) I(R3736t2113) I(R3737t1637) I(R3737t1381) I(R3738t1822) I(R3738t2710) I(R3738t1917) I(R3738t1384) I(R3739t1671) I(R3739t3453) I(R3740t765) I(R3740t140) I(R3740t2493) I(R3741t1816) I(R3741t1697) I(R3741t1220) I(R3741t559) I(R3741t950) I(R3742t2841) I(R3742t2144) I(R3743t1020) I(R3743t2134) I(R3743t2559) I(R3744t626) I(R3744t3574) I(R3745t2013) I(R3745t3080) I(R3745t2762) I(R3746t1138) I(R3747t686) I(R3747t745) I(R3747t548) I(R3747t2473) I(R3748t846) I(R3748t2495) I(R3748t239) I(R3748t533) I(R3748t3501) I(R3749t2787) I(R3750t3012) I(R3750t1491) I(R3750t2648) I(R3751t1718) I(R3751t2562) I(R3752t1246) I(R3752t847) I(R3753t1067) I(R3754t3172) I(R3755t1414) I(R3755t3558) I(R3756t1699) I(R3756t2515) I(R3756t714) I(R3756t41) I(R3757t1069) I(R3757t1530) I(R3757t2448) I(R3757t787) I(R3758t2677) I(R3758t1575) I(R3758t3095) I(R3758t3608) I(R3759t1825) I(R3759t3345) I(R3759t461) I(R3759t475) I(R3759t362) I(R3760t2073) I(R3760t3648) I(R3761t2165) I(R3761t3046) I(R3762t146) I(R3762t2106) I(R3762t3175) I(R3763t1984) I(R3763t2352) I(R3763t563) I(R3764t1737) I(R3765t2718) I(R3765t556) I(R3766t1459) I(R3767t1212) I(R3767t2870) I(R3767t2142) I(R3767t1760) I(R3769t2886) I(R3769t1745) I(R3770t1284) I(R3770t2297) I(R3770t1880) I(R3771t2045) I(R3771t871) I(R3771t2616) I(R3772t2731) I(R3773t1973) I(R3774t3451) I(R3774t2249) I(R3774t1672) I(R3774t3163) I(R3775t2274) I(R3775t2230) I(R3776t3695) I(R3776t778) I(R3776t3067) I(R3776t427) I(R3777t332) I(R3777t829) I(R3779t1124) I(R3779t1174) I(R3779t3107) I(R3779t232) I(R3779t1580) I(R3780t1083) I(R3780t1791) I(R3780t1343) I(R3780t1607) I(R3781t2884) I(R3781t1559) I(R3782t1255) I(R3783t109) I(R3783t2423) I(R3783t546) I(R3784t1314) I(R3784t2967) I(R3785t737) I(R3785t1725) I(R3785t82) I(R3785t583) I(R3786t2831) I(R3786t2326) I(R3786t337) I(R3786t3493) I(R3787t743) I(R3787t2615) I(R3787t198) I(R3788t535) I(R3788t3419) I(R3788t1594) I(R3788t2912) I(R3788t759) I(R3789t376) I(R3789t1920) I(R3790t2196) I(R3791t2836) I(R3791t3482) I(R3791t1597) I(R3791t69) I(R3791t194) I(R3791t3131) I(R3793t1909) I(R3794t122) I(R3795t1379) I(R3796t1271) I(R3796t1650) I(R3797t1572) I(R3797t1881) I(R3797t3731) I(R3798t300) I(R3798t3597) I(R3798t1642) I(R3798t328) I(R3798t752) I(R3798t3732) I(R3798t3189) I(R3799t3069) I(R3799t1030) I(R3799t3724) I(R3800t2925) I(R3801t464) I(R3801t1217) I(R3802t2988) I(R3802t8) I(R3803t2105) I(R3803t3175) I(R3803t3762) I(R3803t2106) I(R3804t3511) I(R3804t1157) I(R3804t3794) I(R3805t543) I(R3805t418) I(R3806t2094) I(R3806t1373) I(R3807t1850) I(R3807t2344) I(R3807t1449) I(R3808t1955) I(R3808t1049) I(R3808t2221) I(R3809t74) I(R3809t1584) I(R3809t3503) I(R3810t1693) I(R3810t3499) I(R3811t1450) I(R3811t1092) I(R3812t688) I(R3812t813) I(R3813t3619) I(R3813t3807) I(R3813t1997) I(R3814t1204) I(R3814t1678) I(R3814t3255) I(R3815t3761) I(R3816t2285) I(R3816t2482) I(R3816t3576) I(R3817t2277) I(R3817t2014) I(R3818t1139) I(R3819t2964) I(R3820t520) I(R3820t566) I(R3821t3075) I(R3821t3291) I(R3821t61) I(R3821t91) I(R3822t129) I(R3822t465) I(R3823t2339) I(R3823t99) I(R3824t1184) I(R3824t3818) I(R3824t1307) I(R3825t2130) I(R3826t2235) I(R3826t1907) I(R3827t748) I(R3828t339) I(R3828t1834) I(R3828t455) I(R3828t1888) I(R3829t2334) I(R3829t1713) I(R3829t1401) I(R3829t1968) I(R3830t464) I(R3830t1819) I(R3831t701) I(R3832t313) I(R3833t2342) I(R3834t1900) I(R3834t2265) I(R3834t581) I(R3835t1150) I(R3835t2934) I(R3835t723) I(R3836t2499) I(R3836t348) I(R3836t3473) I(R3837t818) I(R3838t3272) I(R3838t3050) I(R3838t3490) I(R3839t650) I(R3839t2039) I(R3840t577) I(R3840t1989) I(R3840t2194) I(R3840t2997) I(R3840t3041) I(R3841t1191) I(R3841t3350) I(R3841t2599) I(R3841t2762) I(R3841t820) I(R3842t710) I(R3842t3044) I(R3842t2159) I(R3843t539) I(R3843t1842) I(R3844t3030) I(R3844t1029) I(R3844t1925) I(R3845t1908) I(R3846t852) I(R3846t2613) I(R3846t2258) I(R3847t3452) I(R3848t1131) I(R3848t2836) I(R3848t3482) I(R3848t1661) I(R3848t3112) I(R3848t2652) I(R3849t2683) I(R3850t740) I(R3850t2008) I(R3851t2143) I(R3851t65) I(R3853t3094) I(R3853t907) I(R3853t3698) I(R3854t2604) I(R3854t1931) I(R3854t2744) I(R3855t2972) I(R3855t3466) I(R3856t467) I(R3856t1198) I(R3857t1245) I(R3858t1077) I(R3858t3322) I(R3859t3076) I(R3859t104) I(R3859t1291) I(R3860t1713) I(R3860t1814) I(R3860t2975) I(R3861t3141) I(R3861t1574) I(R3861t835) I(R3863t1327) I(R3863t2992) I(R3864t687) I(R3865t896) I(R3865t460) I(R3865t823) I(R3866t2057) I(R3866t254) I(R3867t1840) I(R3868t32) I(R3868t3093) I(R3868t3595) I(R3869t2872) I(R3869t2568) I(R3869t1846) I(R3870t36) I(R3871t1098) I(R3871t3208) I(R3871t3030) I(R3871t2125) I(R3872t1539) I(R3873t121) I(R3873t2784) I(R3873t2158) I(R3874t1776) I(R3874t1925) I(R3875t1349) I(R3875t2874) I(R3875t258) I(R3876t125) I(R3877t2172) I(R3879t1891) I(R3879t2557) I(R3879t2535) I(R3879t822) I(R3879t17) I(R3879t3583) I(R3880t1147) I(R3880t2483) I(R3881t406) I(R3881t473) I(R3881t1133) I(R3881t2487) I(R3882t2833) I(R3882t3633) I(R3883t2823) I(R3883t466) I(R3884t3431) I(R3884t2386) I(R3885t1806) I(R3885t1247) I(R3886t97) I(R3886t3618) I(R3888t1046) I(R3890t2595) I(R3891t1797) I(R3891t1519) I(R3891t631) I(R3892t3396) I(R3892t43) I(R3892t1524) I(R3893t2333) I(R3893t2576) I(R3894t1211) I(R3894t1677) I(R3894t1548) I(R3895t2331) I(R3895t108) I(R3895t1836) I(R3895t964) I(R3896t658) I(R3896t454) I(R3896t3852) I(R3897t88) I(R3897t1476) I(R3898t552) I(R3898t2763) I(R3898t1924) I(R3898t3225) I(R3899t3103) I(R3899t1830) I(R3899t1077) I(R3900t60) I(R3900t2258) I(R3900t3397) I(R3901t1983) I(R3901t1487) I(R3902t1240) I(R3902t2821) I(R3903t955) I(R3903t1837) I(R3904t920) I(R3904t2145) I(R3905t1960) I(R3905t2138) I(R3905t716) I(R3906t464) I(R3906t3830) I(R3906t2755) I(R3906t1819) I(R3907t2478) I(R3907t3347) I(R3907t2917) I(R3908t836) I(R3909t3203) I(R3910t2273) I(R3910t851) I(R3911t287) I(R3911t2547) I(R3911t2178) I(R3912t1922) I(R3912t1813) I(R3913t1707) I(R3913t3908) I(R3914t3152) I(R3915t31) I(R3915t2617) I(R3915t2098) I(R3916t698) I(R3916t1091) I(R3916t497) I(R3916t1847) I(R3916t1628) I(R3916t1094) I(R3917t2941) I(R3917t1146) I(R3917t1760) I(R3917t3767) I(R3918t542) I(R3919t3514) I(R3919t1880) I(R3920t1803) I(R3920t1716) I(R3922t1711) I(R3922t672) I(R3923t3632) I(R3923t874) I(R3924t2964) I(R3924t3819) I(R3924t2522) I(R3925t2887) I(R3925t2527) I(R3925t1511) I(R3926t3897) I(R3926t1476) I(R3927t895) I(R3928t1375) I(R3928t3656) I(R3929t710) I(R3929t3842) I(R3929t2159) I(R3929t2733) I(R3930t3443) I(R3930t29) I(R3930t811) I(R3931t806) I(R3931t756) I(R3931t3681) I(R3932t401) I(R3932t2719) I(R3933t1240) I(R3933t3902) I(R3934t1582) I(R3936t2562) I(R3937t2146) I(R3937t2218) I(R3937t2797) I(R3937t913) I(R3938t1088) I(R3939t646) I(R3939t1916) I(R3939t3686) I(R3939t1251) I(R3940t1875) I(R3940t2261) I(R3941t562) I(R3941t3173) I(R3942t1783) I(R3942t165) I(R3943t3900) I(R3943t60) I(R3943t1353) I(R3943t920) I(R3944t661) I(R3944t798) I(R3945t3530) I(R3945t3051) I(R3945t2639) I(R3946t2895) I(R3946t826) I(R3947t2154) I(R3948t2358) I(R3948t2764) I(R3949t3191) I(R3949t2780) I(R3949t2844) I(R3950t612) I(R3952t459) I(R3952t2701) I(R3952t1649) I(R3952t788) I(R3952t2231) I(R3953t3652) I(R3953t3195) I(R3954t2659) I(R3954t3653) I(R3954t1569) I(R3954t2706) I(R3955t2228) I(R3955t1111) I(R3956t1811) I(R3956t1443) I(R3957t348) I(R3958t132) I(R3959t1328) I(R3959t2022) I(R3959t3105) I(R3959t3641) I(R3960t198) I(R3961t2268) I(R3962t965) I(R3963t1454) I(R3963t1067) I(R3963t396) I(R3963t293) I(R3964t705) I(R3964t2216) I(R3965t1130) I(R3965t2338) I(R3965t3307) I(R3965t863) I(R3966t1354) I(R3966t1420) I(R3966t1244) I(R3967t2162) I(R3967t2160) I(R3967t3275) I(R3967t2088) I(R3969t900) I(R3969t3599) I(R3970t3274) I(R3971t720) I(R3971t1549) I(R3971t567) I(R3971t2957) I(R3972t2156) I(R3972t255) I(R3972t2608) I(R3973t1477) I(R3973t1001) I(R3973t3425) I(R3974t2815) I(R3975t3915) I(R3975t31) I(R3975t2613) I(R3975t3846) I(R3976t512) I(R3977t538) I(R3978t49) I(R3978t443) I(R3979t1020) I(R3979t3235) I(R3980t3175) I(R3980t1602) I(R3981t517) I(R3982t3749) I(R3983t2544) I(R3983t2781) I(R3983t1626) I(R3983t1708) I(R3984t489) I(R3984t2524) I(R3984t109) I(R3984t3783) I(R3984t92) I(R3985t773) I(R3985t961) I(R3985t732) I(R3986t140) I(R3987t1761) I(R3988t2309) I(R3988t3313) I(R3988t2032) I(R3989t3236) I(R3990t629) I(R3990t1630) I(R3991t1653) I(R3991t2537) I(R3991t2877) I(R3991t3068) I(R3991t712) I(R3992t276) I(R3992t1733) I(R3993t2930) I(R3993t3423) I(R3993t3573) I(R3994t1029) I(R3994t803) I(R3994t858) I(R3995t3228) I(R3995t2783) I(R3997t95) I(R3997t699) I(R3997t2160) I(R3997t3275) I(R3998t2802) I(R3999t2989) I(R4000t187) I(R4000t2590) I(R4000t3382) I(R4001t3453) I(R4001t726) I(R4001t2825) I(R4002t2789) I(R4003t344) I(R4003t176) I(R4004t68) I(R4004t2554) I(R4004t3493) I(R4005t2784) I(R4006t765) I(R4007t87) I(R4007t411) I(R4007t566) I(R4007t3820) I(R4008t1765) I(R4008t3843) I(R4008t1842) I(R4009t2043) I(R4009t1270) I(R4009t268) I(R4010t693) I(R4010t1143) I(R4010t1023) I(R4011t1676) I(R4011t2062) I(R4011t1252) I(R4014t874) I(R4015t1077) I(R4015t3899) I(R4015t1393) I(R4015t3508) I(R4015t1830) I(R4016t2936) I(R4016t1873) I(R4016t1256) I(R4017t405) I(R4018t3477) I(R4018t2728) I(R4019t3755) I(R4019t696) I(R4019t1414) I(R4020t2634) I(R4020t2643) I(R4020t1186) I(R4021t402) I(R4021t1439) I(R4021t1445) I(R4022t1247) I(R4022t1304) I(R4023t1331) I(R4023t1579) I(R4026t2776) I(R4026t1312) I(R4027t1564) I(R4028t3228) I(R4028t3676) I(R4028t2150) I(R4028t1198) I(R4029t1344) I(R4029t1825) I(R4029t3345) I(R4029t461) I(R4029t1483) I(R4029t2834) I(R4030t3343) I(R4031t2457) I(R4031t2150) I(R4032t1912) I(R4033t155) I(R4033t2796) I(R4033t3665) I(R4034t1827) I(R4034t2306) I(R4034t1419) I(R4035t3040) I(R4035t1004) I(R4035t1306) I(R4036t3024) I(R4036t829) I(R4037t978) I(R4038t807) I(R4038t753) I(R4038t1565) I(R4038t3323) I(R4040t1000) I(R4040t3601) I(R4041t1318) I(R4041t1621) I(R4042t3476) I(R4042t2734) I(R4043t3454) I(R4044t498) I(R4044t3986) I(R4045t3352) I(R4046t1078) I(R4046t3095) I(R4046t1685) I(R4048t1957) I(R4048t3059) I(R4048t962) I(R4049t717) I(R4050t2024) I(R4050t954) I(R4051t1281) I(R4051t738) I(R4051t3049) I(R4052t2814) I(R4052t3340) I(R4052t3194) I(R4052t1123) I(R4052t3605) I(R4053t958) I(R4054t44) I(R4054t3352) I(R4055t816) I(R4055t2381) I(R4055t607) I(R4057t1456) I(R4057t3088) I(R4057t1511) I(R4058t3823) I(R4058t2390) I(R4059t186) I(R4059t990) I(R4059t2071) I(R4059t2950) I(R4060t3259) I(R4060t3052) I(R4061t1262) I(R4063t339) I(R4063t1888) I(R4063t3828) I(R4064t3411) I(R4064t808) I(R4065t1207) I(R4066t486) I(R4066t1465) I(R4066t1710) I(R4067t3618) I(R4067t3608) I(R4067t1078) I(R4068t1890) I(R4068t3411) I(R4068t4064) I(R4069t2423) I(R4070t1411) I(R4070t3921) I(R4071t1798) I(R4071t3380) I(R4071t799) I(R4072t1495) I(R4072t1041) I(R4072t1542) I(R4073t118) I(R4073t839) I(R4073t1348) I(R4074t3091) I(R4075t879) I(R4075t3120) I(R4076t317) I(R4077t3112) I(R4077t2424) I(R4077t549) I(R4078t2809) I(R4078t3811) I(R4078t1092) I(R4078t1331) I(R4078t4023) I(R4078t1588) I(R4079t1076) I(R4079t2844) I(R4079t3949) I(R4080t1842) I(R4080t1349) I(R4081t2276) I(R4081t611) I(R4082t1110) I(R4082t1648) I(R4082t1096) I(R4082t3479) I(R4083t1958) I(R4084t596) I(R4084t938) I(R4084t100) I(R4084t1430) I(R4085t1126) I(R4085t3027) I(R4086t1021) I(R4087t1117) I(R4088t3677) I(R4088t2253) I(R4088t1265) I(R4088t522) I(R4089t2574) I(R4090t158) I(R4090t236) I(R4090t1540) I(R4091t2525) I(R4091t2860) I(R4091t2002) I(R4091t1892) I(R4092t2591) I(R4092t2054) I(R4092t394) I(R4093t1287) I(R4093t2116) I(R4093t1317) I(R4093t892) I(R4094t941) I(R4094t3187) I(R4094t1025) I(R4095t2676) I(R4095t2193) I(R4096t2938) I(R4096t1929) I(R4096t2191) I(R4096t3973) I(R4096t1477) I(R4097t1750) I(R4097t760) I(R4097t2695) I(R4097t3233) I(R4098t425) I(R4099t3450) I(R4099t307) I(R4100t3623) I(R4101t2956) I(R4101t2341) I(R4102t643) I(R4102t3614) I(R4102t943) I(R4102t990) I(R4102t4059) I(R4102t2071) I(R4103t1270) I(R4104t2740) I(R4105t1415) I(R4105t3519) I(R4105t204) I(R4106t1351) I(R4106t3910) I(R4106t851) I(R4107t2015) I(R4107t1577) I(R4107t2560) I(R4108t459) I(R4108t3602) I(R4108t793) I(R4108t2036) I(R4109t468) I(R4109t1132) I(R4109t1619) I(R4110t397) I(R4110t2305) I(R4111t2155) I(R4111t2440) I(R4111t3461) I(R4111t3242) I(R4112t83) I(R4112t2525) I(R4112t1288) I(R4112t2860) I(R4113t2657) I(R4113t2545) I(R4113t219) I(R4114t1144) I(R4115t3237) I(R4115t918) I(R4115t336) I(R4116t1440) I(R4116t1338) I(R4116t471) I(R4117t1561) I(R4118t4067) I(R4119t401) I(R4119t3040) I(R4119t4035) I(R4119t1004) I(R4120t382) I(R4120t3503) I(R4120t3809) I(R4121t2819) I(R4121t1196) I(R4122t795) I(R4122t1447) I(R4122t2158) I(R4123t916) I(R4123t523) I(R4123t2320) I(R4124t89) I(R4124t154) I(R4124t2100) I(R4124t1777) I(R4124t176) I(R4125t1147) I(R4125t3880) I(R4126t1605) I(R4126t334) I(R4126t1166) I(R4127t583) I(R4127t3785) I(R4127t82) I(R4127t3150) I(R4128t1513) I(R4129t1123) I(R4129t1566) I(R4129t925) I(R4129t2372) I(R4130t383) I(R4130t2532) I(R4131t4100) I(R4131t1702) I(R4132t3742) I(R4132t2144) I(R4132t3162) I(R4133t2681) I(R4133t3164) I(R4133t1511) I(R4133t4057) I(R4133t3088) I(R4134t2922) I(R4134t146) I(R4134t164) I(R4135t1870) I(R4136t2002) I(R4136t4091) I(R4136t1892) I(R4136t2243) I(R4136t1485) I(R4137t921) I(R4137t3087) I(R4137t1173) I(R4137t923) I(R4137t3564) I(R4138t2523) I(R4138t2418) I(R4138t102) I(R4138t1466) I(R4139t2606) I(R4139t1040) I(R4140t2318) I(R4140t1918) I(R4141t3296) I(R4141t1734) I(R4142t536) I(R4142t2724) I(R4142t2888) I(R4142t3457) I(R4143t1247) I(R4143t3885) I(R4143t2003) I(R4143t2969) I(R4144t410) I(R4144t3581) I(R4145t1780) I(R4146t3294) I(R4146t2044) I(R4146t1521) I(R4147t1076) I(R4147t2575) I(R4147t3903) I(R4147t1837) I(R4147t3949) I(R4147t4079) I(R4148t312) I(R4148t3477) I(R4148t467) I(R4148t3856) I(R4148t2728) I(R4149t2965) I(R4149t676) I(R4149t2158) I(R4150t1619) I(R4151t237) I(R4152t1654) I(R4152t109) I(R4153t2682) I(R4153t3246) I(R4154t197) I(R4155t1038) I(R4155t2545) I(R4155t4113) I(R4156t1910) I(R4156t2963) I(R4156t1455) I(R4156t1647) I(R4157t262) I(R4157t2738) I(R4158t2807) I(R4158t3213) I(R4158t3145) I(R4158t3502) I(R4158t1510) I(R4159t390) I(R4159t418) I(R4159t3805) I(R4160t3290) I(R4160t4044) I(R4161t2048) I(R4161t2579) I(R4161t526) I(R4162t3442) I(R4162t2047) I(R4162t1812) I(R4162t3634) I(R4163t103) I(R4164t2624) I(R4164t3047) I(R4164t2255) I(R4165t2505) I(R4165t3258) I(R4165t1172) I(R4165t2375) I(R4166t2553) I(R4166t132) I(R4166t1249) I(R4167t344) I(R4167t756) I(R4167t4003) I(R4168t2569) I(R4168t354) I(R4169t1870) I(R4169t3693) I(R4170t3874) I(R4170t1925) I(R4170t3844) I(R4170t3030) I(R4171t2069) I(R4171t2137) I(R4172t363) I(R4173t2464) I(R4173t2660) I(R4173t3602) I(R4174t3886) I(R4174t3758) I(R4174t3608) I(R4174t3618) I(R4175t1509) I(R4175t1417) I(R4176t3155) I(R4176t1262) I(R4176t3410) I(R4176t2867) I(R4177t397) I(R4177t2728) I(R4177t2305) I(R4178t4127) I(R4178t583) I(R4178t857) I(R4178t1231) I(R4178t2864) I(R4179t854) I(R4179t2543) I(R4180t544) I(R4180t1953) I(R4181t2210) I(R4181t502) I(R4181t1729) I(R4182t3350) I(R4183t832) I(R4183t2509) I(R4183t3503) I(R4183t1586) I(R4184t1897) I(R4184t416) I(R4184t3546) I(R4185t3883) I(R4186t1956) I(R4186t3994) I(R4187t1125) I(R4187t2316) I(R4187t2814) I(R4188t3314) I(R4189t3156) I(R4189t3435) I(R4189t3232) I(R4190t115) I(R4190t24) I(R4191t2456) I(R4191t4105) I(R4191t4185) I(R4192t613) I(R4192t2389) I(R4192t247) I(R4192t869) I(R4193t2146) I(R4193t2218) I(R4193t2471) I(R4194t3233) I(R4194t1441) I(R4195t1178) I(R4195t1227) I(R4196t527) I(R4196t4062) I(R4197t107) I(R4197t1199) I(R4197t2812) I(R4197t4169) I(R4197t3693) I(R4198t3116) I(R4198t3460) I(R4198t2720) I(R4199t2224) I(R4200t336) I(R4200t4115) I(R4200t918) I(R4200t2127) I(R4201t32) I(R4201t3868) I(R4202t3039) I(R4202t1037) I(R4202t2980) I(R4202t1500) I(R4203t2978) I(R4204t217) I(R4204t933) I(R4204t1442) I(R4205t363) I(R4206t2632) I(R4207t453) I(R4207t1908) I(R4208t4043) I(R4208t3454) I(R4209t593) I(R4209t1321) I(R4210t1082) I(R4210t2486) I(R4210t2280) I(R4211t1522) I(R4211t1754) I(R4211t2031) I(R4212t3269) I(R4213t3525) I(R4213t2271) I(R4214t3709) I(R4215t888) I(R4215t3321) I(R4216t3941) I(R4216t562) I(R4216t3403) I(R4217t779) I(R4217t2454) I(R4218t4081) I(R4218t611) I(R4218t1389) I(R4219t2902) I(R4220t1652) I(R4220t3674) I(R4221t3755) I(R4221t3558) I(R4221t170) I(R4221t2227) I(R4221t33) I(R4222t3281) I(R4223t903) I(R4223t2552) I(R4224t1136) I(R4224t2476) I(R4225t205) I(R4226t442) I(R4226t2793) I(R4227t1403) I(R4227t1400) I(R4227t1583) I(R4228t1863) I(R4228t2010) I(R4228t2097) I(R4229t1436) I(R4229t3031) I(R4230t1717) I(R4230t4207) I(R4230t1319) I(R4231t1307) I(R4232t478) I(R4233t3182) I(R4233t248) I(R4234t1617) I(R4234t2661) I(R4235t3590) I(R4235t2406) I(R4235t773) I(R4236t3684) I(R4236t260) I(R4236t4193) I(R4237t2670) I(R4237t957) I(R4237t3264) I(R4237t2211) I(R4238t3760) I(R4238t1600) I(R4239t3781) I(R4239t835) I(R4240t2328) I(R4240t1149) I(R4240t807) I(R4240t1899) I(R4241t3710) I(R4241t3692) I(R4241t1613) I(R4243t2772) I(R4244t2766) I(R4244t3251) I(R4244t3390) I(R4245t751) I(R4245t2691) I(R4246t3154) I(R4246t1704) I(R4247t2882) I(R4247t1188) I(R4247t178) I(R4248t1431) I(R4248t3300) I(R4248t1353) I(R4248t1318) I(R4248t4041) I(R4249t1261) I(R4249t3302) I(R4250t3253) I(R4250t3441) I(R4250t3127) I(R4251t2212) I(R4251t2566) I(R4251t2795) I(R4252t1504) I(R4252t197) I(R4252t4154) I(R4253t3032) I(R4253t3414) I(R4254t1371) I(R4254t2761) I(R4255t1793) I(R4256t96) I(R4256t1599) I(R4256t2792) I(R4256t1763) I(R4257t1603) I(R4257t1758) I(R4257t1079) I(R4257t696) I(R4258t95) I(R4258t2160) I(R4258t2703) I(R4259t1614) I(R4260t3330) I(R4260t268) I(R4260t1270) I(R4260t899) I(R4261t2268) I(R4261t3961) I(R4261t3486) I(R4262t587) I(R4262t100) I(R4263t146) I(R4263t4134) I(R4263t164) I(R4264t1661) I(R4264t2513) I(R4264t438) I(R4264t549) I(R4265t1980) I(R4265t1716) I(R4265t3920) I(R4267t936) I(R4267t1987) I(R4268t3445) I(R4269t1459) I(R4269t3766) I(R4270t282) I(R4270t1050) I(R4271t1886) I(R4271t4195) I(R4272t3913) I(R4272t3908) I(R4272t836) I(R4272t377) I(R4273t3888) I(R4273t1046) I(R4275t1216) I(R4275t955) I(R4275t462) I(R4276t2629) I(R4276t3901) I(R4277t1109) I(R4278t963) I(R4278t1106) I(R4279t2380) I(R4280t3203) I(R4280t3909) I(R4280t3385) I(R4280t1923) I(R4280t885) I(R4281t553) I(R4282t3921) I(R4282t1411) I(R4282t4070) I(R4283t1505) I(R4283t4065) I(R4284t2938) I(R4284t1477) I(R4284t4070) I(R4285t1805) I(R4285t4) I(R4286t426) I(R4287t1250) I(R4289t2718) I(R4290t682) I(R4291t815) I(R4291t2788) I(R4291t2440) I(R4291t3461) I(R4292t3817) I(R4292t2854) I(R4293t2602) I(R4294t2051) I(R4294t3269) I(R4294t4212) I(R4295t1788) I(R4295t156) I(R4296t2805) I(R4297t2709) I(R4297t2777) I(R4297t2942) I(R4297t2954) I(R4298t1881) I(R4298t3797) I(R4299t2061) I(R4299t2821) I(R4299t446) I(R4300t3018) I(R4300t956) I(R4301t3202) I(R4301t1186) I(R4302t1310) I(R4302t1518) I(R4302t1465) I(R4303t2467) I(R4303t3713) I(R4303t2599) I(R4303t2041) I(R4304t3624) I(R4304t2624) I(R4305t2558) I(R4305t1927) I(R4305t3658) I(R4306t1068) I(R4306t2999) I(R4306t2556) I(R4307t545) I(R4307t3498) I(R4307t697) I(R4307t1986) I(R4308t3821) I(R4308t61) I(R4308t3291) I(R4309t2115) I(R4310t898) I(R4310t2053) I(R4311t780) I(R4311t2924) I(R4312t578) I(R4312t1879) I(R4312t1781) I(R4313t2909) I(R4313t3868) I(R4314t3717) I(R4314t279) I(R4314t3553) I(R4314t1526) I(R4314t120) I(R4315t561) I(R4315t931) I(R4315t3299) I(R4316t790) I(R4316t1434) I(R4317t3507) I(R4317t538) I(R4317t1143) I(R4317t1023) I(R4318t1825) I(R4318t4029) I(R4318t1344) I(R4319t1624) I(R4320t1580) I(R4320t2713) I(R4321t2406) I(R4321t4235) I(R4321t3590) I(R4321t1544) I(R4321t53) I(R4322t1353) I(R4322t4248) I(R4322t1318) I(R4322t2258) I(R4322t60) I(R4323t1478) I(R4323t905) I(R4325t3004) I(R4325t493) I(R4326t1265) I(R4326t3724) I(R4326t1433) I(R4326t1030) I(R4326t3799) I(R4327t898) I(R4327t2053) I(R4327t4284) I(R4327t2938) I(R4327t428) I(R4327t656) I(R4328t2270) I(R4328t519) I(R4329t1941) I(R4329t1390) I(R4329t2418) I(R4329t322) I(R4331t3091) I(R4331t4074) I(R4332t1145) I(R4332t3797) I(R4333t3623) I(R4334t4123) I(R4334t523) I(R4335t2958) I(R4336t404) I(R4336t1725) I(R4336t3867) I(R4337t4141) I(R4337t2807) I(R4338t3455) I(R4339t2512) I(R4339t1752) I(R4340t1500) I(R4340t2442) I(R4340t4202) I(R4340t2614) I(R4340t2214) I(R4341t781) I(R4342t3446) I(R4343t3364) I(R4343t4314) I(R4344t228) I(R4344t4138) I(R4344t1466) I(R4344t2949) I(R4345t3449) I(R4345t1949) I(R4345t3006) I(R4345t2357) I(R4346t429) I(R4346t3643) I(R4346t2279) I(R4346t3357) I(R4346t1832) I(R4347t3157) I(R4348t1371) I(R4348t4267) I(R4348t936) I(R4348t4254) I(R4349t3946) I(R4350t1284) I(R4350t3770) I(R4350t683) I(R4351t1075) I(R4351t3297) I(R4351t3651) I(R4352t3094) I(R4352t3853) I(R4353t982) I(R4353t3364) I(R4353t4343) I(R4353t4314) I(R4353t120) I(R4353t1823) I(R4354t3077) I(R4354t3701) I(R4354t3776) I(R4354t3695) I(R4355t4082) I(R4356t1063) I(R4357t907) I(R4357t2802) I(R4358t1377) I(R4358t2474) I(R4358t1969) I(R4359t3646) I(R4359t903) I(R4359t4223) I(R4360t2466) I(R4360t3467) I(R4360t2190) I(R4362t2046) I(R4362t1889) I(R4362t3890) I(R4362t2595) I(R4363t1145) I(R4363t1227) I(R4363t1233) I(R4363t331) I(R4364t1726) I(R4365t3161) I(R4365t3882) I(R4366t1462) I(R4367t1377) I(R4367t4358) I(R4367t1969) I(R4367t2619) I(R4368t1721) I(R4369t2258) I(R4369t3846) I(R4369t3975) I(R4370t1205) I(R4370t1833) I(R4371t1633) I(R4371t3146) I(R4371t2868) I(R4371t2641) I(R4372t2310) I(R4372t4246) I(R4372t3056) I(R4373t317) I(R4373t4076) I(R4374t1649) I(R4374t1958) I(R4375t2553) I(R4375t4166) I(R4375t132) I(R4375t3958) I(R4375t2594) I(R4376t1032) I(R4376t3161) I(R4376t1988) I(R4376t4365) I(R4377t355) I(R4377t1083) I(R4377t3780) I(R4377t4265) I(R4378t813) I(R4378t1902) I(R4378t617) I(R4378t3421) I(R4378t1541) I(R4378t470) I(R4378t999) I(R4379t551) I(R4379t2596) I(R4379t605) I(R4380t229) I(R4380t3637) I(R4380t3100) I(R4380t3567) I(R4381t3145) I(R4381t4158) I(R4381t3502) I(R4382t2281) I(R4382t257) I(R4382t3694) I(R4383t298) I(R4383t4103) I(R4383t902) I(R4384t1122) I(R4386t1973) I(R4386t50) I(R4386t2257) I(R4387t2635) I(R4387t2880) I(R4388t628) I(R4388t3418) I(R4388t2412) I(R4388t256) I(R4388t3393) I(R4389t4132) I(R4389t3742) I(R4390t2737) I(R4391t2962) I(R4392t4389) I(R4392t708) I(R4393t579) I(R4393t414) I(R4394t610) I(R4394t2744) I(R4394t141) I(R4395t2566) I(R4395t3610) I(R4395t1457) I(R4395t2883) I(R4396t4308) I(R4396t61) I(R4397t1232) I(R4397t333) I(R4398t1502) I(R4398t78) I(R4398t256) I(R4399t1293) I(R4399t472) I(R4399t988) I(R4399t1335) I(R4400t1457) I(R4400t4395) I(R4400t1324) I(R4401t3056) I(R4401t4372) I(R4401t1445) I(R4401t4021) I(R4401t3154) I(R4401t4246) I(R4402t2162) I(R4402t2517) I(R4402t2054) I(R4402t1293) I(R4402t2280) I(R4402t2109) I(R4403t72) I(R4403t1019) I(R4404t2522) I(R4405t1276) I(R4406t1138) I(R4407t186) I(R4407t990) I(R4407t4059) I(R4408t3247) I(R4408t2742) I(R4408t1490) I(R4409t1574) I(R4409t2758) I(R4410t2007) I(R4412t3514) I(R4412t3942) I(R4413t2427) I(R4413t3725) I(R4414t3312) I(R4415t2988) I(R4415t3597) I(R4415t300) I(R4415t3802) I(R4416t3620) I(R4416t1646) I(R4416t110) I(R4416t3009) I(R4418t2772) I(R4418t4243) I(R4419t2651) I(R4419t3287) I(R4419t1665) I(R4419t192) I(R4419t3570) I(R4419t565) I(R4420t11) I(R4420t1819) I(R4420t3830) I(R4420t304) I(R4420t1015) I(R4421t900) I(R4421t3969) I(R4421t757) I(R4421t50) I(R4421t1973) I(R4421t3773) I(R4422t3114) I(R4423t355) I(R4423t2567) I(R4424t2623) I(R4424t3434) I(R4425t4215) I(R4425t888) I(R4426t2607) I(R4426t1599) I(R4427t2066) I(R4427t1459) I(R4428t1505) I(R4428t4283) I(R4428t4065) I(R4429t4005) I(R4429t1619) I(R4430t3331) I(R4430t404) I(R4431t3427) I(R4432t3556) I(R4432t2908) I(R4432t2) I(R4433t3772) I(R4433t2342) I(R4433t3833) I(R4434t2281) I(R4435t3047) I(R4435t4164) I(R4435t2255) I(R4436t1687) I(R4436t2191) I(R4437t4393) I(R4437t1135) I(R4438t906) I(R4438t2290) I(R4438t3659) I(R4438t3585) I(R4438t569) I(R4439t2782) I(R4439t741) I(R4439t3413) I(R4439t1197) I(R4440t1940) I(R4440t3187) I(R4441t3395) I(R4441t1351) I(R4441t4106) I(R4443t1240) I(R4443t3933) I(R4443t3734) I(R4444t630) I(R4444t3619) I(R4444t3813) I(R4445t4226) I(R4445t107) I(R4445t2858) I(R4445t2793) I(R4446t1705) I(R4446t2055) I(R4447t821) I(R4447t1877) I(R4447t2804) I(R4448t1865) I(R4449t3681) I(R4449t3931) I(R4449t806) I(R4450t2761) I(R4450t834) I(R4451t3968) I(R4451t3349) I(R4451t4333) I(R4451t3623) I(R4452t1087) I(R4452t2850) I(R4453t1994) I(R4453t3206) I(R4453t3384) I(R4454t1944) I(R4454t1919) I(R4454t2734) I(R4454t4042) I(R4455t1994) I(R4455t4453) I(R4456t4284) I(R4456t4327) I(R4456t898) I(R4457t1704) I(R4457t4246) I(R4457t4372) I(R4457t2310) I(R4458t545) I(R4458t3304) I(R4458t1418) I(R4458t633) I(R4458t3706) I(R4459t1983) I(R4459t3901) I(R4459t4276) I(R4459t2629) I(R4459t2935) I(R4459t2293) I(R4460t1304) I(R4460t2969) I(R4460t4143) I(R4460t1247) I(R4460t4022) I(R4461t116) I(R4461t1134) I(R4462t2298) I(R4462t3595) I(R4462t3093) I(R4462t2678) I(R4462t2093) I(R4463t621) I(R4463t3731) I(R4463t75) I(R4463t3517) I(R4464t2714) I(R4464t1274) I(R4464t2221) I(R4465t416) I(R4465t3546) I(R4466t2611) I(R4466t1878) I(R4467t41) I(R4467t1699) I(R4467t3317) I(R4468t4312) I(R4468t2582) I(R4469t2501) I(R4469t3149) I(R4469t1113) I(R4470t363) I(R4470t4172) I(R4470t4205) I(R4471t2265) I(R4471t2801) I(R4471t1992) I(R4471t1749) I(R4471t3834) I(R4472t3951) I(R4472t4224) I(R4472t2476) I(R4472t987) I(R4472t3325) I(R4473t454) I(R4473t1352) I(R4473t133) I(R4473t3852) I(R4473t3896) I(R4474t298) I(R4474t899) I(R4474t4260) I(R4474t1270) I(R4474t4103) I(R4474t4383) I(R4475t2070) I(R4475t1425) I(R4475t3326) I(R4476t1705) I(R4476t2039) I(R4476t3839) I(R4477t189) I(R4477t2674) I(R4478t1186) I(R4478t3268) I(R4479t3188) I(R4480t2941) I(R4480t2859) I(R4481t3504) I(R4482t1090) I(R4482t1848) I(R4482t768) I(R4483t138) I(R4483t2650) I(R4483t46) I(R4483t849) I(R4484t1438) I(R4484t2697) I(R4484t2420) I(R4484t4188) I(R4484t3314) I(R4485t3014) I(R4485t309) I(R4485t1194) I(R4485t372) I(R4486t131) I(R4486t1995) I(R4486t990) I(R4486t4407) I(R4487t3255) I(R4487t3814) I(R4487t4290) I(R4488t1156) I(R4488t3510) I(R4488t3351) I(R4488t2607) I(R4489t1296) I(R4489t4114) I(R4489t330) I(R4490t612) I(R4490t1668) I(R4490t3019) I(R4491t2857) I(R4491t1809) I(R4492t2594) I(R4493t3472) I(R4493t1459) I(R4493t2066) I(R4494t3951) I(R4494t4472) I(R4494t3325) I(R4494t398) I(R4495t1206) I(R4495t2890) I(R4495t2426) I(R4495t554) I(R4496t3794) I(R4496t3804) I(R4496t1157) I(R4496t3736) I(R4497t3109) I(R4498t2431) I(R4498t3473) I(R4498t3836) I(R4499t3227) I(R4499t1392) I(R4499t1591) I(R4500t2483) I(R4500t3880) I(R4500t2984) I(R4501t538) I(R4501t4317) I(R4502t3591) I(R4502t1108) I(R4503t341) I(R4503t3439) I(R4503t1775) I(R4503t201) I(R4504t1552) I(R4504t2502) I(R4505t4037) I(R4505t3992) I(R4506t1878) I(R4506t4466) I(R4506t3263) I(R4507t3893) I(R4507t2576) I(R4507t3394) I(R4507t1379) I(R4507t3795) I(R4508t615) I(R4508t4479) I(R4509t171) I(R4509t2482) I(R4510t4134) I(R4510t164) I(R4510t863) I(R4510t487) I(R4510t2207) I(R4511t1720) I(R4511t3636) I(R4512t1654) I(R4512t4152) I(R4513t24) I(R4514t3109) I(R4514t4497) I(R4514t2399) I(R4515t943) I(R4515t1812) I(R4516t3374) I(R4516t4225) I(R4517t3825) I(R4517t994) I(R4518t401) I(R4518t4119) I(R4518t2089) I(R4519t1407) I(R4519t3415) I(R4520t765) I(R4520t3740) I(R4520t2493) I(R4520t3516) I(R4520t4006) I(R4521t1968) I(R4521t3672) I(R4522t1268) I(R4522t1787) I(R4523t3513) I(R4523t3448) I(R4524t160) I(R4524t285) I(R4525t665) I(R4525t1326) I(R4525t3508) I(R4526t3401) I(R4526t1999) I(R4526t1214) I(R4526t98) I(R4526t2331) I(R4527t3508) I(R4527t4525) I(R4527t665) I(R4527t325) I(R4528t1079) I(R4528t64) I(R4528t460) I(R4529t1797) I(R4529t1579) I(R4529t3135) I(R4530t1195) I(R4530t1084) I(R4531t2518) I(R4531t2205) I(R4532t2626) I(R4532t2561) I(R4532t3133) I(R4533t2217) I(R4533t2257) I(R4534t3449) I(R4534t1949) I(R4534t4345) I(R4535t2260) I(R4535t1397) I(R4536t3494) I(R4536t3509) I(R4536t4145) I(R4536t1780) I(R4537t1064) I(R4537t1043) I(R4537t1432) I(R4538t1532) I(R4538t2855) I(R4539t3182) I(R4539t4233) I(R4540t4447) I(R4541t1894) I(R4541t2729) I(R4541t357) I(R4542t2744) I(R4542t3854) I(R4542t1755) I(R4542t4394) I(R4543t1116) I(R4544t468) I(R4544t507) I(R4544t4109) I(R4545t3173) I(R4545t4044) I(R4545t3986) I(R4547t167) I(R4547t2753) I(R4547t3579) I(R4548t4540) I(R4548t4447) I(R4548t2804) I(R4549t3489) I(R4550t1094) I(R4550t1628) I(R4550t3565) I(R4550t3959) I(R4550t2022) I(R4550t3627) I(R4551t1905) I(R4551t294) I(R4552t3512) I(R4552t3628) I(R4552t1555) I(R4553t1182) I(R4553t3667) I(R4554t652) I(R4554t673) I(R4554t758) I(R4554t4221) I(R4554t33) I(R4555t1745) I(R4556t1292) I(R4556t1427) I(R4556t1616) I(R4557t1959) I(R4557t3973) I(R4558t2334) I(R4558t2388) I(R4559t2635) I(R4559t729) I(R4559t359) I(R4560t254) I(R4560t3866) I(R4560t4162) I(R4561t546) I(R4561t3705) I(R4561t1225) I(R4562t1303) I(R4562t1299) I(R4563t4199) I(R4564t1318) I(R4564t2258) I(R4564t4041) I(R4564t3846) I(R4565t2968) I(R4565t3670) I(R4565t2393) I(R4566t432) I(R4566t3461) I(R4566t4111) I(R4566t3242) I(R4566t4390) I(R4567t4222) I(R4568t3507) I(R4568t4317) I(R4568t4501) I(R4569t1155) I(R4569t2232) I(R4570t10) I(R4570t4465) I(R4571t1098) I(R4571t3936) I(R4571t2562) I(R4571t3751) I(R4571t1718) I(R4571t1332) I(R4571t3208) I(R4572t3718) I(R4572t3726) I(R4572t30) I(R4572t1796) I(R4573t3433) I(R4573t991) I(R4574t2295) I(R4574t43) I(R4575t1835) I(R4575t3329) I(R4575t116) I(R4575t2185) I(R4576t264) I(R4576t2906) I(R4576t3207) I(R4577t173) I(R4577t2803) I(R4577t1093) I(R4577t627) I(R4578t3193) I(R4579t4072) I(R4579t1542) I(R4579t2365) I(R4579t2641) I(R4580t4203) I(R4581t2329) I(R4581t917) I(R4582t3543) I(R4582t4060) I(R4582t3259) I(R4582t86) I(R4583t3806) I(R4583t1373) I(R4583t2955) I(R4583t3109) I(R4584t834) I(R4584t4450) I(R4584t2175) I(R4584t1780) I(R4585t1192) I(R4585t1630) I(R4585t629) I(R4586t1774) I(R4587t2515) I(R4587t1699) I(R4587t1310) I(R4588t2070) I(R4589t2829) I(R4589t3723) I(R4589t2946) I(R4590t2178) I(R4590t1813) I(R4590t3912) I(R4591t4180) I(R4591t544) I(R4592t514) I(R4592t1264) I(R4592t1278) I(R4592t1461) I(R4592t2366) I(R4592t3631) I(R4593t3040) I(R4593t2855) I(R4593t2586) I(R4593t3262) I(R4594t3508) I(R4594t4527) I(R4594t4015) I(R4594t1393) I(R4594t521) I(R4594t325) I(R4595t2483) I(R4595t2984) I(R4595t3259) I(R4595t484) I(R4596t2195) I(R4596t3249) I(R4596t2503) I(R4596t3370) I(R4597t1146) I(R4597t3917) I(R4597t1875) I(R4597t3344) I(R4598t3565) I(R4598t1979) I(R4598t856) I(R4599t4361) I(R4599t1672) I(R4599t2249) I(R4599t2466) I(R4599t3889) I(R4601t1633) I(R4601t2901) I(R4602t1734) I(R4602t3296) I(R4602t310) I(R4602t1869) I(R4603t740) I(R4603t3850) I(R4604t1659) I(R4605t4097) I(R4606t2543) I(R4606t4245) I(R4606t850) I(R4608t3292) I(R4609t327) I(R4610t2076) I(R4610t657) I(R4611t903) I(R4611t314) I(R4611t492) I(R4612t3657) I(R4612t1517) I(R4613t3643) I(R4613t4346) I(R4613t1832) I(R4613t2370) I(R4613t800) I(R4614t1256) I(R4614t4016) I(R4614t2936) I(R4615t1027) I(R4615t1756) I(R4615t2760) I(R4616t1271) I(R4616t2046) I(R4616t4362) I(R4616t3796) I(R4617t160) I(R4617t3293) I(R4617t1236) I(R4618t1180) I(R4618t117) I(R4618t878) I(R4618t1316) I(R4618t2400) I(R4619t4445) I(R4619t2878) I(R4619t107) I(R4620t3962) I(R4621t985) I(R4621t251) I(R4621t2802) I(R4621t3998) I(R4622t952) I(R4622t2714) I(R4622t3504) I(R4622t1901) I(R4622t2099) I(R4623t1491) I(R4623t1345) I(R4623t3012) I(R4624t1659) I(R4624t579) I(R4625t2591) I(R4625t4006) I(R4626t4504) I(R4626t2502) I(R4626t2610) I(R4627t2526) I(R4627t20) I(R4628t1102) I(R4628t395) I(R4628t895) I(R4629t1364) I(R4629t2915) I(R4629t2333) I(R4630t3945) I(R4630t2385) I(R4630t767) I(R4631t1301) I(R4631t3078) I(R4631t3265) I(R4632t1759) I(R4632t1654) I(R4632t2886) I(R4632t3769) I(R4632t1745) I(R4632t4555) I(R4633t1697) I(R4633t1220) I(R4634t1890) I(R4634t4068) I(R4634t4175) I(R4635t1165) I(R4635t1937) I(R4635t2035) I(R4635t3385) I(R4636t4141) I(R4636t4337) I(R4636t2807) I(R4636t3213) I(R4638t3447) I(R4638t3806) I(R4639t4515) I(R4639t943) I(R4639t4296) I(R4639t2805) I(R4640t1847) I(R4640t1628) I(R4640t3565) I(R4640t4598) I(R4641t1488) I(R4642t4510) I(R4642t2207) I(R4642t3355) I(R4643t1062) I(R4644t1761) I(R4644t2662) I(R4645t1460) I(R4645t1520) I(R4645t2773) I(R4646t687) I(R4646t2939) I(R4646t2945) I(R4647t3202) I(R4647t4045) I(R4647t3352) I(R4647t1715) I(R4648t447) I(R4648t1321) I(R4649t382) I(R4649t4120) I(R4649t4053) I(R4649t958) I(R4650t2646) I(R4650t4638) I(R4650t3806) I(R4651t621) I(R4651t3517) I(R4651t2006) I(R4652t3704) I(R4652t317) I(R4652t1644) I(R4653t241) I(R4653t660) I(R4654t2641) I(R4654t3644) I(R4654t2365) I(R4655t4219) I(R4655t2902) I(R4655t979) I(R4656t2309) I(R4656t3988) I(R4656t2032) I(R4658t1371) I(R4658t215) I(R4658t4254) I(R4659t2607) I(R4659t4426) I(R4659t4488) I(R4659t96) I(R4659t4256) I(R4659t1599) I(R4660t2623) I(R4660t994) I(R4660t4517) I(R4660t3825) I(R4661t4299) I(R4661t1358) I(R4661t590) I(R4662t1000) I(R4662t1354) I(R4662t3601) I(R4662t1244) I(R4662t3966) I(R4663t3970) I(R4663t3274) I(R4663t403) I(R4663t1044) I(R4664t983) I(R4664t2625) I(R4664t2138) I(R4664t994) I(R4664t4517) I(R4664t3825) I(R4664t2130) I(R4664t1570) I(R4665t2001) I(R4665t996) I(R4666t4042) I(R4667t588) I(R4667t946) I(R4667t2024) I(R4667t4050) I(R4668t1406) I(R4668t3391) I(R4668t1206) I(R4668t3566) I(R4668t1473) I(R4669t922) I(R4669t392) I(R4669t883) I(R4669t370) I(R4669t3661) I(R4670t2222) I(R4670t2864) I(R4670t4178) I(R4670t4192) I(R4670t247) I(R4670t869) I(R4671t2829) I(R4672t4667) I(R4672t3381) I(R4672t946) I(R4673t1831) I(R4673t950) I(R4673t1688) I(R4674t35) I(R4674t125) I(R4674t3876) I(R4674t3424) I(R4675t3525) I(R4675t4213) I(R4676t310) I(R4676t4651) I(R4676t949) I(R4676t2562) I(R4677t2817) I(R4677t3802) I(R4678t1213) I(R4678t21) I(R4679t815) I(R4680t129) I(R4680t868) I(R4680t2851) I(R4680t1638) I(R4681t983) I(R4681t2507) I(R4681t1960) I(R4681t2993) I(R4682t3307) I(R4682t1492) I(R4682t1130) I(R4683t1895) I(R4683t3185) I(R4683t3367) I(R4684t4380) I(R4684t3100) I(R4685t4573) I(R4685t3433) I(R4685t1601) I(R4685t824) I(R4685t367) I(R4686t527) I(R4687t710) I(R4687t3929) I(R4687t734) I(R4687t150) I(R4688t3694) I(R4688t3944) I(R4688t798) I(R4688t500) I(R4689t3122) I(R4690t1516) I(R4691t717) I(R4691t1667) I(R4691t4049) I(R4692t4411) I(R4692t3888) I(R4692t4273) I(R4693t958) I(R4693t4649) I(R4693t479) I(R4694t74) I(R4694t4433) I(R4694t3772) I(R4695t3721) I(R4695t2695) I(R4695t1427) I(R4695t3099) I(R4697t1986) I(R4697t697) I(R4697t3621) I(R4698t1184) I(R4698t3824) I(R4699t3516) I(R4699t4006) I(R4699t70) I(R4699t528) I(R4699t680) I(R4699t3670) I(R4700t3575) I(R4700t3707) I(R4700t2398) I(R4700t502) I(R4701t2008) I(R4702t2323) I(R4702t1681) I(R4702t1969) I(R4702t2474) I(R4703t2354) I(R4703t3535) I(R4703t1526) I(R4703t4314) I(R4703t3553) I(R4704t2757) I(R4704t1809) I(R4704t3688) I(R4704t2465) I(R4704t805) I(R4705t1148) I(R4705t4437) I(R4706t1137) I(R4706t3016) I(R4706t3684) I(R4707t715) I(R4707t4259) I(R4708t792) I(R4708t3351) I(R4708t1264) I(R4708t1278) I(R4709t3024) I(R4709t4036) I(R4709t205) I(R4709t4225) I(R4709t4516) I(R4709t1664) I(R4709t2019) I(R4710t886) I(R4710t4047) I(R4710t1668) I(R4710t4490) I(R4710t612) I(R4711t4110) I(R4711t1198) I(R4711t2305) I(R4712t1890) I(R4712t4634) I(R4712t1608) I(R4712t2923) I(R4713t2023) I(R4713t1061) I(R4714t740) I(R4714t1344) I(R4714t633) I(R4714t3706) I(R4714t1843) I(R4714t2834) I(R4715t4022) I(R4715t1675) I(R4716t1908) I(R4716t4207) I(R4717t2310) I(R4717t4457) I(R4718t746) I(R4718t1218) I(R4718t1056) I(R4719t1061) I(R4719t1643) I(R4719t1793) I(R4720t3182) I(R4720t4539) I(R4720t2736) I(R4720t2960) I(R4721t114) I(R4721t1673) I(R4721t1627) I(R4721t1240) I(R4721t346) I(R4722t2489) I(R4723t232) I(R4724t2468) I(R4724t2173) I(R4725t908) I(R4725t3423) I(R4725t838) I(R4726t4017) I(R4726t4083) I(R4726t2862) I(R4727t2908) I(R4728t1602) I(R4728t2101) I(R4729t81) I(R4729t2533) I(R4729t1000) I(R4729t4040) I(R4730t991) I(R4730t3041) I(R4730t2928) I(R4730t2997) I(R4731t3487) I(R4731t758) I(R4732t1507) I(R4732t3172) I(R4733t1931) I(R4733t3854) I(R4733t4542) I(R4733t1755) I(R4733t4115) I(R4734t1234) I(R4734t1828) I(R4734t4234) I(R4734t1617) I(R4735t2978) I(R4735t4203) I(R4736t2297) I(R4736t3770) I(R4736t683) I(R4736t4350) I(R4737t1734) I(R4737t4141) I(R4737t3936) I(R4738t1059) I(R4738t601) I(R4738t159) I(R4739t4160) I(R4739t252) I(R4739t3333) I(R4739t3290) I(R4740t2958) I(R4741t833) I(R4741t2899) I(R4742t2437) I(R4743t635) I(R4743t2370) I(R4743t540) I(R4743t2640) I(R4744t4074) I(R4744t172) I(R4744t718) I(R4745t80) I(R4746t1200) I(R4746t957) I(R4746t4237) I(R4746t1637) I(R4747t1228) I(R4748t4024) I(R4748t2279) I(R4748t560) I(R4749t23) I(R4749t1013) I(R4749t1338) I(R4750t401) I(R4750t2089) I(R4750t2719) I(R4750t3932) I(R4751t841) I(R4751t2368) I(R4752t153) I(R4753t1816) I(R4753t3741) I(R4754t4277) I(R4754t1063) I(R4755t1378) I(R4755t2976) I(R4755t3412) I(R4755t2867) I(R4755t4176) I(R4755t3155) I(R4756t2086) I(R4756t3081) I(R4756t3544) I(R4756t338) I(R4756t1893) I(R4757t1089) I(R4757t90) I(R4757t736) I(R4758t4074) I(R4758t4331) I(R4758t3437) I(R4759t3927) I(R4760t4411) I(R4760t1543) I(R4760t1348) I(R4760t4273) I(R4760t4692) I(R4761t2371) I(R4761t1671) I(R4761t3739) I(R4761t3453) I(R4762t2311) I(R4762t1205) I(R4763t136) I(R4763t1331) I(R4763t3495) I(R4763t2077) I(R4764t3467) I(R4764t4360) I(R4764t2190) I(R4765t1732) I(R4766t3014) I(R4766t4485) I(R4766t309) I(R4766t2044) I(R4766t4146) I(R4766t1521) I(R4767t4423) I(R4767t2567) I(R4768t3632) I(R4768t3923) I(R4768t2591) I(R4768t394) I(R4768t3022) I(R4769t2425) I(R4770t4318) I(R4770t1344) I(R4770t740) I(R4770t3850) I(R4770t2008) I(R4770t4701) I(R4771t4404) I(R4771t4504) I(R4772t3232) I(R4772t4189) I(R4772t3435) I(R4773t3699) I(R4773t550) I(R4773t373) I(R4773t1253) I(R4774t806) I(R4774t1224) I(R4774t433) I(R4774t4082) I(R4774t4355) I(R4775t2475) I(R4775t1562) I(R4776t4590) I(R4776t4383) I(R4776t1757) I(R4777t4583) I(R4777t4310) I(R4779t198) I(R4779t3787) I(R4781t1811) I(R4781t3956) I(R4782t4740) I(R4782t1651) I(R4783t3780) I(R4783t4377) I(R4783t4265) I(R4783t1980) I(R4783t1607) I(R4784t2) I(R4784t4432) I(R4784t3086) I(R4784t2782) I(R4784t2908) I(R4785t777) I(R4785t1509) I(R4786t1404) I(R4787t46) I(R4787t289) I(R4787t2996) I(R4787t1559) I(R4787t3781) I(R4788t444) I(R4788t779) I(R4788t632) I(R4788t508) I(R4788t2454) I(R4788t4217) I(R4789t3176) I(R4789t4537) I(R4789t2232) I(R4790t2988) I(R4790t3802) I(R4790t4677) I(R4790t2817) I(R4791t580) I(R4791t852) I(R4791t1476) I(R4791t1658) I(R4791t1239) I(R4792t573) I(R4792t1612) I(R4793t3113) I(R4793t1649) I(R4793t4374) I(R4794t1627) I(R4794t1240) I(R4795t2941) I(R4795t3917) I(R4796t2756) I(R4797t2977) I(R4797t3255) I(R4797t3708) I(R4797t682) I(R4797t4290) I(R4797t4487) I(R4798t4103) I(R4798t4383) I(R4798t1270) I(R4798t902) I(R4799t3273) I(R4800t1099) I(R4800t3017) I(R4800t2325) I(R4800t3887) I(R4801t254) I(R4801t4560) I(R4801t243) I(R4801t2581) I(R4801t678) I(R4801t3442) I(R4801t4162) I(R4802t689) I(R4802t2856) I(R4802t1222) I(R4803t4118) I(R4803t930) I(R4803t2833) I(R4803t1380) I(R4804t4451) I(R4804t3623) I(R4804t4100) I(R4805t2841) I(R4805t3742) I(R4805t4389) I(R4805t4392) I(R4805t3491) I(R4805t603) I(R4806t985) I(R4806t3444) I(R4806t1589) I(R4808t3761) I(R4808t1180) I(R4808t3709) I(R4810t1821) I(R4810t144) I(R4810t780) I(R4811t423) I(R4812t444) I(R4812t779) I(R4812t1083) I(R4812t1791) I(R4813t689) I(R4813t4802) I(R4813t2856) I(R4813t708) I(R4814t877) I(R4814t894) I(R4814t3612) I(R4814t3524) I(R4815t2693) I(R4815t4555) I(R4816t52) I(R4816t823) I(R4817t3292) I(R4817t4608) I(R4817t2944) I(R4818t3084) I(R4818t1600) I(R4819t1363) I(R4819t1587) I(R4820t86) I(R4820t3543) I(R4820t3375) I(R4821t3331) I(R4821t3867) I(R4821t4336) I(R4821t404) I(R4821t4430) I(R4822t590) I(R4823t4765) I(R4823t1732) I(R4823t985) I(R4823t251) I(R4824t3116) I(R4824t3460) I(R4824t2068) I(R4824t1950) I(R4825t51) I(R4826t4100) I(R4826t4131) I(R4826t3623) I(R4826t4333) I(R4826t1702) I(R4827t4427) I(R4827t1706) I(R4828t2759) I(R4828t1685) I(R4828t1575) I(R4828t2605) I(R4829t3471) I(R4829t1297) I(R4829t3346) I(R4829t3466) I(R4829t34) I(R4830t4584) I(R4830t3268) I(R4831t579) I(R4831t4393) I(R4831t414) I(R4832t948) I(R4832t4632) I(R4832t4555) I(R4832t4815) I(R4832t2693) I(R4833t1268) I(R4833t957) I(R4833t351) I(R4833t3232) I(R4835t1054) I(R4836t177) I(R4836t2981) I(R4836t3639) I(R4836t3068) I(R4836t2877) I(R4837t1974) I(R4837t2845) I(R4837t2172) I(R4837t3284) I(R4838t602) I(R4838t3664) I(R4838t3117) I(R4838t3083) I(R4839t1765) I(R4839t4008) I(R4839t1349) I(R4839t4080) I(R4839t1842) I(R4840t2021) I(R4840t4313) I(R4840t2909) I(R4840t1261) I(R4841t1287) I(R4841t2365) I(R4841t409) I(R4842t2606) I(R4842t3429) I(R4842t2882) I(R4843t88) I(R4843t817) I(R4844t4686) I(R4844t4790) I(R4845t4289) I(R4846t812) I(R4847t19) I(R4847t2313) I(R4847t2824) I(R4848t1184) I(R4849t3406) I(R4850t412) I(R4850t731) I(R4850t3108) I(R4850t1308) I(R4851t1685) I(R4851t4828) I(R4851t2759) I(R4852t3023) I(R4852t2683) I(R4852t3849) I(R4853t727) I(R4853t1458) I(R4853t2771) I(R4853t2304) I(R4854t986) I(R4854t4002) I(R4855t4384) I(R4855t1404) I(R4855t4786) I(R4856t2145) I(R4856t3904) I(R4856t476) I(R4856t3596) I(R4856t2508) I(R4856t1353) I(R4856t920) I(R4857t1304) I(R4857t2969) I(R4857t2634) I(R4857t4020) I(R4857t4022) I(R4858t1470) I(R4858t2516) I(R4858t3450) I(R4859t3900) I(R4859t709) I(R4860t3200) I(R4860t3104) I(R4860t3557) I(R4861t4404) I(R4861t2121) I(R4861t2522) I(R4862t4404) I(R4862t4771) I(R4862t2522) I(R4863t3312) I(R4863t4544) I(R4863t4005) I(R4863t4414) I(R4864t4089) I(R4864t2574) I(R4864t2230) I(R4864t1289) I(R4864t1681) I(R4865t2055) I(R4865t4446) I(R4865t250) I(R4865t3729) I(R4865t1705) I(R4866t2288) I(R4866t3533) I(R4866t237) I(R4866t4151) I(R4866t1138) I(R4867t3061) I(R4868t2722) I(R4868t3667) I(R4869t2975) I(R4869t3860) I(R4870t4642) I(R4870t4510) I(R4871t2611) I(R4872t643) I(R4872t3118) I(R4872t1785) I(R4872t2950) I(R4872t2071) I(R4873t262) I(R4873t4157) I(R4874t2429) I(R4874t1160) I(R4874t2324) I(R4875t4457) I(R4875t4717) I(R4875t2872) I(R4875t3869) I(R4875t1846) I(R4876t2620) I(R4876t1719) I(R4876t3930) I(R4876t811) I(R4876t3577) I(R4877t1991) I(R4877t1033) I(R4877t4325) I(R4878t3127) I(R4878t2630) I(R4878t1904) I(R4878t3563) I(R4879t4074) I(R4879t4744) I(R4880t1118) I(R4881t4698) I(R4881t1184) I(R4882t2891) I(R4882t2324) I(R4882t862) I(R4883t4873) I(R4883t4425) I(R4883t4215) I(R4884t1994) I(R4884t3206) I(R4884t1175) I(R4885t3412) I(R4885t3555) I(R4886t2886) I(R4886t3769) I(R4886t1745) I(R4887t2556) I(R4887t2897) I(R4888t2075) I(R4888t3264) I(R4888t210) I(R4888t4522) I(R4889t774) I(R4889t2481) I(R4890t3847) I(R4891t2092) I(R4891t2688) I(R4891t125) I(R4891t1858) I(R4892t2758) I(R4892t3299) I(R4892t2819) I(R4893t2494) I(R4893t79) I(R4894t875) I(R4894t2729) I(R4894t826) I(R4895t4461) I(R4895t627) I(R4895t292) I(R4896t378) I(R4896t272) I(R4896t584) I(R4896t1424) I(R4897t4312) I(R4897t4468) I(R4897t1781) I(R4897t2904) I(R4897t2582) I(R4898t1818) I(R4899t3243) I(R4899t2716) I(R4899t1012) I(R4900t2766) I(R4900t2539) I(R4901t2457) I(R4901t2299) I(R4901t3047) I(R4901t4435) I(R4902t3334) I(R4903t4270) I(R4903t4580) I(R4903t424) I(R4904t3511) I(R4905t2536) I(R4905t2717) I(R4906t2646) I(R4906t188) I(R4906t656) I(R4907t4047) I(R4908t3440) I(R4908t1834) I(R4908t3417) I(R4909t1238) I(R4909t3096) I(R4909t3048) I(R4910t1189) I(R4910t2448) I(R4910t137) I(R4910t2379) I(R4911t3604) I(R4912t4342) I(R4912t481) I(R4912t1977) I(R4912t1481) I(R4912t1849) I(R4912t2973) I(R4913t2708) I(R4913t281) I(R4913t1660) I(R4915t465) I(R4915t1494) I(R4916t4453) I(R4916t4455) I(R4916t32) I(R4916t4201) I(R4917t69) I(R4917t4238) I(R4917t1600) I(R4918t453) I(R4918t3845) I(R4918t1908) I(R4919t1376) I(R4920t4025) I(R4920t1065) I(R4921t688) I(R4921t3812) I(R4922t404) I(R4922t4430) I(R4923t916) I(R4923t2552) I(R4923t4223) I(R4923t4359) I(R4923t3646) I(R4923t4334) I(R4923t4123) I(R4924t4266) I(R4925t3904) I(R4925t920) I(R4925t3943) I(R4925t3900) I(R4925t4859) I(R4926t3477) I(R4926t4018) I(R4926t2728) I(R4926t166) I(R4926t1578) I(R4926t312) I(R4927t3283) I(R4927t2846) I(R4927t295) I(R4928t1080) I(R4928t1057) I(R4928t3241) I(R4928t3063) I(R4929t59) I(R4929t1405) I(R4929t463) I(R4929t275) I(R4930t2310) I(R4930t4717) I(R4930t2460) I(R4930t2971) I(R4931t2566) I(R4931t4251) I(R4931t2341) I(R4931t2883) I(R4933t790) I(R4933t4316) I(R4933t4242) I(R4934t4752) I(R4935t1463) I(R4935t2001) I(R4935t3680) I(R4935t996) I(R4935t4665) I(R4936t649) I(R4936t3204) I(R4936t404) I(R4936t4922) I(R4937t3385) I(R4937t1165) I(R4937t184) I(R4938t2264) I(R4938t2889) I(R4938t2998) I(R4939t2014) I(R4939t3817) I(R4939t2112) I(R4940t2290) I(R4940t3659) I(R4940t4378) I(R4940t617) I(R4941t987) I(R4941t3542) I(R4941t3847) I(R4941t3452) I(R4942t2321) I(R4942t2805) I(R4942t4639) I(R4942t3634) I(R4943t1535) I(R4943t2186) I(R4944t4417) I(R4945t1675) I(R4945t655) I(R4946t4794) I(R4946t1627) I(R4946t3260) I(R4946t4600) I(R4948t973) I(R4948t2403) I(R4949t2223) I(R4949t3588) I(R4949t3864) I(R4950t2885) I(R4950t2131) I(R4951t4231) I(R4951t4848) I(R4952t3649) I(R4952t2644) I(R4953t3682) I(R4953t3755) I(R4953t4221) I(R4954t78) I(R4954t3393) I(R4954t4388) I(R4954t256) I(R4954t4398) I(R4955t1483) I(R4955t4029) I(R4955t1843) I(R4955t2834) I(R4956t3596) I(R4956t4856) I(R4956t476) I(R4956t3650) I(R4957t2586) I(R4957t4593) I(R4957t2855) I(R4957t2101) I(R4957t14) I(R4958t1462) I(R4958t4366) I(R4958t2118) I(R4958t4166) I(R4958t132) I(R4959t2282) I(R4959t1972) I(R4959t2136) I(R4959t2208) I(R4960t1347) I(R4960t3355) I(R4960t1319) I(R4961t3218) I(R4961t2295) I(R4961t2699) I(R4961t4440) I(R4962t2292) I(R4962t106) I(R4962t3236) I(R4963t4004) I(R4963t2554) I(R4963t119) I(R4963t1151) I(R4963t3493) I(R4964t4323) I(R4964t1478) I(R4965t1812) I(R4965t4515) I(R4965t943) I(R4965t4102) I(R4965t3614) I(R4966t3289) I(R4967t1610) I(R4967t3664) I(R4968t3310) I(R4968t381) I(R4968t2512) I(R4969t4862) I(R4969t2522) I(R4969t3924) I(R4970t162) I(R4970t1772) I(R4970t2751) I(R4970t2679) I(R4971t3747) I(R4971t4477) I(R4971t2674) I(R4971t2473) I(R4972t2361) I(R4972t4532) I(R4972t2626) I(R4973t3857) I(R4973t887) I(R4973t3328) I(R4974t1381) I(R4974t1935) I(R4975t174) I(R4975t1322) I(R4975t3236) I(R4975t1727) I(R4976t3234) I(R4976t3651) I(R4976t1076) I(R4976t2575) I(R4977t874) I(R4977t1496) I(R4977t1845) I(R4977t3211) I(R4978t2251) I(R4978t2785) I(R4978t4809) I(R4979t832) I(R4979t2731) I(R4979t3438) I(R4980t3539) I(R4980t677) I(R4981t4104) I(R4981t2871) I(R4981t2538) I(R4981t371) I(R4981t3152) I(R4981t2740) I(R4982t1161) I(R4982t1728) I(R4982t2356) I(R4982t2387) I(R4982t706) I(R4983t1192) I(R4983t1630) I(R4983t4585) I(R4984t1177) I(R4984t3337) I(R4985t1720) I(R4985t2104) I(R4986t4069) I(R4986t903) I(R4986t4223) I(R4987t3347) I(R4987t2726) I(R4987t1621) I(R4987t1166) I(R4988t1712) I(R4988t2498) I(R4989t71) I(R4989t1380) I(R4989t4803) I(R4989t4118) I(R4989t4067) I(R4990t2756) I(R4990t4711) I(R4990t1198) I(R4990t3676) I(R4990t1764) I(R4991t3189) I(R4991t3798) I(R4991t3732) I(R4992t4367) I(R4992t2619) I(R4992t1381) I(R4993t175) I(R4993t3490) I(R4993t7) I(R4993t751) I(R4994t1216) I(R4994t3584) I(R4994t354) I(R4994t3903) I(R4995t3179) I(R4995t2749) I(R4996t2417) I(R4997t4570) I(R4997t4465) I(R4998t1997) I(R4998t3813) I(R4998t4444) I(R4999t534) I(R4999t2183) I(R4999t185) I(R5000t230) I(R5000t2947) I(R5000t3153) I(R5001t3726) I(R5001t2337) I(R5001t4615) I(R5001t2760) I(R5002t3398) I(R5002t700) I(R5002t2555) I(R5003t4915) I(R5003t4203) I(R5003t4580) I(R5004t4199) I(R5004t2215) I(R5005t107) I(R5005t4619) I(R5005t1199) I(R5005t2812) I(R5005t2878) I(R5006t3305) I(R5006t2070) I(R5006t2643) I(R5006t1186) I(R5006t530) I(R5007t2593) I(R5007t3422) I(R5008t2346) I(R5008t3538) I(R5008t651) I(R5008t1461) I(R5009t152) I(R5009t1542) I(R5009t1495) I(R5009t3089) I(R5010t2430) I(R5010t3106) I(R5010t526) I(R5010t4161) I(R5010t2048) I(R5011t3679) I(R5011t2113) I(R5011t3736) I(R5012t222) I(R5012t1844) I(R5012t3469) I(R5012t2911) I(R5012t3412) I(R5013t1449) I(R5013t264) I(R5013t4576) I(R5013t3207) I(R5013t1007) I(R5014t1391) I(R5014t1486) I(R5014t3599) I(R5015t1416) I(R5015t2906) I(R5016t4365) I(R5016t4376) I(R5016t1988) I(R5017t2146) I(R5017t4193) I(R5018t3388) I(R5018t1956) I(R5018t4186) I(R5018t1120) I(R5019t2919) I(R5019t115) I(R5020t2990) I(R5020t1399) I(R5020t2531) I(R5020t130) I(R5020t726) I(R5021t4279) I(R5021t2806) I(R5022t2386) I(R5022t3884) I(R5022t430) I(R5022t1546) I(R5022t3431) I(R5023t519) I(R5024t1560) I(R5024t4019) I(R5024t3755) I(R5024t4953) I(R5024t3682) I(R5025t111) I(R5026t4871) I(R5026t3354) I(R5027t770) I(R5027t2335) I(R5027t3023) I(R5027t3689) I(R5028t784) I(R5028t1602) I(R5028t3980) I(R5029t4218) I(R5029t4081) I(R5030t3914) I(R5030t3152) I(R5030t2740) I(R5031t1411) I(R5031t4282) I(R5031t2880) I(R5032t2659) I(R5033t290) I(R5033t1238) I(R5033t3252) I(R5033t1340) I(R5034t118) I(R5034t3515) I(R5034t144) I(R5034t4810) I(R5034t1821) I(R5035t450) I(R5035t3918) I(R5036t997) I(R5036t80) I(R5037t346) I(R5037t4721) I(R5037t1240) I(R5037t4443) I(R5037t3734) I(R5038t179) I(R5039t531) I(R5039t2857) I(R5039t101) I(R5040t1258) I(R5040t3240) I(R5040t1506) I(R5040t124) I(R5041t718) I(R5041t2459) I(R5041t1248) I(R5042t2648) I(R5042t910) I(R5042t1851) I(R5042t3448) I(R5043t2162) I(R5043t2517) I(R5043t1740) I(R5043t2088) I(R5044t4752) I(R5044t153) I(R5045t1544) I(R5045t3361) I(R5045t2712) I(R5046t1696) I(R5046t3339) I(R5047t3450) I(R5047t4099) I(R5047t3315) I(R5048t4157) I(R5048t3134) I(R5049t263) I(R5049t3212) I(R5049t3237) I(R5049t702) I(R5049t2363) I(R5050t1387) I(R5051t698) I(R5051t3974) I(R5051t1094) I(R5052t1624) I(R5052t2854) I(R5052t4292) I(R5052t4319) I(R5053t4843) I(R5053t14) I(R5053t817) I(R5054t1896) I(R5054t4056) I(R5054t25) I(R5055t1333) I(R5055t1685) I(R5055t1988) I(R5055t1032) I(R5056t3231) I(R5056t417) I(R5056t3144) I(R5057t1706) I(R5057t4827) I(R5057t4427) I(R5057t1459) I(R5057t3766) I(R5058t744) I(R5058t2631) I(R5059t1360) I(R5059t4128) I(R5060t3599) I(R5060t3969) I(R5060t5014) I(R5060t3773) I(R5060t4421) I(R5061t265) I(R5061t1558) I(R5061t1684) I(R5062t1955) I(R5062t1049) I(R5062t2499) I(R5062t3836) I(R5062t4498) I(R5063t2990) I(R5063t3134) I(R5063t283) I(R5064t3870) I(R5064t2894) I(R5064t2897) I(R5064t4887) I(R5065t2505) I(R5065t1080) I(R5065t4928) I(R5066t421) I(R5066t1219) I(R5066t616) I(R5067t2703) I(R5067t4258) I(R5067t2486) I(R5067t2160) I(R5068t1274) I(R5068t2221) I(R5068t4101) I(R5069t4366) I(R5069t4958) I(R5069t132) I(R5070t3927) I(R5070t895) I(R5071t446) I(R5071t4299) I(R5071t4661) I(R5071t1800) I(R5071t1982) I(R5072t1721) I(R5072t4368) I(R5072t1576) I(R5073t1183) I(R5073t3239) I(R5074t3764) I(R5074t159) I(R5075t541) I(R5075t2573) I(R5075t859) I(R5075t3321) I(R5075t1503) I(R5075t2011) I(R5076t1769) I(R5076t3456) I(R5077t1891) I(R5077t3270) I(R5077t2557) I(R5078t110) I(R5078t4854) I(R5078t4002) I(R5079t4090) I(R5079t1540) I(R5080t548) I(R5080t2843) I(R5080t891) I(R5080t2473) I(R5081t4162) I(R5081t4560) I(R5081t3634) I(R5081t3348) I(R5081t2057) I(R5081t3866) I(R5082t3320) I(R5082t2081) I(R5083t305) I(R5083t2449) I(R5083t1934) I(R5084t3205) I(R5084t11) I(R5084t1015) I(R5084t3987) I(R5085t3737) I(R5085t1381) I(R5085t4992) I(R5086t3833) I(R5086t4433) I(R5087t2585) I(R5087t965) I(R5088t416) I(R5088t4465) I(R5088t1057) I(R5088t1897) I(R5089t4031) I(R5089t2150) I(R5089t3995) I(R5090t2993) I(R5090t4681) I(R5090t267) I(R5090t2371) I(R5090t4761) I(R5090t3905) I(R5090t1960) I(R5091t3318) I(R5091t1043) I(R5091t4537) I(R5091t4789) I(R5091t3176) I(R5091t2504) I(R5092t4794) I(R5092t1240) I(R5092t1034) I(R5093t2399) I(R5095t2914) I(R5095t4696) I(R5095t606) I(R5096t1951) I(R5096t3031) I(R5096t4229) I(R5097t113) I(R5097t2621) I(R5098t1739) I(R5099t329) I(R5099t2284) I(R5100t847) I(R5100t1715) I(R5100t3509) I(R5100t3752) I(R5101t1298) I(R5101t788) I(R5101t1649) I(R5101t4793) I(R5102t2924) I(R5102t4311) I(R5102t1821) I(R5102t1795) I(R5103t5059) I(R5103t1616) I(R5103t4556) I(R5103t1292) I(R5103t4128) I(R5104t1712) I(R5104t1349) I(R5104t4080) I(R5104t4988) I(R5105t2045) I(R5105t3343) I(R5105t3771) I(R5107t3114) I(R5107t4422) I(R5108t842) I(R5108t3554) I(R5108t1466) I(R5108t102) I(R5109t1257) I(R5109t2910) I(R5109t3832) I(R5110t3534) I(R5110t818) I(R5110t3837) I(R5110t2546) I(R5111t3126) I(R5112t1496) I(R5112t4977) I(R5112t4014) I(R5113t1582) I(R5113t771) I(R5113t3735) I(R5113t2067) I(R5114t1906) I(R5114t913) I(R5115t2161) I(R5117t3921) I(R5117t4070) I(R5117t4284) I(R5118t1014) I(R5118t2666) I(R5118t511) I(R5118t1241) I(R5118t557) I(R5119t1416) I(R5119t3267) I(R5119t5015) I(R5120t3486) I(R5121t2447) I(R5122t414) I(R5123t955) I(R5123t4275) I(R5123t809) I(R5123t2521) I(R5123t1357) I(R5124t1105) I(R5124t3377) I(R5125t3450) I(R5125t4099) I(R5125t307) I(R5126t3447) I(R5126t2094) I(R5126t3806) I(R5126t4638) I(R5127t4269) I(R5127t3766) I(R5127t358) I(R5128t4283) I(R5129t2743) I(R5130t2970) I(R5130t2968) I(R5130t3055) I(R5130t3098) I(R5131t2672) I(R5131t3596) I(R5131t1170) I(R5131t269) I(R5131t3119) I(R5132t178) I(R5132t4781) I(R5132t1811) I(R5133t4722) I(R5133t2489) I(R5133t2488) I(R5134t2262) I(R5134t2602) I(R5134t356) I(R5134t4293) I(R5135t4535) I(R5135t1397) I(R5135t2813) I(R5135t476) I(R5136t2733) I(R5137t1203) I(R5138t1786) I(R5138t4628) I(R5138t1102) I(R5139t2442) I(R5139t2935) I(R5139t2214) I(R5139t4340) I(R5140t989) I(R5141t1071) I(R5141t2927) I(R5142t2209) I(R5142t2578) I(R5142t3025) I(R5142t1766) I(R5142t1127) I(R5142t94) I(R5143t2737) I(R5143t717) I(R5143t1667) I(R5143t1106) I(R5143t4278) I(R5143t963) I(R5144t1604) I(R5144t1680) I(R5144t2114) I(R5145t4679) I(R5145t4500) I(R5146t2705) I(R5146t4025) I(R5146t4265) I(R5147t1182) I(R5147t2722) I(R5147t4868) I(R5147t3667) I(R5148t1095) I(R5148t319) I(R5149t2417) I(R5149t3983) I(R5149t2544) I(R5150t371) I(R5150t3152) I(R5151t3338) I(R5152t2306) I(R5152t1827) I(R5152t4034) I(R5153t3928) I(R5153t2673) I(R5153t2921) I(R5153t3656) I(R5154t1991) I(R5154t4877) I(R5154t4325) I(R5155t2612) I(R5155t2644) I(R5155t1861) I(R5156t625) I(R5156t818) I(R5157t2436) I(R5157t449) I(R5158t1470) I(R5158t4858) I(R5159t3431) I(R5159t2587) I(R5159t2263) I(R5159t217) I(R5160t1013) I(R5160t4749) I(R5160t4116) I(R5160t1338) I(R5161t4204) I(R5161t217) I(R5161t5159) I(R5162t642) I(R5162t2082) I(R5162t1088) I(R5162t3938) I(R5162t3082) I(R5163t761) I(R5163t2840) I(R5163t1421) I(R5164t3698) I(R5164t3853) I(R5164t907) I(R5164t4357) I(R5164t2802) I(R5164t251) I(R5164t4823) I(R5165t2733) I(R5165t451) I(R5166t129) I(R5166t3822) I(R5166t2330) I(R5167t1168) I(R5167t2608) I(R5167t3972) I(R5167t2156) I(R5168t4324) I(R5169t2996) I(R5169t1965) I(R5170t294) I(R5170t4551) I(R5170t2359) I(R5171t372) I(R5171t4424) I(R5171t3434) I(R5171t318) I(R5172t3280) I(R5172t2093) I(R5172t2678) I(R5173t1038) I(R5173t4155) I(R5174t598) I(R5174t790) I(R5174t635) I(R5174t1113) I(R5174t1434) I(R5175t1524) I(R5175t3485) I(R5175t43) I(R5175t3892) I(R5176t2062) I(R5176t1676) I(R5177t1140) I(R5177t2945) I(R5177t3376) I(R5178t2710) I(R5178t1384) I(R5178t654) I(R5179t2233) I(R5179t2757) I(R5179t4704) I(R5179t1809) I(R5180t3504) I(R5180t4481) I(R5180t1901) I(R5181t4881) I(R5181t128) I(R5181t3818) I(R5182t1109) I(R5182t2995) I(R5182t2690) I(R5183t1899) I(R5183t4947) I(R5184t727) I(R5184t2702) I(R5184t1458) I(R5184t4853) I(R5185t1693) I(R5185t2332) I(R5185t2226) I(R5185t2336) I(R5186t2421) I(R5186t3032) I(R5186t4408) I(R5186t3247) I(R5187t2315) I(R5187t2094) I(R5188t4962) I(R5188t3236) I(R5188t3989) I(R5189t3935) I(R5190t978) I(R5190t4505) I(R5190t4037) I(R5191t1351) I(R5191t4106) I(R5191t25) I(R5193t1487) I(R5193t3901) I(R5193t4276) I(R5194t4303) I(R5194t3713) I(R5195t2025) I(R5195t691) I(R5195t1115) I(R5195t1150) I(R5196t3429) I(R5196t891) I(R5196t2473) I(R5196t4971) I(R5196t2674) I(R5196t1187) I(R5196t1623) I(R5197t2035) I(R5197t4635) I(R5198t2349) I(R5198t3996) I(R5199t2169) I(R5199t4334) I(R5199t523) I(R5200t81) I(R5200t311) I(R5200t2180) I(R5201t1128) I(R5201t1469) I(R5202t3069) I(R5202t801) I(R5202t3724) I(R5203t2825) I(R5203t2531) I(R5203t1730) I(R5203t794) I(R5203t1784) I(R5204t2845) I(R5204t4837) I(R5204t1615) I(R5204t2172) I(R5205t1444) I(R5205t653) I(R5206t3896) I(R5206t3852) I(R5207t182) I(R5207t2705) I(R5207t5146) I(R5207t4025) I(R5208t3343) I(R5208t4030) I(R5210t1514) I(R5210t2416) I(R5210t1140) I(R5210t3633) I(R5211t1554) I(R5211t3313) I(R5211t3988) I(R5212t2527) I(R5212t1711) I(R5212t2549) I(R5213t3542) I(R5213t4941) I(R5213t3452) I(R5214t717) I(R5214t4049) I(R5214t4390) I(R5214t2737) I(R5214t5143) I(R5215t274) I(R5215t892) I(R5215t3914) I(R5215t3152) I(R5216t1955) I(R5216t3126) I(R5216t5111) I(R5216t4464) I(R5217t250) I(R5217t2055) I(R5217t3241) I(R5217t3063) I(R5217t448) I(R5217t3523) I(R5218t285) I(R5218t2132) I(R5218t1611) I(R5218t4524) I(R5219t2376) I(R5220t4273) I(R5220t5034) I(R5220t118) I(R5220t4073) I(R5221t4502) I(R5221t2383) I(R5221t3715) I(R5221t1108) I(R5222t1913) I(R5222t3377) I(R5222t5124) I(R5222t1105) I(R5222t3470) I(R5222t1618) I(R5223t1145) I(R5223t4332) I(R5223t1388) I(R5223t1572) I(R5223t3797) I(R5224t2621) I(R5224t507) I(R5224t4544) I(R5225t1403) I(R5226t1013) I(R5226t516) I(R5227t1444) I(R5227t5205) I(R5228t997) I(R5228t4966) I(R5229t1750) I(R5229t4811) I(R5230t424) I(R5230t4903) I(R5230t4580) I(R5230t4203) I(R5230t4735) I(R5231t1965) I(R5231t5169) I(R5232t2159) I(R5232t3842) I(R5232t451) I(R5232t3964) I(R5233t1483) I(R5233t4955) I(R5233t1843) I(R5233t2689) I(R5233t691) I(R5234t1740) I(R5234t2517) I(R5234t2054) I(R5234t4402) I(R5235t1296) I(R5235t5004) I(R5235t2215) I(R5235t330) I(R5236t555) I(R5236t3397) I(R5237t4552) I(R5237t1555) I(R5237t670) I(R5238t3611) I(R5238t4276) I(R5238t5193) I(R5239t3422) I(R5239t2816) I(R5239t542) I(R5240t3139) I(R5240t3061) I(R5241t1669) I(R5241t2494) I(R5241t4893) I(R5241t4212) I(R5242t2273) I(R5242t93) I(R5242t3500) I(R5243t2980) I(R5245t2164) I(R5245t2828) I(R5245t3197) I(R5245t3413) I(R5246t1139) I(R5246t4927) I(R5246t1350) I(R5246t3818) I(R5247t4538) I(R5247t3040) I(R5247t4119) I(R5248t1367) I(R5248t3590) I(R5248t1237) I(R5249t2309) I(R5249t3313) I(R5249t3800) I(R5249t4656) I(R5250t2505) I(R5250t3258) I(R5250t5065) I(R5250t10) I(R5251t1982) I(R5251t5071) I(R5251t988) I(R5252t2521) I(R5252t1357) I(R5253t561) I(R5253t2919) I(R5253t3205) I(R5253t5084) I(R5253t11) I(R5254t3699) I(R5255t1151) I(R5255t4963) I(R5255t580) I(R5255t271) I(R5255t119) I(R5256t4083) I(R5256t4726) I(R5256t2862) I(R5256t4947) I(R5257t2618) I(R5258t830) I(R5259t277) I(R5259t1538) I(R5260t620) I(R5260t933) I(R5261t4944) I(R5262t3970) I(R5262t26) I(R5262t2409) I(R5263t2322) I(R5263t227) I(R5264t907) I(R5264t2802) I(R5264t3998) I(R5264t1948) I(R5264t638) I(R5264t1181) I(R5265t3909) I(R5265t3203) I(R5265t2369) I(R5266t2664) I(R5266t96) I(R5266t3527) I(R5267t5261) I(R5267t4944) I(R5268t4567) I(R5268t4222) I(R5269t2591) I(R5269t4625) I(R5269t4006) I(R5269t4699) I(R5269t70) I(R5269t4092) I(R5270t2414) I(R5270t1291) I(R5270t1737) I(R5270t3363) I(R5270t1936) I(R5271t2357) I(R5271t3006) I(R5272t407) I(R5272t4311) I(R5272t2924) I(R5273t904) I(R5273t2323) I(R5274t55) I(R5274t613) I(R5274t4192) I(R5274t4670) I(R5274t4178) I(R5274t2102) I(R5275t4753) I(R5276t4131) I(R5276t3522) I(R5276t4100) I(R5277t2379) I(R5277t1689) I(R5278t1710) I(R5278t1952) I(R5278t486) I(R5278t1465) I(R5278t4302) I(R5278t3387) I(R5278t3696) I(R5279t4255) I(R5279t2665) I(R5279t2189) I(R5280t369) I(R5280t4279) I(R5280t1561) I(R5281t2825) I(R5281t5203) I(R5281t1784) I(R5282t2015) I(R5282t1082) I(R5282t4210) I(R5282t1577) I(R5283t5231) I(R5283t1559) I(R5283t1965) I(R5284t772) I(R5284t385) I(R5285t2180) I(R5285t5200) I(R5285t81) I(R5286t3724) I(R5286t1265) I(R5286t4088) I(R5286t2253) I(R5287t2013) I(R5287t2307) I(R5287t3745) I(R5287t2762) I(R5287t2866) I(R5288t2631) I(R5288t5058) I(R5288t4098) I(R5289t1337) I(R5290t452) I(R5290t2853) I(R5290t762) I(R5291t3847) I(R5291t3325) I(R5291t987) I(R5291t4941) I(R5293t4324) I(R5293t3390) I(R5294t4039) I(R5294t1810) I(R5294t1539) I(R5294t3872) I(R5295t1183) I(R5295t5073) I(R5295t2570) I(R5295t3239) I(R5296t1611) I(R5296t2327) I(R5296t771) I(R5296t969) I(R5296t2132) I(R5297t3887) I(R5297t4800) I(R5298t1493) I(R5298t3522) I(R5298t1563) I(R5299t4398) I(R5299t256) I(R5300t4406) I(R5300t1138) I(R5301t2856) I(R5302t2410) I(R5302t1410) I(R5302t253) I(R5303t1721) I(R5303t4368) I(R5303t2942) I(R5304t205) I(R5304t2893) I(R5304t3777) I(R5305t1939) I(R5305t3327) I(R5305t3654) I(R5306t2373) I(R5306t2081) I(R5306t2363) I(R5306t263) I(R5307t915) I(R5307t1254) I(R5307t917) I(R5308t2752) I(R5308t585) I(R5308t1355) I(R5309t4244) I(R5309t2766) I(R5310t4849) I(R5310t3406) I(R5310t2583) I(R5310t2115) I(R5311t1070) I(R5311t537) I(R5311t1634) I(R5311t865) I(R5312t4675) I(R5312t3636) I(R5313t3751) I(R5314t2334) I(R5314t3671) I(R5314t4558) I(R5315t2963) I(R5315t1455) I(R5315t4156) I(R5316t470) I(R5316t5038) I(R5316t179) I(R5316t3715) I(R5316t2383) I(R5317t2970) I(R5317t532) I(R5317t1569) I(R5317t3635) I(R5318t529) I(R5318t2051) I(R5318t4011) I(R5318t2062) I(R5318t5176) I(R5318t242) I(R5319t2513) I(R5319t4264) I(R5319t3719) I(R5319t438) I(R5320t3612) I(R5320t65) I(R5320t3851) I(R5321t183) I(R5321t1235) I(R5322t2323) I(R5322t5273) I(R5322t2474) I(R5322t4702) I(R5323t2117) I(R5323t664) I(R5324t3026) I(R5324t4848) I(R5325t3106) I(R5326t1824) I(R5326t3720) I(R5326t4683) I(R5326t3367) I(R5327t2826) I(R5327t2083) I(R5327t3109) I(R5327t4310) I(R5328t2239) I(R5328t2366) I(R5328t2920) I(R5328t3631) I(R5329t187) I(R5329t3382) I(R5329t4924) I(R5330t1787) I(R5330t3232) I(R5330t4189) I(R5331t2431) I(R5332t2854) I(R5333t21) I(R5333t4678) I(R5333t2699) I(R5333t2295) I(R5334t2634) I(R5334t4020) I(R5334t1186) I(R5334t4478) I(R5335t1747) I(R5335t3615) I(R5336t1712) I(R5336t5104) I(R5336t1349) I(R5336t258) I(R5337t1325) I(R5337t2078) I(R5337t1915) I(R5338t2919) I(R5338t5253) I(R5338t11) I(R5338t115) I(R5338t5019) I(R5339t4086) I(R5339t4983) I(R5340t640) I(R5340t1571) I(R5340t3603) I(R5341t2501) I(R5341t3020) I(R5341t1113) I(R5341t4469) I(R5342t3815) I(R5342t5290) I(R5342t762) I(R5342t436) I(R5343t588) I(R5343t2490) I(R5344t1937) I(R5344t193) I(R5345t1552) I(R5345t4504) I(R5345t4771) I(R5346t3802) I(R5346t4677) I(R5346t8) I(R5347t180) I(R5347t4027) I(R5347t1564) I(R5348t1563) I(R5348t4868) I(R5349t5315) I(R5349t1455) I(R5349t4274) I(R5350t4497) I(R5350t4514) I(R5352t4759) I(R5352t2792) I(R5353t1621) I(R5353t4041) I(R5353t4564) I(R5353t3846) I(R5354t1436) I(R5354t4229) I(R5355t2642) I(R5355t7) I(R5355t4993) I(R5355t5023) I(R5356t1948) I(R5356t3998) I(R5356t5264) I(R5357t2787) I(R5357t2994) I(R5357t3059) I(R5357t962) I(R5358t2643) I(R5358t4020) I(R5358t1675) I(R5359t3405) I(R5359t3054) I(R5359t3572) I(R5360t3924) I(R5360t2522) I(R5361t1492) I(R5362t3086) I(R5362t741) I(R5362t3814) I(R5362t1204) I(R5363t3565) I(R5363t4550) I(R5363t3959) I(R5363t1979) I(R5364t3575) I(R5364t3707) I(R5364t2926) I(R5364t2093) I(R5364t1423) I(R5365t4822) I(R5365t4397) I(R5365t1232) I(R5366t1695) I(R5366t1041) I(R5368t971) I(R5368t2552) I(R5368t4223) I(R5368t4986) I(R5369t1364) I(R5369t2915) I(R5370t2051) I(R5370t2595) I(R5370t1252) I(R5370t4011) I(R5370t5318) I(R5371t2114) I(R5372t4149) I(R5372t4150) I(R5372t3873) I(R5372t2158) I(R5373t2131) I(R5373t3978) I(R5374t1836) I(R5374t3895) I(R5374t998) I(R5374t76) I(R5374t2975) I(R5374t4869) I(R5374t3860) I(R5374t3672) I(R5374t108) I(R5375t696) I(R5375t1079) I(R5375t4019) I(R5375t64) I(R5375t4528) I(R5377t214) I(R5377t3537) I(R5377t3474) I(R5378t5261) I(R5379t3715) I(R5379t5316) I(R5379t1313) I(R5379t236) I(R5379t179) I(R5380t3689) I(R5380t3002) I(R5380t1626) I(R5381t882) I(R5381t4696) I(R5381t2034) I(R5382t2994) I(R5382t2563) I(R5383t3188) I(R5383t3452) I(R5383t4479) I(R5384t2213) I(R5384t339) I(R5384t4063) I(R5385t1243) I(R5385t748) I(R5385t3550) I(R5386t1261) I(R5386t4249) I(R5387t3348) I(R5387t1018) I(R5387t2057) I(R5387t5081) I(R5388t826) I(R5388t3946) I(R5388t2508) I(R5388t2278) I(R5388t4349) I(R5389t3196) I(R5389t3203) I(R5389t4280) I(R5389t885) I(R5390t3720) I(R5390t646) I(R5390t1644) I(R5391t1228) I(R5391t2465) I(R5391t3688) I(R5391t2519) I(R5392t2208) I(R5392t2622) I(R5393t3767) I(R5393t3917) I(R5394t1005) I(R5394t3379) I(R5394t1885) I(R5395t943) I(R5395t4639) I(R5395t4296) I(R5395t2805) I(R5395t3445) I(R5395t4268) I(R5396t4385) I(R5396t210) I(R5397t2994) I(R5397t5382) I(R5397t3059) I(R5397t5357) I(R5398t497) I(R5399t423) I(R5399t1360) I(R5399t65) I(R5399t2929) I(R5399t3336) I(R5400t1039) I(R5400t3074) I(R5400t2163) I(R5400t3655) I(R5400t674) I(R5401t2298) I(R5401t3595) I(R5401t3868) I(R5402t5360) I(R5402t3924) I(R5402t3819) I(R5402t4104) I(R5403t74) I(R5403t841) I(R5403t3809) I(R5404t4253) I(R5404t3563) I(R5404t939) I(R5404t3414) I(R5405t371) I(R5405t2538) I(R5405t5150) I(R5405t2901) I(R5406t1801) I(R5406t2768) I(R5406t1631) I(R5406t1214) I(R5407t605) I(R5407t4379) I(R5407t2297) I(R5407t4736) I(R5407t683) I(R5407t551) I(R5408t1952) I(R5408t4013) I(R5408t326) I(R5409t1333) I(R5409t5055) I(R5409t2759) I(R5409t4851) I(R5409t1685) I(R5410t5169) I(R5410t1965) I(R5410t4723) I(R5410t5106) I(R5411t2646) I(R5411t4650) I(R5411t3806) I(R5411t4583) I(R5411t656) I(R5411t4906) I(R5412t408) I(R5412t3888) I(R5413t2215) I(R5413t5004) I(R5413t4199) I(R5413t2224) I(R5414t139) I(R5414t1747) I(R5414t3974) I(R5414t2815) I(R5415t3145) I(R5415t4381) I(R5416t3633) I(R5416t3882) I(R5417t2013) I(R5417t3745) I(R5417t3080) I(R5418t2634) I(R5418t4857) I(R5418t4143) I(R5418t834) I(R5418t1874) I(R5419t3935) I(R5419t5189) I(R5419t2857) I(R5420t1636) I(R5420t3013) I(R5420t2812) I(R5420t5005) I(R5420t2878) I(R5421t3082) I(R5421t5162) I(R5421t3938) I(R5421t1088) I(R5422t1372) I(R5422t2954) I(R5422t3129) I(R5423t1369) I(R5423t1993) I(R5423t2612) I(R5423t1365) I(R5424t2137) I(R5424t3354) I(R5424t5026) I(R5425t939) I(R5425t1230) I(R5426t2462) I(R5428t3414) I(R5428t4253) I(R5428t3032) I(R5429t2394) I(R5430t2240) I(R5430t694) I(R5430t2105) I(R5431t1803) I(R5431t3920) I(R5431t1716) I(R5431t3240) I(R5431t5040) I(R5432t3933) I(R5432t4443) I(R5432t3981) I(R5433t2889) I(R5433t4938) I(R5434t2273) I(R5434t3910) I(R5434t851) I(R5434t3500) I(R5435t2941) I(R5435t4480) I(R5435t2859) I(R5435t4795) I(R5436t1366) I(R5436t5245) I(R5436t3413) I(R5436t4439) I(R5436t741) I(R5437t40) I(R5437t1688) I(R5438t1268) I(R5438t4522) I(R5438t1787) I(R5438t2598) I(R5438t3232) I(R5438t4833) I(R5439t1135) I(R5441t111) I(R5441t5025) I(R5442t2747) I(R5442t2982) I(R5442t704) I(R5442t1212) I(R5442t3767) I(R5443t1089) I(R5443t4757) I(R5443t736) I(R5443t2920) I(R5444t1024) I(R5444t2985) I(R5444t1036) I(R5444t2199) I(R5444t19) I(R5445t3933) I(R5445t2593) I(R5445t5007) I(R5445t3981) I(R5445t5432) I(R5446t1362) I(R5446t2790) I(R5446t2636) I(R5447t2684) I(R5447t915) I(R5447t4950) I(R5448t2097) I(R5448t893) I(R5448t2010) I(R5448t4228) I(R5449t1116) I(R5449t4543) I(R5449t2896) I(R5450t782) I(R5450t4914) I(R5451t848) I(R5451t1769) I(R5451t4718) I(R5451t1056) I(R5451t3301) I(R5451t2287) I(R5452t4151) I(R5452t2585) I(R5452t4866) I(R5453t5041) I(R5453t3142) I(R5453t1220) I(R5453t2080) I(R5453t1248) I(R5454t3298) I(R5454t5324) I(R5454t4848) I(R5454t1184) I(R5454t4881) I(R5455t262) I(R5455t4873) I(R5455t3638) I(R5455t4425) I(R5455t4883) I(R5456t3172) I(R5456t2711) I(R5456t3592) I(R5456t3782) I(R5456t4732) I(R5457t1859) I(R5457t4239) I(R5457t835) I(R5457t135) I(R5458t2843) I(R5459t3548) I(R5459t5019) I(R5460t815) I(R5460t4679) I(R5461t3387) I(R5461t3696) I(R5461t2069) I(R5461t4171) I(R5461t2137) I(R5462t4452) I(R5463t5309) I(R5463t2766) I(R5463t4900) I(R5463t4012) I(R5464t5173) I(R5464t4155) I(R5464t3314) I(R5464t4188) I(R5465t2083) I(R5465t5327) I(R5465t2399) I(R5466t699) I(R5466t2913) I(R5466t532) I(R5466t3997) I(R5467t766) I(R5467t1579) I(R5467t2065) I(R5467t3495) I(R5467t4023) I(R5468t447) I(R5468t4648) I(R5468t1321) I(R5468t4209) I(R5469t4482) I(R5469t1090) I(R5470t2675) I(R5470t3465) I(R5470t2713) I(R5470t5106) I(R5470t775) I(R5471t408) I(R5471t5412) I(R5471t3888) I(R5471t1046) I(R5472t89) I(R5472t3416) I(R5472t1648) I(R5472t1110) I(R5473t1859) I(R5473t5457) I(R5473t4239) I(R5474t4226) I(R5474t4445) I(R5474t442) I(R5475t3872) I(R5475t1539) I(R5475t662) I(R5476t992) I(R5476t3192) I(R5476t5387) I(R5477t515) I(R5477t3823) I(R5477t4058) I(R5478t1095) I(R5478t4407) I(R5478t4486) I(R5479t5422) I(R5479t2954) I(R5479t4297) I(R5479t2942) I(R5479t5303) I(R5480t4300) I(R5480t1072) I(R5480t3018) I(R5481t922) I(R5481t4669) I(R5481t5423) I(R5481t3661) I(R5482t3316) I(R5483t1670) I(R5483t2247) I(R5483t2871) I(R5483t1084) I(R5483t2506) I(R5484t3367) I(R5484t4683) I(R5484t3185) I(R5485t4267) I(R5485t4762) I(R5486t322) I(R5486t4329) I(R5487t5137) I(R5488t4461) I(R5488t1087) I(R5488t1134) I(R5489t459) I(R5489t3602) I(R5489t4173) I(R5489t2660) I(R5490t4362) I(R5490t4616) I(R5490t3796) I(R5490t1650) I(R5491t305) I(R5491t5083) I(R5491t570) I(R5491t3531) I(R5492t4082) I(R5492t3479) I(R5492t2628) I(R5493t5300) I(R5493t1531) I(R5493t1609) I(R5494t3571) I(R5494t3289) I(R5495t4511) I(R5495t2637) I(R5495t3636) I(R5496t26) I(R5496t819) I(R5496t5262) I(R5496t3970) I(R5496t3208) I(R5497t456) I(R5497t3569) I(R5497t457) I(R5497t58) I(R5498t4907) I(R5498t4047) I(R5498t4128) I(R5499t3213) I(R5499t4158) I(R5499t3145) I(R5499t2172) I(R5499t3877) I(R5500t3221) I(R5500t4184) I(R5500t3546) I(R5501t1319) I(R5501t4087) I(R5502t1841) I(R5502t774) I(R5502t4889) I(R5502t2481) I(R5503t1037) I(R5503t4202) I(R5504t2720) I(R5504t4198) I(R5504t329) I(R5504t3474) I(R5504t214) I(R5506t2881) I(R5506t2936) I(R5506t3614) I(R5507t3581) I(R5507t3071) I(R5507t1369) I(R5508t2322) I(R5508t5263) I(R5508t518) I(R5508t1762) I(R5509t1099) I(R5509t3017) I(R5510t3159) I(R5510t368) I(R5511t3062) I(R5511t3629) I(R5512t2463) I(R5512t4633) I(R5512t1697) I(R5512t3741) I(R5512t4753) I(R5512t5275) I(R5513t1068) I(R5513t2556) I(R5513t4887) I(R5513t5064) I(R5513t3870) I(R5514t3393) I(R5514t4585) I(R5514t2875) I(R5515t2783) I(R5515t3995) I(R5515t5089) I(R5515t4031) I(R5515t2255) I(R5515t4164) I(R5515t2624) I(R5515t4304) I(R5516t152) I(R5516t5009) I(R5516t1542) I(R5516t4579) I(R5517t4563) I(R5517t2065) I(R5517t5467) I(R5517t3495) I(R5518t5097) I(R5518t113) I(R5518t1355) I(R5518t585) I(R5519t4312) I(R5519t4468) I(R5519t578) I(R5519t4503) I(R5519t341) I(R5519t2582) I(R5520t2658) I(R5520t1714) I(R5520t4903) I(R5521t500) I(R5521t1829) I(R5521t2119) I(R5522t2914) I(R5522t382) I(R5522t606) I(R5523t1376) I(R5524t2958) I(R5524t4335) I(R5525t410) I(R5525t4144) I(R5525t4952) I(R5526t4007) I(R5526t3820) I(R5527t733) I(R5527t2007) I(R5527t3458) I(R5527t564) I(R5527t6) I(R5527t799) I(R5527t2016) I(R5528t4328) I(R5528t1043) I(R5528t5091) I(R5528t3318) I(R5528t519) I(R5529t1213) I(R5529t2712) I(R5529t5045) I(R5529t2699) I(R5529t5333) I(R5529t4678) I(R5530t4240) I(R5530t807) I(R5530t4947) I(R5531t4104) I(R5531t4981) I(R5531t2871) I(R5531t2247) I(R5531t3819) I(R5531t5402) I(R5532t722) I(R5532t4796) I(R5533t2367) I(R5533t676) I(R5534t3081) I(R5534t2086) I(R5535t970) I(R5535t2455) I(R5536t1341) I(R5536t2864) I(R5536t1231) I(R5536t5121) I(R5537t852) I(R5537t3846) I(R5537t2613) I(R5537t31) I(R5537t589) I(R5538t667) I(R5539t667) I(R5539t1220) I(R5539t3142) I(R5539t5453) I(R5540t2217) I(R5540t2940) I(R5540t663) I(R5540t984) I(R5540t4533) I(R5541t2832) I(R5541t3507) I(R5541t4568) I(R5541t4501) I(R5542t2165) I(R5542t782) I(R5542t5450) I(R5542t4808) I(R5542t3761) I(R5543t3012) I(R5543t1277) I(R5543t4341) I(R5544t3968) I(R5544t4804) I(R5544t2152) I(R5544t3578) I(R5544t3033) I(R5545t3253) I(R5545t757) I(R5545t3127) I(R5545t4250) I(R5546t3714) I(R5547t687) I(R5547t4646) I(R5548t888) I(R5549t1760) I(R5549t1962) I(R5549t2142) I(R5550t447) I(R5550t3184) I(R5550t1121) I(R5550t4648) I(R5551t4508) I(R5551t3049) I(R5552t606) I(R5552t2437) I(R5552t4742) I(R5552t382) I(R5554t1941) I(R5554t2228) I(R5554t3077) I(R5555t1319) I(R5555t5501) I(R5555t4960) I(R5555t1117) I(R5555t4087) I(R5556t3348) I(R5556t5387) I(R5556t1018) I(R5556t2444) I(R5557t4879) I(R5557t4744) I(R5557t718) I(R5557t1248) I(R5557t2080) I(R5557t327) I(R5558t4104) I(R5558t1281) I(R5559t4434) I(R5559t5521) I(R5559t2119) I(R5560t3298) I(R5560t5454) I(R5560t3222) I(R5560t3026) I(R5560t5324) I(R5561t2672) I(R5561t1851) I(R5562t3271) I(R5562t614) I(R5563t4261) I(R5563t3486) I(R5563t5120) I(R5564t15) I(R5564t2264) I(R5564t4938) I(R5564t2231) I(R5564t1975) I(R5565t5151) I(R5566t310) I(R5566t1472) I(R5566t1869) I(R5566t4602) I(R5567t4745) I(R5567t945) I(R5567t2059) I(R5568t1112) I(R5568t1168) I(R5568t2458) I(R5568t5482) I(R5569t3782) I(R5569t3592) I(R5569t5456) I(R5571t1701) I(R5571t2989) I(R5571t2947) I(R5572t4932) I(R5572t4032) I(R5572t1389) I(R5572t4218) I(R5573t1167) I(R5574t2754) I(R5574t4607) I(R5575t4826) I(R5575t2732) I(R5575t1553) I(R5576t3445) I(R5576t4268) I(R5576t3178) I(R5577t3200) I(R5577t4860) I(R5577t2654) I(R5578t4997) I(R5578t4570) I(R5579t2374) I(R5579t1479) I(R5580t1926) I(R5580t1396) I(R5580t636) I(R5580t3538) I(R5581t3101) I(R5581t5138) I(R5581t4628) I(R5581t395) I(R5581t1011) I(R5582t4397) I(R5582t3651) I(R5582t4351) I(R5582t1075) I(R5582t333) I(R5583t2340) I(R5583t341) I(R5583t3439) I(R5584t5035) I(R5584t3918) I(R5584t542) I(R5584t690) I(R5584t1356) I(R5585t3265) I(R5585t3078) I(R5585t1346) I(R5585t2922) I(R5586t648) I(R5586t272) I(R5587t5192) I(R5587t4950) I(R5587t2131) I(R5588t1545) I(R5588t2823) I(R5588t2948) I(R5588t339) I(R5588t5384) I(R5589t5361) I(R5589t4551) I(R5589t5170) I(R5590t1928) I(R5590t337) I(R5591t175) I(R5591t3463) I(R5591t4993) I(R5591t3490) I(R5591t501) I(R5591t1051) I(R5592t4053) I(R5592t5498) I(R5593t3218) I(R5593t4961) I(R5594t1800) I(R5594t3211) I(R5595t1310) I(R5595t4302) I(R5595t1518) I(R5596t1423) I(R5596t3707) I(R5597t2174) I(R5597t255) I(R5598t807) I(R5598t4038) I(R5598t5530) I(R5598t3334) I(R5598t3323) I(R5599t3171) I(R5599t3580) I(R5599t1252) I(R5600t2258) I(R5600t3900) I(R5600t4369) I(R5600t555) I(R5600t5236) I(R5600t3397) I(R5601t451) I(R5601t5232) I(R5602t3796) I(R5603t225) I(R5603t4765) I(R5603t1732) I(R5604t2319) I(R5605t3188) I(R5605t5383) I(R5605t3452) I(R5605t3847) I(R5605t4890) I(R5606t2218) I(R5606t4193) I(R5606t2797) I(R5606t787) I(R5606t2471) I(R5607t3062) I(R5607t2033) I(R5607t1962) I(R5607t1746) I(R5608t812) I(R5608t3279) I(R5609t94) I(R5609t5142) I(R5609t2978) I(R5609t1127) I(R5610t1916) I(R5610t3939) I(R5610t646) I(R5610t5390) I(R5611t4076) I(R5611t4373) I(R5612t4182) I(R5613t4480) I(R5613t1779) I(R5613t2727) I(R5614t355) I(R5614t4423) I(R5614t1083) I(R5614t4377) I(R5615t2931) I(R5615t2881) I(R5615t5506) I(R5615t2936) I(R5616t2312) I(R5616t3200) I(R5616t5078) I(R5616t110) I(R5616t3104) I(R5617t3128) I(R5617t3669) I(R5617t2172) I(R5617t3365) I(R5618t606) I(R5618t2437) I(R5618t2743) I(R5618t5129) I(R5618t4696) I(R5618t5095) I(R5620t3976) I(R5620t2974) I(R5620t4288) I(R5621t812) I(R5621t4846) I(R5622t1536) I(R5622t4645) I(R5622t1520) I(R5622t2184) I(R5623t617) I(R5623t4940) I(R5623t2290) I(R5623t4422) I(R5624t4258) I(R5624t95) I(R5624t1789) I(R5625t4492) I(R5625t2594) I(R5626t2201) I(R5627t3875) I(R5627t1247) I(R5627t4022) I(R5627t4715) I(R5627t258) I(R5628t3964) I(R5628t5232) I(R5628t3842) I(R5628t3044) I(R5629t1194) I(R5629t2983) I(R5629t1736) I(R5630t1205) I(R5630t4370) I(R5631t490) I(R5631t1040) I(R5632t500) I(R5632t4688) I(R5632t3694) I(R5632t4382) I(R5633t5292) I(R5633t5419) I(R5634t178) I(R5634t5132) I(R5634t4781) I(R5634t5371) I(R5634t2114) I(R5634t5144) I(R5635t4914) I(R5635t4214) I(R5635t3709) I(R5635t2443) I(R5636t3768) I(R5636t1202) I(R5638t1059) I(R5638t4383) I(R5638t4776) I(R5640t5408) I(R5641t2741) I(R5641t5421) I(R5641t1088) I(R5641t1409) I(R5642t4384) I(R5642t2977) I(R5642t3255) I(R5642t1122) I(R5643t4212) I(R5643t5241) I(R5643t4893) I(R5644t2671) I(R5644t811) I(R5644t3577) I(R5644t3687) I(R5644t2197) I(R5645t497) I(R5645t1091) I(R5645t3447) I(R5645t4638) I(R5645t4650) I(R5646t1915) I(R5647t52) I(R5647t4816) I(R5647t3682) I(R5647t2296) I(R5647t823) I(R5648t2384) I(R5648t2783) I(R5648t2932) I(R5648t769) I(R5648t1683) I(R5649t49) I(R5649t3978) I(R5649t5373) I(R5650t3172) I(R5650t1507) I(R5650t1580) I(R5651t63) I(R5651t3487) I(R5651t2750) I(R5651t4731) I(R5652t235) I(R5652t2673) I(R5653t2182) I(R5653t2235) I(R5653t3826) I(R5653t1907) I(R5653t399) I(R5653t2584) I(R5654t739) I(R5654t1474) I(R5655t3821) I(R5655t1704) I(R5655t4246) I(R5655t3154) I(R5656t1188) I(R5656t1187) I(R5656t1320) I(R5657t3114) I(R5657t3420) I(R5658t3204) I(R5658t227) I(R5658t1762) I(R5659t2312) I(R5659t2812) I(R5660t2846) I(R5660t2528) I(R5660t671) I(R5660t2487) I(R5661t3611) I(R5661t5238) I(R5661t1907) I(R5661t3826) I(R5661t5193) I(R5662t4523) I(R5662t1345) I(R5663t2872) I(R5663t4875) I(R5663t3075) I(R5664t574) I(R5664t4024) I(R5665t5332) I(R5665t618) I(R5666t4775) I(R5667t49) I(R5667t934) I(R5667t2665) I(R5668t1299) I(R5668t2219) I(R5668t1516) I(R5668t4690) I(R5669t2549) I(R5669t5212) I(R5669t2680) I(R5669t672) I(R5670t1993) I(R5670t2612) I(R5670t2644) I(R5670t3071) I(R5671t5367) I(R5671t2906) I(R5671t2126) I(R5671t2344) I(R5671t246) I(R5672t4584) I(R5672t4830) I(R5672t834) I(R5672t1874) I(R5672t3268) I(R5673t3870) I(R5673t36) I(R5674t2018) I(R5674t1660) I(R5674t4913) I(R5674t281) I(R5674t477) I(R5675t1236) I(R5675t1611) I(R5675t3288) I(R5675t3293) I(R5676t1622) I(R5676t3332) I(R5676t571) I(R5677t586) I(R5677t3179) I(R5677t981) I(R5677t3497) I(R5678t2789) I(R5678t2972) I(R5678t2475) I(R5679t3421) I(R5679t3659) I(R5679t4940) I(R5679t4378) I(R5680t5534) I(R5680t3081) I(R5680t84) I(R5681t1073) I(R5681t4688) I(R5681t3944) I(R5681t661) I(R5682t5678) I(R5682t2475) I(R5682t644) I(R5682t1129) I(R5682t2254) I(R5683t26) I(R5683t803) I(R5683t1501) I(R5684t4107) I(R5684t4144) I(R5684t410) I(R5685t3994) I(R5685t858) I(R5686t4866) I(R5686t5452) I(R5686t1138) I(R5686t3746) I(R5686t2842) I(R5686t2585) I(R5687t5597) I(R5688t421) I(R5688t5066) I(R5688t1219) I(R5688t3660) I(R5689t2337) I(R5689t5001) I(R5689t4615) I(R5689t469) I(R5690t260) I(R5690t3642) I(R5690t890) I(R5691t4511) I(R5691t4675) I(R5691t5312) I(R5691t3636) I(R5692t882) I(R5692t5095) I(R5692t4696) I(R5692t5381) I(R5693t4345) I(R5693t3449) I(R5693t576) I(R5693t747) I(R5694t2353) I(R5694t4295) I(R5694t1788) I(R5694t2905) I(R5695t2360) I(R5695t1990) I(R5695t2839) I(R5695t1339) I(R5695t3534) I(R5696t5010) I(R5696t2430) I(R5696t2268) I(R5696t2048) I(R5697t2166) I(R5697t3186) I(R5697t2058) I(R5698t386) I(R5698t4142) I(R5698t1953) I(R5699t1450) I(R5699t4967) I(R5700t3609) I(R5700t828) I(R5701t2458) I(R5701t2771) I(R5701t1196) I(R5701t5482) I(R5701t5568) I(R5702t640) I(R5702t3663) I(R5702t567) I(R5702t1571) I(R5702t5340) I(R5703t871) I(R5703t3771) I(R5703t4917) I(R5703t69) I(R5704t1540) I(R5704t2518) I(R5705t782) I(R5705t5450) I(R5705t4914) I(R5706t5665) I(R5706t4292) I(R5706t2854) I(R5706t5332) I(R5707t3789) I(R5707t1920) I(R5708t4074) I(R5708t4879) I(R5709t2023) I(R5709t3174) I(R5709t3626) I(R5710t1109) I(R5710t5182) I(R5710t303) I(R5711t4934) I(R5712t2343) I(R5712t1795) I(R5712t1821) I(R5712t5034) I(R5712t5220) I(R5712t4273) I(R5713t2057) I(R5713t3866) I(R5713t66) I(R5713t860) I(R5713t2433) I(R5713t254) I(R5714t3197) I(R5714t2205) I(R5714t2225) I(R5715t3778) I(R5715t746) I(R5716t828) I(R5716t3609) I(R5716t291) I(R5716t3645) I(R5716t259) I(R5717t1858) I(R5717t125) I(R5717t4674) I(R5717t35) I(R5718t3296) I(R5718t4141) I(R5718t4636) I(R5718t3213) I(R5718t5499) I(R5718t1869) I(R5719t386) I(R5719t5698) I(R5719t1953) I(R5720t3849) I(R5720t1068) I(R5720t2999) I(R5721t4170) I(R5721t2125) I(R5721t3871) I(R5721t3030) I(R5722t1282) I(R5722t793) I(R5722t2036) I(R5722t2701) I(R5722t1649) I(R5722t4374) I(R5722t1958) I(R5723t1987) I(R5723t4267) I(R5724t3863) I(R5724t3853) I(R5724t3698) I(R5724t2992) I(R5725t1972) I(R5725t3251) I(R5725t128) I(R5725t5181) I(R5726t3466) I(R5726t4829) I(R5726t3855) I(R5727t62) I(R5727t2681) I(R5727t1711) I(R5728t1360) I(R5728t5059) I(R5728t1480) I(R5728t2811) I(R5729t4844) I(R5729t4790) I(R5729t2988) I(R5730t2113) I(R5730t3057) I(R5730t3736) I(R5730t3160) I(R5730t672) I(R5730t2680) I(R5731t1894) I(R5731t4541) I(R5731t1431) I(R5731t357) I(R5732t5099) I(R5732t3630) I(R5733t3015) I(R5733t3554) I(R5733t5108) I(R5733t842) I(R5734t782) I(R5734t5705) I(R5734t512) I(R5734t3976) I(R5734t5620) I(R5734t4914) I(R5735t5709) I(R5735t1003) I(R5735t443) I(R5735t3626) I(R5736t4952) I(R5737t2260) I(R5737t2813) I(R5737t476) I(R5737t4956) I(R5737t3650) I(R5738t1630) I(R5738t3990) I(R5739t191) I(R5739t2192) I(R5739t1753) I(R5740t1930) I(R5740t302) I(R5741t1342) I(R5742t832) I(R5742t2509) I(R5742t2540) I(R5743t536) I(R5744t3982) I(R5745t4040) I(R5745t5284) I(R5745t772) I(R5745t194) I(R5746t1829) I(R5746t5521) I(R5746t1583) I(R5746t2751) I(R5746t2679) I(R5746t2128) I(R5746t2119) I(R5747t5428) I(R5747t3518) I(R5747t1230) I(R5748t5227) I(R5748t1444) I(R5748t2454) I(R5748t508) I(R5749t2165) I(R5749t5630) I(R5749t452) I(R5749t3046) I(R5750t56) I(R5750t3226) I(R5750t1964) I(R5750t474) I(R5750t2103) I(R5750t1482) I(R5751t1741) I(R5751t1072) I(R5751t5480) I(R5752t868) I(R5752t909) I(R5752t4680) I(R5752t1638) I(R5752t1766) I(R5753t1022) I(R5753t3370) I(R5753t422) I(R5754t2180) I(R5755t4842) I(R5755t2435) I(R5756t5169) I(R5756t1150) I(R5756t3835) I(R5756t2934) I(R5756t134) I(R5757t2115) I(R5757t3170) I(R5758t1703) I(R5758t3064) I(R5758t851) I(R5758t5434) I(R5758t3500) I(R5758t2867) I(R5759t3682) I(R5759t4953) I(R5759t5647) I(R5759t52) I(R5759t758) I(R5759t4554) I(R5759t4221) I(R5760t1926) I(R5760t5580) I(R5760t328) I(R5761t1709) I(R5761t3108) I(R5761t412) I(R5761t641) I(R5761t85) I(R5762t2208) I(R5762t5392) I(R5762t901) I(R5763t2056) I(R5763t1749) I(R5764t293) I(R5764t2739) I(R5765t466) I(R5765t521) I(R5765t4594) I(R5765t1393) I(R5766t3529) I(R5766t2913) I(R5767t1692) I(R5767t3396) I(R5767t3892) I(R5767t1524) I(R5768t1852) I(R5768t5711) I(R5768t4934) I(R5768t4752) I(R5768t5044) I(R5769t190) I(R5769t3379) I(R5770t734) I(R5770t4687) I(R5770t1690) I(R5770t1790) I(R5771t4562) I(R5771t1299) I(R5771t2219) I(R5772t1266) I(R5772t3529) I(R5772t5766) I(R5773t1958) I(R5773t4374) I(R5774t5135) I(R5774t4535) I(R5774t558) I(R5775t4062) I(R5776t3754) I(R5776t3194) I(R5777t825) I(R5777t853) I(R5777t1656) I(R5778t1789) I(R5778t3215) I(R5778t3529) I(R5778t5766) I(R5778t2913) I(R5778t5624) I(R5779t4055) I(R5779t816) I(R5780t4160) I(R5780t3290) I(R5781t925) I(R5782t5267) I(R5782t4944) I(R5782t4417) I(R5783t832) I(R5783t4979) I(R5783t5742) I(R5784t5510) I(R5784t3624) I(R5785t1473) I(R5785t2577) I(R5785t3391) I(R5785t3113) I(R5785t1751) I(R5786t3977) I(R5786t2412) I(R5786t3418) I(R5786t2461) I(R5786t538) I(R5787t3308) I(R5787t1787) I(R5787t4522) I(R5787t5396) I(R5787t4385) I(R5788t1098) I(R5788t5553) I(R5788t4737) I(R5788t3936) I(R5788t4571) I(R5789t2196) I(R5789t3790) I(R5789t1489) I(R5789t1430) I(R5790t381) I(R5790t5136) I(R5790t2266) I(R5791t4104) I(R5791t5558) I(R5791t2740) I(R5791t5030) I(R5792t3504) I(R5792t4481) I(R5792t2714) I(R5792t4464) I(R5792t1274) I(R5792t5180) I(R5793t101) I(R5793t1550) I(R5793t5593) I(R5793t4961) I(R5793t4440) I(R5793t3187) I(R5794t5494) I(R5794t3571) I(R5795t876) I(R5795t3602) I(R5795t4173) I(R5795t2464) I(R5796t978) I(R5796t1487) I(R5796t2124) I(R5797t3488) I(R5797t616) I(R5797t974) I(R5797t576) I(R5798t2766) I(R5798t3251) I(R5798t3254) I(R5798t2539) I(R5798t4900) I(R5799t5630) I(R5799t5749) I(R5799t1205) I(R5799t940) I(R5799t452) I(R5800t323) I(R5800t2734) I(R5801t5415) I(R5801t501) I(R5801t3490) I(R5801t3050) I(R5801t3502) I(R5801t4381) I(R5802t695) I(R5802t1576) I(R5802t2609) I(R5802t3129) I(R5803t2328) I(R5803t4240) I(R5803t1899) I(R5804t3116) I(R5804t272) I(R5804t5586) I(R5804t648) I(R5804t1906) I(R5805t1679) I(R5805t1619) I(R5805t2367) I(R5806t1951) I(R5806t5096) I(R5806t3229) I(R5806t2084) I(R5806t3031) I(R5807t4022) I(R5807t4715) I(R5807t4857) I(R5807t4020) I(R5807t5358) I(R5807t1675) I(R5808t1185) I(R5808t3683) I(R5808t4809) I(R5808t4978) I(R5809t5332) I(R5809t2369) I(R5810t1959) I(R5810t4557) I(R5810t3973) I(R5810t3425) I(R5811t4548) I(R5811t2804) I(R5811t2452) I(R5811t67) I(R5811t3337) I(R5811t4984) I(R5812t1803) I(R5813t2300) I(R5813t4660) I(R5813t2623) I(R5813t3434) I(R5814t2041) I(R5814t73) I(R5815t4643) I(R5815t1062) I(R5815t986) I(R5815t4854) I(R5815t4002) I(R5816t381) I(R5816t157) I(R5816t5136) I(R5816t5790) I(R5817t1922) I(R5817t601) I(R5817t2564) I(R5818t44) I(R5818t1450) I(R5818t2809) I(R5819t3720) I(R5819t5326) I(R5819t4683) I(R5820t62) I(R5820t2529) I(R5820t5727) I(R5820t1711) I(R5820t3922) I(R5821t3193) I(R5821t2099) I(R5822t4067) I(R5822t4118) I(R5822t1078) I(R5822t4046) I(R5822t930) I(R5822t4803) I(R5823t3332) I(R5823t5676) I(R5823t571) I(R5823t208) I(R5823t124) I(R5824t3437) I(R5824t888) I(R5824t4425) I(R5825t2414) I(R5825t5270) I(R5825t1291) I(R5826t3588) I(R5826t2965) I(R5826t2380) I(R5826t240) I(R5826t380) I(R5827t1371) I(R5827t4658) I(R5827t215) I(R5828t3781) I(R5828t4239) I(R5829t4605) I(R5829t3449) I(R5830t1017) I(R5830t3083) I(R5831t2092) I(R5831t2688) I(R5831t3398) I(R5831t5002) I(R5831t1858) I(R5832t2899) I(R5832t5277) I(R5833t38) I(R5833t2733) I(R5833t3929) I(R5833t4687) I(R5833t734) I(R5834t4745) I(R5834t2059) I(R5834t5567) I(R5835t3710) I(R5835t4241) I(R5836t4513) I(R5836t4211) I(R5836t1522) I(R5836t1859) I(R5836t5457) I(R5836t24) I(R5837t2748) I(R5837t2637) I(R5837t5495) I(R5838t1786) I(R5838t5138) I(R5838t1102) I(R5838t895) I(R5838t5070) I(R5839t1976) I(R5839t661) I(R5840t3359) I(R5840t3512) I(R5841t1142) I(R5841t1773) I(R5841t3000) I(R5841t831) I(R5841t1367) I(R5841t1237) I(R5842t1659) I(R5842t4604) I(R5842t579) I(R5842t4624) I(R5843t1805) I(R5844t4607) I(R5844t524) I(R5845t2475) I(R5845t1635) I(R5845t439) I(R5845t2009) I(R5845t1562) I(R5845t4775) I(R5846t4867) I(R5846t914) I(R5847t5665) I(R5847t618) I(R5847t1412) I(R5847t3214) I(R5847t1221) I(R5848t1171) I(R5848t3331) I(R5848t4936) I(R5848t649) I(R5849t1159) I(R5849t1488) I(R5849t196) I(R5849t3576) I(R5849t2775) I(R5850t2992) I(R5850t3698) I(R5850t4823) I(R5850t5164) I(R5851t628) I(R5851t195) I(R5851t2461) I(R5852t5312) I(R5853t310) I(R5853t4676) I(R5853t2562) I(R5853t3936) I(R5853t4737) I(R5853t1734) I(R5854t1079) I(R5854t4257) I(R5854t3031) I(R5854t4229) I(R5855t1765) I(R5855t3480) I(R5855t4839) I(R5855t1349) I(R5855t3875) I(R5855t2874) I(R5856t4467) I(R5856t112) I(R5856t3317) I(R5857t608) I(R5857t142) I(R5857t3092) I(R5858t4053) I(R5858t5592) I(R5858t5498) I(R5858t4907) I(R5858t4693) I(R5858t958) I(R5859t4512) I(R5860t2940) I(R5860t5439) I(R5860t4386) I(R5861t675) I(R5861t1340) I(R5861t3324) I(R5861t112) I(R5861t3317) I(R5862t2290) I(R5862t5623) I(R5862t906) I(R5862t5657) I(R5862t3114) I(R5862t4422) I(R5863t5295) I(R5863t1183) I(R5863t3064) I(R5863t3410) I(R5864t4026) I(R5864t1312) I(R5864t220) I(R5864t2761) I(R5864t1882) I(R5864t5775) I(R5865t103) I(R5865t3714) I(R5865t5546) I(R5866t639) I(R5866t354) I(R5866t4168) I(R5867t1098) I(R5867t5788) I(R5867t5553) I(R5869t4852) I(R5869t5673) I(R5869t5720) I(R5869t3849) I(R5870t143) I(R5871t3282) I(R5871t3055) I(R5871t2968) I(R5872t423) I(R5872t4811) I(R5872t4194) I(R5873t1540) I(R5873t5704) I(R5873t3459) I(R5873t2518) I(R5874t459) I(R5874t3952) I(R5874t2231) I(R5874t1975) I(R5875t2835) I(R5875t5700) I(R5876t2015) I(R5876t3649) I(R5876t4952) I(R5877t5639) I(R5877t3727) I(R5878t2470) I(R5878t1124) I(R5878t3779) I(R5879t1109) I(R5879t5182) I(R5879t4277) I(R5880t2601) I(R5880t3295) I(R5881t1624) I(R5881t5244) I(R5881t3583) I(R5882t219) I(R5882t3560) I(R5882t2657) I(R5882t2682) I(R5882t4153) I(R5882t3246) I(R5882t3526) I(R5883t1252) I(R5883t2139) I(R5884t1924) I(R5884t3898) I(R5884t2763) I(R5884t1222) I(R5885t1315) I(R5885t2487) I(R5885t3881) I(R5886t324) I(R5886t3058) I(R5886t2898) I(R5886t3190) I(R5887t5757) I(R5887t3239) I(R5888t5116) I(R5888t5257) I(R5889t1618) I(R5889t1669) I(R5889t5222) I(R5889t3592) I(R5890t2049) I(R5890t3197) I(R5890t3413) I(R5891t2120) I(R5892t1480) I(R5892t631) I(R5892t2811) I(R5892t5728) I(R5893t3746) I(R5893t2669) I(R5894t407) I(R5894t2924) I(R5894t1795) I(R5894t1173) I(R5894t4137) I(R5894t923) I(R5895t1593) I(R5895t3027) I(R5895t4691) I(R5895t1667) I(R5896t5761) I(R5896t641) I(R5896t754) I(R5896t1035) I(R5897t1301) I(R5897t88) I(R5897t817) I(R5897t2101) I(R5898t4759) I(R5898t5352) I(R5898t3927) I(R5898t5070) I(R5899t1899) I(R5899t5183) I(R5899t2201) I(R5899t5626) I(R5899t5256) I(R5899t4947) I(R5900t5261) I(R5900t3287) I(R5900t3245) I(R5901t5176) I(R5901t1162) I(R5902t2221) I(R5902t2795) I(R5902t2499) I(R5902t1049) I(R5903t2590) I(R5903t3382) I(R5903t5329) I(R5903t1387) I(R5903t5050) I(R5905t5367) I(R5905t877) I(R5905t4814) I(R5906t368) I(R5906t5510) I(R5906t2325) I(R5906t3180) I(R5906t3159) I(R5907t812) I(R5907t5608) I(R5907t498) I(R5907t2655) I(R5908t819) I(R5908t3208) I(R5908t3030) I(R5909t4758) I(R5911t1077) I(R5911t3858) I(R5912t906) I(R5912t2225) I(R5912t569) I(R5913t16) I(R5913t1072) I(R5913t1855) I(R5913t5751) I(R5914t3971) I(R5914t567) I(R5914t3248) I(R5915t4094) I(R5915t5039) I(R5915t2719) I(R5916t5437) I(R5916t1688) I(R5916t4673) I(R5916t1660) I(R5916t4913) I(R5917t691) I(R5917t2689) I(R5918t1345) I(R5918t5662) I(R5918t4523) I(R5918t3513) I(R5918t3650) I(R5918t739) I(R5918t5654) I(R5919t3542) I(R5919t932) I(R5919t3452) I(R5919t5213) I(R5920t2526) I(R5920t4627) I(R5920t20) I(R5920t306) I(R5920t2026) I(R5921t1034) I(R5921t4210) I(R5921t1082) I(R5922t1783) I(R5922t3048) I(R5922t4909) I(R5922t1238) I(R5922t290) I(R5922t308) I(R5922t165) I(R5922t3942) I(R5923t970) I(R5923t5843) I(R5923t1805) I(R5924t2814) I(R5924t4187) I(R5924t4052) I(R5924t3194) I(R5925t2683) I(R5925t166) I(R5925t1578) I(R5925t2484) I(R5926t5386) I(R5926t4249) I(R5926t3584) I(R5927t4269) I(R5927t1459) I(R5928t2027) I(R5928t3700) I(R5929t1229) I(R5929t1983) I(R5929t3901) I(R5930t4337) I(R5930t2807) I(R5930t1510) I(R5930t572) I(R5931t1792) I(R5931t1444) I(R5931t2937) I(R5932t1920) I(R5932t701) I(R5932t3831) I(R5933t951) I(R5934t2343) I(R5934t5712) I(R5934t1046) I(R5934t4273) I(R5935t2001) I(R5935t2003) I(R5935t4665) I(R5936t3282) I(R5936t5871) I(R5936t937) I(R5936t919) I(R5936t3055) I(R5937t5927) I(R5937t1459) I(R5937t4493) I(R5937t3469) I(R5938t2817) I(R5938t4677) I(R5939t2765) I(R5939t2168) I(R5940t4949) I(R5940t4095) I(R5941t574) I(R5941t1257) I(R5941t313) I(R5942t3292) I(R5942t4608) I(R5942t2179) I(R5942t1674) I(R5942t2659) I(R5943t978) I(R5943t5190) I(R5943t5796) I(R5944t379) I(R5944t5532) I(R5944t4796) I(R5944t5124) I(R5945t875) I(R5945t2729) I(R5945t5427) I(R5946t3115) I(R5946t66) I(R5947t2698) I(R5947t2842) I(R5948t1831) I(R5948t4634) I(R5948t4712) I(R5949t1946) I(R5949t2769) I(R5950t4822) I(R5950t5365) I(R5950t1232) I(R5950t3167) I(R5950t690) I(R5950t3593) I(R5950t2816) I(R5951t4597) I(R5951t2727) I(R5952t3267) I(R5952t5119) I(R5952t5015) I(R5952t4023) I(R5952t1579) I(R5952t4529) I(R5952t3135) I(R5953t4512) I(R5953t4152) I(R5953t109) I(R5953t3675) I(R5954t4384) I(R5954t1122) I(R5955t4509) I(R5955t2775) I(R5956t420) I(R5956t1478) I(R5956t4323) I(R5956t905) I(R5957t1032) I(R5957t3703) I(R5957t5055) I(R5957t1333) I(R5958t1669) I(R5958t5889) I(R5958t3592) I(R5959t5619) I(R5959t84) I(R5960t61) I(R5960t4396) I(R5960t5885) I(R5961t973) I(R5961t4948) I(R5961t2396) I(R5962t4127) I(R5962t4178) I(R5962t3150) I(R5962t480) I(R5962t551) I(R5962t2596) I(R5962t2102) I(R5962t5274) I(R5963t1755) I(R5963t4733) I(R5963t4115) I(R5963t3237) I(R5963t702) I(R5963t3622) I(R5964t725) I(R5964t1445) I(R5965t4732) I(R5965t3782) I(R5965t5456) I(R5966t1203) I(R5966t5137) I(R5966t5487) I(R5967t2178) I(R5967t3551) I(R5967t1813) I(R5967t4590) I(R5968t2550) I(R5968t213) I(R5968t677) I(R5969t1603) I(R5969t4257) I(R5969t3404) I(R5969t1436) I(R5969t4229) I(R5969t5854) I(R5970t3192) I(R5970t1370) I(R5970t992) I(R5971t2060) I(R5971t3289) I(R5971t4966) I(R5972t4248) I(R5972t4126) I(R5972t1166) I(R5973t812) I(R5973t928) I(R5973t4846) I(R5974t1336) I(R5974t5603) I(R5974t225) I(R5974t1261) I(R5974t4840) I(R5975t4251) I(R5975t5068) I(R5975t4101) I(R5975t2341) I(R5975t4931) I(R5976t964) I(R5976t3401) I(R5976t5743) I(R5977t4588) I(R5978t1358) I(R5978t2837) I(R5979t2060) I(R5979t5971) I(R5979t3679) I(R5979t122) I(R5980t654) I(R5980t2129) I(R5980t1384) I(R5980t3727) I(R5980t5877) I(R5981t4411) I(R5981t4692) I(R5981t3888) I(R5981t5412) I(R5981t865) I(R5982t2382) I(R5982t2831) I(R5983t4412) I(R5983t308) I(R5984t1814) I(R5984t3860) I(R5984t2975) I(R5984t1242) I(R5985t553) I(R5986t2351) I(R5986t938) I(R5986t3381) I(R5987t1900) I(R5987t3834) I(R5987t581) I(R5987t3582) I(R5988t2921) I(R5988t5153) I(R5989t1686) I(R5989t2031) I(R5989t3053) I(R5989t2316) I(R5989t3605) I(R5990t3131) I(R5990t194) I(R5990t385) I(R5990t2615) I(R5991t5639) I(R5991t5877) I(R5992t2825) I(R5992t5281) I(R5993t4375) I(R5993t1260) I(R5994t2008) I(R5994t5631) I(R5994t1040) I(R5994t4139) I(R5995t4724) I(R5996t2180) I(R5996t5754) I(R5997t1087) I(R5997t4452) I(R5997t2838) I(R5998t2632) I(R5998t2861) I(R5998t3559) I(R5998t4206) I(R5999t3459) I(R5999t1540) I(R5999t4090) I(R5999t236) I(R6000t2928) I(R6000t4730) I(R6000t5933) I(R6001t3932) I(R6001t3079) I(R6001t3590) I(R6001t5248) I(R6002t2595) I(R6003t4461) I(R6003t4895) I(R6003t627) I(R6003t2497) I(R6003t2827) I(R6003t1087) I(R6003t5488) I(R6004t956) I(R6004t3001) I(R6004t3018) I(R6005t2322) I(R6005t364) I(R6005t2535) I(R6005t3879) I(R6005t822) I(R6006t719) I(R6006t1223) I(R6007t177) I(R6007t2981) I(R6007t1404) I(R6007t4786) I(R6008t1560) I(R6008t5024) I(R6008t3682) I(R6008t2296) I(R6008t245) I(R6009t4017) I(R6009t405) I(R6009t2668) I(R6009t1206) I(R6009t1406) I(R6010t1466) I(R6010t3554) I(R6010t1515) I(R6010t2949) I(R6011t426) I(R6011t3957) I(R6011t1047) I(R6011t3341) I(R6012t4074) I(R6012t4744) I(R6012t3437) I(R6012t4758) I(R6013t2726) I(R6013t352) I(R6013t4987) I(R6014t3945) I(R6014t4630) I(R6014t2385) I(R6014t2639) I(R6015t757) I(R6015t5545) I(R6015t3563) I(R6015t4878) I(R6015t3127) I(R6016t3412) I(R6016t5012) I(R6016t2911) I(R6016t3555) I(R6016t4885) I(R6017t2252) I(R6017t3774) I(R6018t1284) I(R6018t4350) I(R6018t683) I(R6018t1840) I(R6018t3867) I(R6019t3283) I(R6019t3402) I(R6019t5392) I(R6019t2622) I(R6020t5509) I(R6020t3835) I(R6020t2934) I(R6020t2325) I(R6020t3017) I(R6021t5685) I(R6021t4186) I(R6021t3994) I(R6022t4540) I(R6022t708) I(R6022t4392) I(R6023t2728) I(R6023t4177) I(R6023t4926) I(R6023t166) I(R6023t2683) I(R6023t3849) I(R6024t410) I(R6024t5876) I(R6024t4952) I(R6024t5525) I(R6025t1673) I(R6025t114) I(R6025t47) I(R6026t2248) I(R6026t3753) I(R6026t2484) I(R6026t5925) I(R6027t4840) I(R6027t4313) I(R6027t3868) I(R6027t5401) I(R6028t3) I(R6028t3552) I(R6028t4470) I(R6028t4172) I(R6029t575) I(R6029t2276) I(R6029t4130) I(R6030t1725) I(R6030t4336) I(R6030t1700) I(R6030t1840) I(R6030t3867) I(R6031t1132) I(R6031t3479) I(R6031t1096) I(R6031t3416) I(R6031t1619) I(R6031t4109) I(R6032t2609) I(R6032t3129) I(R6032t5422) I(R6032t5479) I(R6033t1737) I(R6033t2564) I(R6034t1954) I(R6034t1093) I(R6034t4577) I(R6035t3610) I(R6035t4395) I(R6035t4400) I(R6035t3339) I(R6035t2212) I(R6036t1401) I(R6036t1968) I(R6036t4521) I(R6036t3672) I(R6036t5374) I(R6036t3860) I(R6036t1713) I(R6037t3287) I(R6037t5900) I(R6037t5378) I(R6037t5261) I(R6038t3966) I(R6038t1420) I(R6039t485) I(R6039t829) I(R6039t5042) I(R6039t910) I(R6040t1151) I(R6040t4963) I(R6040t3493) I(R6040t3786) I(R6040t337) I(R6040t5590) I(R6040t1928) I(R6042t4726) I(R6042t5773) I(R6042t1958) I(R6042t4083) I(R6043t461) I(R6043t1483) I(R6044t2392) I(R6044t1936) I(R6044t2653) I(R6045t401) I(R6045t4119) I(R6045t2420) I(R6045t3932) I(R6046t3400) I(R6046t669) I(R6046t2106) I(R6046t3762) I(R6047t363) I(R6047t4172) I(R6047t1655) I(R6047t2982) I(R6047t704) I(R6047t1212) I(R6048t656) I(R6048t2053) I(R6048t5411) I(R6048t4583) I(R6048t4777) I(R6048t4310) I(R6049t1379) I(R6049t3795) I(R6049t2017) I(R6049t2213) I(R6049t1053) I(R6049t2576) I(R6049t3394) I(R6050t3012) I(R6050t4623) I(R6050t1345) I(R6050t4341) I(R6050t5543) I(R6051t5408) I(R6051t4013) I(R6052t1028) I(R6052t2974) I(R6052t5620) I(R6053t5814) I(R6053t2041) I(R6053t4281) I(R6053t553) I(R6053t3481) I(R6054t5361) I(R6054t5589) I(R6055t5000) I(R6055t3153) I(R6055t3386) I(R6055t1517) I(R6055t4612) I(R6056t4187) I(R6056t3172) I(R6056t3754) I(R6056t5776) I(R6056t3194) I(R6056t5924) I(R6057t3704) I(R6057t1211) I(R6057t1677) I(R6057t317) I(R6057t4652) I(R6058t2563) I(R6058t5382) I(R6058t5397) I(R6058t3059) I(R6058t3683) I(R6059t3313) I(R6059t662) I(R6059t3800) I(R6059t5249) I(R6060t3151) I(R6060t4841) I(R6061t2008) I(R6061t3850) I(R6061t4603) I(R6062t5206) I(R6062t3852) I(R6062t469) I(R6062t1594) I(R6063t1238) I(R6063t4909) I(R6063t3096) I(R6063t3324) I(R6063t5861) I(R6063t1340) I(R6063t5033) I(R6064t347) I(R6064t3270) I(R6064t2557) I(R6064t5077) I(R6065t152) I(R6065t5009) I(R6065t3151) I(R6065t2752) I(R6065t794) I(R6065t3378) I(R6066t2459) I(R6066t5041) I(R6066t3157) I(R6066t3142) I(R6066t5453) I(R6067t1028) I(R6067t2974) I(R6067t1596) I(R6067t4288) I(R6067t5620) I(R6068t4592) I(R6068t3631) I(R6069t2494) I(R6069t3470) I(R6069t2556) I(R6069t4887) I(R6070t173) I(R6070t4577) I(R6070t627) I(R6070t292) I(R6071t2141) I(R6071t3169) I(R6071t365) I(R6071t2422) I(R6072t1266) I(R6072t3529) I(R6072t597) I(R6073t4799) I(R6074t4222) I(R6074t4567) I(R6074t5056) I(R6074t3231) I(R6074t3281) I(R6075t479) I(R6075t4693) I(R6075t5858) I(R6075t4907) I(R6075t2688) I(R6076t5073) I(R6076t3395) I(R6076t5887) I(R6077t1712) I(R6077t4607) I(R6077t2498) I(R6077t4988) I(R6078t2200) I(R6078t2903) I(R6078t4985) I(R6079t880) I(R6079t2385) I(R6079t3569) I(R6080t2157) I(R6080t3381) I(R6080t4672) I(R6080t946) I(R6081t20) I(R6081t4627) I(R6081t963) I(R6082t3331) I(R6082t5344) I(R6082t1171) I(R6083t2197) I(R6083t3687) I(R6083t3577) I(R6084t4932) I(R6084t5029) I(R6085t96) I(R6085t3665) I(R6085t4659) I(R6085t4488) I(R6085t1264) I(R6086t555) I(R6087t3337) I(R6087t67) I(R6087t59) I(R6087t4929) I(R6087t463) I(R6088t4422) I(R6088t5623) I(R6088t5107) I(R6088t2064) I(R6089t3199) I(R6089t4591) I(R6090t3168) I(R6091t183) I(R6091t5321) I(R6091t1235) I(R6091t2778) I(R6092t216) I(R6092t3521) I(R6092t1384) I(R6092t3738) I(R6092t1917) I(R6093t2895) I(R6093t3946) I(R6093t229) I(R6093t5388) I(R6093t4349) I(R6094t922) I(R6094t5481) I(R6094t392) I(R6094t1365) I(R6094t5423) I(R6095t846) I(R6095t2495) I(R6095t3748) I(R6096t1153) I(R6096t1865) I(R6096t4448) I(R6096t170) I(R6097t5877) I(R6097t4557) I(R6097t2085) I(R6097t3727) I(R6098t217) I(R6098t2401) I(R6099t4479) I(R6099t5383) I(R6099t3452) I(R6099t932) I(R6100t3471) I(R6100t5888) I(R6100t1297) I(R6100t4829) I(R6101t653) I(R6101t1805) I(R6101t4285) I(R6102t1176) I(R6102t881) I(R6102t3029) I(R6103t2498) I(R6103t2169) I(R6103t523) I(R6103t3506) I(R6103t3085) I(R6104t4779) I(R6104t3787) I(R6104t2615) I(R6104t5990) I(R6105t23) I(R6105t3491) I(R6105t603) I(R6105t4805) I(R6105t2841) I(R6106t2248) I(R6106t3753) I(R6106t6026) I(R6107t1883) I(R6107t3402) I(R6107t901) I(R6107t5762) I(R6107t5392) I(R6107t6019) I(R6108t5332) I(R6108t2369) I(R6108t3666) I(R6109t2448) I(R6109t3757) I(R6109t4910) I(R6109t137) I(R6109t1069) I(R6110t3604) I(R6110t4911) I(R6111t991) I(R6111t4231) I(R6111t1307) I(R6112t1252) I(R6112t5599) I(R6112t2244) I(R6112t1943) I(R6113t4198) I(R6113t5804) I(R6113t3116) I(R6114t2842) I(R6114t2585) I(R6115t4939) I(R6115t3991) I(R6115t2112) I(R6116t1699) I(R6116t4587) I(R6116t2028) I(R6116t1518) I(R6116t5595) I(R6116t1310) I(R6117t3200) I(R6117t5577) I(R6117t3013) I(R6117t2654) I(R6118t4141) I(R6118t4337) I(R6118t5553) I(R6118t5788) I(R6118t4737) I(R6119t1195) I(R6119t2901) I(R6120t885) I(R6120t3096) I(R6120t3464) I(R6120t2012) I(R6121t4144) I(R6121t5684) I(R6121t3529) I(R6121t597) I(R6121t3581) I(R6122t5562) I(R6122t3271) I(R6122t2408) I(R6122t2148) I(R6122t6083) I(R6123t4417) I(R6123t4944) I(R6123t1745) I(R6123t4555) I(R6123t647) I(R6124t4950) I(R6124t5587) I(R6124t2885) I(R6124t5192) I(R6125t5562) I(R6125t614) I(R6125t1208) I(R6125t2339) I(R6125t2520) I(R6126t1457) I(R6126t560) I(R6126t429) I(R6127t3625) I(R6127t3691) I(R6127t1573) I(R6127t369) I(R6127t1945) I(R6128t2013) I(R6128t5417) I(R6128t163) I(R6128t2916) I(R6128t2721) I(R6129t68) I(R6129t4004) I(R6129t4690) I(R6129t1516) I(R6129t3493) I(R6130t2707) I(R6130t1095) I(R6130t605) I(R6130t2297) I(R6131t2789) I(R6131t4002) I(R6131t5078) I(R6131t5616) I(R6131t2312) I(R6132t1798) I(R6132t3444) I(R6132t1589) I(R6132t2016) I(R6132t5527) I(R6132t799) I(R6133t375) I(R6133t686) I(R6134t1471) I(R6134t1770) I(R6134t5201) I(R6135t3518) I(R6135t3561) I(R6135t320) I(R6135t3515) I(R6136t2029) I(R6136t2798) I(R6136t5722) I(R6136t1958) I(R6137t826) I(R6137t1353) I(R6137t3300) I(R6138t2634) I(R6138t5334) I(R6138t1874) I(R6138t5672) I(R6138t3268) I(R6138t4478) I(R6139t1737) I(R6139t3764) I(R6139t5074) I(R6139t6033) I(R6140t3061) I(R6140t3766) I(R6140t5240) I(R6142t1412) I(R6142t5847) I(R6142t1653) I(R6143t3718) I(R6143t3726) I(R6143t5001) I(R6143t2760) I(R6144t1871) I(R6144t600) I(R6145t3456) I(R6145t5076) I(R6145t1769) I(R6146t4801) I(R6146t678) I(R6146t1140) I(R6147t4876) I(R6147t2918) I(R6147t2114) I(R6147t5371) I(R6147t1719) I(R6148t464) I(R6148t3801) I(R6149t2388) I(R6149t818) I(R6150t5039) I(R6150t5179) I(R6150t2233) I(R6150t5915) I(R6151t1243) I(R6151t5385) I(R6151t2209) I(R6151t3550) I(R6152t1456) I(R6152t1709) I(R6153t5273) I(R6153t904) I(R6153t116) I(R6153t4575) I(R6154t530) I(R6154t3038) I(R6154t703) I(R6155t3241) I(R6155t1897) I(R6156t3349) I(R6156t533) I(R6156t239) I(R6156t2245) I(R6157t1121) I(R6157t3184) I(R6157t447) I(R6157t2250) I(R6158t4879) I(R6158t5557) I(R6158t327) I(R6158t5708) I(R6159t590) I(R6159t4397) I(R6160t205) I(R6160t5304) I(R6160t4709) I(R6160t4036) I(R6160t829) I(R6160t3777) I(R6161t552) I(R6161t3225) I(R6161t3898) I(R6162t5314) I(R6162t4558) I(R6162t2388) I(R6163t784) I(R6163t5028) I(R6163t1602) I(R6163t4728) I(R6164t151) I(R6164t2323) I(R6165t1140) I(R6165t5177) I(R6165t5210) I(R6165t3633) I(R6165t2945) I(R6166t3417) I(R6166t4908) I(R6166t2403) I(R6166t1933) I(R6166t1834) I(R6167t4364) I(R6167t1527) I(R6168t1702) I(R6168t4131) I(R6168t1169) I(R6168t2698) I(R6168t5947) I(R6168t3522) I(R6168t5276) I(R6169t2682) I(R6169t2626) I(R6169t4972) I(R6169t2361) I(R6170t3380) I(R6170t1410) I(R6171t3556) I(R6171t4432) I(R6171t1404) I(R6171t4855) I(R6171t4384) I(R6171t5954) I(R6172t650) I(R6172t5610) I(R6172t3704) I(R6172t721) I(R6173t491) I(R6173t3702) I(R6174t5613) I(R6175t911) I(R6175t30) I(R6175t1796) I(R6176t3014) I(R6176t4485) I(R6176t413) I(R6176t3691) I(R6176t827) I(R6177t5486) I(R6177t4138) I(R6177t2418) I(R6177t4329) I(R6178t4802) I(R6178t689) I(R6178t3285) I(R6178t1862) I(R6178t338) I(R6178t1209) I(R6179t694) I(R6179t525) I(R6180t1596) I(R6180t6067) I(R6180t1028) I(R6181t1320) I(R6181t1898) I(R6181t5641) I(R6182t1790) I(R6182t5770) I(R6183t1897) I(R6183t5088) I(R6183t6155) I(R6183t3241) I(R6184t3426) I(R6184t2294) I(R6185t5359) I(R6185t3054) I(R6185t5702) I(R6185t1571) I(R6186t1854) I(R6186t2467) I(R6186t4303) I(R6186t2041) I(R6187t126) I(R6187t2488) I(R6187t3695) I(R6187t494) I(R6188t4262) I(R6188t4769) I(R6189t4144) I(R6189t6121) I(R6189t3581) I(R6190t663) I(R6190t248) I(R6190t984) I(R6190t5540) I(R6191t2198) I(R6192t4914) I(R6192t5635) I(R6192t1028) I(R6192t6052) I(R6192t5620) I(R6192t5734) I(R6193t2707) I(R6193t6130) I(R6193t131) I(R6194t1868) I(R6195t3573) I(R6195t3993) I(R6195t2930) I(R6196t3421) I(R6196t5679) I(R6196t3659) I(R6196t4438) I(R6196t3585) I(R6196t2600) I(R6197t226) I(R6197t3165) I(R6197t4154) I(R6197t4252) I(R6198t3450) I(R6198t5125) I(R6198t4858) I(R6198t5158) I(R6199t232) I(R6199t1580) I(R6199t4320) I(R6199t2713) I(R6200t3568) I(R6200t3878) I(R6200t6017) I(R6200t2252) I(R6201t2626) I(R6201t2657) I(R6201t6179) I(R6202t3132) I(R6202t2963) I(R6202t5315) I(R6202t5349) I(R6203t2040) I(R6203t3948) I(R6203t2358) I(R6204t5219) I(R6204t5441) I(R6204t111) I(R6205t886) I(R6205t2820) I(R6205t3398) I(R6205t5831) I(R6205t2688) I(R6206t5219) I(R6206t4291) I(R6207t235) I(R6207t2748) I(R6207t5837) I(R6208t5729) I(R6208t1642) I(R6208t3798) I(R6208t3597) I(R6208t2988) I(R6209t415) I(R6209t1908) I(R6209t3845) I(R6210t5323) I(R6210t3807) I(R6211t208) I(R6211t1460) I(R6211t2773) I(R6212t1685) I(R6212t4046) I(R6212t1988) I(R6212t5016) I(R6213t63) I(R6213t3487) I(R6213t2690) I(R6213t5182) I(R6213t5710) I(R6213t303) I(R6213t13) I(R6213t758) I(R6214t1793) I(R6214t4719) I(R6215t2546) I(R6215t3090) I(R6215t2360) I(R6216t1540) I(R6216t3918) I(R6216t5035) I(R6216t450) I(R6217t92) I(R6217t3984) I(R6217t3783) I(R6218t265) I(R6218t5145) I(R6218t4679) I(R6219t3238) I(R6219t286) I(R6219t2574) I(R6219t2230) I(R6220t3264) I(R6220t4888) I(R6220t4237) I(R6220t957) I(R6220t4833) I(R6220t1268) I(R6220t4522) I(R6221t1733) I(R6221t4835) I(R6222t2193) I(R6222t1873) I(R6223t1963) I(R6223t646) I(R6223t437) I(R6223t948) I(R6224t873) I(R6224t1989) I(R6224t2432) I(R6225t1336) I(R6225t3444) I(R6225t4806) I(R6225t5603) I(R6225t5974) I(R6226t1723) I(R6226t2692) I(R6226t2391) I(R6227t1155) I(R6227t4569) I(R6227t2962) I(R6227t2232) I(R6228t2618) I(R6228t5292) I(R6229t4114) I(R6229t1610) I(R6229t1591) I(R6229t4499) I(R6229t3227) I(R6230t1100) I(R6230t1938) I(R6230t914) I(R6231t4074) I(R6231t5708) I(R6231t3091) I(R6232t1063) I(R6232t4356) I(R6233t590) I(R6233t4822) I(R6233t5365) I(R6233t4397) I(R6233t6159) I(R6234t3587) I(R6234t3130) I(R6234t356) I(R6235t4050) I(R6235t4667) I(R6236t4882) I(R6236t862) I(R6237t1286) I(R6237t2128) I(R6237t2119) I(R6237t4769) I(R6237t6188) I(R6238t460) I(R6238t3865) I(R6238t1330) I(R6238t1279) I(R6238t2500) I(R6238t3209) I(R6239t138) I(R6239t3498) I(R6239t929) I(R6239t1986) I(R6239t4307) I(R6240t4898) I(R6240t84) I(R6240t5680) I(R6241t5063) I(R6241t3089) I(R6241t1495) I(R6241t4072) I(R6241t1695) I(R6241t283) I(R6242t310) I(R6242t5566) I(R6242t1472) I(R6242t1615) I(R6242t3353) I(R6242t4676) I(R6243t829) I(R6243t4036) I(R6243t6039) I(R6243t3024) I(R6244t1243) I(R6244t5385) I(R6244t3310) I(R6244t3827) I(R6244t748) I(R6245t3343) I(R6245t4030) I(R6245t1244) I(R6245t634) I(R6246t282) I(R6246t2156) I(R6246t297) I(R6246t255) I(R6246t3972) I(R6247t2949) I(R6247t4344) I(R6247t5337) I(R6248t3979) I(R6248t1020) I(R6248t5640) I(R6249t5779) I(R6249t981) I(R6249t816) I(R6250t4962) I(R6250t5188) I(R6250t3989) I(R6250t1633) I(R6250t3146) I(R6251t689) I(R6251t3285) I(R6251t4813) I(R6251t708) I(R6251t4392) I(R6251t4805) I(R6251t3491) I(R6252t1559) I(R6252t5283) I(R6252t3107) I(R6252t3779) I(R6252t232) I(R6252t4723) I(R6252t5410) I(R6252t1965) I(R6253t731) I(R6253t840) I(R6253t1164) I(R6253t412) I(R6254t3238) I(R6254t6219) I(R6254t1553) I(R6254t5575) I(R6254t4826) I(R6254t2230) I(R6255t5921) I(R6255t4210) I(R6255t2280) I(R6256t4635) I(R6256t1165) I(R6256t4937) I(R6256t3385) I(R6257t2043) I(R6257t902) I(R6257t4383) I(R6257t4776) I(R6257t1757) I(R6258t2187) I(R6258t2474) I(R6258t5322) I(R6258t5273) I(R6258t6153) I(R6259t325) I(R6259t4594) I(R6259t5961) I(R6260t122) I(R6260t5979) I(R6260t3679) I(R6260t5011) I(R6261t1405) I(R6261t59) I(R6261t2452) I(R6262t870) I(R6262t1879) I(R6263t1314) I(R6263t1529) I(R6263t3784) I(R6263t981) I(R6264t1866) I(R6264t4281) I(R6264t5985) I(R6265t5926) I(R6265t5386) I(R6265t1261) I(R6266t1856) I(R6266t2759) I(R6266t1647) I(R6268t5140) I(R6269t1455) I(R6269t1856) I(R6269t1647) I(R6270t407) I(R6270t5272) I(R6270t780) I(R6270t4311) I(R6271t1052) I(R6271t2487) I(R6271t1698) I(R6272t3246) I(R6272t3526) I(R6272t5069) I(R6272t4153) I(R6273t2154) I(R6273t3536) I(R6274t1085) I(R6274t2079) I(R6274t700) I(R6274t5002) I(R6274t3950) I(R6274t612) I(R6275t2729) I(R6275t5945) I(R6275t1605) I(R6275t1894) I(R6276t383) I(R6276t1474) I(R6277t3260) I(R6277t47) I(R6277t6025) I(R6277t1673) I(R6278t4106) I(R6278t5191) I(R6278t3910) I(R6278t2273) I(R6278t5242) I(R6278t93) I(R6278t3462) I(R6279t1482) I(R6279t400) I(R6279t887) I(R6279t3328) I(R6280t1229) I(R6280t5781) I(R6280t925) I(R6281t291) I(R6281t2569) I(R6281t4168) I(R6281t5866) I(R6282t2514) I(R6282t1277) I(R6282t5543) I(R6283t1750) I(R6283t5229) I(R6283t4811) I(R6283t5872) I(R6283t4194) I(R6283t3233) I(R6284t5195) I(R6284t1115) I(R6284t2996) I(R6284t46) I(R6285t3772) I(R6285t4433) I(R6285t2342) I(R6285t3438) I(R6285t2731) I(R6286t1514) I(R6286t2581) I(R6286t243) I(R6286t2902) I(R6286t4219) I(R6287t2704) I(R6287t915) I(R6287t5447) I(R6287t4950) I(R6287t2885) I(R6288t2733) I(R6288t5136) I(R6288t38) I(R6289t1726) I(R6289t4364) I(R6290t4207) I(R6290t4716) I(R6290t4230) I(R6291t5229) I(R6291t4605) I(R6291t2404) I(R6291t423) I(R6291t4811) I(R6292t4070) I(R6292t4284) I(R6292t1001) I(R6292t3973) I(R6292t1477) I(R6293t1944) I(R6293t4454) I(R6293t2897) I(R6293t2894) I(R6294t331) I(R6294t4363) I(R6294t1233) I(R6295t125) I(R6295t4891) I(R6295t3876) I(R6295t2688) I(R6296t3761) I(R6296t3815) I(R6296t5342) I(R6296t436) I(R6296t4808) I(R6297t950) I(R6297t1831) I(R6297t5948) I(R6297t4634) I(R6297t4175) I(R6297t1417) I(R6298t2665) I(R6298t5279) I(R6298t4713) I(R6299t4610) I(R6299t4549) I(R6300t1216) I(R6300t4994) I(R6300t3903) I(R6300t955) I(R6300t462) I(R6302t1079) I(R6302t3031) I(R6302t5806) I(R6302t4528) I(R6303t737) I(R6303t969) I(R6303t3220) I(R6303t404) I(R6303t4936) I(R6303t771) I(R6304t3234) I(R6304t2575) I(R6304t4976) I(R6305t2415) I(R6306t2060) I(R6306t5971) I(R6306t4966) I(R6306t5228) I(R6307t5092) I(R6307t1034) I(R6307t5921) I(R6308t1059) I(R6308t4738) I(R6308t601) I(R6308t496) I(R6309t4974) I(R6310t5197) I(R6310t4635) I(R6311t5319) I(R6311t3719) I(R6311t3648) I(R6311t1886) I(R6311t4271) I(R6312t5367) I(R6312t5671) I(R6312t246) I(R6312t3524) I(R6312t4814) I(R6312t5905) I(R6313t4945) I(R6313t258) I(R6313t5336) I(R6313t655) I(R6314t113) I(R6314t5097) I(R6314t2621) I(R6314t5224) I(R6314t507) I(R6314t3540) I(R6314t2108) I(R6315t4198) I(R6315t5504) I(R6315t214) I(R6315t3460) I(R6316t1805) I(R6316t5843) I(R6317t235) I(R6317t2104) I(R6317t4985) I(R6318t2965) I(R6318t4149) I(R6318t5826) I(R6318t2380) I(R6318t1945) I(R6318t4122) I(R6318t2158) I(R6319t2446) I(R6319t1625) I(R6319t2614) I(R6319t1) I(R6320t4027) I(R6320t4163) I(R6321t1116) I(R6321t4543) I(R6321t2565) I(R6321t4607) I(R6321t5844) I(R6321t524) I(R6322t1088) I(R6322t2082) I(R6322t1409) I(R6323t430) I(R6323t1546) I(R6323t147) I(R6323t604) I(R6324t4985) I(R6324t6078) I(R6324t3525) I(R6324t3163) I(R6325t521) I(R6325t4594) I(R6325t6259) I(R6325t947) I(R6326t3790) I(R6326t5789) I(R6326t1489) I(R6327t1731) I(R6327t5780) I(R6327t5907) I(R6327t5608) I(R6328t2512) I(R6329t701) I(R6329t2739) I(R6329t1454) I(R6329t293) I(R6330t579) I(R6330t4831) I(R6331t424) I(R6331t1752) I(R6331t2978) I(R6331t4735) I(R6332t1782) I(R6332t2635) I(R6332t3054) I(R6332t3405) I(R6333t2772) I(R6333t4243) I(R6334t1216) I(R6334t4275) I(R6334t5123) I(R6334t1357) I(R6334t5252) I(R6334t543) I(R6334t3584) I(R6335t4309) I(R6335t4056) I(R6335t5054) I(R6335t25) I(R6336t6126) I(R6337t206) I(R6337t1022) I(R6337t5753) I(R6337t5733) I(R6337t842) I(R6338t896) I(R6338t2750) I(R6338t3865) I(R6338t6322) I(R6338t2082) I(R6339t2510) I(R6339t6279) I(R6339t1482) I(R6339t56) I(R6340t156) I(R6340t5487) I(R6341t2606) I(R6341t4247) I(R6341t2882) I(R6342t1670) I(R6342t2506) I(R6343t5035) I(R6343t5584) I(R6343t1356) I(R6344t4446) I(R6344t776) I(R6344t2780) I(R6345t5396) I(R6345t210) I(R6346t6320) I(R6346t4163) I(R6346t3589) I(R6346t1901) I(R6346t5180) I(R6347t3351) I(R6347t4488) I(R6347t1264) I(R6347t6085) I(R6348t6055) I(R6348t4612) I(R6348t3657) I(R6348t1887) I(R6348t1489) I(R6349t3568) I(R6349t5910) I(R6350t5979) I(R6350t3121) I(R6351t4849) I(R6351t5310) I(R6351t4056) I(R6351t6335) I(R6351t4309) I(R6351t2115) I(R6352t646) I(R6352t1251) I(R6352t335) I(R6353t4252) I(R6353t3778) I(R6354t3166) I(R6355t2277) I(R6355t403) I(R6355t2112) I(R6356t1934) I(R6356t2753) I(R6357t5961) I(R6357t2396) I(R6357t1512) I(R6357t3261) I(R6358t2125) I(R6358t670) I(R6358t2355) I(R6359t5439) I(R6359t1973) I(R6360t2312) I(R6360t3471) I(R6360t6131) I(R6360t2789) I(R6360t34) I(R6361t1619) I(R6361t4109) I(R6361t4429) I(R6362t160) I(R6362t4524) I(R6363t5207) I(R6363t554) I(R6363t4495) I(R6364t470) I(R6364t5316) I(R6364t1541) I(R6364t179) I(R6364t5038) I(R6365t1447) I(R6365t795) I(R6365t4122) I(R6365t1521) I(R6366t1722) I(R6366t2011) I(R6367t282) I(R6367t4270) I(R6367t6246) I(R6367t5003) I(R6367t4580) I(R6367t4903) I(R6368t5824) I(R6368t2395) I(R6368t5455) I(R6368t4425) I(R6369t427) I(R6369t2072) I(R6370t2668) I(R6370t6363) I(R6370t5207) I(R6370t4025) I(R6370t4920) I(R6371t414) I(R6371t4831) I(R6371t5122) I(R6371t6330) I(R6372t2497) I(R6372t2827) I(R6372t1087) I(R6372t5997) I(R6372t2838) I(R6373t458) I(R6373t599) I(R6373t1927) I(R6373t2005) I(R6373t3407) I(R6374t3977) I(R6374t5786) I(R6374t1159) I(R6374t4641) I(R6375t4177) I(R6375t6023) I(R6375t3849) I(R6375t5720) I(R6376t2497) I(R6376t6372) I(R6376t2838) I(R6376t1484) I(R6376t3244) I(R6376t4577) I(R6376t627) I(R6377t2676) I(R6377t2193) I(R6377t2806) I(R6378t5764) I(R6378t396) I(R6378t3963) I(R6378t293) I(R6379t1898) I(R6379t6181) I(R6379t1320) I(R6379t5656) I(R6379t2314) I(R6380t943) I(R6380t1995) I(R6380t131) I(R6381t3521) I(R6381t1426) I(R6381t6092) I(R6382t1720) I(R6382t4511) I(R6382t4985) I(R6382t6324) I(R6383t5173) I(R6383t5464) I(R6383t4538) I(R6383t4188) I(R6384t100) I(R6384t4084) I(R6384t4262) I(R6384t5789) I(R6384t1430) I(R6385t4772) I(R6385t2018) I(R6385t2387) I(R6385t3435) I(R6386t3211) I(R6386t3148) I(R6387t785) I(R6387t859) I(R6387t2786) I(R6387t786) I(R6387t5636) I(R6387t1202) I(R6387t541) I(R6388t4393) I(R6388t4437) I(R6388t1135) I(R6388t414) I(R6389t2019) I(R6389t5619) I(R6389t5289) I(R6389t1337) I(R6389t2514) I(R6390t2431) I(R6390t3126) I(R6390t5331) I(R6391t6280) I(R6391t1487) I(R6391t3901) I(R6391t5929) I(R6392t3105) I(R6392t845) I(R6393t3350) I(R6393t3841) I(R6393t2599) I(R6393t3713) I(R6393t5612) I(R6393t4182) I(R6394t377) I(R6394t2170) I(R6394t4033) I(R6394t155) I(R6395t1073) I(R6395t5681) I(R6395t3250) I(R6396t1751) I(R6397t2821) I(R6397t1280) I(R6397t4299) I(R6398t2340) I(R6398t3218) I(R6398t3439) I(R6398t2374) I(R6398t5579) I(R6398t1479) I(R6399t1855) I(R6399t6198) I(R6400t5623) I(R6400t6088) I(R6400t2064) I(R6401t3399) I(R6402t3352) I(R6402t44) I(R6403t781) I(R6403t4341) I(R6403t5543) I(R6403t1277) I(R6404t5620) I(R6404t3976) I(R6404t512) I(R6404t905) I(R6404t5956) I(R6405t4830) I(R6405t3202) I(R6405t4301) I(R6405t1186) I(R6405t4478) I(R6405t3268) I(R6406t3923) I(R6406t874) I(R6406t4014) I(R6407t5085) I(R6407t2670) I(R6407t4237) I(R6407t4746) I(R6407t1637) I(R6407t3737) I(R6408t745) I(R6408t548) I(R6408t5458) I(R6408t5742) I(R6408t5783) I(R6409t3188) I(R6409t5360) I(R6409t4479) I(R6410t3583) I(R6410t184) I(R6410t4937) I(R6411t5880) I(R6412t4413) I(R6412t3725) I(R6412t658) I(R6412t3424) I(R6413t331) I(R6413t4363) I(R6414t1125) I(R6414t3053) I(R6414t5989) I(R6414t2316) I(R6415t3001) I(R6415t6004) I(R6415t2120) I(R6415t2364) I(R6416t5960) I(R6416t5885) I(R6416t3881) I(R6416t473) I(R6417t1867) I(R6418t298) I(R6418t4474) I(R6418t899) I(R6418t2824) I(R6419t1844) I(R6419t4755) I(R6419t2867) I(R6419t3408) I(R6420t1386) I(R6420t730) I(R6420t1311) I(R6421t1167) I(R6421t5573) I(R6421t1896) I(R6421t3996) I(R6422t4289) I(R6422t3226) I(R6422t1964) I(R6423t1295) I(R6423t1031) I(R6423t2459) I(R6423t6066) I(R6423t3157) I(R6424t912) I(R6424t1576) I(R6424t3550) I(R6425t2721) I(R6425t3615) I(R6426t1285) I(R6426t2050) I(R6426t1554) I(R6426t4342) I(R6426t3446) I(R6427t1386) I(R6427t833) I(R6427t724) I(R6428t4584) I(R6428t4830) I(R6428t1780) I(R6428t4536) I(R6428t3494) I(R6428t1715) I(R6428t4647) I(R6428t3202) I(R6428t6405) I(R6429t3294) I(R6429t4146) I(R6429t1771) I(R6430t1367) I(R6430t3590) I(R6430t4235) I(R6431t228) I(R6431t804) I(R6431t3699) I(R6431t5254) I(R6432t882) I(R6432t2034) I(R6432t5381) I(R6433t2197) I(R6433t5562) I(R6433t6122) I(R6433t6083) I(R6434t5116) I(R6434t4169) I(R6434t5659) I(R6435t421) I(R6435t5688) I(R6435t3660) I(R6436t4673) I(R6436t5916) I(R6436t1660) I(R6436t1816) I(R6436t3741) I(R6436t950) I(R6437t4873) I(R6437t4883) I(R6437t4215) I(R6438t5928) I(R6438t5406) I(R6438t1214) I(R6439t981) I(R6439t6263) I(R6439t3784) I(R6439t3497) I(R6440t6352) I(R6440t335) I(R6440t1172) I(R6441t1548) I(R6441t1677) I(R6441t4497) I(R6441t4076) I(R6441t317) I(R6442t215) I(R6442t4658) I(R6442t2175) I(R6442t4584) I(R6442t4450) I(R6442t2761) I(R6442t4254) I(R6443t3800) I(R6443t4039) I(R6444t768) I(R6444t2099) I(R6444t4622) I(R6444t1901) I(R6445t3168) I(R6445t6090) I(R6445t4778) I(R6445t2850) I(R6446t846) I(R6446t6095) I(R6446t3035) I(R6446t2732) I(R6446t3501) I(R6447t4643) I(R6447t5815) I(R6448t900) I(R6448t3969) I(R6448t5260) I(R6449t6194) I(R6449t1868) I(R6449t1341) I(R6449t5536) I(R6449t1382) I(R6450t195) I(R6450t5851) I(R6450t3399) I(R6450t6401) I(R6451t3230) I(R6451t3406) I(R6451t1440) I(R6452t1864) I(R6452t149) I(R6453t1651) I(R6453t3066) I(R6453t2712) I(R6453t3361) I(R6454t6175) I(R6454t30) I(R6455t909) I(R6455t5003) I(R6455t4203) I(R6455t2978) I(R6455t1127) I(R6456t6323) I(R6456t604) I(R6456t3136) I(R6457t2530) I(R6458t5044) I(R6458t153) I(R6459t5694) I(R6459t4295) I(R6460t4415) I(R6460t3189) I(R6460t1435) I(R6460t3026) I(R6460t3802) I(R6461t1987) I(R6461t5723) I(R6461t5485) I(R6461t4267) I(R6462t5593) I(R6462t5189) I(R6462t5419) I(R6462t2857) I(R6462t101) I(R6462t5793) I(R6463t2786) I(R6463t859) I(R6464t3932) I(R6464t6045) I(R6464t6001) I(R6464t5248) I(R6464t1237) I(R6464t1773) I(R6464t2697) I(R6464t2420) I(R6465t1997) I(R6465t4998) I(R6466t1446) I(R6466t1590) I(R6466t2572) I(R6466t2542) I(R6466t195) I(R6466t2461) I(R6467t2955) I(R6467t5187) I(R6467t2094) I(R6467t1373) I(R6468t2281) I(R6468t4434) I(R6468t257) I(R6468t761) I(R6470t3542) I(R6470t5919) I(R6470t4835) I(R6471t5505) I(R6471t3198) I(R6471t87) I(R6472t1968) I(R6472t2388) I(R6472t4521) I(R6472t3672) I(R6472t3837) I(R6473t864) I(R6473t3430) I(R6474t3876) I(R6474t5351) I(R6474t6075) I(R6475t2817) I(R6475t5938) I(R6475t3680) I(R6476t6000) I(R6476t5933) I(R6477t2979) I(R6477t2026) I(R6477t5145) I(R6477t4679) I(R6477t815) I(R6478t1881) I(R6478t3353) I(R6478t6242) I(R6478t4298) I(R6479t6148) I(R6479t4505) I(R6479t5190) I(R6479t5943) I(R6480t4040) I(R6480t5745) I(R6480t3601) I(R6480t1606) I(R6481t1122) I(R6481t5954) I(R6481t3086) I(R6481t5362) I(R6481t1204) I(R6482t6034) I(R6482t1954) I(R6482t3244) I(R6483t2686) I(R6483t3843) I(R6483t539) I(R6483t2863) I(R6484t2903) I(R6484t6078) I(R6484t4985) I(R6484t6317) I(R6484t1249) I(R6484t1260) I(R6485t2099) I(R6485t5111) I(R6485t5216) I(R6485t4464) I(R6486t735) I(R6486t4550) I(R6486t3627) I(R6487t1297) I(R6487t2462) I(R6487t5426) I(R6487t5888) I(R6487t6100) I(R6488t2032) I(R6488t2702) I(R6488t6452) I(R6488t1864) I(R6488t1458) I(R6489t711) I(R6489t3034) I(R6489t350) I(R6489t3343) I(R6489t6245) I(R6489t634) I(R6490t3722) I(R6490t3186) I(R6490t2058) I(R6491t2960) I(R6491t4720) I(R6491t4539) I(R6491t3792) I(R6492t3792) I(R6492t414) I(R6493t886) I(R6493t3398) I(R6493t5002) I(R6493t6274) I(R6493t3950) I(R6493t612) I(R6493t4710) I(R6494t973) I(R6494t4948) I(R6494t324) I(R6494t5886) I(R6494t3190) I(R6494t3417) I(R6494t2403) I(R6495t6132) I(R6496t1498) I(R6496t2774) I(R6496t2337) I(R6496t3726) I(R6496t2639) I(R6496t1794) I(R6497t763) I(R6497t816) I(R6497t6249) I(R6497t981) I(R6497t586) I(R6498t2455) I(R6498t3052) I(R6498t4418) I(R6499t2234) I(R6499t366) I(R6499t869) I(R6499t4192) I(R6499t2389) I(R6499t2300) I(R6499t5813) I(R6499t4660) I(R6500t3760) I(R6500t4238) I(R6500t2073) I(R6501t5114) I(R6502t4809) I(R6502t5808) I(R6502t3683) I(R6502t6058) I(R6502t3059) I(R6503t1334) I(R6503t3002) I(R6503t5380) I(R6503t3689) I(R6503t5027) I(R6503t3023) I(R6503t4852) I(R6503t5869) I(R6503t5673) I(R6503t36) I(R6503t755) I(R6504t4252) I(R6504t1504) I(R6504t647) I(R6504t1872) I(R6505t555) I(R6505t6086) I(R6505t5600) I(R6505t4369) I(R6505t3975) I(R6506t3211) I(R6506t6386) I(R6506t6159) I(R6506t1800) I(R6507t2243) I(R6507t4136) I(R6507t1892) I(R6507t3065) I(R6507t3730) I(R6508t3722) I(R6508t3186) I(R6508t2166) I(R6508t1820) I(R6509t730) I(R6509t1386) I(R6509t6427) I(R6509t724) I(R6509t2617) I(R6509t3915) I(R6509t2098) I(R6510t442) I(R6510t2465) I(R6512t4437) I(R6512t4705) I(R6512t5439) I(R6512t1135) I(R6513t4752) I(R6513t4934) I(R6513t3532) I(R6513t1966) I(R6514t1178) I(R6514t1388) I(R6514t549) I(R6514t4077) I(R6514t2424) I(R6515t5357) I(R6515t962) I(R6515t1810) I(R6515t6061) I(R6516t3420) I(R6516t1197) I(R6517t5638) I(R6517t496) I(R6517t6308) I(R6517t1059) I(R6518t1705) I(R6518t4446) I(R6518t2780) I(R6518t6344) I(R6519t1876) I(R6519t3008) I(R6519t1537) I(R6520t780) I(R6521t830) I(R6521t5226) I(R6521t516) I(R6521t2153) I(R6522t5615) I(R6522t2931) I(R6522t2193) I(R6522t6222) I(R6523t4642) I(R6523t4870) I(R6523t365) I(R6523t2422) I(R6523t3355) I(R6524t4199) I(R6524t4563) I(R6524t2077) I(R6524t136) I(R6524t5235) I(R6524t5004) I(R6525t5058) I(R6525t4867) I(R6525t5846) I(R6525t914) I(R6526t625) I(R6526t5036) I(R6526t80) I(R6526t4745) I(R6527t4601) I(R6527t3223) I(R6527t6119) I(R6527t2901) I(R6528t178) I(R6528t4247) I(R6528t1320) I(R6528t5656) I(R6528t1188) I(R6529t5000) I(R6529t2947) I(R6529t5571) I(R6530t2481) I(R6530t2849) I(R6530t1663) I(R6531t1471) I(R6531t417) I(R6531t5056) I(R6532t421) I(R6532t6435) I(R6533t147) I(R6533t435) I(R6533t1546) I(R6533t5022) I(R6534t348) I(R6534t3957) I(R6534t6011) I(R6534t1047) I(R6534t3102) I(R6535t464) I(R6535t3906) I(R6535t2755) I(R6535t1359) I(R6535t6479) I(R6535t6148) I(R6536t167) I(R6536t1629) I(R6536t1861) I(R6536t5155) I(R6536t2612) I(R6536t1365) I(R6537t318) I(R6537t592) I(R6537t2389) I(R6537t613) I(R6537t55) I(R6538t2129) I(R6538t5980) I(R6538t1571) I(R6538t3603) I(R6539t4354) I(R6539t3695) I(R6539t3070) I(R6540t372) I(R6540t5171) I(R6540t5629) I(R6540t1194) I(R6540t4485) I(R6541t4608) I(R6541t5942) I(R6541t2179) I(R6541t1674) I(R6541t2913) I(R6541t5766) I(R6542t4945) I(R6542t6313) I(R6542t258) I(R6542t5627) I(R6543t1712) I(R6543t5336) I(R6543t6313) I(R6543t3326) I(R6543t2565) I(R6543t6321) I(R6543t4607) I(R6543t6077) I(R6544t2206) I(R6544t1776) I(R6545t2551) I(R6546t3276) I(R6546t5680) I(R6547t1896) I(R6547t6421) I(R6547t5054) I(R6547t4056) I(R6547t5573) I(R6548t828) I(R6548t5716) I(R6548t259) I(R6548t1356) I(R6548t3167) I(R6549t3305) I(R6549t4588) I(R6549t5977) I(R6550t2741) I(R6550t3483) I(R6550t5641) I(R6550t5421) I(R6550t3082) I(R6550t2314) I(R6551t377) I(R6551t270) I(R6551t1089) I(R6551t6188) I(R6552t2848) I(R6552t2944) I(R6552t4817) I(R6552t5032) I(R6553t1405) I(R6553t3716) I(R6553t600) I(R6554t4157) I(R6554t5048) I(R6554t4873) I(R6554t6437) I(R6554t4215) I(R6555t306) I(R6555t1807) I(R6556t2935) I(R6556t5139) I(R6556t2293) I(R6557t4411) I(R6557t5981) I(R6558t1440) I(R6558t1475) I(R6558t3011) I(R6558t471) I(R6558t4116) I(R6559t1891) I(R6559t5077) I(R6559t3270) I(R6560t3331) I(R6560t5344) I(R6561t2756) I(R6561t4796) I(R6561t5944) I(R6561t5124) I(R6561t3377) I(R6561t2149) I(R6562t1064) I(R6562t1432) I(R6562t2962) I(R6562t6227) I(R6562t1155) I(R6563t4054) I(R6563t5100) I(R6563t1715) I(R6563t4647) I(R6563t3352) I(R6564t110) I(R6564t4416) I(R6564t1646) I(R6564t986) I(R6564t4854) I(R6564t5078) I(R6565t2403) I(R6565t6166) I(R6566t4482) I(R6566t2099) I(R6566t1848) I(R6567t2529) I(R6567t5740) I(R6567t302) I(R6568t5416) I(R6568t3633) I(R6568t2945) I(R6568t4646) I(R6569t1859) I(R6569t2588) I(R6569t5473) I(R6569t4239) I(R6569t3781) I(R6569t2884) I(R6570t317) I(R6570t4373) I(R6570t5611) I(R6570t3720) I(R6571t3548) I(R6571t135) I(R6572t1798) I(R6572t4071) I(R6572t4700) I(R6573t5440) I(R6573t3744) I(R6574t17) I(R6574t822) I(R6574t3204) I(R6574t649) I(R6575t3179) I(R6576t814) I(R6576t2411) I(R6576t3921) I(R6577t2070) I(R6577t4475) I(R6577t1468) I(R6578t113) I(R6578t6314) I(R6578t2108) I(R6578t1742) I(R6578t4093) I(R6578t2116) I(R6579t1841) I(R6579t5502) I(R6579t2481) I(R6579t6530) I(R6580t3851) I(R6580t5320) I(R6580t3612) I(R6581t3075) I(R6581t3821) I(R6581t2872) I(R6581t1883) I(R6581t91) I(R6582t5803) I(R6582t1663) I(R6582t2201) I(R6582t1899) I(R6583t517) I(R6583t3981) I(R6584t6340) I(R6584t5487) I(R6584t5137) I(R6584t3311) I(R6585t2243) I(R6585t5484) I(R6585t3185) I(R6586t2294) I(R6586t2286) I(R6587t1121) I(R6587t5904) I(R6587t2333) I(R6587t2915) I(R6588t2688) I(R6588t2820) I(R6588t6075) I(R6588t4907) I(R6589t1870) I(R6589t4135) I(R6589t4747) I(R6590t5955) I(R6591t5408) I(R6591t5640) I(R6591t6248) I(R6591t1838) I(R6592t5947) I(R6592t6168) I(R6592t3522) I(R6593t3414) I(R6593t5428) I(R6593t5747) I(R6593t1230) I(R6594t1759) I(R6594t1172) I(R6594t6440) I(R6595t98) I(R6595t4526) I(R6595t3090) I(R6595t2546) I(R6595t5110) I(R6595t108) I(R6595t2331) I(R6596t3230) I(R6596t6451) I(R6596t1854) I(R6596t4056) I(R6596t6351) I(R6596t4849) I(R6596t3406) I(R6598t139) I(R6598t972) I(R6598t1592) I(R6598t2815) I(R6599t1391) I(R6599t1486) I(R6600t5805) I(R6600t2367) I(R6600t5533) I(R6600t676) I(R6600t4150) I(R6601t4675) I(R6601t4361) I(R6601t4599) I(R6601t1672) I(R6602t74) I(R6602t2692) I(R6602t841) I(R6602t5403) I(R6603t4639) I(R6603t4942) I(R6603t1812) I(R6603t3634) I(R6604t4177) I(R6604t6375) I(R6605t872) I(R6605t6476) I(R6605t5933) I(R6605t951) I(R6606t1507) I(R6606t5650) I(R6606t2713) I(R6606t4320) I(R6606t1580) I(R6607t5542) I(R6607t4808) I(R6607t3709) I(R6607t4214) I(R6607t5635) I(R6607t4914) I(R6608t911) I(R6608t6175) I(R6608t6454) I(R6608t6079) I(R6608t880) I(R6609t4772) I(R6609t6385) I(R6609t2018) I(R6609t3478) I(R6610t2567) I(R6610t968) I(R6611t28) I(R6611t2042) I(R6611t5425) I(R6611t1230) I(R6612t5431) I(R6612t5040) I(R6612t1506) I(R6612t3587) I(R6612t6234) I(R6613t575) I(R6613t6029) I(R6613t2276) I(R6613t1694) I(R6613t57) I(R6613t393) I(R6613t977) I(R6614t6590) I(R6614t2832) I(R6614t5541) I(R6614t3507) I(R6615t5928) I(R6615t6438) I(R6615t3700) I(R6615t1801) I(R6615t5406) I(R6616t727) I(R6616t2702) I(R6616t2032) I(R6616t4656) I(R6616t3800) I(R6616t2925) I(R6617t1276) I(R6617t4405) I(R6618t4503) I(R6618t5519) I(R6618t201) I(R6618t578) I(R6619t1483) I(R6619t6043) I(R6619t3166) I(R6619t6354) I(R6619t5233) I(R6620t620) I(R6620t900) I(R6620t939) I(R6620t5425) I(R6620t6611) I(R6620t2042) I(R6621t3676) I(R6621t3228) I(R6621t3995) I(R6622t5947) I(R6622t6592) I(R6622t2038) I(R6623t3930) I(R6623t4876) I(R6623t3443) I(R6623t995) I(R6623t2918) I(R6623t6147) I(R6624t2424) I(R6624t3112) I(R6624t2652) I(R6624t1368) I(R6625t1729) I(R6625t4181) I(R6625t1423) I(R6625t2238) I(R6626t5176) I(R6626t5318) I(R6626t5901) I(R6626t1162) I(R6626t242) I(R6627t3309) I(R6627t140) I(R6627t3740) I(R6627t765) I(R6627t1808) I(R6628t208) I(R6628t1460) I(R6628t5823) I(R6628t571) I(R6628t4645) I(R6629t287) I(R6629t3106) I(R6630t1532) I(R6630t4538) I(R6630t6383) I(R6630t4188) I(R6630t4484) I(R6630t2420) I(R6631t1511) I(R6631t4057) I(R6631t1456) I(R6631t1942) I(R6631t2348) I(R6632t117) I(R6632t2346) I(R6632t5008) I(R6632t1461) I(R6632t2366) I(R6632t878) I(R6633t2368) I(R6633t4751) I(R6633t5498) I(R6633t5592) I(R6634t5683) I(R6634t26) I(R6634t819) I(R6634t5908) I(R6635t944) I(R6635t2707) I(R6635t131) I(R6635t4412) I(R6635t3514) I(R6636t1838) I(R6636t6591) I(R6636t6248) I(R6636t1020) I(R6636t3743) I(R6636t2559) I(R6637t3302) I(R6637t6267) I(R6637t639) I(R6637t5866) I(R6638t5423) I(R6638t5481) I(R6638t1369) I(R6638t5507) I(R6638t6301) I(R6639t6169) I(R6639t4153) I(R6639t2682) I(R6640t3868) I(R6640t4201) I(R6640t1770) I(R6641t3412) I(R6641t4885) I(R6641t3555) I(R6641t358) I(R6641t671) I(R6641t2487) I(R6641t6271) I(R6641t1052) I(R6641t1378) I(R6642t4614) I(R6642t1645) I(R6642t1812) I(R6642t3614) I(R6642t5506) I(R6642t2936) I(R6643t1418) I(R6643t4603) I(R6643t740) I(R6644t5973) I(R6644t2399) I(R6644t4514) I(R6644t5350) I(R6644t4846) I(R6645t2689) I(R6645t5917) I(R6645t46) I(R6645t4483) I(R6645t849) I(R6647t3505) I(R6647t3776) I(R6648t1922) I(R6648t5817) I(R6648t4234) I(R6649t2538) I(R6649t5405) I(R6649t1195) I(R6649t1084) I(R6649t5483) I(R6649t2871) I(R6650t467) I(R6650t213) I(R6650t5968) I(R6650t2550) I(R6650t783) I(R6650t244) I(R6651t305) I(R6651t5491) I(R6651t5469) I(R6651t4482) I(R6651t3531) I(R6652t2791) I(R6652t5335) I(R6652t3080) I(R6652t2762) I(R6653t5856) I(R6653t2028) I(R6653t6116) I(R6654t3900) I(R6654t4859) I(R6654t709) I(R6654t977) I(R6654t3397) I(R6655t991) I(R6655t4730) I(R6655t6111) I(R6655t6000) I(R6656t1375) I(R6656t3928) I(R6656t5868) I(R6656t3656) I(R6657t1306) I(R6657t2663) I(R6657t337) I(R6657t2326) I(R6658t919) I(R6658t5936) I(R6658t1557) I(R6659t4908) I(R6659t3417) I(R6659t3190) I(R6659t2329) I(R6659t3673) I(R6660t1028) I(R6660t6192) I(R6660t5635) I(R6660t2443) I(R6660t1403) I(R6660t4227) I(R6660t1400) I(R6660t6180) I(R6661t1531) I(R6661t5493) I(R6661t5300) I(R6661t4406) I(R6661t2323) I(R6662t197) I(R6662t4815) I(R6662t4555) I(R6662t6123) I(R6662t647) I(R6663t2659) I(R6663t3653) I(R6663t5032) I(R6663t2188) I(R6663t1305) I(R6664t3357) I(R6664t4346) I(R6664t2279) I(R6664t4748) I(R6664t4024) I(R6665t1986) I(R6665t4697) I(R6665t3141) I(R6665t2925) I(R6666t78) I(R6666t1097) I(R6666t1192) I(R6666t4585) I(R6666t5514) I(R6666t3393) I(R6666t4954) I(R6667t51) I(R6667t367) I(R6667t3409) I(R6668t1674) I(R6668t2913) I(R6668t5466) I(R6668t532) I(R6668t5317) I(R6668t1569) I(R6668t3954) I(R6669t1970) I(R6669t58) I(R6670t5172) I(R6670t3280) I(R6670t3121) I(R6671t1547) I(R6671t2764) I(R6672t6362) I(R6672t285) I(R6672t4524) I(R6673t1450) I(R6673t5818) I(R6673t5699) I(R6673t1152) I(R6673t44) I(R6674t1443) I(R6674t3956) I(R6674t2148) I(R6674t6122) I(R6674t2620) I(R6675t2810) I(R6675t417) I(R6675t5056) I(R6676t2133) I(R6676t1865) I(R6677t666) I(R6677t311) I(R6677t5745) I(R6677t5284) I(R6678t3704) I(R6678t4652) I(R6678t1644) I(R6678t5390) I(R6678t5610) I(R6678t6172) I(R6679t365) I(R6679t2441) I(R6679t6523) I(R6680t1404) I(R6680t2981) I(R6680t3639) I(R6681t1336) I(R6681t3444) I(R6681t2021) I(R6681t4840) I(R6681t5974) I(R6682t2876) I(R6682t5238) I(R6682t3611) I(R6683t202) I(R6683t2647) I(R6683t3586) I(R6684t4731) I(R6684t52) I(R6684t758) I(R6685t225) I(R6685t1261) I(R6685t5603) I(R6685t4249) I(R6686t408) I(R6686t5412) I(R6686t5981) I(R6686t3195) I(R6687t6154) I(R6687t530) I(R6687t1186) I(R6687t4301) I(R6688t1027) I(R6688t1756) I(R6688t2555) I(R6688t4615) I(R6689t3622) I(R6689t2363) I(R6689t5306) I(R6690t5852) I(R6691t3767) I(R6691t5442) I(R6691t5393) I(R6692t497) I(R6692t5398) I(R6692t4640) I(R6693t579) I(R6693t4624) I(R6693t5122) I(R6693t6371) I(R6693t6330) I(R6694t2687) I(R6694t1241) I(R6694t6273) I(R6695t2419) I(R6695t4440) I(R6695t1940) I(R6696t3804) I(R6696t3794) I(R6696t2839) I(R6697t3115) I(R6697t5946) I(R6697t3700) I(R6697t2027) I(R6697t3124) I(R6697t66) I(R6698t1180) I(R6698t4618) I(R6698t2400) I(R6698t2991) I(R6698t3709) I(R6698t4808) I(R6699t4287) I(R6699t37) I(R6700t1894) I(R6700t4541) I(R6700t6275) I(R6700t2729) I(R6701t985) I(R6701t2007) I(R6701t733) I(R6701t2016) I(R6702t23) I(R6702t4749) I(R6702t1013) I(R6702t5226) I(R6702t6521) I(R6703t1048) I(R6703t6197) I(R6703t226) I(R6703t168) I(R6704t1959) I(R6704t4557) I(R6704t6097) I(R6705t6508) I(R6705t3722) I(R6705t924) I(R6705t694) I(R6706t3312) I(R6706t4414) I(R6707t4767) I(R6707t5146) I(R6707t2705) I(R6707t2567) I(R6708t1073) I(R6708t2404) I(R6708t419) I(R6709t670) I(R6709t5237) I(R6709t2723) I(R6709t2355) I(R6710t6344) I(R6710t6155) I(R6710t1897) I(R6710t4184) I(R6710t3191) I(R6710t2780) I(R6710t776) I(R6711t5620) I(R6711t6404) I(R6711t5956) I(R6711t4288) I(R6712t369) I(R6712t6127) I(R6712t1945) I(R6712t2380) I(R6712t4279) I(R6712t5280) I(R6713t2038) I(R6713t6622) I(R6713t6592) I(R6713t1408) I(R6714t5017) I(R6714t4193) I(R6714t4236) I(R6714t3684) I(R6715t1939) I(R6715t2873) I(R6715t2358) I(R6715t2764) I(R6715t6671) I(R6715t1547) I(R6715t3327) I(R6716t546) I(R6716t3281) I(R6716t3144) I(R6717t25) I(R6717t5191) I(R6718t3621) I(R6718t6643) I(R6718t1418) I(R6718t697) I(R6719t4125) I(R6719t3862) I(R6719t2026) I(R6719t5920) I(R6720t6081) I(R6720t5143) I(R6720t963) I(R6721t4072) I(R6721t4579) I(R6721t2641) I(R6721t1041) I(R6722t1678) I(R6722t4290) I(R6722t4487) I(R6722t3814) I(R6723t5281) I(R6723t143) I(R6723t121) I(R6723t1784) I(R6724t162) I(R6724t1772) I(R6724t736) I(R6725t2792) I(R6725t5352) I(R6725t1599) I(R6726t5626) I(R6726t2029) I(R6726t2798) I(R6726t774) I(R6726t4889) I(R6727t5637) I(R6727t4477) I(R6727t189) I(R6728t1252) I(R6728t5883) I(R6728t2139) I(R6728t1943) I(R6728t6112) I(R6729t3536) I(R6729t560) I(R6729t4748) I(R6730t754) I(R6730t1164) I(R6730t6253) I(R6730t412) I(R6730t641) I(R6731t5538) I(R6731t667) I(R6731t5539) I(R6731t3142) I(R6732t494) I(R6732t6187) I(R6732t2488) I(R6732t5133) I(R6733t1657) I(R6733t1676) I(R6733t1162) I(R6733t3194) I(R6733t4052) I(R6733t1123) I(R6734t1377) I(R6734t4358) I(R6734t2211) I(R6735t2693) I(R6735t948) I(R6735t437) I(R6736t770) I(R6736t5027) I(R6736t1163) I(R6736t2335) I(R6737t583) I(R6737t857) I(R6737t3785) I(R6738t625) I(R6738t6526) I(R6738t5036) I(R6739t3179) I(R6739t5677) I(R6739t2749) I(R6739t3497) I(R6740t6096) I(R6740t170) I(R6740t2227) I(R6741t6362) I(R6741t6672) I(R6741t285) I(R6742t5699) I(R6742t4114) I(R6742t1144) I(R6743t5332) I(R6743t6108) I(R6743t2369) I(R6743t5809) I(R6744t2252) I(R6744t6349) I(R6745t5508) I(R6745t518) I(R6746t3439) I(R6746t4503) I(R6746t2374) I(R6746t3396) I(R6746t1775) I(R6747t2020) I(R6747t6170) I(R6748t2388) I(R6748t6149) I(R6748t6162) I(R6748t6526) I(R6748t625) I(R6748t5156) I(R6748t818) I(R6749t4098) I(R6749t5288) I(R6749t2631) I(R6749t2432) I(R6750t1624) I(R6750t1863) I(R6750t223) I(R6750t3817) I(R6750t4292) I(R6750t5052) I(R6750t4319) I(R6751t2876) I(R6751t5238) I(R6751t4276) I(R6751t2629) I(R6752t1978) I(R6752t3028) I(R6752t2317) I(R6753t812) I(R6753t5608) I(R6753t3279) I(R6753t928) I(R6753t5973) I(R6754t6204) I(R6754t5219) I(R6754t2376) I(R6754t3574) I(R6754t3744) I(R6755t3166) I(R6755t3728) I(R6755t461) I(R6755t6043) I(R6755t6619) I(R6756t5659) I(R6756t6434) I(R6756t2812) I(R6756t4197) I(R6756t4169) I(R6757t1324) I(R6757t2501) I(R6757t4400) I(R6757t6035) I(R6757t3339) I(R6757t5046) I(R6757t4469) I(R6758t1536) I(R6758t1549) I(R6758t3663) I(R6758t640) I(R6758t2184) I(R6758t5622) I(R6759t2107) I(R6759t639) I(R6759t291) I(R6759t3645) I(R6760t640) I(R6760t6758) I(R6760t2184) I(R6760t3603) I(R6760t5340) I(R6761t5090) I(R6761t3905) I(R6761t716) I(R6762t3495) I(R6762t5467) I(R6762t1331) I(R6762t4023) I(R6763t224) I(R6763t2511) I(R6763t3358) I(R6763t1402) I(R6764t560) I(R6764t3536) I(R6764t2154) I(R6764t1620) I(R6765t1143) I(R6765t4317) I(R6765t4010) I(R6765t1023) I(R6766t4531) I(R6766t2225) I(R6766t5714) I(R6766t2205) I(R6767t4968) I(R6767t157) I(R6767t451) I(R6767t5601) I(R6767t6328) I(R6767t2512) I(R6768t6723) I(R6768t4414) I(R6768t4863) I(R6768t4005) I(R6768t2784) I(R6768t121) I(R6769t2328) I(R6769t5803) I(R6769t2551) I(R6769t6530) I(R6769t1663) I(R6769t6582) I(R6770t1400) I(R6770t1583) I(R6770t3484) I(R6770t661) I(R6770t798) I(R6770t1829) I(R6771t2284) I(R6771t3436) I(R6771t5099) I(R6771t5732) I(R6771t3630) I(R6771t2203) I(R6771t340) I(R6772t3830) I(R6772t4420) I(R6772t956) I(R6772t3001) I(R6772t2662) I(R6772t304) I(R6773t200) I(R6773t875) I(R6773t2353) I(R6773t3100) I(R6773t3637) I(R6774t228) I(R6774t4344) I(R6774t6431) I(R6774t5254) I(R6774t5646) I(R6774t1915) I(R6775t2157) I(R6775t6080) I(R6775t3381) I(R6775t5986) I(R6775t938) I(R6776t1290) I(R6776t3037) I(R6776t3245) I(R6776t1665) I(R6776t4419) I(R6776t192) I(R6777t3067) I(R6777t1793) I(R6777t126) I(R6777t3695) I(R6777t778) I(R6778t3012) I(R6778t3750) I(R6778t5543) I(R6778t6282) I(R6778t3024) I(R6778t2648) I(R6779t1426) I(R6779t6381) I(R6779t866) I(R6779t3105) I(R6779t845) I(R6779t753) I(R6779t1565) I(R6779t1361) I(R6780t2285) I(R6780t449) I(R6780t5157) I(R6780t4911) I(R6781t5953) I(R6781t5859) I(R6781t4512) I(R6782t4061) I(R6782t1262) I(R6783t1343) I(R6783t3780) I(R6783t6693) I(R6783t5122) I(R6783t2937) I(R6784t1733) I(R6784t6221) I(R6784t4835) I(R6784t1054) I(R6785t2121) I(R6785t2522) I(R6785t5360) I(R6786t3893) I(R6786t4507) I(R6787t2481) I(R6787t4889) I(R6787t6726) I(R6788t244) I(R6788t3857) I(R6788t4973) I(R6788t6279) I(R6789t2425) I(R6789t3999) I(R6789t2989) I(R6789t3790) I(R6789t2196) I(R6789t4769) I(R6790t1538) I(R6790t2421) I(R6790t5186) I(R6790t3247) I(R6790t668) I(R6791t854) I(R6791t2691) I(R6791t4245) I(R6791t751) I(R6791t5023) I(R6791t519) I(R6791t3318) I(R6791t2504) I(R6792t2530) I(R6792t233) I(R6793t4375) I(R6793t5993) I(R6793t2594) I(R6793t2347) I(R6794t616) I(R6794t5066) I(R6794t1219) I(R6795t5791) I(R6795t3914) I(R6795t5030) I(R6796t5191) I(R6796t6717) I(R6796t3462) I(R6796t6278) I(R6797t5289) I(R6797t4220) I(R6797t5619) I(R6797t6389) I(R6798t2998) I(R6799t5547) I(R6799t4095) I(R6799t5940) I(R6800t582) I(R6800t1016) I(R6800t389) I(R6801t160) I(R6801t1236) I(R6801t5675) I(R6801t1611) I(R6801t5218) I(R6801t4524) I(R6802t1769) I(R6802t5076) I(R6802t3456) I(R6802t1872) I(R6802t3037) I(R6802t1290) I(R6802t1706) I(R6803t5254) I(R6803t375) I(R6803t1055) I(R6803t2078) I(R6803t1915) I(R6804t459) I(R6804t5489) I(R6804t2660) I(R6804t15) I(R6804t5564) I(R6804t1975) I(R6805t3253) I(R6805t963) I(R6805t4278) I(R6805t3441) I(R6805t4250) I(R6806t1815) I(R6806t3535) I(R6807t5724) I(R6807t3853) I(R6807t2319) I(R6808t2105) I(R6808t3803) I(R6808t3175) I(R6808t1537) I(R6808t6519) I(R6808t1876) I(R6808t1903) I(R6809t1615) I(R6809t5204) I(R6809t2172) I(R6809t3877) I(R6810t3733) I(R6810t1012) I(R6810t2716) I(R6810t3295) I(R6810t1860) I(R6811t3197) I(R6811t5714) I(R6811t2205) I(R6811t3094) I(R6811t2828) I(R6811t5245) I(R6812t3753) I(R6812t1748) I(R6812t1454) I(R6812t1067) I(R6813t2551) I(R6813t6545) I(R6813t163) I(R6813t6128) I(R6813t2013) I(R6814t2995) I(R6814t5182) I(R6814t2597) I(R6814t5879) I(R6815t763) I(R6815t1446) I(R6815t659) I(R6815t3010) I(R6816t1121) I(R6816t6587) I(R6816t2915) I(R6816t5369) I(R6817t2594) I(R6817t5625) I(R6817t4375) I(R6817t3958) I(R6818t374) I(R6818t6501) I(R6818t5114) I(R6819t4311) I(R6819t5102) I(R6819t780) I(R6819t4810) I(R6819t1821) I(R6820t644) I(R6820t1635) I(R6820t5845) I(R6820t2475) I(R6820t5682) I(R6821t3401) I(R6821t5976) I(R6821t4526) I(R6821t1999) I(R6821t5743) I(R6822t2020) I(R6822t6747) I(R6823t1846) I(R6823t3869) I(R6823t2568) I(R6823t1104) I(R6823t4930) I(R6824t298) I(R6824t4383) I(R6824t5638) I(R6824t1059) I(R6824t4738) I(R6825t3258) I(R6825t5250) I(R6825t4152) I(R6825t2375) I(R6825t4165) I(R6826t1418) I(R6826t6643) I(R6826t740) I(R6826t633) I(R6827t10) I(R6827t92) I(R6827t4780) I(R6828t1371) I(R6828t4348) I(R6828t4267) I(R6828t2110) I(R6829t5107) I(R6829t6088) I(R6829t6544) I(R6830t1257) I(R6830t5109) I(R6830t5941) I(R6830t313) I(R6830t3832) I(R6831t632) I(R6831t2865) I(R6832t2862) I(R6832t3334) I(R6832t5598) I(R6832t5256) I(R6833t44) I(R6833t4054) I(R6833t3352) I(R6833t6402) I(R6834t6731) I(R6834t3142) I(R6834t2204) I(R6834t1417) I(R6834t6297) I(R6835t5116) I(R6835t2618) I(R6835t5257) I(R6835t5888) I(R6836t5689) I(R6836t469) I(R6836t3419) I(R6836t3788) I(R6836t535) I(R6837t3559) I(R6837t5998) I(R6837t2893) I(R6837t2861) I(R6838t2181) I(R6838t2492) I(R6839t423) I(R6839t1360) I(R6839t1441) I(R6839t1427) I(R6839t4556) I(R6839t1616) I(R6840t5381) I(R6840t5777) I(R6840t853) I(R6840t2843) I(R6840t2034) I(R6841t3234) I(R6841t1232) I(R6841t4397) I(R6842t2015) I(R6842t3649) I(R6842t3432) I(R6842t5282) I(R6843t6386) I(R6843t6506) I(R6843t6159) I(R6843t3148) I(R6844t1951) I(R6844t5096) I(R6844t4229) I(R6845t2183) I(R6845t4999) I(R6845t1801) I(R6845t2768) I(R6845t302) I(R6846t4718) I(R6846t5451) I(R6846t746) I(R6846t5715) I(R6846t6145) I(R6846t1769) I(R6847t1229) I(R6847t6280) I(R6847t5781) I(R6847t1943) I(R6847t2244) I(R6847t1983) I(R6848t527) I(R6848t4062) I(R6848t4196) I(R6849t446) I(R6849t5071) I(R6849t5251) I(R6849t988) I(R6850t3665) I(R6850t6085) I(R6850t1264) I(R6850t514) I(R6851t152) I(R6851t6065) I(R6851t6060) I(R6851t3151) I(R6852t1081) I(R6852t5079) I(R6852t1540) I(R6852t6216) I(R6852t3918) I(R6853t3257) I(R6853t1857) I(R6853t4045) I(R6853t3352) I(R6853t6402) I(R6854t728) I(R6854t1563) I(R6854t2415) I(R6854t5348) I(R6855t2328) I(R6855t1149) I(R6855t3959) I(R6855t1328) I(R6856t2904) I(R6856t1323) I(R6856t5189) I(R6856t3935) I(R6857t277) I(R6857t5259) I(R6857t6135) I(R6857t3561) I(R6857t1538) I(R6858t5650) I(R6858t3172) I(R6858t2470) I(R6858t5878) I(R6859t3532) I(R6859t1966) I(R6859t4845) I(R6859t4289) I(R6859t2718) I(R6860t705) I(R6860t2229) I(R6860t2216) I(R6860t424) I(R6860t4903) I(R6860t5520) I(R6860t1714) I(R6861t145) I(R6861t1528) I(R6861t1771) I(R6861t6429) I(R6862t173) I(R6862t2803) I(R6862t292) I(R6862t904) I(R6862t2715) I(R6863t6798) I(R6863t343) I(R6864t1451) I(R6864t5) I(R6865t5631) I(R6865t3982) I(R6865t3749) I(R6865t3138) I(R6865t1040) I(R6865t490) I(R6866t2614) I(R6866t4340) I(R6866t1625) I(R6866t3039) I(R6866t4202) I(R6867t3696) I(R6867t5461) I(R6867t2069) I(R6867t4013) I(R6867t6051) I(R6868t3019) I(R6868t1668) I(R6868t4710) I(R6868t4047) I(R6869t1695) I(R6869t5366) I(R6869t3134) I(R6869t5048) I(R6870t2741) I(R6870t3483) I(R6870t5641) I(R6870t6181) I(R6870t1898) I(R6871t4951) I(R6871t1998) I(R6871t4231) I(R6872t4051) I(R6872t5402) I(R6872t4104) I(R6872t5558) I(R6872t1281) I(R6873t2254) I(R6873t6447) I(R6873t5815) I(R6873t4002) I(R6874t1203) I(R6874t2246) I(R6874t1117) I(R6874t4087) I(R6874t5966) I(R6875t2301) I(R6875t2933) I(R6875t5740) I(R6875t1930) I(R6876t4939) I(R6876t6115) I(R6876t2014) I(R6876t1653) I(R6876t3991) I(R6877t1226) I(R6877t2050) I(R6877t1285) I(R6878t2292) I(R6878t4962) I(R6878t1041) I(R6878t3146) I(R6878t6250) I(R6879t1759) I(R6879t6594) I(R6879t4632) I(R6879t4832) I(R6879t948) I(R6879t1963) I(R6879t6440) I(R6880t2322) I(R6880t5508) I(R6880t6745) I(R6881t317) I(R6881t1644) I(R6881t5390) I(R6881t3720) I(R6881t6570) I(R6882t379) I(R6882t5944) I(R6882t5124) I(R6882t1105) I(R6883t3463) I(R6883t1051) I(R6884t4324) I(R6884t5293) I(R6884t3266) I(R6885t209) I(R6885t873) I(R6885t6224) I(R6885t2432) I(R6886t2096) I(R6886t2533) I(R6887t3518) I(R6887t5747) I(R6887t6135) I(R6887t3561) I(R6887t2421) I(R6887t3032) I(R6887t5428) I(R6888t4519) I(R6888t6583) I(R6888t3981) I(R6888t5445) I(R6888t5007) I(R6889t2817) I(R6889t4790) I(R6889t4844) I(R6889t6475) I(R6890t1613) I(R6890t4241) I(R6890t1921) I(R6890t3403) I(R6890t3547) I(R6891t3257) I(R6891t1103) I(R6891t1242) I(R6891t5984) I(R6891t1857) I(R6891t6853) I(R6892t3822) I(R6892t5166) I(R6892t465) I(R6893t2992) I(R6893t3863) I(R6893t5850) I(R6893t6267) I(R6894t882) I(R6894t4120) I(R6894t382) I(R6894t5522) I(R6894t5692) I(R6895t2790) I(R6895t5446) I(R6895t2636) I(R6895t2735) I(R6896t4354) I(R6896t4637) I(R6896t3701) I(R6897t1521) I(R6897t3014) I(R6897t827) I(R6898t4834) I(R6898t685) I(R6898t488) I(R6899t4089) I(R6899t4864) I(R6899t2619) I(R6899t1681) I(R6900t2695) I(R6900t4097) I(R6900t760) I(R6901t2018) I(R6901t706) I(R6901t2387) I(R6902t6647) I(R6902t3505) I(R6903t2277) I(R6903t6355) I(R6903t5313) I(R6904t6221) I(R6904t5919) I(R6904t6470) I(R6904t4835) I(R6905t4288) I(R6905t6711) I(R6905t6067) I(R6905t1596) I(R6905t5956) I(R6906t2603) I(R6906t3068) I(R6906t3639) I(R6906t5262) I(R6906t3970) I(R6906t4663) I(R6906t1044) I(R6907t611) I(R6907t4218) I(R6907t2460) I(R6907t4930) I(R6907t2971) I(R6907t1389) I(R6908t3468) I(R6909t1475) I(R6909t6558) I(R6909t3230) I(R6910t3937) I(R6911t1276) I(R6911t6617) I(R6911t1250) I(R6911t2716) I(R6912t2310) I(R6912t4930) I(R6912t2460) I(R6912t1474) I(R6912t725) I(R6913t2475) I(R6913t4775) I(R6913t5666) I(R6913t2656) I(R6914t1883) I(R6914t2872) I(R6914t2568) I(R6914t3254) I(R6914t750) I(R6915t4255) I(R6915t5279) I(R6915t6298) I(R6915t4713) I(R6915t1061) I(R6915t4719) I(R6916t686) I(R6916t6133) I(R6916t4979) I(R6917t6864) I(R6917t2638) I(R6917t1592) I(R6917t681) I(R6917t5) I(R6918t3449) I(R6918t4534) I(R6918t1949) I(R6918t3712) I(R6918t5829) I(R6919t238) I(R6919t1877) I(R6919t2804) I(R6919t5811) I(R6919t2452) I(R6920t1215) I(R6920t3571) I(R6920t5494) I(R6920t3289) I(R6920t5971) I(R6920t3074) I(R6920t1039) I(R6921t200) I(R6921t875) I(R6921t826) I(R6921t4894) I(R6922t923) I(R6922t5894) I(R6923t4287) I(R6923t6699) I(R6923t1325) I(R6923t2511) I(R6924t5914) I(R6924t3971) I(R6925t1358) I(R6925t5978) I(R6926t2825) I(R6926t5203) I(R6926t2531) I(R6926t130) I(R6926t726) I(R6927t474) I(R6927t1964) I(R6927t6422) I(R6927t4289) I(R6927t4845) I(R6928t1292) I(R6928t4556) I(R6928t3099) I(R6928t4695) I(R6929t866) I(R6929t1426) I(R6929t2191) I(R6930t974) I(R6930t576) I(R6930t5693) I(R6930t3449) I(R6930t5829) I(R6931t6822) I(R6931t6867) I(R6931t2069) I(R6931t4171) I(R6932t5010) I(R6932t5696) I(R6932t2430) I(R6933t2498) I(R6933t6077) I(R6933t4607) I(R6933t5574) I(R6933t3085) I(R6934t3405) I(R6934t5359) I(R6935t344) I(R6935t4167) I(R6935t756) I(R6935t3681) I(R6935t1110) I(R6936t2750) I(R6936t6338) I(R6936t2082) I(R6936t642) I(R6936t1499) I(R6936t63) I(R6936t5651) I(R6937t4653) I(R6937t241) I(R6937t2397) I(R6937t681) I(R6937t5198) I(R6938t5424) I(R6938t3387) I(R6938t4466) I(R6938t4871) I(R6938t5026) I(R6939t1811) I(R6939t3956) I(R6939t1443) I(R6939t1409) I(R6940t4) I(R6940t970) I(R6940t4285) I(R6940t1805) I(R6940t5923) I(R6941t5314) I(R6941t6162) I(R6941t3671) I(R6941t945) I(R6941t2059) I(R6942t395) I(R6942t4628) I(R6942t137) I(R6942t4910) I(R6942t2379) I(R6943t2929) I(R6943t894) I(R6943t3612) I(R6943t5320) I(R6943t65) I(R6944t2463) I(R6944t4657) I(R6944t1273) I(R6944t5209) I(R6944t301) I(R6945t4149) I(R6945t5372) I(R6945t4150) I(R6945t6600) I(R6945t676) I(R6946t468) I(R6946t507) I(R6946t3540) I(R6946t433) I(R6946t2628) I(R6946t3479) I(R6947t4300) I(R6948t5378) I(R6948t6037) I(R6948t3287) I(R6948t2651) I(R6949t400) I(R6949t887) I(R6949t1394) I(R6949t4973) I(R6950t1290) I(R6950t6776) I(R6950t192) I(R6950t1706) I(R6951t28) I(R6951t3562) I(R6951t118) I(R6951t839) I(R6951t266) I(R6952t5863) I(R6952t4061) I(R6952t1262) I(R6953t6415) I(R6953t2120) I(R6953t5891) I(R6954t4519) I(R6954t6888) I(R6954t5007) I(R6954t3422) I(R6954t3415) I(R6955t1223) I(R6955t719) I(R6955t2576) I(R6955t6049) I(R6955t1053) I(R6956t2390) I(R6956t2299) I(R6956t4901) I(R6956t3047) I(R6957t5655) I(R6957t3154) I(R6958t1287) I(R6958t4841) I(R6958t1355) I(R6958t2116) I(R6959t2107) I(R6959t2319) I(R6959t5604) I(R6959t6343) I(R6959t1356) I(R6959t3645) I(R6959t6759) I(R6960t1929) I(R6960t2191) I(R6960t1687) I(R6960t3641) I(R6960t3959) I(R6960t5363) I(R6960t1979) I(R6961t565) I(R6961t3570) I(R6961t3139) I(R6962t2317) I(R6962t6794) I(R6962t616) I(R6962t5797) I(R6963t1099) I(R6963t5509) I(R6963t29) I(R6963t3443) I(R6963t3166) I(R6963t6354) I(R6964t4026) I(R6964t4062) I(R6964t5775) I(R6964t5864) I(R6965t4259) I(R6965t1614) I(R6965t2763) I(R6965t552) I(R6967t2341) I(R6967t2883) I(R6967t4931) I(R6968t1015) I(R6968t4644) I(R6968t1761) I(R6968t3987) I(R6968t5084) I(R6969t171) I(R6969t4509) I(R6969t5955) I(R6969t6590) I(R6969t2288) I(R6970t2321) I(R6970t4942) I(R6970t2805) I(R6970t3445) I(R6970t3178) I(R6970t5556) I(R6970t2444) I(R6971t2060) I(R6971t6306) I(R6971t997) I(R6971t5228) I(R6972t517) I(R6972t1497) I(R6972t261) I(R6972t3734) I(R6972t4443) I(R6972t5432) I(R6972t3981) I(R6973t590) I(R6973t6159) I(R6973t6506) I(R6973t1800) I(R6973t5071) I(R6973t4661) I(R6974t1177) I(R6974t4540) I(R6974t6022) I(R6974t4392) I(R6975t2278) I(R6975t5388) I(R6975t269) I(R6975t3567) I(R6975t4380) I(R6975t229) I(R6975t6093) I(R6976t2451) I(R6976t3306) I(R6976t154) I(R6976t1679) I(R6976t1721) I(R6976t5072) I(R6977t3221) I(R6977t1128) I(R6977t1469) I(R6978t2626) I(R6978t6201) I(R6978t4532) I(R6978t2561) I(R6978t6705) I(R6978t694) I(R6978t6179) I(R6979t6948) I(R6979t492) I(R6979t314) I(R6979t2986) I(R6980t3003) I(R6980t3315) I(R6980t5047) I(R6981t2248) I(R6981t6106) I(R6982t2823) I(R6982t2213) I(R6982t5384) I(R6982t5588) I(R6983t4099) I(R6983t5047) I(R6983t3315) I(R6984t4301) I(R6984t6687) I(R6984t6154) I(R6984t4045) I(R6985t6947) I(R6985t6221) I(R6985t6904) I(R6986t5936) I(R6986t6658) I(R6986t1557) I(R6986t937) I(R6987t502) I(R6987t4700) I(R6987t1423) I(R6987t6625) I(R6987t4181) I(R6988t3460) I(R6988t4824) I(R6988t2068) I(R6989t509) I(R6989t2384) I(R6989t4304) I(R6989t775) I(R6990t906) I(R6990t5912) I(R6990t2225) I(R6990t5714) I(R6991t10) I(R6991t5250) I(R6991t5065) I(R6991t4928) I(R6991t1057) I(R6992t2241) I(R6992t3677) I(R6992t1329) I(R6992t5050) I(R6992t1387) I(R6993t3892) I(R6993t43) I(R6994t6229) I(R6994t6454) I(R6994t3227) I(R6995t1679) I(R6995t5805) I(R6995t1619) I(R6995t6031) I(R6995t3416) I(R6996t4146) I(R6996t143) I(R6997t2669) I(R6997t5893) I(R6997t3746) I(R6997t5686) I(R6997t2842) I(R6997t5947) I(R6997t2698) I(R6998t3207) I(R6999t891) I(R6999t3429) I(R6999t4842) I(R6999t5755) I(R6999t2435) I(R7000t253) I(R7000t2559) I(R7000t3743) I(R7000t2134) I(R7000t2536) I(R7001t2848) I(R7001t6552) I(R7001t5032) I(R7001t1568) I(R7002t4567) I(R7002t4780) I(R7002t5578) I(R7002t4997) I(R7002t6977) I(R7003t3380) I(R7003t4071) I(R7004t4762) I(R7004t5485) I(R7004t2110) I(R7004t6828) I(R7004t4267) I(R7005t870) I(R7005t3654) I(R7005t3327) I(R7006t1871) I(R7006t1309) I(R7006t2264) I(R7006t600) I(R7006t6144) I(R7007t142) I(R7007t3690) I(R7007t2822) I(R7008t5819) I(R7009t4731) I(R7009t4816) I(R7009t52) I(R7009t6684) I(R7010t5550) I(R7010t3486) I(R7010t4261) I(R7010t3961) I(R7010t5904) I(R7010t6587) I(R7010t1121) I(R7011t364) I(R7011t4549) I(R7011t6745) I(R7011t6880) I(R7012t3588) I(R7012t2367) I(R7012t5533) I(R7012t676) I(R7012t2965) I(R7012t5826) I(R7013t2324) I(R7013t862) I(R7013t3198) I(R7013t3125) I(R7014t1825) I(R7014t4318) I(R7014t362) I(R7014t1680) I(R7014t4701) I(R7014t4770) I(R7015t854) I(R7015t4179) I(R7015t2691) I(R7015t4245) I(R7015t4606) I(R7015t2543) I(R7016t6229) I(R7016t330) I(R7016t4489) I(R7016t4114) I(R7017t1105) I(R7017t2556) I(R7017t6069) I(R7017t3470) I(R7018t93) I(R7018t2147) I(R7018t3462) I(R7018t6796) I(R7018t6717) I(R7018t25) I(R7019t39) I(R7019t1748) I(R7019t1464) I(R7019t701) I(R7019t6329) I(R7019t1454) I(R7020t4208) I(R7020t5937) I(R7020t4493) I(R7020t3472) I(R7020t3454) I(R7021t411) I(R7021t862) I(R7021t6236) I(R7021t6838) I(R7021t2181) I(R7022t2411) I(R7022t6576) I(R7022t814) I(R7023t5144) I(R7023t5634) I(R7023t178) I(R7023t4247) I(R7023t6341) I(R7024t4685) I(R7024t367) I(R7025t4268) I(R7026t1390) I(R7026t2418) I(R7026t102) I(R7026t2489) I(R7026t4722) I(R7027t4898) I(R7027t1818) I(R7028t403) I(R7028t4663) I(R7028t3274) I(R7029t3956) I(R7029t4781) I(R7029t1719) I(R7029t2620) I(R7029t6674) I(R7030t285) I(R7030t5218) I(R7030t5763) I(R7030t2132) I(R7031t5205) I(R7031t5227) I(R7031t5748) I(R7032t3395) I(R7032t4441) I(R7032t4106) I(R7032t851) I(R7033t6084) I(R7033t4088) I(R7033t522) I(R7033t2276) I(R7033t4081) I(R7033t5029) I(R7034t72) I(R7034t4995) I(R7034t3179) I(R7034t6575) I(R7035t2823) I(R7035t3883) I(R7035t6982) I(R7036t1693) I(R7036t5185) I(R7036t2226) I(R7036t6406) I(R7037t2065) I(R7037t2224) I(R7037t5517) I(R7037t4563) I(R7037t4199) I(R7038t4033) I(R7038t6394) I(R7038t270) I(R7038t377) I(R7039t6429) I(R7039t4146) I(R7039t6996) I(R7039t143) I(R7039t5870) I(R7040t128) I(R7040t4324) I(R7041t3320) I(R7041t5082) I(R7041t6689) I(R7041t5306) I(R7041t2081) I(R7042t4339) I(R7042t424) I(R7042t6860) I(R7042t2216) I(R7042t6328) I(R7042t2512) I(R7043t3795) I(R7043t3702) I(R7043t268) I(R7043t3330) I(R7043t3143) I(R7043t2017) I(R7043t6049) I(R7044t2448) I(R7044t77) I(R7044t1689) I(R7045t478) I(R7045t1223) I(R7045t6955) I(R7045t1053) I(R7046t3054) I(R7046t3710) I(R7046t5835) I(R7047t1770) I(R7047t6640) I(R7047t3868) I(R7047t4313) I(R7048t4587) I(R7048t1310) I(R7048t4302) I(R7048t5278) I(R7048t3387) I(R7049t280) I(R7049t2243) I(R7049t6585) I(R7049t5484) I(R7049t3367) I(R7049t2094) I(R7050t5870) I(R7051t6473) I(R7051t6426) I(R7051t1554) I(R7051t3430) I(R7052t3557) I(R7052t3606) I(R7052t3009) I(R7052t4416) I(R7052t110) I(R7052t4860) I(R7053t3522) I(R7053t5298) I(R7053t6592) I(R7053t6713) I(R7053t5348) I(R7053t1563) I(R7054t1596) I(R7054t6905) I(R7054t419) I(R7055t5576) I(R7055t6730) I(R7055t754) I(R7055t3178) I(R7056t872) I(R7056t6605) I(R7056t1350) I(R7056t951) I(R7057t5151) I(R7057t5565) I(R7057t3338) I(R7057t2035) I(R7058t5475) I(R7058t662) I(R7058t6059) I(R7058t3800) I(R7059t864) I(R7059t481) I(R7059t4912) I(R7059t4342) I(R7060t2646) I(R7060t4650) I(R7060t5645) I(R7060t497) I(R7060t5398) I(R7060t4906) I(R7061t1538) I(R7061t6790) I(R7061t3561) I(R7061t2421) I(R7062t1360) I(R7062t5059) I(R7062t1616) I(R7062t5103) I(R7063t1368) I(R7063t3353) I(R7064t4819) I(R7064t6599) I(R7064t3136) I(R7064t3692) I(R7064t1981) I(R7065t2535) I(R7065t2557) I(R7065t6064) I(R7065t364) I(R7066t3562) I(R7066t118) I(R7067t435) I(R7067t1557) I(R7067t6986) I(R7067t937) I(R7067t604) I(R7067t6323) I(R7067t147) I(R7068t2162) I(R7068t5043) I(R7068t2088) I(R7068t3967) I(R7069t2710) I(R7069t5178) I(R7069t1822) I(R7069t2485) I(R7069t2773) I(R7069t1520) I(R7069t2184) I(R7069t6760) I(R7069t3603) I(R7069t654) I(R7070t4573) I(R7070t4685) I(R7070t991) I(R7070t6111) I(R7070t7024) I(R7071t1241) I(R7071t6694) I(R7071t5664) I(R7071t557) I(R7072t6444) I(R7072t2373) I(R7072t5306) I(R7072t263) I(R7072t1901) I(R7073t6279) I(R7073t6788) I(R7073t3328) I(R7073t4973) I(R7074t6234) I(R7075t5959) I(R7075t6546) I(R7075t5680) I(R7075t84) I(R7076t2259) I(R7076t2810) I(R7076t6675) I(R7076t953) I(R7077t5285) I(R7078t1531) I(R7078t1609) I(R7078t171) I(R7078t2288) I(R7079t233) I(R7079t2155) I(R7079t6792) I(R7079t4111) I(R7080t187) I(R7080t5329) I(R7080t4924) I(R7080t4266) I(R7081t2876) I(R7081t6751) I(R7081t5238) I(R7081t6682) I(R7082t705) I(R7082t1226) I(R7082t2229) I(R7082t1864) I(R7082t6452) I(R7082t149) I(R7083t5945) I(R7083t875) I(R7083t6773) I(R7083t2353) I(R7084t4540) I(R7084t6974) I(R7084t4548) I(R7084t5811) I(R7084t4984) I(R7084t1177) I(R7085t5661) I(R7085t2124) I(R7085t1487) I(R7085t5193) I(R7086t3071) I(R7086t5670) I(R7086t3581) I(R7086t4144) I(R7086t5525) I(R7086t4952) I(R7086t2644) I(R7087t249) I(R7087t1751) I(R7087t6396) I(R7087t1298) I(R7088t569) I(R7088t3585) I(R7088t3459) I(R7089t2051) I(R7089t4294) I(R7089t5370) I(R7089t2595) I(R7089t3890) I(R7090t2494) I(R7090t4893) I(R7090t4887) I(R7090t6069) I(R7091t2242) I(R7091t3774) I(R7091t3163) I(R7091t2347) I(R7092t3157) I(R7092t4347) I(R7093t6350) I(R7093t1423) I(R7093t3121) I(R7094t383) I(R7094t4130) I(R7094t2460) I(R7094t1474) I(R7094t6276) I(R7095t3505) I(R7095t6902) I(R7096t2987) I(R7096t1255) I(R7097t1675) I(R7097t4945) I(R7097t4715) I(R7097t5627) I(R7097t6542) I(R7098t4358) I(R7098t2185) I(R7098t2187) I(R7098t2474) I(R7099t2049) I(R7099t6990) I(R7099t5714) I(R7099t3197) I(R7100t763) I(R7100t1446) I(R7100t6497) I(R7100t586) I(R7100t1590) I(R7100t6466) I(R7101t331) I(R7101t657) I(R7101t2076) I(R7101t6294) I(R7102t3530) I(R7102t3945) I(R7102t4630) I(R7103t6099) I(R7103t6904) I(R7103t5919) I(R7103t932) I(R7104t178) I(R7104t5132) I(R7104t1811) I(R7104t6939) I(R7104t1409) I(R7104t5641) I(R7104t6181) I(R7104t1320) I(R7105t848) I(R7105t2287) I(R7105t3454) I(R7105t3472) I(R7106t2008) I(R7106t5994) I(R7106t5631) I(R7106t6865) I(R7106t3982) I(R7106t5744) I(R7107t1228) I(R7107t5391) I(R7107t2090) I(R7107t4747) I(R7108t1190) I(R7108t3420) I(R7108t5657) I(R7108t5862) I(R7108t906) I(R7108t6990) I(R7109t51) I(R7109t367) I(R7109t2003) I(R7109t5935) I(R7109t2001) I(R7109t4825) I(R7110t1042) I(R7110t2537) I(R7110t6142) I(R7111t2417) I(R7111t5149) I(R7111t3983) I(R7112t1576) I(R7112t5802) I(R7112t5072) I(R7112t6032) I(R7112t2609) I(R7113t4639) I(R7113t6603) I(R7113t4515) I(R7113t1812) I(R7114t5087) I(R7114t2585) I(R7114t6114) I(R7115t5311) I(R7115t3195) I(R7115t3953) I(R7115t3652) I(R7116t5323) I(R7116t6210) I(R7116t4964) I(R7116t4323) I(R7117t1396) I(R7117t5580) I(R7117t796) I(R7117t1642) I(R7117t328) I(R7117t5760) I(R7118t322) I(R7118t1691) I(R7118t2523) I(R7118t199) I(R7118t373) I(R7119t646) I(R7119t6352) I(R7119t1251) I(R7119t3939) I(R7120t2540) I(R7120t5742) I(R7120t6408) I(R7120t6432) I(R7121t1182) I(R7121t4553) I(R7121t2073) I(R7121t1886) I(R7122t3450) I(R7122t4858) I(R7122t5047) I(R7122t6980) I(R7122t2516) I(R7123t5957) I(R7123t1333) I(R7124t1362) I(R7124t2794) I(R7124t5446) I(R7124t2636) I(R7124t1269) I(R7125t2340) I(R7125t5583) I(R7125t2904) I(R7125t341) I(R7126t5978) I(R7126t6925) I(R7126t4822) I(R7127t2076) I(R7127t7101) I(R7127t3033) I(R7127t1233) I(R7127t6294) I(R7128t1679) I(R7128t1721) I(R7128t2942) I(R7128t5303) I(R7129t5237) I(R7129t6709) I(R7129t2723) I(R7129t1257) I(R7130t820) I(R7130t1006) I(R7130t2791) I(R7130t6652) I(R7130t5335) I(R7131t6895) I(R7131t2790) I(R7131t2831) I(R7132t889) I(R7132t975) I(R7132t56) I(R7132t3226) I(R7132t6422) I(R7133t1512) I(R7133t3733) I(R7133t3261) I(R7133t1860) I(R7133t6810) I(R7134t2852) I(R7134t419) I(R7135t6299) I(R7135t4610) I(R7135t2076) I(R7135t797) I(R7136t5880) I(R7136t3261) I(R7137t3422) I(R7137t6954) I(R7137t3415) I(R7138t3476) I(R7138t2734) I(R7138t323) I(R7138t3342) I(R7139t1705) I(R7139t4476) I(R7139t2039) I(R7139t6518) I(R7140t2340) I(R7140t7125) I(R7140t1323) I(R7140t6856) I(R7140t2904) I(R7141t1246) I(R7141t3752) I(R7141t847) I(R7141t4998) I(R7142t4406) I(R7142t6661) I(R7142t1289) I(R7142t2230) I(R7142t3775) I(R7143t3534) I(R7143t5110) I(R7143t5695) I(R7143t2360) I(R7143t6215) I(R7143t2546) I(R7144t921) I(R7144t1173) I(R7144t2343) I(R7144t5934) I(R7144t1046) I(R7144t408) I(R7144t3364) I(R7145t2770) I(R7145t1786) I(R7145t5838) I(R7145t1156) I(R7145t5329) I(R7145t5903) I(R7145t1387) I(R7146t4904) I(R7146t672) I(R7146t3160) I(R7147t46) I(R7147t6645) I(R7147t6284) I(R7147t5195) I(R7147t691) I(R7147t5917) I(R7148t6838) I(R7148t2181) I(R7148t566) I(R7148t520) I(R7149t2165) I(R7149t5749) I(R7149t3761) I(R7149t3046) I(R7150t2405) I(R7150t3131) I(R7150t1302) I(R7150t2745) I(R7150t4779) I(R7150t6104) I(R7150t5990) I(R7151t855) I(R7151t3214) I(R7151t1412) I(R7151t960) I(R7152t4277) I(R7152t4754) I(R7152t5879) I(R7152t1063) I(R7153t1633) I(R7153t4371) I(R7153t6250) I(R7153t3146) I(R7154t2007) I(R7154t4410) I(R7154t3458) I(R7154t5527) I(R7155t2492) I(R7155t6838) I(R7155t7148) I(R7156t3624) I(R7156t4304) I(R7156t6989) I(R7156t775) I(R7157t534) I(R7157t4999) I(R7157t2183) I(R7157t1370) I(R7158t4242) I(R7158t1043) I(R7158t5528) I(R7158t4328) I(R7159t5200) I(R7159t4729) I(R7159t4040) I(R7159t5745) I(R7159t6677) I(R7159t311) I(R7160t4286) I(R7160t3957) I(R7161t4442) I(R7161t5931) I(R7161t1444) I(R7161t653) I(R7162t1410) I(R7162t6170) I(R7162t5302) I(R7162t2410) I(R7163t2960) I(R7163t161) I(R7164t1178) I(R7164t4195) I(R7164t4271) I(R7164t6311) I(R7164t5319) I(R7164t438) I(R7165t6610) I(R7165t968) I(R7165t608) I(R7165t5857) I(R7165t182) I(R7166t5643) I(R7166t323) I(R7166t5800) I(R7167t4776) I(R7167t1757) I(R7167t2043) I(R7167t3702) I(R7168t4975) I(R7169t6433) I(R7169t3180) I(R7169t2520) I(R7169t6125) I(R7169t5562) I(R7170t1398) I(R7170t4516) I(R7170t4225) I(R7171t1480) I(R7171t2929) I(R7171t6943) I(R7172t4099) I(R7172t6983) I(R7172t307) I(R7173t2960) I(R7173t7163) I(R7173t3792) I(R7173t6491) I(R7174t1502) I(R7174t2261) I(R7174t3940) I(R7174t2345) I(R7174t78) I(R7174t4398) I(R7175t863) I(R7175t3307) I(R7175t487) I(R7175t1717) I(R7176t1275) I(R7176t5570) I(R7176t3366) I(R7177t3797) I(R7177t4298) I(R7177t6478) I(R7178t581) I(R7178t619) I(R7178t2056) I(R7178t5763) I(R7178t7030) I(R7178t2132) I(R7178t1382) I(R7179t1191) I(R7179t3350) I(R7179t3996) I(R7179t5198) I(R7179t6937) I(R7179t681) I(R7179t1640) I(R7180t2787) I(R7180t3138) I(R7180t6865) I(R7180t3749) I(R7181t4146) I(R7181t6996) I(R7181t143) I(R7181t6723) I(R7182t4897) I(R7182t5257) I(R7182t5426) I(R7182t1781) I(R7183t3024) I(R7183t6778) I(R7183t6282) I(R7183t2514) I(R7184t669) I(R7184t2105) I(R7184t1141) I(R7185t454) I(R7185t658) I(R7185t3424) I(R7185t4674) I(R7185t35) I(R7185t445) I(R7185t133) I(R7186t20) I(R7186t2737) I(R7186t1807) I(R7186t6555) I(R7186t306) I(R7187t6305) I(R7187t2415) I(R7187t4195) I(R7187t4271) I(R7188t6928) I(R7188t4751) I(R7188t841) I(R7188t2391) I(R7188t1978) I(R7188t3099) I(R7189t269) I(R7189t6975) I(R7189t3119) I(R7190t1891) I(R7190t6559) I(R7190t3270) I(R7190t1624) I(R7190t5881) I(R7190t3583) I(R7191t4822) I(R7191t7126) I(R7191t5978) I(R7191t2837) I(R7191t3422) I(R7191t5239) I(R7191t2816) I(R7191t5950) I(R7192t4724) I(R7192t5995) I(R7193t4239) I(R7193t5828) I(R7193t835) I(R7193t3045) I(R7194t312) I(R7194t1578) I(R7194t244) I(R7194t6650) I(R7194t467) I(R7195t5332) I(R7195t5665) I(R7195t5847) I(R7195t1221) I(R7195t3496) I(R7195t6108) I(R7196t3723) I(R7196t4589) I(R7196t3962) I(R7197t2442) I(R7197t3697) I(R7197t5243) I(R7197t2980) I(R7197t1500) I(R7198t1171) I(R7198t6082) I(R7198t884) I(R7198t193) I(R7198t5344) I(R7199t1325) I(R7199t6923) I(R7199t4287) I(R7199t2949) I(R7199t6247) I(R7199t5337) I(R7200t3188) I(R7200t6409) I(R7200t5360) I(R7200t6785) I(R7200t2121) I(R7201t604) I(R7201t3547) I(R7202t188) I(R7202t4906) I(R7202t6692) I(R7202t5398) I(R7202t7060) I(R7203t1161) I(R7203t1728) I(R7203t4982) I(R7204t4921) I(R7204t2154) I(R7204t3812) I(R7205t3101) I(R7205t1030) I(R7206t3221) I(R7206t6977) I(R7206t5500) I(R7206t4997) I(R7206t7002) I(R7207t4741) I(R7207t2899) I(R7207t5832) I(R7207t1433) I(R7208t982) I(R7208t1568) I(R7208t7001) I(R7208t2848) I(R7208t1823) I(R7208t4353) I(R7209t5313) I(R7209t2352) I(R7209t5448) I(R7209t893) I(R7210t391) I(R7210t2355) I(R7210t6358) I(R7210t2125) I(R7210t3871) I(R7211t5812) I(R7211t7074) I(R7211t6234) I(R7211t6612) I(R7211t5431) I(R7211t1803) I(R7212t2336) I(R7212t3309) I(R7212t5185) I(R7212t2226) I(R7212t1808) I(R7212t6627) I(R7213t6229) I(R7213t7016) I(R7213t330) I(R7213t3718) I(R7213t4572) I(R7213t30) I(R7213t6454) I(R7213t6994) I(R7214t769) I(R7214t2932) I(R7214t1764) I(R7215t5756) I(R7215t134) I(R7215t7156) I(R7216t446) I(R7216t6849) I(R7216t988) I(R7216t472) I(R7217t2684) I(R7217t3978) I(R7217t5373) I(R7217t5447) I(R7218t4117) I(R7218t4279) I(R7218t5280) I(R7218t1561) I(R7219t3403) I(R7219t4216) I(R7219t6890) I(R7219t3547) I(R7219t7201) I(R7220t3563) I(R7220t4878) I(R7220t5404) I(R7220t4253) I(R7220t3032) I(R7220t5186) I(R7220t4408) I(R7220t2742) I(R7220t1904) I(R7221t3402) I(R7221t6019) I(R7221t1133) I(R7221t3881) I(R7221t406) I(R7222t1708) I(R7222t3455) I(R7222t1827) I(R7222t4034) I(R7223t1339) I(R7223t3534) I(R7223t818) I(R7223t5156) I(R7223t625) I(R7223t27) I(R7224t2843) I(R7224t5080) I(R7224t2435) I(R7224t891) I(R7225t4877) I(R7225t207) I(R7225t1481) I(R7225t1033) I(R7226t1155) I(R7226t1064) I(R7226t4537) I(R7226t4789) I(R7227t2240) I(R7227t5430) I(R7227t694) I(R7227t525) I(R7227t2685) I(R7228t542) I(R7228t1081) I(R7228t3918) I(R7228t6852) I(R7229t1461) I(R7229t5008) I(R7229t713) I(R7229t2202) I(R7229t651) I(R7230t5743) I(R7230t5976) I(R7230t536) I(R7230t3457) I(R7230t2951) I(R7230t58) I(R7230t6669) I(R7231t322) I(R7231t5486) I(R7231t7118) I(R7231t2523) I(R7231t4138) I(R7231t6177) I(R7232t2789) I(R7232t5678) I(R7232t4002) I(R7232t6873) I(R7232t2254) I(R7232t5682) I(R7233t7114) I(R7233t5087) I(R7233t965) I(R7233t3962) I(R7233t7196) I(R7233t3723) I(R7234t2295) I(R7234t4574) I(R7234t2374) I(R7234t5579) I(R7234t1479) I(R7235t2971) I(R7235t4930) I(R7235t6823) I(R7235t1104) I(R7235t1389) I(R7236t5830) I(R7236t1103) I(R7236t6891) I(R7237t504) I(R7237t2202) I(R7237t1926) I(R7237t1867) I(R7238t2765) I(R7238t1375) I(R7238t5939) I(R7239t4384) I(R7239t5642) I(R7239t6007) I(R7239t4786) I(R7239t4855) I(R7240t1726) I(R7240t6289) I(R7240t7080) I(R7240t187) I(R7241t6352) I(R7241t6440) I(R7241t646) I(R7241t6223) I(R7241t1963) I(R7241t6879) I(R7242t6766) I(R7242t2225) I(R7242t5912) I(R7242t569) I(R7242t7088) I(R7242t3459) I(R7242t5873) I(R7242t2518) I(R7243t638) I(R7243t1948) I(R7243t2134) I(R7243t7000) I(R7243t2536) I(R7243t2717) I(R7243t3458) I(R7243t7154) I(R7243t5356) I(R7244t1971) I(R7244t2856) I(R7244t5301) I(R7245t1536) I(R7245t4604) I(R7245t5842) I(R7245t802) I(R7246t1045) I(R7246t3066) I(R7246t2799) I(R7247t1951) I(R7247t5354) I(R7247t218) I(R7247t3229) I(R7248t4875) I(R7248t5663) I(R7248t4457) I(R7248t1704) I(R7248t5655) I(R7248t3821) I(R7248t3075) I(R7249t3261) I(R7249t7136) I(R7249t6357) I(R7250t3941) I(R7250t3173) I(R7250t4545) I(R7250t252) I(R7250t1921) I(R7251t1691) I(R7251t6102) I(R7251t3029) I(R7251t373) I(R7252t806) I(R7252t4774) I(R7252t4449) I(R7252t4355) I(R7253t1566) I(R7253t3392) I(R7253t3605) I(R7253t5989) I(R7253t1686) I(R7254t2261) I(R7254t3940) I(R7254t3344) I(R7254t1875) I(R7255t441) I(R7255t909) I(R7255t6455) I(R7255t5003) I(R7255t4915) I(R7255t465) I(R7255t868) I(R7256t338) I(R7256t1862) I(R7256t4756) I(R7256t3544) I(R7256t1263) I(R7257t2664) I(R7257t1763) I(R7257t2471) I(R7257t260) I(R7257t3642) I(R7258t6186) I(R7258t6909) I(R7258t1475) I(R7258t73) I(R7258t5814) I(R7258t2041) I(R7259t4162) I(R7259t3442) I(R7259t4801) I(R7259t678) I(R7260t1422) I(R7260t6566) I(R7260t4482) I(R7260t6651) I(R7261t1057) I(R7261t5088) I(R7261t4928) I(R7261t3241) I(R7261t6183) I(R7262t3667) I(R7262t4553) I(R7262t4868) I(R7262t5348) I(R7262t7053) I(R7262t6713) I(R7262t1408) I(R7263t4492) I(R7263t5625) I(R7264t2310) I(R7264t6912) I(R7264t4372) I(R7264t3056) I(R7264t725) I(R7265t2972) I(R7265t5678) I(R7265t2475) I(R7265t6913) I(R7265t2656) I(R7265t2873) I(R7265t127) I(R7265t3466) I(R7265t3855) I(R7266t1095) I(R7266t5478) I(R7266t6130) I(R7266t6193) I(R7266t131) I(R7266t4486) I(R7267t3234) I(R7267t2835) I(R7267t5875) I(R7267t5700) I(R7267t6841) I(R7268t1523) I(R7268t5610) I(R7268t1916) I(R7268t3523) I(R7269t19) I(R7269t4847) I(R7269t2005) I(R7269t5444) I(R7270t4446) I(R7270t6344) I(R7270t6710) I(R7270t6155) I(R7270t3241) I(R7270t5217) I(R7270t2055) I(R7271t1073) I(R7271t7054) I(R7271t419) I(R7271t6708) I(R7272t2165) I(R7272t5749) I(R7272t5630) I(R7272t4370) I(R7272t1833) I(R7272t782) I(R7272t5542) I(R7273t281) I(R7273t477) I(R7273t351) I(R7274t1334) I(R7274t2544) I(R7274t2894) I(R7274t5064) I(R7274t3870) I(R7274t36) I(R7274t755) I(R7275t1010) I(R7275t1949) I(R7276t1463) I(R7276t3409) I(R7276t5938) I(R7276t6475) I(R7276t3680) I(R7277t2886) I(R7277t3675) I(R7277t4986) I(R7278t2143) I(R7278t6580) I(R7278t3851) I(R7279t4082) I(R7279t5492) I(R7279t4774) I(R7279t433) I(R7279t2628) I(R7280t5427) I(R7280t5945) I(R7280t6275) I(R7280t1605) I(R7281t180) I(R7281t6336) I(R7281t6126) I(R7281t1457) I(R7281t4395) I(R7281t2883) I(R7281t6967) I(R7281t2341) I(R7282t3007) I(R7282t3686) I(R7282t3063) I(R7283t1121) I(R7283t6816) I(R7283t5369) I(R7283t2250) I(R7284t5151) I(R7284t5565) I(R7284t3338) I(R7284t1880) I(R7284t3919) I(R7284t3514) I(R7284t3464) I(R7285t2718) I(R7285t3765) I(R7285t6859) I(R7285t3532) I(R7285t556) I(R7286t6800) I(R7286t2010) I(R7286t5448) I(R7286t7209) I(R7286t2352) I(R7286t563) I(R7287t1639) I(R7287t483) I(R7287t4969) I(R7288t6591) I(R7288t2559) I(R7288t7000) I(R7288t253) I(R7288t2410) I(R7289t915) I(R7289t5307) I(R7289t5447) I(R7289t2684) I(R7289t917) I(R7290t996) I(R7290t4935) I(R7290t1312) I(R7291t1038) I(R7291t1876) I(R7291t4155) I(R7291t2545) I(R7291t2685) I(R7291t1903) I(R7292t5900) I(R7292t6504) I(R7292t1872) I(R7292t3245) I(R7293t5369) I(R7293t1364) I(R7293t1517) I(R7293t4612) I(R7293t3657) I(R7294t909) I(R7294t6455) I(R7294t1127) I(R7294t1766) I(R7294t5752) I(R7295t4418) I(R7295t6498) I(R7295t2772) I(R7295t6333) I(R7295t3052) I(R7296t3909) I(R7296t5265) I(R7296t2369) I(R7296t5809) I(R7297t5966) I(R7297t6874) I(R7297t4230) I(R7297t1319) I(R7297t5501) I(R7297t4087) I(R7298t728) I(R7298t3578) I(R7298t1961) I(R7299t207) I(R7299t1598) I(R7299t2427) I(R7299t9) I(R7299t1991) I(R7300t6244) I(R7300t381) I(R7300t4968) I(R7300t3310) I(R7301t2795) I(R7301t4251) I(R7301t5902) I(R7301t2221) I(R7301t5068) I(R7301t5975) I(R7302t4452) I(R7302t5997) I(R7302t2838) I(R7303t3969) I(R7303t6448) I(R7303t5260) I(R7303t933) I(R7303t1442) I(R7303t2272) I(R7303t3599) I(R7304t5082) I(R7304t1967) I(R7304t2081) I(R7305t3699) I(R7305t4773) I(R7305t550) I(R7306t6182) I(R7306t1594) I(R7307t4586) I(R7307t2708) I(R7307t4913) I(R7307t5916) I(R7307t5437) I(R7308t4347) I(R7308t777) I(R7309t6783) I(R7309t7161) I(R7309t5122) I(R7310t5458) I(R7310t6408) I(R7310t7120) I(R7310t6432) I(R7310t2034) I(R7310t2843) I(R7311t3524) I(R7311t4814) I(R7311t7134) I(R7311t2852) I(R7311t3383) I(R7312t6910) I(R7312t3937) I(R7312t913) I(R7313t234) I(R7313t1153) I(R7313t1603) I(R7313t1758) I(R7314t985) I(R7314t6701) I(R7314t4621) I(R7314t3998) I(R7314t4410) I(R7315t4325) I(R7315t4877) I(R7315t3004) I(R7315t1977) I(R7315t1033) I(R7316t1852) I(R7316t5768) I(R7316t5044) I(R7316t18) I(R7317t3004) I(R7317t7315) I(R7317t1977) I(R7317t481) I(R7317t493) I(R7318t4366) I(R7318t831) I(R7318t4235) I(R7318t773) I(R7318t3985) I(R7319t1419) I(R7319t3689) I(R7319t770) I(R7319t2306) I(R7319t4034) I(R7320t7277) I(R7320t4986) I(R7320t903) I(R7320t4611) I(R7321t439) I(R7321t2009) I(R7321t810) I(R7322t3296) I(R7322t5718) I(R7322t1869) I(R7322t4602) I(R7323t7246) I(R7323t3485) I(R7324t1100) I(R7324t6230) I(R7324t2846) I(R7324t872) I(R7324t6605) I(R7324t914) I(R7325t189) I(R7325t2674) I(R7325t5196) I(R7325t1187) I(R7326t6673) I(R7326t602) I(R7326t1017) I(R7326t1152) I(R7327t2968) I(R7327t5130) I(R7327t532) I(R7328t327) I(R7328t1273) I(R7328t6944) I(R7328t4657) I(R7329t1434) I(R7329t4316) I(R7329t1113) I(R7329t3149) I(R7329t4391) I(R7330t97) I(R7330t381) I(R7330t5790) I(R7330t2266) I(R7331t6980) I(R7331t5321) I(R7331t1235) I(R7331t2778) I(R7331t1224) I(R7332t6355) I(R7332t6903) I(R7332t5313) I(R7332t3751) I(R7332t7028) I(R7332t403) I(R7333t180) I(R7333t1564) I(R7333t6336) I(R7333t7281) I(R7334t1824) I(R7334t5326) I(R7334t3367) I(R7335t3429) I(R7335t5196) I(R7335t2882) I(R7335t1623) I(R7336t2662) I(R7336t3001) I(R7336t6415) I(R7336t6953) I(R7337t4605) I(R7337t3250) I(R7337t2404) I(R7337t6291) I(R7338t1657) I(R7338t6733) I(R7338t1123) I(R7338t5781) I(R7338t6847) I(R7338t1943) I(R7338t2139) I(R7339t4017) I(R7339t6009) I(R7339t4726) I(R7339t6042) I(R7339t1406) I(R7340t7278) I(R7340t7311) I(R7340t4814) I(R7340t3612) I(R7340t6580) I(R7341t4086) I(R7341t1021) I(R7342t1114) I(R7342t3591) I(R7342t5546) I(R7343t2298) I(R7343t2926) I(R7343t5401) I(R7344t2970) I(R7344t837) I(R7344t3635) I(R7345t4126) I(R7345t1605) I(R7345t1894) I(R7345t5731) I(R7345t1431) I(R7346t675) I(R7346t1340) I(R7346t1164) I(R7346t6253) I(R7346t840) I(R7346t714) I(R7347t2013) I(R7347t2307) I(R7347t2849) I(R7347t1385) I(R7348t4248) I(R7348t5972) I(R7348t1166) I(R7349t4453) I(R7349t5574) I(R7349t2163) I(R7349t32) I(R7349t4916) I(R7350t3015) I(R7350t3243) I(R7350t422) I(R7350t5753) I(R7351t1835) I(R7351t3329) I(R7351t1087) I(R7351t2850) I(R7351t6445) I(R7351t2407) I(R7352t3357) I(R7352t6664) I(R7352t4024) I(R7352t5664) I(R7352t574) I(R7353t1853) I(R7353t5502) I(R7353t774) I(R7353t2798) I(R7353t1282) I(R7353t793) I(R7353t3602) I(R7354t1922) I(R7354t3912) I(R7354t1813) I(R7355t3335) I(R7355t3574) I(R7355t1684) I(R7355t5061) I(R7355t265) I(R7356t1254) I(R7356t5307) I(R7356t1024) I(R7356t3440) I(R7356t789) I(R7356t917) I(R7357t6556) I(R7357t1581) I(R7358t4504) I(R7358t4626) I(R7358t4771) I(R7358t4862) I(R7358t4969) I(R7358t7287) I(R7359t1491) I(R7359t4623) I(R7359t1345) I(R7359t5662) I(R7359t2648) I(R7360t593) I(R7360t4209) I(R7360t5099) I(R7360t329) I(R7360t5504) I(R7360t2720) I(R7361t3917) I(R7361t5393) I(R7361t5435) I(R7361t4795) I(R7362t2325) I(R7362t4800) I(R7362t5906) I(R7362t3180) I(R7362t3887) I(R7363t1956) I(R7363t3556) I(R7363t6680) I(R7363t1404) I(R7363t6171) I(R7364t2222) I(R7364t2864) I(R7364t1341) I(R7364t1868) I(R7364t366) I(R7364t869) I(R7365t1849) I(R7365t4912) I(R7365t1481) I(R7365t2151) I(R7366t5720) I(R7366t5869) I(R7366t1068) I(R7366t5513) I(R7366t3870) I(R7366t5673) I(R7367t2941) I(R7367t3917) I(R7367t4597) I(R7367t5951) I(R7367t5613) I(R7367t4480) I(R7368t6783) I(R7368t7309) I(R7368t2937) I(R7368t5931) I(R7368t7161) I(R7369t924) I(R7369t6705) I(R7369t2496) I(R7369t2561) I(R7369t6978) I(R7370t3886) I(R7370t4174) I(R7370t4274) I(R7370t2266) I(R7370t97) I(R7371t45) I(R7371t2888) I(R7371t767) I(R7371t4630) I(R7372t2319) I(R7372t5604) I(R7373t4024) I(R7373t4748) I(R7373t6729) I(R7373t5664) I(R7374t5214) I(R7374t4390) I(R7375t2327) I(R7375t5113) I(R7376t5268) I(R7376t4780) I(R7376t6827) I(R7376t92) I(R7377t1531) I(R7377t2715) I(R7377t151) I(R7377t6164) I(R7378t2330) I(R7378t5166) I(R7378t3217) I(R7378t6892) I(R7379t2370) I(R7379t540) I(R7379t3832) I(R7379t313) I(R7379t1832) I(R7380t5676) I(R7380t1622) I(R7381t1634) I(R7381t865) I(R7381t5981) I(R7381t6557) I(R7382t4707) I(R7382t6161) I(R7383t7323) I(R7383t2295) I(R7383t4574) I(R7383t43) I(R7384t3977) I(R7384t6374) I(R7384t4641) I(R7384t4501) I(R7384t538) I(R7385t1385) I(R7385t1866) I(R7385t4281) I(R7385t6264) I(R7386t6309) I(R7386t4689) I(R7386t3122) I(R7386t3035) I(R7386t6446) I(R7386t6095) I(R7387t716) I(R7387t994) I(R7387t2138) I(R7387t3905) I(R7388t6490) I(R7388t3722) I(R7388t3617) I(R7389t3204) I(R7389t4936) I(R7389t6303) I(R7389t771) I(R7389t3735) I(R7389t2067) I(R7390t2735) I(R7390t2719) I(R7390t4750) I(R7390t2089) I(R7390t4518) I(R7391t6744) I(R7391t3273) I(R7391t4799) I(R7391t5910) I(R7391t6349) I(R7392t1006) I(R7392t1985) I(R7392t139) I(R7392t5414) I(R7392t1747) I(R7392t5335) I(R7392t7130) I(R7393t3804) I(R7393t2933) I(R7393t6696) I(R7394t2076) I(R7394t2491) I(R7394t7135) I(R7394t797) I(R7394t1762) I(R7394t2667) I(R7394t181) I(R7395t99) I(R7395t2084) I(R7396t3551) I(R7396t5967) I(R7396t1234) I(R7396t4734) I(R7396t4234) I(R7396t6648) I(R7396t1922) I(R7396t7354) I(R7396t1813) I(R7397t7025) I(R7397t4268) I(R7397t5395) I(R7397t943) I(R7397t6380) I(R7398t4014) I(R7398t5112) I(R7398t4977) I(R7398t874) I(R7399t6133) I(R7399t1055) I(R7399t3360) I(R7399t4979) I(R7399t6916) I(R7400t5449) I(R7400t2896) I(R7400t3571) I(R7400t5794) I(R7401t3301) I(R7401t5451) I(R7401t660) I(R7401t3454) I(R7401t2287) I(R7402t1994) I(R7402t4884) I(R7402t1471) I(R7402t1770) I(R7402t6640) I(R7403t2228) I(R7403t7152) I(R7403t5879) I(R7404t2919) I(R7404t5019) I(R7404t5459) I(R7404t931) I(R7404t4315) I(R7404t561) I(R7405t6341) I(R7405t7023) I(R7405t5144) I(R7405t1604) I(R7405t1680) I(R7406t93) I(R7406t5242) I(R7406t3500) I(R7406t222) I(R7407t2) I(R7407t5954) I(R7407t6481) I(R7407t3086) I(R7408t4818) I(R7408t2616) I(R7408t2000) I(R7409t1951) I(R7409t6844) I(R7409t7247) I(R7409t5354) I(R7409t4229) I(R7410t3173) I(R7410t3941) I(R7411t2109) I(R7411t2162) I(R7411t5067) I(R7411t2160) I(R7411t3967) I(R7412t1380) I(R7412t2833) I(R7412t6568) I(R7412t5416) I(R7412t3882) I(R7413t6289) I(R7413t6884) I(R7413t3266) I(R7414t19) I(R7414t2199) I(R7414t1036) I(R7414t2313) I(R7415t5106) I(R7415t5470) I(R7415t5410) I(R7415t4723) I(R7415t232) I(R7415t6199) I(R7415t2713) I(R7416t301) I(R7416t6944) I(R7416t5209) I(R7416t2900) I(R7417t3088) I(R7417t3164) I(R7417t4057) I(R7417t1456) I(R7417t6152) I(R7417t1709) I(R7417t85) I(R7418t6486) I(R7418t3974) I(R7418t5051) I(R7418t1094) I(R7418t4550) I(R7419t3559) I(R7419t5998) I(R7419t1893) I(R7419t1209) I(R7419t4206) I(R7420t1984) I(R7420t2352) I(R7421t61) I(R7421t91) I(R7421t5960) I(R7421t6416) I(R7421t473) I(R7422t3145) I(R7422t5415) I(R7422t3128) I(R7422t1051) I(R7422t501) I(R7422t5801) I(R7423t2030) I(R7423t2299) I(R7423t6956) I(R7423t4980) I(R7424t944) I(R7424t2707) I(R7424t506) I(R7424t1880) I(R7424t3919) I(R7424t3514) I(R7425t1289) I(R7425t1681) I(R7425t7142) I(R7425t6661) I(R7425t2323) I(R7425t4702) I(R7426t3069) I(R7426t5202) I(R7426t3724) I(R7426t3799) I(R7427t2825) I(R7427t5992) I(R7427t4001) I(R7428t4) I(R7428t148) I(R7428t970) I(R7428t2237) I(R7428t3219) I(R7428t54) I(R7429t5794) I(R7429t5494) I(R7429t3289) I(R7429t4966) I(R7429t5228) I(R7429t997) I(R7429t6184) I(R7429t3426) I(R7430t1120) I(R7430t6829) I(R7430t6544) I(R7430t1776) I(R7431t6463) I(R7431t5548) I(R7431t859) I(R7432t3050) I(R7432t3272) I(R7432t2135) I(R7432t1009) I(R7433t3202) I(R7433t4045) I(R7433t4647) I(R7434t440) I(R7434t961) I(R7434t3985) I(R7434t773) I(R7434t53) I(R7434t2548) I(R7435t982) I(R7435t3953) I(R7436t3428) I(R7436t748) I(R7436t5385) I(R7436t3550) I(R7436t912) I(R7437t5615) I(R7437t6522) I(R7437t6222) I(R7437t1873) I(R7437t2936) I(R7438t6396) I(R7438t2171) I(R7438t1751) I(R7439t2718) I(R7439t556) I(R7439t3539) I(R7439t677) I(R7440t3278) I(R7440t7103) I(R7440t6904) I(R7440t6985) I(R7441t3751) I(R7441t7420) I(R7441t5313) I(R7442t3889) I(R7442t4599) I(R7442t4361) I(R7443t443) I(R7443t3978) I(R7443t4581) I(R7443t2329) I(R7443t3626) I(R7444t5808) I(R7444t1185) I(R7444t493) I(R7444t7317) I(R7444t481) I(R7445t87) I(R7445t6459) I(R7445t4295) I(R7445t156) I(R7445t5526) I(R7445t4007) I(R7446t4160) I(R7446t5780) I(R7446t6327) I(R7446t5907) I(R7446t498) I(R7446t4044) I(R7447t2490) I(R7447t2250) I(R7447t6157) I(R7447t447) I(R7447t5468) I(R7448t1345) I(R7448t5918) I(R7448t5654) I(R7448t1474) I(R7448t6912) I(R7448t725) I(R7449t3302) I(R7449t6267) I(R7449t6637) I(R7450t904) I(R7450t5273) I(R7450t2323) I(R7450t6164) I(R7451t4389) I(R7451t4392) I(R7451t6974) I(R7451t1177) I(R7451t3337) I(R7451t6087) I(R7451t463) I(R7451t1429) I(R7452t2188) I(R7452t3652) I(R7452t1305) I(R7453t4055) I(R7453t5779) I(R7453t6249) I(R7453t981) I(R7453t6263) I(R7453t1529) I(R7453t2381) I(R7454t4785) I(R7454t1947) I(R7455t7408) I(R7455t4818) I(R7455t3084) I(R7455t2381) I(R7455t1529) I(R7455t959) I(R7456t212) I(R7456t3052) I(R7456t4060) I(R7456t3259) I(R7457t200) I(R7457t6921) I(R7457t6773) I(R7457t3637) I(R7457t2895) I(R7457t3946) I(R7457t826) I(R7458t1620) I(R7459t87) I(R7459t7445) I(R7459t6471) I(R7459t5505) I(R7459t6459) I(R7460t2402) I(R7460t2667) I(R7461t1285) I(R7461t6877) I(R7461t5628) I(R7461t3044) I(R7461t710) I(R7462t5464) I(R7462t4113) I(R7462t219) I(R7462t3000) I(R7462t1142) I(R7462t3314) I(R7463t3204) I(R7463t5658) I(R7463t1582) I(R7463t3934) I(R7464t3514) I(R7464t7284) I(R7464t3464) I(R7464t1783) I(R7464t3942) I(R7464t4412) I(R7465t546) I(R7465t4561) I(R7465t6716) I(R7465t3144) I(R7465t5056) I(R7465t6675) I(R7465t7076) I(R7465t953) I(R7465t1225) I(R7466t1123) I(R7466t7338) I(R7466t5781) I(R7466t925) I(R7467t1621) I(R7467t2726) I(R7467t5353) I(R7467t3846) I(R7467t852) I(R7468t3415) I(R7468t1081) I(R7468t1313) I(R7469t2113) I(R7469t3057) I(R7469t3679) I(R7469t2238) I(R7470t3876) I(R7470t6295) I(R7470t2688) I(R7470t6075) I(R7470t6474) I(R7471t1117) I(R7471t5427) I(R7472t1130) I(R7472t4682) I(R7472t1492) I(R7472t5361) I(R7473t7027) I(R7473t1818) I(R7473t3170) I(R7473t1508) I(R7473t2153) I(R7473t830) I(R7474t3511) I(R7474t4904) I(R7474t3804) I(R7474t7393) I(R7474t2933) I(R7475t1390) I(R7475t1941) I(R7475t3070) I(R7475t6539) I(R7475t5554) I(R7476t2025) I(R7476t5195) I(R7476t1150) I(R7476t3835) I(R7476t723) I(R7477t1041) I(R7477t6878) I(R7477t5366) I(R7477t2738) I(R7478t622) I(R7478t3469) I(R7479t3305) I(R7479t5006) I(R7479t2070) I(R7479t4588) I(R7479t6549) I(R7480t379) I(R7480t5944) I(R7480t5532) I(R7480t2999) I(R7481t478) I(R7481t3386) I(R7481t4232) I(R7482t5168) I(R7482t128) I(R7482t7040) I(R7482t4324) I(R7483t6467) I(R7483t4076) I(R7483t5611) I(R7483t5187) I(R7484t4333) I(R7484t5575) I(R7484t533) I(R7485t1783) I(R7485t3048) I(R7485t4909) I(R7485t3096) I(R7485t6120) I(R7485t3464) I(R7485t7464) I(R7486t3176) I(R7486t2504) I(R7487t6127) I(R7487t1945) I(R7487t6318) I(R7487t4122) I(R7488t4325) I(R7488t5154) I(R7488t1991) I(R7488t7299) I(R7489t5986) I(R7489t7447) I(R7489t2250) I(R7490t1650) I(R7490t3580) I(R7490t6002) I(R7491t1152) I(R7491t7326) I(R7491t1017) I(R7491t5830) I(R7491t7236) I(R7491t1103) I(R7492t4904) I(R7492t7146) I(R7492t5820) I(R7493t3253) I(R7493t2257) I(R7493t4533) I(R7493t6805) I(R7494t877) I(R7494t1519) I(R7494t894) I(R7494t6943) I(R7494t7171) I(R7495t1534) I(R7495t3299) I(R7495t2819) I(R7495t3316) I(R7496t4506) I(R7496t3263) I(R7496t3108) I(R7496t1308) I(R7497t2586) I(R7497t3262) I(R7497t288) I(R7497t5053) I(R7497t14) I(R7498t1276) I(R7498t2601) I(R7498t6411) I(R7498t616) I(R7498t4405) I(R7499t2739) I(R7499t6378) I(R7499t5764) I(R7500t23) I(R7500t6702) I(R7500t6521) I(R7500t3491) I(R7500t6105) I(R7502t1896) I(R7502t5198) I(R7502t2349) I(R7502t2147) I(R7502t25) I(R7502t5054) I(R7503t4731) I(R7503t3865) I(R7503t896) I(R7503t2750) I(R7503t5651) I(R7504t1371) I(R7504t5827) I(R7504t2110) I(R7504t6828) I(R7505t4333) I(R7505t4451) I(R7505t7484) I(R7505t533) I(R7505t6156) I(R7505t3349) I(R7506t4904) I(R7506t7146) I(R7506t3160) I(R7506t1157) I(R7506t3804) I(R7506t3511) I(R7507t3306) I(R7507t2100) I(R7507t3025) I(R7507t2209) I(R7508t3061) I(R7508t4867) I(R7508t3139) I(R7509t2809) I(R7509t5818) I(R7509t4078) I(R7509t3811) I(R7509t1450) I(R7510t1176) I(R7510t2176) I(R7510t2177) I(R7510t2690) I(R7510t2995) I(R7510t2597) I(R7510t6814) I(R7510t3955) I(R7510t1111) I(R7511t1782) I(R7511t2635) I(R7511t5639) I(R7512t5031) I(R7512t4387) I(R7512t2880) I(R7513t1896) I(R7513t6421) I(R7513t7502) I(R7513t5198) I(R7513t3996) I(R7514t6231) I(R7514t5708) I(R7515t3456) I(R7515t6145) I(R7515t6353) I(R7515t3778) I(R7515t5715) I(R7515t6846) I(R7516t7376) I(R7516t6217) I(R7516t92) I(R7517t4605) I(R7517t3712) I(R7517t6918) I(R7517t5829) I(R7518t2226) I(R7518t1808) I(R7519t4937) I(R7519t5244) I(R7519t5881) I(R7520t2319) I(R7520t6807) I(R7520t7372) I(R7521t5254) I(R7521t7305) I(R7521t3699) I(R7522t4397) I(R7522t5582) I(R7522t6841) I(R7522t3234) I(R7522t3651) I(R7523t1587) I(R7523t3054) I(R7523t6185) I(R7523t5702) I(R7524t2529) I(R7524t5820) I(R7524t7492) I(R7524t6875) I(R7524t5740) I(R7524t6567) I(R7525t34) I(R7525t2972) I(R7525t4829) I(R7525t5726) I(R7525t3855) I(R7526t826) I(R7526t6137) I(R7526t2729) I(R7526t4541) I(R7526t357) I(R7526t3300) I(R7527t408) I(R7527t6686) I(R7527t7144) I(R7527t3953) I(R7527t3195) I(R7528t3723) I(R7528t7233) I(R7528t7114) I(R7528t6114) I(R7528t2038) I(R7529t3331) I(R7529t6082) I(R7529t6560) I(R7529t5344) I(R7530t4629) I(R7530t6006) I(R7530t1364) I(R7531t4066) I(R7531t682) I(R7531t4290) I(R7531t1710) I(R7532t5325) I(R7532t3106) I(R7532t6629) I(R7532t287) I(R7532t3911) I(R7532t2547) I(R7532t3620) I(R7533t4607) I(R7533t5844) I(R7533t5574) I(R7533t524) I(R7534t6019) I(R7534t7221) I(R7534t3283) I(R7534t2846) I(R7534t5660) I(R7535t5926) I(R7535t3584) I(R7535t543) I(R7535t1735) I(R7536t4259) I(R7536t6965) I(R7536t4707) I(R7536t7382) I(R7536t6161) I(R7536t552) I(R7537t4511) I(R7537t5691) I(R7537t4675) I(R7537t3525) I(R7537t6324) I(R7537t6382) I(R7538t8) I(R7538t5346) I(R7538t6871) I(R7538t4951) I(R7539t6782) I(R7540t1436) I(R7540t5969) I(R7541t1423) I(R7541t5364) I(R7541t7093) I(R7541t3121) I(R7541t3280) I(R7541t5172) I(R7541t2093) I(R7542t3169) I(R7542t7471) I(R7542t5427) I(R7542t7280) I(R7543t7216) I(R7543t446) I(R7543t4299) I(R7543t2061) I(R7543t1034) I(R7543t5921) I(R7544t3195) I(R7544t6686) I(R7544t7115) I(R7544t5311) I(R7544t865) I(R7544t5981) I(R7545t4656) I(R7545t6616) I(R7545t5249) I(R7545t3800) I(R7546t3830) I(R7546t6772) I(R7546t1217) I(R7546t3801) I(R7546t464) I(R7547t594) I(R7547t2150) I(R7547t4028) I(R7547t1198) I(R7548t4456) I(R7548t898) I(R7548t4310) I(R7549t291) I(R7549t6281) I(R7549t5866) I(R7549t639) I(R7549t6759) I(R7550t6798) I(R7550t6863) I(R7550t2998) I(R7550t4938) I(R7550t5564) I(R7550t2231) I(R7550t343) I(R7551t94) I(R7551t5609) I(R7551t3310) I(R7551t2512) I(R7551t1752) I(R7551t6331) I(R7551t2978) I(R7552t6074) I(R7552t4567) I(R7552t7002) I(R7552t6977) I(R7552t1469) I(R7553t2027) I(R7553t3700) I(R7553t6697) I(R7554t7328) I(R7554t2080) I(R7554t4657) I(R7555t5282) I(R7555t6842) I(R7555t1082) I(R7555t3303) I(R7555t3432) I(R7556t4687) I(R7556t5770) I(R7556t150) I(R7557t2896) I(R7557t1272) I(R7557t3655) I(R7557t2754) I(R7557t524) I(R7558t1927) I(R7558t2392) I(R7558t2005) I(R7558t6373) I(R7559t272) I(R7559t378) I(R7559t1303) I(R7559t1950) I(R7560t3572) I(R7560t5359) I(R7560t6185) I(R7560t1571) I(R7561t9) I(R7561t1826) I(R7562t3878) I(R7563t879) I(R7563t1128) I(R7563t5201) I(R7563t4075) I(R7564t2505) I(R7564t3007) I(R7564t4165) I(R7564t335) I(R7564t1251) I(R7564t3686) I(R7565t3215) I(R7565t2560) I(R7565t2703) I(R7565t4258) I(R7565t5624) I(R7565t1789) I(R7566t495) I(R7566t3537) I(R7566t5377) I(R7566t214) I(R7566t1556) I(R7567t5252) I(R7567t6334) I(R7567t543) I(R7567t4159) I(R7567t390) I(R7567t2521) I(R7568t411) I(R7568t862) I(R7568t7013) I(R7568t3198) I(R7569t1660) I(R7570t1203) I(R7570t2246) I(R7570t3311) I(R7570t6584) I(R7570t5137) I(R7571t4905) I(R7571t7003) I(R7572t3207) I(R7572t4576) I(R7572t1588) I(R7572t4078) I(R7572t4023) I(R7572t5952) I(R7572t5015) I(R7573t2526) I(R7573t4627) I(R7573t6081) I(R7574t1912) I(R7574t4032) I(R7574t5572) I(R7574t1389) I(R7574t1104) I(R7575t809) I(R7575t5500) I(R7575t4184) I(R7576t828) I(R7576t6548) I(R7576t1232) I(R7576t5950) I(R7576t3167) I(R7577t2694) I(R7577t3304) I(R7577t849) I(R7577t6645) I(R7577t2689) I(R7577t1843) I(R7577t4714) I(R7577t3706) I(R7578t1382) I(R7578t7178) I(R7579t1835) I(R7579t4575) I(R7579t2185) I(R7579t7098) I(R7579t2140) I(R7579t2407) I(R7580t1361) I(R7580t1565) I(R7580t3334) I(R7580t4902) I(R7580t7074) I(R7581t6895) I(R7581t7131) I(R7581t4518) I(R7581t7390) I(R7581t2735) I(R7582t1462) I(R7582t3985) I(R7582t732) I(R7582t2118) I(R7583t4519) I(R7583t6888) I(R7583t6583) I(R7583t517) I(R7583t3607) I(R7583t3715) I(R7583t1407) I(R7584t780) I(R7584t6857) I(R7584t6135) I(R7584t320) I(R7584t144) I(R7584t4810) I(R7585t1693) I(R7585t3810) I(R7585t5621) I(R7586t6072) I(R7586t1266) I(R7587t1942) I(R7587t6631) I(R7587t387) I(R7587t2348) I(R7588t3530) I(R7588t3594) I(R7588t7102) I(R7588t544) I(R7589t1275) I(R7589t3366) I(R7589t1827) I(R7589t39) I(R7590t4884) I(R7590t7402) I(R7590t1471) I(R7590t1175) I(R7591t4333) I(R7591t4826) I(R7591t7484) I(R7591t5575) I(R7592t742) I(R7592t1587) I(R7592t3054) I(R7592t7046) I(R7592t5835) I(R7592t4241) I(R7592t3692) I(R7592t1981) I(R7593t6326) I(R7593t3790) I(R7593t6789) I(R7593t2989) I(R7593t1701) I(R7593t5571) I(R7593t6529) I(R7594t2782) I(R7594t5362) I(R7594t3086) I(R7594t4784) I(R7595t301) I(R7595t2463) I(R7595t6901) I(R7595t5275) I(R7595t5512) I(R7596t4291) I(R7596t6206) I(R7596t5219) I(R7596t6204) I(R7596t6792) I(R7596t7079) I(R7596t4111) I(R7596t2440) I(R7597t1160) I(R7597t2891) I(R7597t3777) I(R7597t332) I(R7598t1578) I(R7598t2484) I(R7598t7194) I(R7598t244) I(R7598t6788) I(R7599t4342) I(R7599t4912) I(R7599t2973) I(R7599t1690) I(R7599t150) I(R7599t3446) I(R7600t1761) I(R7600t4644) I(R7600t2662) I(R7600t7336) I(R7601t687) I(R7601t5547) I(R7601t6799) I(R7601t5940) I(R7601t4949) I(R7601t3864) I(R7602t39) I(R7602t1748) I(R7602t7589) I(R7602t1827) I(R7602t5152) I(R7603t2043) I(R7603t4009) I(R7603t3702) I(R7603t7167) I(R7604t4434) I(R7604t6468) I(R7604t761) I(R7604t2947) I(R7604t5571) I(R7604t2989) I(R7605t498) I(R7605t2655) I(R7605t4044) I(R7605t3986) I(R7605t349) I(R7606t7342) I(R7606t3947) I(R7606t5865) I(R7606t5546) I(R7607t1741) I(R7607t2364) I(R7607t5751) I(R7607t5480) I(R7607t3018) I(R7608t377) I(R7608t2170) I(R7608t4272) I(R7608t836) I(R7608t890) I(R7608t155) I(R7609t6618) I(R7609t967) I(R7609t2168) I(R7609t201) I(R7610t2970) I(R7610t5317) I(R7610t532) I(R7610t7327) I(R7610t5130) I(R7611t6556) I(R7611t7357) I(R7611t1581) I(R7611t5599) I(R7611t6112) I(R7611t2244) I(R7611t2293) I(R7612t6141) I(R7612t7486) I(R7612t3176) I(R7613t935) I(R7613t1636) I(R7613t2878) I(R7613t4619) I(R7614t843) I(R7614t2651) I(R7614t209) I(R7614t6749) I(R7614t4098) I(R7614t425) I(R7615t664) I(R7615t5323) I(R7615t2311) I(R7615t4762) I(R7615t7004) I(R7615t2110) I(R7615t2117) I(R7616t2619) I(R7616t6899) I(R7616t4992) I(R7616t4089) I(R7617t1266) I(R7617t5772) I(R7617t5766) I(R7617t6541) I(R7617t4608) I(R7617t4817) I(R7617t2944) I(R7618t436) I(R7618t762) I(R7618t3538) I(R7618t636) I(R7618t5290) I(R7619t7408) I(R7619t1600) I(R7619t4818) I(R7620t6379) I(R7620t881) I(R7620t3029) I(R7621t248) I(R7621t3182) I(R7621t984) I(R7621t7573) I(R7621t2526) I(R7621t2736) I(R7622t408) I(R7622t5471) I(R7622t1046) I(R7623t1872) I(R7623t3456) I(R7623t6504) I(R7623t4252) I(R7623t6353) I(R7623t7515) I(R7624t4740) I(R7624t235) I(R7624t6317) I(R7624t6484) I(R7625t103) I(R7625t5865) I(R7625t7606) I(R7625t3947) I(R7626t3591) I(R7626t4943) I(R7626t1535) I(R7626t1738) I(R7626t1108) I(R7627t4496) I(R7627t3794) I(R7627t6260) I(R7627t5011) I(R7628t274) I(R7628t3644) I(R7628t4654) I(R7628t2641) I(R7628t5150) I(R7628t3152) I(R7629t4492) I(R7629t2594) I(R7629t6793) I(R7629t2347) I(R7629t2242) I(R7630t1160) I(R7630t4874) I(R7630t6975) I(R7630t7189) I(R7630t3119) I(R7630t3647) I(R7630t332) I(R7631t3934) I(R7631t7463) I(R7631t2953) I(R7632t997) I(R7632t5036) I(R7632t80) I(R7632t2294) I(R7632t6184) I(R7632t7429) I(R7633t1806) I(R7633t3885) I(R7633t1247) I(R7633t5627) I(R7633t3875) I(R7633t2874) I(R7634t1148) I(R7634t579) I(R7634t5842) I(R7634t7245) I(R7634t2111) I(R7635t4277) I(R7635t4754) I(R7635t1063) I(R7635t6232) I(R7636t1530) I(R7636t137) I(R7636t6109) I(R7636t1069) I(R7637t1860) I(R7637t7133) I(R7637t1585) I(R7637t3295) I(R7637t5880) I(R7637t7136) I(R7637t3261) I(R7638t2466) I(R7638t3362) I(R7638t3774) I(R7638t3451) I(R7639t1136) I(R7639t3611) I(R7639t6682) I(R7639t4224) I(R7640t4911) I(R7640t3604) I(R7640t2033) I(R7640t196) I(R7641t2601) I(R7641t7498) I(R7641t5880) I(R7641t6411) I(R7642t4789) I(R7642t2232) I(R7643t2384) I(R7643t2783) I(R7643t5515) I(R7643t4304) I(R7643t6989) I(R7644t5097) I(R7644t5518) I(R7644t5224) I(R7644t2621) I(R7645t3198) I(R7645t6471) I(R7645t5505) I(R7645t4684) I(R7645t4380) I(R7645t3567) I(R7645t296) I(R7645t3125) I(R7645t7013) I(R7646t1282) I(R7646t5722) I(R7646t2798) I(R7646t6136) I(R7647t434) I(R7647t1448) I(R7647t1442) I(R7647t4204) I(R7648t5059) I(R7648t5728) I(R7648t2811) I(R7648t1513) I(R7648t4128) I(R7649t1292) I(R7649t6928) I(R7649t7188) I(R7649t4751) I(R7650t5116) I(R7650t6434) I(R7650t5888) I(R7650t6100) I(R7650t5659) I(R7651t1362) I(R7651t3319) I(R7651t5446) I(R7651t2790) I(R7651t2831) I(R7651t2382) I(R7651t2794) I(R7652t347) I(R7652t6064) I(R7652t3489) I(R7652t4549) I(R7652t7065) I(R7653t5736) I(R7653t3320) I(R7653t1755) I(R7653t4542) I(R7653t4394) I(R7654t1798) I(R7654t6132) I(R7654t799) I(R7654t4071) I(R7655t1645) I(R7655t678) I(R7655t7259) I(R7656t2356) I(R7656t1728) I(R7656t4982) I(R7657t1692) I(R7657t5767) I(R7658t3110) I(R7658t2534) I(R7658t3212) I(R7658t3714) I(R7659t4806) I(R7659t6225) I(R7659t985) I(R7659t1732) I(R7659t5603) I(R7660t3386) I(R7660t7481) I(R7660t3883) I(R7660t4185) I(R7660t4191) I(R7660t4105) I(R7660t204) I(R7661t3305) I(R7661t3426) I(R7661t2294) I(R7661t6586) I(R7661t2286) I(R7661t3038) I(R7661t530) I(R7663t2649) I(R7663t876) I(R7663t5795) I(R7663t3277) I(R7664t5440) I(R7664t6573) I(R7664t3744) I(R7664t6754) I(R7664t6204) I(R7664t111) I(R7665t5824) I(R7665t6368) I(R7665t4758) I(R7665t3437) I(R7666t859) I(R7666t7431) I(R7666t5548) I(R7666t888) I(R7666t4215) I(R7666t3321) I(R7667t711) I(R7667t3784) I(R7667t1314) I(R7667t959) I(R7668t2200) I(R7668t2903) I(R7668t2347) I(R7668t6793) I(R7668t5993) I(R7668t1260) I(R7669t543) I(R7669t3805) I(R7669t7567) I(R7669t4159) I(R7670t6173) I(R7670t6629) I(R7670t3702) I(R7671t3091) I(R7671t6231) I(R7672t2185) I(R7672t2187) I(R7672t4575) I(R7672t6153) I(R7672t6258) I(R7673t2466) I(R7673t7638) I(R7673t4360) I(R7673t2190) I(R7674t5794) I(R7674t5977) I(R7675t3801) I(R7675t6148) I(R7675t6479) I(R7675t4505) I(R7676t1328) I(R7676t163) I(R7676t2916) I(R7676t735) I(R7677t1048) I(R7677t3778) I(R7677t5715) I(R7677t746) I(R7678t4782) I(R7678t4740) I(R7679t3021) I(R7679t3284) I(R7679t3365) I(R7679t2745) I(R7680t3661) I(R7680t3717) I(R7680t4314) I(R7680t279) I(R7680t370) I(R7681t1038) I(R7681t5173) I(R7681t2855) I(R7681t4538) I(R7681t6383) I(R7682t4897) I(R7682t7182) I(R7682t5292) I(R7683t2451) I(R7683t6976) I(R7683t5072) I(R7683t1576) I(R7683t6424) I(R7684t1959) I(R7684t3425) I(R7684t1001) I(R7685t1861) I(R7685t5155) I(R7685t2644) I(R7685t4952) I(R7685t5736) I(R7686t919) I(R7686t3055) I(R7686t3098) I(R7686t537) I(R7686t861) I(R7686t1557) I(R7687t2962) I(R7687t6562) I(R7688t4877) I(R7688t7225) I(R7688t207) I(R7688t1598) I(R7688t1991) I(R7689t4726) I(R7689t2862) I(R7690t3649) I(R7690t4952) I(R7691t435) I(R7691t6533) I(R7691t5022) I(R7691t3431) I(R7691t2587) I(R7691t1634) I(R7691t861) I(R7692t4461) I(R7692t4895) I(R7692t292) I(R7692t904) I(R7692t116) I(R7693t4234) I(R7693t6648) I(R7693t5817) I(R7694t2706) I(R7694t3653) I(R7694t1569) I(R7694t1305) I(R7694t6663) I(R7695t684) I(R7695t6530) I(R7695t6579) I(R7696t1370) I(R7696t5896) I(R7696t1035) I(R7697t3094) I(R7697t4352) I(R7697t6811) I(R7697t2205) I(R7698t3061) I(R7698t914) I(R7698t5846) I(R7698t4867) I(R7699t1661) I(R7699t4264) I(R7699t3848) I(R7699t3112) I(R7699t4077) I(R7699t549) I(R7700t4887) I(R7700t7090) I(R7700t2897) I(R7700t1744) I(R7700t79) I(R7700t4893) I(R7701t2463) I(R7701t2080) I(R7701t7554) I(R7701t4657) I(R7701t6944) I(R7702t372) I(R7702t5171) I(R7702t838) I(R7702t3423) I(R7702t592) I(R7702t318) I(R7703t2867) I(R7703t6419) I(R7703t3500) I(R7703t222) I(R7703t3408) I(R7704t3141) I(R7704t6665) I(R7704t3861) I(R7704t1574) I(R7704t4409) I(R7704t2925) I(R7705t3193) I(R7705t5821) I(R7705t2099) I(R7705t6566) I(R7705t7260) I(R7705t1422) I(R7706t3253) I(R7706t7493) I(R7706t2257) I(R7706t4386) I(R7706t5545) I(R7707t4465) I(R7707t4997) I(R7707t7206) I(R7707t5500) I(R7707t3546) I(R7708t4153) I(R7708t3958) I(R7708t132) I(R7708t5069) I(R7708t6272) I(R7709t5063) I(R7709t1399) I(R7709t3089) I(R7709t6241) I(R7710t1633) I(R7710t6250) I(R7710t3989) I(R7710t4807) I(R7710t3223) I(R7710t6527) I(R7710t4601) I(R7711t4731) I(R7711t7009) I(R7711t4816) I(R7711t823) I(R7711t3865) I(R7711t7503) I(R7712t1912) I(R7712t4032) I(R7712t5572) I(R7712t4012) I(R7712t5463) I(R7712t4900) I(R7712t2539) I(R7713t3751) I(R7713t949) I(R7713t4676) I(R7713t2562) I(R7714t7380) I(R7714t1622) I(R7714t1607) I(R7714t3780) I(R7715t5149) I(R7715t2894) I(R7715t2544) I(R7716t1910) I(R7716t4156) I(R7716t1647) I(R7716t3051) I(R7716t2639) I(R7717t4604) I(R7717t4645) I(R7718t5585) I(R7718t3265) I(R7718t2917) I(R7719t1871) I(R7719t6144) I(R7719t600) I(R7719t6553) I(R7719t1405) I(R7720t3067) I(R7720t427) I(R7721t969) I(R7721t5296) I(R7721t7578) I(R7721t2447) I(R7722t4195) I(R7722t7187) I(R7722t1227) I(R7722t4363) I(R7722t1233) I(R7722t3578) I(R7722t1961) I(R7722t2415) I(R7723t1085) I(R7723t700) I(R7723t5002) I(R7723t2555) I(R7723t6688) I(R7723t5413) I(R7724t367) I(R7724t4685) I(R7724t1551) I(R7724t2450) I(R7724t824) I(R7725t5966) I(R7725t4716) I(R7725t1908) I(R7725t415) I(R7726t2379) I(R7726t5277) I(R7726t1189) I(R7726t2448) I(R7726t7044) I(R7726t1689) I(R7727t2277) I(R7727t893) I(R7728t3384) I(R7728t4453) I(R7729t6717) I(R7729t6796) I(R7729t7018) I(R7730t426) I(R7730t4286) I(R7730t6011) I(R7730t3957) I(R7730t7160) I(R7731t299) I(R7731t1193) I(R7731t5018) I(R7731t3388) I(R7731t221) I(R7731t942) I(R7732t908) I(R7732t4725) I(R7732t838) I(R7732t5769) I(R7733t1081) I(R7733t7468) I(R7733t1313) I(R7733t158) I(R7733t4090) I(R7733t5079) I(R7733t6852) I(R7734t1722) I(R7734t6366) I(R7734t1671) I(R7734t2990) I(R7734t3134) I(R7735t7547) I(R7735t594) I(R7735t2030) I(R7735t7423) I(R7735t4980) I(R7735t677) I(R7735t213) I(R7735t6650) I(R7736t2334) I(R7736t5314) I(R7736t3671) I(R7736t3427) I(R7736t1857) I(R7736t6891) I(R7736t5984) I(R7736t1814) I(R7736t1713) I(R7736t3829) I(R7737t813) I(R7737t3812) I(R7737t7204) I(R7737t2154) I(R7737t6273) I(R7738t1455) I(R7738t6269) I(R7738t4156) I(R7738t1647) I(R7739t2787) I(R7739t2994) I(R7739t5382) I(R7739t825) I(R7740t7478) I(R7740t7406) I(R7740t93) I(R7741t6210) I(R7741t3807) I(R7741t3813) I(R7741t1997) I(R7741t6465) I(R7742t6680) I(R7742t5262) I(R7742t2409) I(R7742t1956) I(R7742t7363) I(R7743t1377) I(R7743t6734) I(R7743t2211) I(R7743t2670) I(R7743t6407) I(R7743t5085) I(R7743t4992) I(R7743t4367) I(R7744t2291) I(R7744t2532) I(R7744t476) I(R7744t4856) I(R7744t2145) I(R7744t709) I(R7744t977) I(R7745t2875) I(R7745t629) I(R7745t1019) I(R7745t6575) I(R7746t4364) I(R7746t1107) I(R7746t1527) I(R7746t6167) I(R7747t5741) I(R7747t3468) I(R7747t1911) I(R7747t3137) I(R7748t1651) I(R7748t6453) I(R7748t440) I(R7748t7434) I(R7748t2548) I(R7748t3361) I(R7749t1480) I(R7749t7171) I(R7749t7494) I(R7749t1519) I(R7749t631) I(R7749t5892) I(R7750t432) I(R7750t4566) I(R7750t1807) I(R7750t2737) I(R7750t4390) I(R7751t10) I(R7751t6827) I(R7751t4780) I(R7751t7002) I(R7751t5578) I(R7751t4570) I(R7752t3138) I(R7752t2435) I(R7752t7224) I(R7752t3369) I(R7753t1788) I(R7753t6340) I(R7753t156) I(R7753t4295) I(R7754t3725) I(R7754t658) I(R7754t3896) I(R7754t5206) I(R7754t926) I(R7755t2832) I(R7755t5541) I(R7755t2775) I(R7755t1488) I(R7755t4641) I(R7755t7384) I(R7755t4501) I(R7756t2070) I(R7756t5006) I(R7756t2643) I(R7756t5358) I(R7757t6761) I(R7757t7050) I(R7757t1528) I(R7757t145) I(R7757t716) I(R7758t331) I(R7758t4610) I(R7758t657) I(R7758t7101) I(R7759t5323) I(R7759t7116) I(R7759t4323) I(R7759t905) I(R7759t6404) I(R7759t512) I(R7759t2311) I(R7759t664) I(R7760t74) I(R7760t1584) I(R7760t4694) I(R7760t3772) I(R7760t2731) I(R7760t1586) I(R7761t621) I(R7761t4463) I(R7761t3731) I(R7761t3797) I(R7761t7177) I(R7762t2618) I(R7762t6228) I(R7762t5257) I(R7762t7182) I(R7762t7682) I(R7762t5292) I(R7763t1036) I(R7763t7414) I(R7763t455) I(R7763t1834) I(R7763t4908) I(R7763t3440) I(R7764t7083) I(R7764t5945) I(R7764t5427) I(R7764t7570) I(R7764t3311) I(R7764t1788) I(R7765t7129) I(R7765t2723) I(R7767t5717) I(R7767t35) I(R7767t445) I(R7768t6957) I(R7768t6782) I(R7768t4061) I(R7768t4401) I(R7768t3154) I(R7769t6701) I(R7769t7314) I(R7769t4410) I(R7769t2007) I(R7770t6670) I(R7770t5971) I(R7770t6920) I(R7770t3074) I(R7770t2678) I(R7771t1881) I(R7771t3353) I(R7771t1368) I(R7771t6624) I(R7772t896) I(R7772t2750) I(R7772t7503) I(R7773t1539) I(R7773t5475) I(R7773t662) I(R7773t2785) I(R7774t3302) I(R7774t4249) I(R7774t5926) I(R7774t3584) I(R7774t354) I(R7774t5866) I(R7774t6637) I(R7775t8) I(R7775t5324) I(R7775t4848) I(R7775t4951) I(R7775t7538) I(R7776t1797) I(R7776t3891) I(R7776t4529) I(R7776t6868) I(R7776t2633) I(R7776t631) I(R7777t2550) I(R7777t5968) I(R7777t2510) I(R7777t975) I(R7777t889) I(R7777t7439) I(R7777t677) I(R7778t3992) I(R7778t1733) I(R7778t1054) I(R7778t3147) I(R7779t911) I(R7779t6175) I(R7779t1796) I(R7779t6014) I(R7779t2385) I(R7779t880) I(R7780t3707) I(R7780t4700) I(R7780t6987) I(R7780t1423) I(R7780t5596) I(R7781t4695) I(R7781t2317) I(R7781t6752) I(R7781t1978) I(R7782t6924) I(R7782t5014) I(R7782t1486) I(R7782t3248) I(R7782t5914) I(R7783t3773) I(R7783t1973) I(R7783t6359) I(R7784t598) I(R7784t2640) I(R7784t4743) I(R7784t635) I(R7785t360) I(R7785t185) I(R7785t4999) I(R7785t6845) I(R7785t302) I(R7785t6567) I(R7786t6412) I(R7786t9) I(R7786t7561) I(R7786t1826) I(R7786t4674) I(R7786t3424) I(R7787t355) I(R7787t4423) I(R7787t4767) I(R7787t6707) I(R7787t5146) I(R7787t4265) I(R7787t4377) I(R7788t1862) I(R7788t3285) I(R7788t6251) I(R7788t3491) I(R7788t7500) I(R7788t1263) I(R7789t513) I(R7789t6631) I(R7789t2348) I(R7790t1216) I(R7790t6300) I(R7790t4275) I(R7790t462) I(R7791t7414) I(R7791t7763) I(R7791t2313) I(R7791t3140) I(R7791t455) I(R7792t1065) I(R7792t4902) I(R7792t2862) I(R7792t7689) I(R7792t405) I(R7793t1403) I(R7793t4227) I(R7793t5225) I(R7794t88) I(R7794t3897) I(R7794t5897) I(R7795t7059) I(R7795t481) I(R7795t7444) I(R7795t5808) I(R7796t4605) I(R7796t7517) I(R7796t3712) I(R7796t1949) I(R7796t7275) I(R7796t7337) I(R7797t1367) I(R7797t6430) I(R7797t5841) I(R7797t831) I(R7797t7318) I(R7797t4235) I(R7798t5344) I(R7798t1937) I(R7798t2035) I(R7798t7057) I(R7798t3338) I(R7799t2876) I(R7799t3697) I(R7799t7197) I(R7800t3392) I(R7800t4513) I(R7800t24) I(R7800t4190) I(R7800t1566) I(R7801t6761) I(R7801t7757) I(R7801t4761) I(R7801t5090) I(R7802t3396) I(R7802t3892) I(R7802t6746) I(R7802t6993) I(R7803t3516) I(R7803t4520) I(R7803t4006) I(R7803t4699) I(R7804t889) I(R7804t7132) I(R7804t6422) I(R7804t4289) I(R7804t2718) I(R7804t7439) I(R7804t7777) I(R7805t3694) I(R7805t4688) I(R7805t5681) I(R7805t6395) I(R7805t3250) I(R7805t7337) I(R7805t7796) I(R7805t7275) I(R7805t1010) I(R7807t3720) I(R7807t5390) I(R7807t646) I(R7807t7008) I(R7807t5819) I(R7808t10) I(R7808t489) I(R7808t6827) I(R7808t92) I(R7808t3984) I(R7809t17) I(R7809t3545) I(R7809t3583) I(R7809t6410) I(R7809t184) I(R7809t884) I(R7810t1292) I(R7810t5103) I(R7810t4128) I(R7810t5498) I(R7810t6633) I(R7810t4751) I(R7810t7649) I(R7811t334) I(R7811t365) I(R7811t3169) I(R7811t7542) I(R7811t7280) I(R7811t1605) I(R7812t7500) I(R7812t7788) I(R7812t1263) I(R7812t3544) I(R7813t5039) I(R7813t6150) I(R7813t4491) I(R7813t2857) I(R7814t1159) I(R7814t6374) I(R7814t1488) I(R7814t4641) I(R7815t825) I(R7815t5777) I(R7816t3077) I(R7816t5554) I(R7816t7475) I(R7816t6539) I(R7816t4354) I(R7817t7459) I(R7817t4684) I(R7817t7645) I(R7817t5505) I(R7818t6235) I(R7818t6910) I(R7818t6501) I(R7818t5343) I(R7819t5277) I(R7819t5832) I(R7819t2379) I(R7819t395) I(R7819t1011) I(R7819t5581) I(R7819t3101) I(R7819t7205) I(R7820t4949) I(R7820t5940) I(R7820t4095) I(R7820t2676) I(R7820t2223) I(R7821t211) I(R7821t2818) I(R7821t1509) I(R7821t4785) I(R7822t862) I(R7822t4882) I(R7822t7013) I(R7822t2324) I(R7823t1838) I(R7823t6591) I(R7823t7288) I(R7823t2559) I(R7824t3932) I(R7824t6001) I(R7824t3079) I(R7824t1025) I(R7825t3455) I(R7826t5709) I(R7826t6298) I(R7826t4713) I(R7826t2023) I(R7827t122) I(R7827t2839) I(R7827t6696) I(R7827t3794) I(R7828t3021) I(R7828t7679) I(R7828t2745) I(R7828t1302) I(R7828t2836) I(R7829t372) I(R7829t838) I(R7829t7732) I(R7829t4485) I(R7830t5281) I(R7830t6723) I(R7830t143) I(R7830t5870) I(R7830t7427) I(R7830t5992) I(R7831t4587) I(R7831t7048) I(R7831t2515) I(R7831t4506) I(R7831t4466) I(R7831t6938) I(R7831t3387) I(R7832t5115) I(R7832t1689) I(R7832t77) I(R7833t1413) I(R7833t2660) I(R7834t1798) I(R7834t3575) I(R7834t4700) I(R7834t6572) I(R7835t1381) I(R7835t4974) I(R7835t4992) I(R7835t7616) I(R7835t6309) I(R7836t74) I(R7836t4694) I(R7836t4433) I(R7836t6226) I(R7836t2692) I(R7836t6602) I(R7837t1826) I(R7837t2437) I(R7837t4742) I(R7837t5351) I(R7838t3928) I(R7838t5524) I(R7838t1375) I(R7839t2050) I(R7839t6426) I(R7839t1554) I(R7839t5211) I(R7839t3988) I(R7839t2032) I(R7839t6488) I(R7839t6452) I(R7839t149) I(R7840t1726) I(R7840t4364) I(R7840t7746) I(R7840t2590) I(R7840t187) I(R7840t7240) I(R7841t6194) I(R7841t1868) I(R7841t808) I(R7842t55) I(R7842t2453) I(R7842t6195) I(R7842t3573) I(R7843t4531) I(R7843t5704) I(R7843t2518) I(R7844t3) I(R7844t3552) I(R7844t1383) I(R7845t6336) I(R7845t7333) I(R7845t1620) I(R7845t6764) I(R7846t4897) I(R7846t7682) I(R7846t5292) I(R7846t2904) I(R7847t7478) I(R7847t7740) I(R7847t7406) I(R7847t222) I(R7847t3469) I(R7848t6017) I(R7848t6200) I(R7848t3774) I(R7848t7638) I(R7848t7673) I(R7848t7562) I(R7848t3878) I(R7849t1743) I(R7849t1335) I(R7849t4399) I(R7849t1293) I(R7850t3987) I(R7850t2608) I(R7850t1761) I(R7851t648) I(R7851t5586) I(R7851t913) I(R7851t3937) I(R7851t2797) I(R7851t5606) I(R7851t787) I(R7852t5618) I(R7852t1656) I(R7852t4325) I(R7852t7488) I(R7852t2743) I(R7852t5129) I(R7853t4094) I(R7853t5915) I(R7853t2719) I(R7853t3932) I(R7853t7824) I(R7853t1025) I(R7854t374) I(R7854t6818) I(R7854t2490) I(R7854t7447) I(R7854t5468) I(R7855t7216) I(R7855t472) I(R7855t2280) I(R7855t6255) I(R7856t2112) I(R7856t6115) I(R7856t712) I(R7856t3991) I(R7857t2908) I(R7857t4727) I(R7857t4784) I(R7857t2782) I(R7857t4439) I(R7857t1197) I(R7857t6516) I(R7858t423) I(R7858t6839) I(R7858t1441) I(R7858t4194) I(R7858t5872) I(R7859t6169) I(R7859t6639) I(R7859t4153) I(R7859t7708) I(R7859t2361) I(R7860t2084) I(R7860t7395) I(R7860t3229) I(R7861t5966) I(R7861t7297) I(R7861t4230) I(R7861t6290) I(R7861t4716) I(R7861t7725) I(R7862t3196) I(R7862t112) I(R7862t3324) I(R7862t5389) I(R7863t2818) I(R7863t7821) I(R7863t1947) I(R7863t7454) I(R7863t4785) I(R7864t916) I(R7864t1283) I(R7864t2552) I(R7864t971) I(R7864t2592) I(R7865t745) I(R7865t6916) I(R7865t4979) I(R7865t5783) I(R7865t6408) I(R7866t2677) I(R7866t1856) I(R7866t6269) I(R7867t2758) I(R7867t1196) I(R7867t2771) I(R7867t4853) I(R7867t2304) I(R7868t1098) I(R7868t5867) I(R7868t5553) I(R7868t2355) I(R7868t391) I(R7869t3817) I(R7869t6750) I(R7869t2277) I(R7869t7727) I(R7869t893) I(R7869t5448) I(R7869t2097) I(R7869t223) I(R7870t4553) I(R7870t7262) I(R7870t1408) I(R7870t3723) I(R7870t3668) I(R7871t6475) I(R7871t6889) I(R7871t4026) I(R7871t4686) I(R7871t4844) I(R7872t5207) I(R7872t6363) I(R7872t182) I(R7872t554) I(R7873t7624) I(R7873t6484) I(R7873t1249) I(R7873t440) I(R7874t1696) I(R7874t3102) I(R7874t1047) I(R7875t2132) I(R7875t7178) I(R7875t5296) I(R7875t7721) I(R7875t7578) I(R7876t1427) I(R7876t4556) I(R7876t4695) I(R7876t6928) I(R7877t4586) I(R7877t1935) I(R7877t1381) I(R7877t3737) I(R7877t1637) I(R7877t1774) I(R7878t5680) I(R7878t6240) I(R7878t3081) I(R7878t4756) I(R7879t3507) I(R7879t6614) I(R7879t1533) I(R7879t237) I(R7880t1761) I(R7880t7600) I(R7880t6953) I(R7880t7336) I(R7881t4761) I(R7881t7801) I(R7881t7757) I(R7881t7050) I(R7881t4001) I(R7881t3453) I(R7882t5585) I(R7882t7718) I(R7882t2922) I(R7883t2048) I(R7883t2579) I(R7883t2268) I(R7883t3961) I(R7884t378) I(R7884t4896) I(R7884t1424) I(R7884t5668) I(R7884t1299) I(R7885t4546) I(R7885t3217) I(R7886t3105) I(R7886t6392) I(R7886t3959) I(R7886t6855) I(R7886t1149) I(R7886t845) I(R7887t244) I(R7887t1060) I(R7887t2510) I(R7887t6339) I(R7887t6279) I(R7887t6788) I(R7888t497) I(R7888t6692) I(R7888t3916) I(R7888t1847) I(R7888t4640) I(R7889t3548) I(R7889t4190) I(R7889t115) I(R7889t5019) I(R7889t5459) I(R7890t1448) I(R7890t6456) I(R7890t3136) I(R7891t992) I(R7891t1018) I(R7891t5387) I(R7891t5476) I(R7892t5885) I(R7892t5960) I(R7892t1315) I(R7892t4396) I(R7893t7227) I(R7893t2657) I(R7893t6201) I(R7893t6179) I(R7893t525) I(R7894t2281) I(R7894t4434) I(R7894t4382) I(R7894t5632) I(R7894t500) I(R7894t5521) I(R7894t5559) I(R7895t5168) I(R7895t4324) I(R7895t6884) I(R7896t4316) I(R7896t7329) I(R7896t4391) I(R7896t2962) I(R7896t7687) I(R7897t3061) I(R7897t6140) I(R7897t3766) I(R7897t5127) I(R7897t358) I(R7897t764) I(R7898t6122) I(R7898t6674) I(R7898t3577) I(R7898t6083) I(R7899t4411) I(R7899t1543) I(R7899t4760) I(R7900t978) I(R7900t4037) I(R7900t3826) I(R7900t5661) I(R7900t7085) I(R7900t2124) I(R7900t5796) I(R7901t968) I(R7901t632) I(R7901t4788) I(R7901t444) I(R7902t2503) I(R7902t3249) I(R7902t1061) I(R7902t4713) I(R7902t2023) I(R7903t2382) I(R7903t5982) I(R7903t2267) I(R7903t3493) I(R7903t3786) I(R7903t2831) I(R7904t5639) I(R7904t5877) I(R7904t1571) I(R7904t6538) I(R7904t5980) I(R7905t3385) I(R7905t5332) I(R7906t3463) I(R7906t6883) I(R7906t1051) I(R7906t5591) I(R7907t605) I(R7907t3286) I(R7907t1095) I(R7907t5148) I(R7907t2453) I(R7908t997) I(R7908t6971) I(R7908t7827) I(R7908t122) I(R7908t2060) I(R7909t1762) I(R7909t7631) I(R7909t2953) I(R7909t2667) I(R7910t3357) I(R7910t7352) I(R7910t313) I(R7910t5941) I(R7910t574) I(R7911t1564) I(R7911t4027) I(R7911t7333) I(R7911t7845) I(R7911t1620) I(R7911t7458) I(R7912t6307) I(R7912t5921) I(R7912t1082) I(R7912t4600) I(R7913t4290) I(R7913t5640) I(R7913t6722) I(R7914t44) I(R7914t4054) I(R7914t7141) I(R7915t6214) I(R7915t6915) I(R7915t4719) I(R7916t4211) I(R7916t5836) I(R7916t4513) I(R7917t6740) I(R7917t4724) I(R7917t2468) I(R7917t2227) I(R7918t411) I(R7918t7568) I(R7918t87) I(R7918t3198) I(R7919t3629) I(R7919t6374) I(R7919t1159) I(R7920t1786) I(R7920t3101) I(R7920t5581) I(R7920t5138) I(R7921t6694) I(R7921t7071) I(R7921t5664) I(R7921t7373) I(R7922t5646) I(R7922t5254) I(R7922t6803) I(R7922t1915) I(R7923t3205) I(R7923t3316) I(R7923t5084) I(R7923t3987) I(R7923t7850) I(R7923t2608) I(R7923t5167) I(R7923t1168) I(R7923t5568) I(R7923t5482) I(R7924t6673) I(R7924t7326) I(R7924t602) I(R7924t3664) I(R7924t4967) I(R7924t5699) I(R7925t2359) I(R7925t5170) I(R7925t5589) I(R7926t533) I(R7926t7484) I(R7926t3501) I(R7926t2732) I(R7926t5575) I(R7927t2214) I(R7927t2614) I(R7927t3171) I(R7927t5599) I(R7927t7611) I(R7927t1581) I(R7928t7196) I(R7928t3962) I(R7928t4620) I(R7928t2829) I(R7929t1403) I(R7929t5225) I(R7929t7793) I(R7929t2751) I(R7930t1074) I(R7930t3488) I(R7930t5797) I(R7930t576) I(R7930t747) I(R7931t5847) I(R7931t6142) I(R7931t1653) I(R7931t618) I(R7932t311) I(R7932t2180) I(R7932t5996) I(R7932t666) I(R7933t2073) I(R7933t3084) I(R7933t6500) I(R7933t4238) I(R7933t1600) I(R7933t4818) I(R7934t285) I(R7934t7030) I(R7934t1992) I(R7934t4471) I(R7934t1749) I(R7934t5763) I(R7935t3941) I(R7935t4216) I(R7935t3403) I(R7935t1921) I(R7935t7250) I(R7936t4553) I(R7936t7121) I(R7936t2073) I(R7936t3668) I(R7936t7870) I(R7937t2513) I(R7937t3719) I(R7937t3648) I(R7937t3760) I(R7937t4238) I(R7937t4917) I(R7937t69) I(R7937t1597) I(R7937t2541) I(R7938t6319) I(R7939t1385) I(R7939t1866) I(R7939t2849) I(R7939t6264) I(R7940t1539) I(R7940t5294) I(R7940t1810) I(R7940t6515) I(R7940t962) I(R7940t1957) I(R7941t1804) I(R7941t5376) I(R7942t6934) I(R7942t3405) I(R7942t1782) I(R7942t7511) I(R7942t5639) I(R7942t3572) I(R7943t6518) I(R7943t7139) I(R7944t2425) I(R7944t3999) I(R7944t6789) I(R7945t4432) I(R7945t6171) I(R7945t5954) I(R7945t7407) I(R7945t2) I(R7946t933) I(R7946t4204) I(R7946t217) I(R7946t6098) I(R7946t620) I(R7946t5260) I(R7947t1363) I(R7947t3248) I(R7947t7782) I(R7947t1486) I(R7947t6599) I(R7948t1021) I(R7948t2345) I(R7948t7341) I(R7948t5128) I(R7949t2333) I(R7949t6587) I(R7949t3893) I(R7949t6786) I(R7949t5904) I(R7950t6492) I(R7950t3792) I(R7951t5031) I(R7951t7512) I(R7951t1411) I(R7951t7684) I(R7951t4387) I(R7952t4531) I(R7952t6766) I(R7952t7242) I(R7952t2518) I(R7953t4665) I(R7953t5935) I(R7953t2003) I(R7953t4143) I(R7953t996) I(R7954t169) I(R7954t1470) I(R7954t4858) I(R7954t2516) I(R7955t1870) I(R7955t6589) I(R7955t3693) I(R7955t2627) I(R7955t2090) I(R7955t7107) I(R7955t4747) I(R7956t91) I(R7956t7421) I(R7956t3402) I(R7956t406) I(R7956t473) I(R7957t1073) I(R7957t5681) I(R7957t5839) I(R7957t661) I(R7958t5349) I(R7958t4274) I(R7958t6288) I(R7958t38) I(R7959t743) I(R7959t6677) I(R7959t5284) I(R7959t385) I(R7959t2615) I(R7960t1002) I(R7960t3322) I(R7960t3858) I(R7960t5911) I(R7960t1077) I(R7960t3899) I(R7961t2481) I(R7961t6530) I(R7961t1663) I(R7961t2201) I(R7961t5626) I(R7961t6726) I(R7961t6787) I(R7962t1498) I(R7962t6496) I(R7962t535) I(R7962t6836) I(R7963t686) I(R7963t6916) I(R7963t7865) I(R7963t745) I(R7964t4335) I(R7964t5524) I(R7964t7838) I(R7964t1375) I(R7965t3710) I(R7965t4241) I(R7965t6890) I(R7965t1921) I(R7965t729) I(R7965t4559) I(R7965t2635) I(R7965t6332) I(R7965t3054) I(R7966t3725) I(R7966t4413) I(R7966t2800) I(R7966t2427) I(R7967t5112) I(R7967t4014) I(R7967t1802) I(R7967t203) I(R7968t647) I(R7968t6504) I(R7968t6123) I(R7968t4417) I(R7968t7292) I(R7969t4227) I(R7969t7793) I(R7969t1583) I(R7969t5746) I(R7969t2751) I(R7969t7929) I(R7970t2274) I(R7970t499) I(R7970t5893) I(R7970t3746) I(R7971t1674) I(R7971t2659) I(R7971t6668) I(R7971t3954) I(R7972t186) I(R7972t321) I(R7972t319) I(R7972t5148) I(R7972t1095) I(R7972t5478) I(R7972t4407) I(R7973t5118) I(R7973t2666) I(R7973t1902) I(R7973t617) I(R7973t6400) I(R7973t2064) I(R7974t7501) I(R7974t5280) I(R7974t1561) I(R7974t1785) I(R7975t2152) I(R7975t7298) I(R7975t3578) I(R7975t5544) I(R7976t1454) I(R7976t3963) I(R7976t6812) I(R7976t1067) I(R7977t1148) I(R7977t4393) I(R7977t4437) I(R7977t4705) I(R7978t4990) I(R7978t3676) I(R7979t509) I(R7979t2675) I(R7979t5470) I(R7979t3465) I(R7980t3598) I(R7980t3704) I(R7980t6057) I(R7980t1211) I(R7981t2068) I(R7982t3853) I(R7982t4352) I(R7982t6807) I(R7982t7520) I(R7982t2696) I(R7982t7697) I(R7983t1391) I(R7984t1676) I(R7984t5176) I(R7984t6733) I(R7984t1162) I(R7984t5901) I(R7985t650) I(R7985t721) I(R7985t203) I(R7986t5985) I(R7986t6264) I(R7986t4281) I(R7986t553) I(R7987t1675) I(R7987t5358) I(R7987t7756) I(R7988t1696) I(R7988t2795) I(R7988t3102) I(R7988t7874) I(R7989t1141) I(R7989t694) I(R7989t5430) I(R7989t2105) I(R7990t3660) I(R7990t5688) I(R7990t3468) I(R7990t3183) I(R7990t1219) I(R7991t1952) I(R7991t5408) I(R7991t6051) I(R7991t6867) I(R7991t3696) I(R7992t1548) I(R7992t5350) I(R7992t6644) I(R7992t4846) I(R7993t5485) I(R7993t6461) I(R7993t4762) I(R7993t1205) I(R7993t5799) I(R7994t5062) I(R7994t4498) I(R7994t2431) I(R7995t4637) I(R7995t3505) I(R7995t6647) I(R7995t3776) I(R7996t255) I(R7996t2608) I(R7996t5597) I(R7996t1761) I(R7996t7850) I(R7997t4064) I(R7997t4068) I(R7997t1509) I(R7997t4175) I(R7997t4634) I(R7998t2684) I(R7998t7289) I(R7998t917) I(R7998t4581) I(R7998t7443) I(R7998t3978) I(R7998t7217) I(R7999t5474) I(R7999t6510) I(R7999t442) I(R8000t927) I(R8000t1658) I(R8000t1239) I(R8001t572) I(R8001t1510) I(R8001t2135) I(R8001t7765) I(R8001t2723) I(R8001t749) I(R8002t693) I(R8002t1446) I(R8002t4010) I(R8002t1143) I(R8002t538) I(R8002t5786) I(R8002t2461) I(R8003t8000) I(R8003t1151) I(R8003t5255) I(R8003t580) I(R8003t1239) I(R8004t513) I(R8004t7789) I(R8004t3925) I(R8004t1511) I(R8004t6631) I(R8005t4995) I(R8005t7034) I(R8005t72) I(R8006t510) I(R8006t1767) I(R8007t55) I(R8007t5274) I(R8007t2102) I(R8007t3286) I(R8007t2453) I(R8007t7842) I(R8008t628) I(R8008t4388) I(R8008t3393) I(R8008t5514) I(R8008t2875) I(R8008t6450) I(R8008t5851) I(R8009t940) I(R8009t5799) I(R8009t452) I(R8009t2853) I(R8009t2445) I(R8010t1859) I(R8010t2588) I(R8010t1522) I(R8010t1754) I(R8011t534) I(R8011t7157) I(R8011t5761) I(R8011t85) I(R8011t3177) I(R8012t4043) I(R8012t4653) I(R8012t660) I(R8012t7401) I(R8012t3454) I(R8013t736) I(R8013t4757) I(R8013t6724) I(R8013t1772) I(R8013t90) I(R8014t1131) I(R8014t1974) I(R8014t3848) I(R8014t2652) I(R8014t2845) I(R8014t4837) I(R8015t1805) I(R8015t5205) I(R8015t653) I(R8016t437) I(R8016t6223) I(R8016t646) I(R8016t7807) I(R8016t7008) I(R8017t177) I(R8017t1042) I(R8017t6007) I(R8017t7239) I(R8017t5642) I(R8017t2977) I(R8017t7110) I(R8018t3347) I(R8018t3907) I(R8018t4987) I(R8019t526) I(R8019t3795) I(R8019t4507) I(R8020t665) I(R8020t1326) I(R8020t482) I(R8020t7136) I(R8020t7249) I(R8020t6357) I(R8021t448) I(R8021t3063) I(R8021t3686) I(R8021t3939) I(R8022t4300) I(R8022t6947) I(R8022t6985) I(R8022t7440) I(R8022t1072) I(R8022t5480) I(R8023t3942) I(R8023t4412) I(R8023t165) I(R8023t308) I(R8023t5983) I(R8024t208) I(R8024t6211) I(R8024t124) I(R8024t1506) I(R8024t2485) I(R8024t7069) I(R8024t2773) I(R8025t281) I(R8025t1200) I(R8025t7273) I(R8025t351) I(R8025t957) I(R8025t4746) I(R8026t7395) I(R8026t6458) I(R8026t4058) I(R8026t3823) I(R8026t99) I(R8027t882) I(R8027t6432) I(R8027t7120) I(R8027t2540) I(R8027t2509) I(R8027t4183) I(R8027t3503) I(R8027t4120) I(R8027t6894) I(R8028t1633) I(R8028t4371) I(R8028t4601) I(R8028t2901) I(R8028t5405) I(R8028t5150) I(R8028t7628) I(R8028t2641) I(R8029t2217) I(R8029t2257) I(R8029t4386) I(R8029t5860) I(R8029t2940) I(R8029t5540) I(R8030t4001) I(R8030t7881) I(R8030t7427) I(R8030t7830) I(R8030t5870) I(R8030t7050) I(R8031t2084) I(R8031t5806) I(R8031t99) I(R8031t3823) I(R8032t7420) I(R8032t7441) I(R8032t949) I(R8032t2006) I(R8032t1984) I(R8033t389) I(R8033t6800) I(R8033t347) I(R8033t2010) I(R8033t7286) I(R8034t5743) I(R8034t6821) I(R8034t1999) I(R8034t5928) I(R8034t2027) I(R8034t536) I(R8035t3928) I(R8035t7838) I(R8035t5524) I(R8035t2958) I(R8035t2673) I(R8035t5153) I(R8036t4391) I(R8036t7329) I(R8037t1707) I(R8037t587) I(R8037t1137) I(R8038t3128) I(R8038t3669) I(R8039t367) I(R8039t7024) I(R8039t6871) I(R8039t7538) I(R8040t1062) I(R8040t3073) I(R8040t1234) I(R8040t6447) I(R8040t4643) I(R8041t5633) I(R8041t5419) I(R8041t3935) I(R8041t6856) I(R8042t636) I(R8042t1396) I(R8042t7618) I(R8042t5290) I(R8042t2853) I(R8042t796) I(R8043t7987) I(R8043t7756) I(R8043t2070) I(R8043t4475) I(R8043t1425) I(R8044t6465) I(R8044t4998) I(R8044t7141) I(R8044t1246) I(R8044t2117) I(R8045t7877) I(R8045t1935) I(R8045t285) I(R8045t1992) I(R8045t40) I(R8046t7083) I(R8046t2353) I(R8046t5694) I(R8046t2905) I(R8047t6265) I(R8047t1261) I(R8047t4840) I(R8047t2909) I(R8047t1735) I(R8048t3592) I(R8048t5889) I(R8048t5569) I(R8048t3782) I(R8048t1255) I(R8048t1913) I(R8048t5222) I(R8049t7092) I(R8049t7308) I(R8049t4347) I(R8050t1345) I(R8050t6050) I(R8050t7448) I(R8050t725) I(R8050t5964) I(R8050t4341) I(R8051t4290) I(R8051t7531) I(R8051t7913) I(R8051t5640) I(R8051t5408) I(R8051t326) I(R8051t1710) I(R8052t547) I(R8052t4105) I(R8052t4191) I(R8052t2456) I(R8052t1393) I(R8053t273) I(R8053t3) I(R8053t7844) I(R8054t723) I(R8055t1334) I(R8055t2544) I(R8055t2781) I(R8055t3002) I(R8055t6503) I(R8056t3279) I(R8056t7022) I(R8056t2411) I(R8056t1731) I(R8056t6327) I(R8056t5608) I(R8057t1147) I(R8057t4125) I(R8057t2736) I(R8057t2960) I(R8057t1682) I(R8058t7832) I(R8058t77) I(R8058t1424) I(R8058t7884) I(R8058t5668) I(R8059t568) I(R8059t3060) I(R8059t319) I(R8059t5148) I(R8059t7907) I(R8060t1708) I(R8060t7222) I(R8060t4034) I(R8060t1419) I(R8060t1626) I(R8061t5115) I(R8061t7832) I(R8061t1689) I(R8061t5277) I(R8061t5832) I(R8062t4866) I(R8062t2288) I(R8062t7078) I(R8062t1609) I(R8063t1816) I(R8063t4753) I(R8063t5275) I(R8064t5863) I(R8064t6952) I(R8064t1262) I(R8064t4176) I(R8064t3410) I(R8065t2555) I(R8065t6688) I(R8066t1125) I(R8066t3053) I(R8066t4187) I(R8066t6056) I(R8066t3172) I(R8066t6858) I(R8066t2470) I(R8066t2031) I(R8067t4050) I(R8067t2146) I(R8067t5017) I(R8067t6714) I(R8067t3684) I(R8067t3016) I(R8067t954) I(R8068t5877) I(R8068t5991) I(R8068t6097) I(R8068t6704) I(R8068t1959) I(R8068t7511) I(R8068t5639) I(R8069t97) I(R8069t7370) I(R8069t2266) I(R8069t7330) I(R8070t3628) I(R8070t1555) I(R8070t4552) I(R8071t7400) I(R8071t5794) I(R8071t7674) I(R8071t5977) I(R8071t4588) I(R8071t2070) I(R8071t6577) I(R8072t339) I(R8072t1739) I(R8072t1933) I(R8072t1834) I(R8072t3828) I(R8073t5652) I(R8073t235) I(R8073t7624) I(R8073t4740) I(R8074t7454) I(R8074t4785) I(R8074t777) I(R8074t7308) I(R8074t8049) I(R8075t1538) I(R8075t5259) I(R8075t6790) I(R8075t668) I(R8076t4109) I(R8076t6361) I(R8076t4429) I(R8076t4863) I(R8076t4544) I(R8077t3193) I(R8077t5821) I(R8077t3126) I(R8077t6390) I(R8077t4578) I(R8078t5378) I(R8078t6948) I(R8078t4886) I(R8078t4611) I(R8078t492) I(R8078t6979) I(R8079t88) I(R8079t4843) I(R8079t5053) I(R8079t1658) I(R8079t4791) I(R8079t1476) I(R8079t3897) I(R8080t6379) I(R8080t7620) I(R8080t881) I(R8080t3082) I(R8080t2314) I(R8081t379) I(R8081t7480) I(R8081t2999) I(R8081t4306) I(R8081t2556) I(R8081t7017) I(R8081t1105) I(R8082t1496) I(R8082t7139) I(R8082t2039) I(R8083t6150) I(R8083t7813) I(R8083t5179) I(R8083t1809) I(R8083t4491) I(R8084t5741) I(R8084t7747) I(R8084t3137) I(R8084t3358) I(R8085t1450) I(R8085t3811) I(R8085t1092) I(R8085t3224) I(R8085t5699) I(R8086t436) I(R8086t6296) I(R8086t3538) I(R8086t2346) I(R8086t117) I(R8086t1180) I(R8086t4808) I(R8087t2779) I(R8087t3374) I(R8087t2086) I(R8087t5534) I(R8088t4260) I(R8088t899) I(R8088t1888) I(R8088t4063) I(R8088t5384) I(R8089t375) I(R8089t6133) I(R8089t686) I(R8089t4477) I(R8089t6727) I(R8090t6769) I(R8090t6530) I(R8090t2849) I(R8090t7347) I(R8090t2013) I(R8090t6813) I(R8091t5313) I(R8091t7209) I(R8091t7441) I(R8091t7420) I(R8091t2352) I(R8092t465) I(R8092t7885) I(R8092t3217) I(R8092t7378) I(R8092t6892) I(R8093t1015) I(R8093t4420) I(R8093t6968) I(R8093t4644) I(R8093t2662) I(R8093t304) I(R8094t1009) I(R8094t7379) I(R8094t3832) I(R8094t5109) I(R8094t2910) I(R8095t3204) I(R8095t7463) I(R8095t2067) I(R8095t5113) I(R8095t1582) I(R8096t97) I(R8096t3886) I(R8097t4139) I(R8097t5994) I(R8097t2606) I(R8098t6106) I(R8098t6981) I(R8098t6812) I(R8099t3562) I(R8099t7066) I(R8099t1230) I(R8099t5747) I(R8099t3518) I(R8100t5791) I(R8100t6795) I(R8100t6091) I(R8100t183) I(R8101t6423) I(R8101t1295) I(R8101t786) I(R8101t6387) I(R8101t5636) I(R8101t3768) I(R8102t1256) I(R8102t4614) I(R8102t3376) I(R8102t5177) I(R8102t1140) I(R8102t678) I(R8102t1645) I(R8102t6642) I(R8103t4107) I(R8103t5684) I(R8103t410) I(R8103t6024) I(R8103t5876) I(R8103t2015) I(R8104t5994) I(R8104t8097) I(R8104t2606) I(R8104t6341) I(R8104t7405) I(R8105t3218) I(R8105t5593) I(R8105t1323) I(R8105t6856) I(R8105t5189) I(R8105t6462) I(R8106t2248) I(R8106t6981) I(R8106t8098) I(R8106t1163) I(R8107t1879) I(R8107t4312) I(R8107t870) I(R8107t3654) I(R8107t7182) I(R8107t1781) I(R8108t1465) I(R8108t4066) I(R8108t3708) I(R8108t682) I(R8108t7531) I(R8109t989) I(R8109t5140) I(R8109t6268) I(R8109t5301) I(R8109t2856) I(R8109t4802) I(R8109t1222) I(R8110t7667) I(R8110t2000) I(R8110t7408) I(R8110t7455) I(R8110t959) I(R8111t128) I(R8111t5181) I(R8111t4881) I(R8111t7482) I(R8112t7565) I(R8112t4210) I(R8112t2486) I(R8112t2703) I(R8113t1687) I(R8113t4436) I(R8113t866) I(R8113t6929) I(R8113t2191) I(R8114t1090) I(R8114t4482) I(R8114t768) I(R8114t2081) I(R8114t1967) I(R8115t4005) I(R8115t4429) I(R8115t8076) I(R8115t4863) I(R8116t1742) I(R8116t2778) I(R8116t6091) I(R8116t8100) I(R8116t6795) I(R8116t1317) I(R8116t4093) I(R8116t6578) I(R8117t655) I(R8117t1675) I(R8117t7987) I(R8117t3326) I(R8117t6543) I(R8117t6313) I(R8118t3139) I(R8118t7508) I(R8118t4867) I(R8118t6525) I(R8118t6961) I(R8119t1032) I(R8119t3161) I(R8119t3703) I(R8119t2416) I(R8119t5210) I(R8119t3633) I(R8119t3882) I(R8119t4365) I(R8120t5996) I(R8120t7932) I(R8120t666) I(R8120t850) I(R8121t1182) I(R8121t2302) I(R8121t6305) I(R8121t7187) I(R8121t4271) I(R8121t1886) I(R8121t7121) I(R8122t7929) I(R8122t1403) I(R8122t2443) I(R8122t2991) I(R8122t2400) I(R8123t353) I(R8123t2890) I(R8123t2426) I(R8123t7007) I(R8123t3690) I(R8123t3042) I(R8124t1093) I(R8124t3244) I(R8124t4577) I(R8124t6376) I(R8125t7278) I(R8125t6708) I(R8125t419) I(R8125t7134) I(R8125t7311) I(R8125t7340) I(R8126t1913) I(R8126t8048) I(R8126t3377) I(R8126t2987) I(R8126t7096) I(R8126t1255) I(R8127t467) I(R8127t3856) I(R8127t6650) I(R8127t7735) I(R8127t7547) I(R8127t1198) I(R8128t6309) I(R8128t7386) I(R8128t6095) I(R8128t6362) I(R8129t505) I(R8129t539) I(R8129t2169) I(R8129t5104) I(R8129t4080) I(R8129t1842) I(R8129t3843) I(R8130t1463) I(R8130t4825) I(R8130t7109) I(R8130t2001) I(R8131t5683) I(R8131t6634) I(R8131t1501) I(R8131t3030) I(R8131t5908) I(R8132t2843) I(R8132t7752) I(R8132t3369) I(R8132t853) I(R8132t6840) I(R8133t1156) I(R8133t4488) I(R8133t6725) I(R8134t5812) I(R8134t7211) I(R8134t7074) I(R8134t7580) I(R8134t4902) I(R8135t989) I(R8135t5140) I(R8135t6268) I(R8135t3225) I(R8135t1924) I(R8136t2648) I(R8136t7359) I(R8136t3448) I(R8136t4523) I(R8136t5662) I(R8137t1707) I(R8137t8037) I(R8137t3913) I(R8137t3908) I(R8137t4706) I(R8137t1137) I(R8138t1871) I(R8138t7719) I(R8138t1405) I(R8138t6261) I(R8139t331) I(R8139t582) I(R8139t75) I(R8139t6413) I(R8140t2985) I(R8140t5444) I(R8140t7269) I(R8140t2005) I(R8140t1086) I(R8141t478) I(R8141t7045) I(R8141t2213) I(R8141t1053) I(R8142t6240) I(R8142t7878) I(R8142t4756) I(R8142t3544) I(R8142t5258) I(R8143t4620) I(R8143t7928) I(R8143t2829) I(R8143t4671) I(R8144t2182) I(R8144t2235) I(R8144t3147) I(R8144t1054) I(R8144t4835) I(R8145t1534) I(R8145t7495) I(R8145t3205) I(R8145t3316) I(R8146t7624) I(R8146t4740) I(R8146t4782) I(R8146t1651) I(R8146t440) I(R8147t2374) I(R8147t7234) I(R8147t6746) I(R8147t7802) I(R8147t6993) I(R8147t43) I(R8147t4574) I(R8148t3379) I(R8148t5394) I(R8148t1885) I(R8148t5769) I(R8149t7216) I(R8149t7543) I(R8149t5921) I(R8149t6255) I(R8149t7855) I(R8150t1072) I(R8150t8022) I(R8150t16) I(R8150t3371) I(R8150t3278) I(R8150t7440) I(R8151t2555) I(R8151t4473) I(R8151t3852) I(R8151t8065) I(R8152t1939) I(R8152t5305) I(R8152t2873) I(R8152t127) I(R8152t2462) I(R8152t5426) I(R8152t7182) I(R8152t8107) I(R8152t3654) I(R8153t129) I(R8153t4680) I(R8153t4003) I(R8153t5166) I(R8154t6694) I(R8154t7921) I(R8154t6273) I(R8154t3536) I(R8154t6729) I(R8154t7373) I(R8155t578) I(R8155t707) I(R8155t967) I(R8155t7609) I(R8156t1507) I(R8156t4732) I(R8156t3465) I(R8156t2713) I(R8156t6606) I(R8157t4216) I(R8157t7219) I(R8157t562) I(R8157t7201) I(R8158t3776) I(R8158t6647) I(R8158t6902) I(R8159t1133) I(R8159t7221) I(R8159t3881) I(R8159t2487) I(R8159t5660) I(R8159t7534) I(R8160t1531) I(R8160t7377) I(R8160t6661) I(R8160t2323) I(R8160t6164) I(R8161t3272) I(R8161t3838) I(R8161t1009) I(R8161t1632) I(R8161t2350) I(R8161t7) I(R8161t3490) I(R8162t5073) I(R8162t6076) I(R8162t5887) I(R8162t3239) I(R8163t604) I(R8163t7201) I(R8163t8157) I(R8163t562) I(R8163t937) I(R8163t7067) I(R8164t1005) I(R8164t5394) I(R8164t7501) I(R8164t7974) I(R8164t1785) I(R8165t3549) I(R8165t3122) I(R8165t4689) I(R8166t2633) I(R8166t7776) I(R8166t6868) I(R8166t4047) I(R8167t722) I(R8167t2305) I(R8168t1660) I(R8168t7569) I(R8168t5674) I(R8168t2018) I(R8168t6901) I(R8169t3499) I(R8169t3810) I(R8169t1802) I(R8169t1932) I(R8169t3598) I(R8169t7980) I(R8170t44) I(R8170t5818) I(R8170t7914) I(R8170t6998) I(R8171t3046) I(R8171t5342) I(R8171t3815) I(R8171t3761) I(R8172t8098) I(R8172t8106) I(R8172t1163) I(R8172t2306) I(R8172t5152) I(R8172t7602) I(R8172t1748) I(R8172t6812) I(R8173t6409) I(R8173t4479) I(R8173t4508) I(R8173t615) I(R8174t381) I(R8174t4968) I(R8174t5816) I(R8174t157) I(R8174t6767) I(R8175t270) I(R8175t1089) I(R8175t7038) I(R8175t4033) I(R8175t5443) I(R8176t6072) I(R8176t7586) I(R8176t1266) I(R8176t7617) I(R8176t6301) I(R8176t597) I(R8177t1725) I(R8177t3785) I(R8177t1700) I(R8177t1840) I(R8177t82) I(R8178t2451) I(R8178t6976) I(R8178t3306) I(R8178t7507) I(R8178t7683) I(R8179t10) I(R8179t489) I(R8179t5250) I(R8179t6825) I(R8179t4152) I(R8179t2524) I(R8180t5953) I(R8180t6781) I(R8180t5859) I(R8180t2886) I(R8180t7277) I(R8180t3675) I(R8181t5083) I(R8181t5491) I(R8181t1934) I(R8181t6356) I(R8181t3210) I(R8181t2220) I(R8181t570) I(R8182t1193) I(R8182t5657) I(R8182t3420) I(R8182t6516) I(R8183t1624) I(R8183t5052) I(R8183t2854) I(R8183t7519) I(R8183t5881) I(R8184t2829) I(R8184t4589) I(R8184t7928) I(R8184t7196) I(R8185t5192) I(R8185t6124) I(R8185t2885) I(R8186t4653) I(R8186t6937) I(R8186t5198) I(R8186t2349) I(R8187t1779) I(R8187t6966) I(R8187t2095) I(R8187t2767) I(R8187t5951) I(R8187t2727) I(R8188t5057) I(R8188t3766) I(R8188t6140) I(R8188t5240) I(R8189t3440) I(R8189t4908) I(R8189t789) I(R8189t3673) I(R8189t6659) I(R8190t59) I(R8190t6261) I(R8190t6087) I(R8190t67) I(R8190t5811) I(R8190t2452) I(R8191t927) I(R8191t1658) I(R8191t8079) I(R8191t5053) I(R8191t7497) I(R8191t288) I(R8192t1398) I(R8192t7170) I(R8192t3374) I(R8192t4516) I(R8193t5477) I(R8193t4058) I(R8193t3159) I(R8193t5906) I(R8193t3180) I(R8194t4094) I(R8194t5915) I(R8194t5039) I(R8194t531) I(R8194t941) I(R8195t394) I(R8195t4092) I(R8195t2054) I(R8195t1293) I(R8195t7849) I(R8195t1743) I(R8195t3022) I(R8196t4193) I(R8196t4236) I(R8196t2471) I(R8197t8142) I(R8197t7027) I(R8197t7473) I(R8197t830) I(R8197t5258) I(R8198t5366) I(R8198t6869) I(R8198t7477) I(R8198t2738) I(R8198t4157) I(R8198t5048) I(R8199t578) I(R8199t8155) I(R8199t707) I(R8199t6262) I(R8199t1879) I(R8200t1931) I(R8200t4733) I(R8200t4115) I(R8201t4802) I(R8201t1222) I(R8201t5884) I(R8201t2763) I(R8201t2632) I(R8201t4206) I(R8202t6597) I(R8202t5285) I(R8202t2180) I(R8202t5754) I(R8202t5996) I(R8202t8120) I(R8203t1854) I(R8203t6186) I(R8203t6596) I(R8203t3230) I(R8203t6909) I(R8203t7258) I(R8204t114) I(R8204t1931) I(R8204t3734) I(R8204t918) I(R8204t4115) I(R8204t8200) I(R8205t5457) I(R8205t5836) I(R8205t24) I(R8205t6571) I(R8205t135) I(R8206t3000) I(R8206t3560) I(R8206t831) I(R8206t7318) I(R8206t4366) I(R8206t5069) I(R8206t6272) I(R8206t3526) I(R8207t5509) I(R8207t6963) I(R8207t8054) I(R8207t723) I(R8207t3835) I(R8207t6020) I(R8208t298) I(R8208t6418) I(R8208t2824) I(R8208t159) I(R8208t4738) I(R8208t6824) I(R8209t548) I(R8209t5080) I(R8209t2843) I(R8209t5458) I(R8209t6408) I(R8210t2135) I(R8210t8001) I(R8210t7765) I(R8210t7129) I(R8210t1257) I(R8210t2910) I(R8211t608) I(R8211t2865) I(R8211t6831) I(R8211t3092) I(R8212t598) I(R8212t5174) I(R8212t7784) I(R8212t635) I(R8213t899) I(R8213t6418) I(R8213t2824) I(R8213t2313) I(R8213t3140) I(R8214t2252) I(R8214t6744) I(R8214t6017) I(R8214t3273) I(R8214t7391) I(R8215t6597) I(R8215t8202) I(R8215t7612) I(R8215t7486) I(R8215t2504) I(R8216t2676) I(R8216t6377) I(R8216t240) I(R8217t6934) I(R8217t7942) I(R8217t5359) I(R8217t3572) I(R8218t3147) I(R8218t8144) I(R8218t7778) I(R8218t3826) I(R8218t2235) I(R8219t4261) I(R8219t5563) I(R8219t3557) I(R8220t6000) I(R8220t6476) I(R8220t6605) I(R8220t7324) I(R8220t914) I(R8220t6525) I(R8221t4174) I(R8221t7370) I(R8221t7866) I(R8221t2677) I(R8221t3758) I(R8222t2033) I(R8222t5607) I(R8222t2870) I(R8222t2142) I(R8222t5549) I(R8222t1962) I(R8223t5106) I(R8223t5470) I(R8223t775) I(R8223t7156) I(R8224t4345) I(R8224t2357) I(R8224t1467) I(R8224t1002) I(R8225t4232) I(R8225t478) I(R8225t8141) I(R8226t1376) I(R8226t4919) I(R8226t2859) I(R8226t4480) I(R8226t5613) I(R8226t6174) I(R8227t3810) I(R8227t7992) I(R8227t4846) I(R8227t5621) I(R8227t7585) I(R8228t374) I(R8228t6818) I(R8228t2490) I(R8228t5343) I(R8228t7818) I(R8228t6501) I(R8229t6265) I(R8229t5926) I(R8229t7535) I(R8229t1735) I(R8230t5271) I(R8230t1421) I(R8230t5163) I(R8230t761) I(R8230t3006) I(R8231t3202) I(R8231t7433) I(R8231t4045) I(R8231t6984) I(R8231t4301) I(R8232t1230) I(R8232t3562) I(R8232t8099) I(R8233t3121) I(R8233t6350) I(R8233t6670) I(R8233t7770) I(R8233t5971) I(R8233t5979) I(R8234t2987) I(R8234t3377) I(R8234t8126) I(R8235t2815) I(R8235t6598) I(R8235t2580) I(R8235t345) I(R8235t1288) I(R8236t5633) I(R8236t8041) I(R8236t5292) I(R8236t7846) I(R8236t2904) I(R8236t6856) I(R8237t3183) I(R8237t7990) I(R8237t2317) I(R8237t6962) I(R8237t6794) I(R8237t1219) I(R8238t6738) I(R8238t27) I(R8238t5036) I(R8239t6018) I(R8239t3338) I(R8239t7798) I(R8239t3867) I(R8240t544) I(R8240t7588) I(R8240t2888) I(R8240t7371) I(R8240t4630) I(R8240t7102) I(R8241t2787) I(R8241t7739) I(R8241t825) I(R8241t3369) I(R8241t7752) I(R8241t3138) I(R8241t7180) I(R8242t2008) I(R8242t7106) I(R8242t5744) I(R8242t6515) I(R8242t6061) I(R8243t3110) I(R8243t7658) I(R8243t2534) I(R8243t103) I(R8243t5865) I(R8243t3714) I(R8244t5352) I(R8244t5898) I(R8244t5070) I(R8244t5838) I(R8244t7145) I(R8244t1156) I(R8244t8133) I(R8244t6725) I(R8245t352) I(R8245t1301) I(R8245t1476) I(R8245t3926) I(R8245t3897) I(R8245t7794) I(R8245t5897) I(R8246t6336) I(R8246t7845) I(R8246t6126) I(R8246t560) I(R8246t6764) I(R8247t3243) I(R8247t4899) I(R8247t2716) I(R8247t431) I(R8248t857) I(R8248t6737) I(R8248t3785) I(R8248t737) I(R8248t969) I(R8248t2447) I(R8248t5121) I(R8248t5536) I(R8248t1231) I(R8249t5770) I(R8249t7556) I(R8249t1690) I(R8249t7599) I(R8249t150) I(R8250t7461) I(R8250t710) I(R8250t4687) I(R8250t150) I(R8250t7599) I(R8250t3446) I(R8251t4819) I(R8251t7064) I(R8251t1587) I(R8251t1981) I(R8252t209) I(R8252t843) I(R8252t2986) I(R8253t6425) I(R8253t5414) I(R8253t1747) I(R8253t3615) I(R8254t1178) I(R8254t4195) I(R8254t1227) I(R8254t2074) I(R8255t5212) I(R8255t5669) I(R8255t1711) I(R8255t3922) I(R8255t672) I(R8256t6877) I(R8256t7461) I(R8256t1226) I(R8256t705) I(R8256t3964) I(R8256t5628) I(R8257t6910) I(R8257t7818) I(R8257t7312) I(R8257t913) I(R8257t5114) I(R8257t6501) I(R8258t2649) I(R8258t7695) I(R8258t684) I(R8259t4053) I(R8259t5403) I(R8259t841) I(R8259t2368) I(R8259t6633) I(R8259t5592) I(R8260t3242) I(R8260t4566) I(R8260t7374) I(R8260t4390) I(R8261t2025) I(R8261t6354) I(R8261t6963) I(R8261t8054) I(R8262t3517) I(R8262t4463) I(R8262t75) I(R8262t582) I(R8262t6800) I(R8262t7286) I(R8262t563) I(R8262t3763) I(R8262t1984) I(R8263t3543) I(R8263t4820) I(R8263t1558) I(R8263t265) I(R8263t6218) I(R8263t3375) I(R8264t7892) I(R8264t4396) I(R8264t6782) I(R8264t7539) I(R8265t290) I(R8265t1164) I(R8265t6730) I(R8266t2110) I(R8266t7504) I(R8266t5827) I(R8266t215) I(R8266t1780) I(R8266t4145) I(R8266t3752) I(R8266t1246) I(R8267t1955) I(R8267t5062) I(R8267t5216) I(R8267t3126) I(R8267t2431) I(R8267t7994) I(R8268t5088) I(R8268t6991) I(R8268t1057) I(R8269t1956) I(R8269t7742) I(R8269t4186) I(R8269t6021) I(R8269t5685) I(R8269t858) I(R8269t2409) I(R8270t4145) I(R8270t4536) I(R8270t3509) I(R8270t5100) I(R8270t3752) I(R8270t8266) I(R8271t3630) I(R8271t3486) I(R8271t5120) I(R8272t2784) I(R8272t3873) I(R8272t4005) I(R8272t4429) I(R8272t1619) I(R8272t4150) I(R8272t5372) I(R8273t2280) I(R8273t2109) I(R8273t7411) I(R8273t5067) I(R8274t301) I(R8274t7595) I(R8274t6901) I(R8274t706) I(R8274t7416) I(R8275t7290) I(R8275t4143) I(R8275t7953) I(R8275t996) I(R8276t4745) I(R8276t5834) I(R8276t6526) I(R8276t6748) I(R8276t6162) I(R8276t6941) I(R8276t2059) I(R8277t482) I(R8277t8020) I(R8277t7136) I(R8277t5880) I(R8277t6411) I(R8278t1678) I(R8278t3979) I(R8278t6248) I(R8279t3754) I(R8279t2711) I(R8279t1162) I(R8279t3194) I(R8279t5776) I(R8280t4184) I(R8280t6710) I(R8280t7575) I(R8280t3191) I(R8281t2894) I(R8281t7715) I(R8281t6293) I(R8282t109) I(R8282t2423) I(R8282t4069) I(R8282t4986) I(R8282t7277) I(R8282t3675) I(R8283t4387) I(R8283t7951) I(R8283t7684) I(R8283t1959) I(R8283t8068) I(R8283t7511) I(R8283t2635) I(R8284t7146) I(R8284t7492) I(R8284t672) I(R8284t3922) I(R8284t5820) I(R8285t7905) I(R8285t3385) I(R8286t3257) I(R8286t1152) I(R8286t6673) I(R8287t864) I(R8287t7059) I(R8287t7795) I(R8287t5808) I(R8287t4978) I(R8287t2251) I(R8287t284) I(R8288t1021) I(R8288t1192) I(R8288t4983) I(R8288t5339) I(R8288t4086) I(R8289t2875) I(R8289t5514) I(R8289t629) I(R8289t4585) I(R8290t1548) I(R8290t7992) I(R8290t6441) I(R8290t4497) I(R8290t5350) I(R8291t4586) I(R8291t7307) I(R8291t1774) I(R8291t1637) I(R8291t1200) I(R8291t2708) I(R8292t2815) I(R8292t3974) I(R8292t5051) I(R8292t698) I(R8293t6228) I(R8293t6835) I(R8293t2618) I(R8294t1339) I(R8294t7223) I(R8294t27) I(R8294t8238) I(R8294t2839) I(R8295t1148) I(R8295t4705) I(R8295t6512) I(R8295t5439) I(R8295t6924) I(R8295t3971) I(R8295t720) I(R8295t2111) I(R8296t2382) I(R8296t7981) I(R8296t2068) I(R8296t1303) I(R8296t2219) I(R8297t1778) I(R8297t7410) I(R8298t588) I(R8298t2490) I(R8298t7447) I(R8298t7489) I(R8298t4672) I(R8298t4667) I(R8299t1652) I(R8299t4220) I(R8299t4792) I(R8299t2570) I(R8300t6086) I(R8300t2617) I(R8300t3915) I(R8300t3975) I(R8300t6505) I(R8301t2590) I(R8301t1058) I(R8301t5050) I(R8301t5903) I(R8302t6301) I(R8302t6638) I(R8302t8176) I(R8302t597) I(R8302t3581) I(R8302t5507) I(R8303t578) I(R8303t6618) I(R8303t8155) I(R8303t7609) I(R8304t2668) I(R8304t6370) I(R8304t405) I(R8304t7792) I(R8304t1065) I(R8304t4920) I(R8305t5125) I(R8305t6198) I(R8305t6399) I(R8305t307) I(R8306t3350) I(R8306t4182) I(R8306t5612) I(R8306t3996) I(R8306t7179) I(R8307t1050) I(R8307t4270) I(R8307t2658) I(R8307t5520) I(R8307t4903) I(R8308t2436) I(R8308t6034) I(R8308t6482) I(R8308t5157) I(R8309t2486) I(R8309t4210) I(R8309t5067) I(R8309t8273) I(R8309t2280) I(R8310t4132) I(R8310t4389) I(R8310t3162) I(R8310t2004) I(R8310t1429) I(R8310t7451) I(R8311t1067) I(R8311t3753) I(R8311t7598) I(R8311t2484) I(R8311t6026) I(R8312t4117) I(R8312t7218) I(R8312t4279) I(R8312t5021) I(R8312t2806) I(R8312t2193) I(R8312t6522) I(R8313t8297) I(R8313t937) I(R8313t562) I(R8313t3941) I(R8313t7410) I(R8314t6260) I(R8314t7627) I(R8314t122) I(R8314t3794) I(R8315t784) I(R8315t2922) I(R8315t4134) I(R8315t146) I(R8315t3762) I(R8316t1761) I(R8316t7880) I(R8316t7996) I(R8316t5891) I(R8316t6953) I(R8317t6302) I(R8317t2339) I(R8317t1119) I(R8318t383) I(R8318t558) I(R8318t5774) I(R8318t6276) I(R8319t931) I(R8319t7404) I(R8319t135) I(R8319t6571) I(R8319t3548) I(R8319t5459) I(R8320t3307) I(R8320t7175) I(R8320t1717) I(R8320t4230) I(R8320t4207) I(R8320t453) I(R8321t6268) I(R8321t8135) I(R8321t7766) I(R8322t1300) I(R8322t6322) I(R8322t1409) I(R8322t1443) I(R8322t1210) I(R8323t1163) I(R8323t2248) I(R8323t2335) I(R8323t2683) I(R8323t5925) I(R8323t6026) I(R8324t1014) I(R8324t5118) I(R8324t7973) I(R8324t2064) I(R8325t2390) I(R8325t556) I(R8325t7439) I(R8325t3539) I(R8325t4980) I(R8325t7423) I(R8325t6956) I(R8326t8175) I(R8326t3631) I(R8326t5328) I(R8326t2920) I(R8326t5443) I(R8327t6406) I(R8327t7036) I(R8327t2226) I(R8327t7518) I(R8327t2591) I(R8327t4768) I(R8327t3923) I(R8328t6089) I(R8328t7123) I(R8329t3880) I(R8329t4500) I(R8329t3862) I(R8329t6719) I(R8329t4125) I(R8330t202) I(R8330t2986) I(R8330t8252) I(R8331t1742) I(R8331t2778) I(R8331t1224) I(R8332t936) I(R8332t4348) I(R8332t1882) I(R8332t5864) I(R8332t2761) I(R8332t4254) I(R8333t2898) I(R8333t3190) I(R8333t6659) I(R8333t2329) I(R8333t7443) I(R8333t3626) I(R8333t3174) I(R8333t342) I(R8334t6518) I(R8334t7943) I(R8334t2780) I(R8334t2844) I(R8334t3297) I(R8334t7139) I(R8335t3156) I(R8336t5604) I(R8336t6959) I(R8336t7372) I(R8336t2696) I(R8336t450) I(R8336t5035) I(R8336t6343) I(R8337t1816) I(R8337t6436) I(R8337t1660) I(R8337t7569) I(R8337t8063) I(R8338t352) I(R8338t1301) I(R8338t8018) I(R8338t3907) I(R8338t2917) I(R8338t3265) I(R8338t4631) I(R8339t7321) I(R8339t439) I(R8340t3046) I(R8340t5749) I(R8340t452) I(R8340t5290) I(R8340t5342) I(R8340t8171) I(R8341t693) I(R8341t4010) I(R8341t1023) I(R8341t965) I(R8341t3962) I(R8341t4620) I(R8341t8143) I(R8341t659) I(R8342t4557) I(R8342t6092) I(R8342t1384) I(R8342t2085) I(R8342t6097) I(R8343t5832) I(R8343t7207) I(R8343t7819) I(R8343t7205) I(R8343t1030) I(R8343t1433) I(R8344t2663) I(R8344t6657) I(R8344t2326) I(R8344t4518) I(R8344t4119) I(R8344t1004) I(R8345t6699) I(R8345t6763) I(R8345t3358) I(R8345t37) I(R8346t1045) I(R8346t7246) I(R8346t7323) I(R8346t7383) I(R8346t2295) I(R8347t5376) I(R8347t1333) I(R8347t2759) I(R8347t6266) I(R8347t3051) I(R8348t6479) I(R8348t6535) I(R8348t5943) I(R8348t2372) I(R8348t1359) I(R8349t825) I(R8349t7815) I(R8349t7739) I(R8349t5382) I(R8350t7325) I(R8350t1187) I(R8350t5656) I(R8350t6379) I(R8350t6511) I(R8351t2969) I(R8351t4143) I(R8351t4857) I(R8351t5418) I(R8352t618) I(R8352t3372) I(R8352t2014) I(R8352t6876) I(R8352t1653) I(R8352t7931) I(R8353t936) I(R8353t2445) I(R8353t1882) I(R8353t5864) I(R8353t5775) I(R8353t4062) I(R8353t8009) I(R8354t6699) I(R8354t6923) I(R8354t2511) I(R8354t6763) I(R8354t8345) I(R8355t7156) I(R8355t7215) I(R8355t3624) I(R8355t5784) I(R8355t134) I(R8356t3669) I(R8356t8038) I(R8356t6883) I(R8356t198) I(R8356t4779) I(R8357t5345) I(R8357t4890) I(R8357t4771) I(R8358t1321) I(R8358t4209) I(R8358t7360) I(R8358t5099) I(R8358t5732) I(R8358t3630) I(R8358t8271) I(R8359t970) I(R8359t5535) I(R8359t2455) I(R8359t6498) I(R8359t4418) I(R8359t4243) I(R8359t5843) I(R8359t5923) I(R8360t4299) I(R8360t4661) I(R8360t1358) I(R8360t2837) I(R8360t1280) I(R8360t6397) I(R8361t160) I(R8361t6362) I(R8361t8128) I(R8361t6095) I(R8361t2495) I(R8361t3293) I(R8361t4617) I(R8362t4807) I(R8362t7710) I(R8362t3989) I(R8362t3236) I(R8362t4975) I(R8362t1322) I(R8363t4003) I(R8363t8153) I(R8363t4680) I(R8363t2851) I(R8363t1777) I(R8363t176) I(R8364t1391) I(R8364t7983) I(R8364t6599) I(R8364t7064) I(R8364t3136) I(R8364t7890) I(R8365t1141) I(R8365t7989) I(R8365t694) I(R8365t6705) I(R8365t6508) I(R8365t1820) I(R8366t1946) I(R8366t7784) I(R8366t2640) I(R8367t1145) I(R8367t4332) I(R8367t4363) I(R8367t6413) I(R8367t8139) I(R8368t3391) I(R8368t5773) I(R8369t1679) I(R8369t7128) I(R8369t2367) I(R8370t2604) I(R8370t2744) I(R8370t141) I(R8370t3649) I(R8370t6842) I(R8370t3432) I(R8370t3260) I(R8371t233) I(R8371t2155) I(R8371t3242) I(R8372t7152) I(R8372t4637) I(R8372t7095) I(R8373t1363) I(R8373t4819) I(R8373t1587) I(R8373t7523) I(R8373t5702) I(R8373t567) I(R8373t5914) I(R8373t3248) I(R8374t1080) I(R8374t3007) I(R8374t4928) I(R8374t3063) I(R8374t7282) I(R8375t3283) I(R8375t4927) I(R8375t6019) I(R8375t2622) I(R8375t1139) I(R8376t4496) I(R8376t7627) I(R8376t3736) I(R8376t5011) I(R8377t499) I(R8377t2274) I(R8377t2230) I(R8377t6254) I(R8377t4826) I(R8377t1702) I(R8378t6134) I(R8378t4075) I(R8378t3120) I(R8378t2909) I(R8378t4313) I(R8378t7047) I(R8378t1770) I(R8379t6829) I(R8379t7430) I(R8379t1120) I(R8380t5175) I(R8380t3485) I(R8380t7678) I(R8380t4740) I(R8380t2958) I(R8380t4335) I(R8381t1296) I(R8381t4489) I(R8381t4114) I(R8381t1144) I(R8381t136) I(R8381t6524) I(R8381t5235) I(R8382t1647) I(R8382t7716) I(R8382t3051) I(R8382t8347) I(R8382t6266) I(R8383t5536) I(R8383t6449) I(R8383t5121) I(R8384t4506) I(R8384t7831) I(R8384t2515) I(R8385t3431) I(R8385t3884) I(R8385t2386) I(R8385t434) I(R8385t7647) I(R8385t4204) I(R8385t5161) I(R8385t5159) I(R8386t8074) I(R8386t3768) I(R8387t6074) I(R8387t7552) I(R8387t5056) I(R8387t6531) I(R8387t1471) I(R8387t6134) I(R8387t5201) I(R8387t1469) I(R8388t2832) I(R8388t6614) I(R8388t2775) I(R8388t5955) I(R8388t6590) I(R8389t299) I(R8389t7731) I(R8389t1193) I(R8389t4727) I(R8390t5857) I(R8390t3690) I(R8390t142) I(R8391t3243) I(R8391t4899) I(R8391t1012) I(R8391t3733) I(R8391t422) I(R8391t7350) I(R8392t6858) I(R8392t5878) I(R8392t3779) I(R8393t5419) I(R8393t1228) I(R8393t4747) I(R8394t5553) I(R8394t7868) I(R8394t572) I(R8394t5930) I(R8394t4337) I(R8394t6118) I(R8395t4274) I(R8395t6288) I(R8395t7958) I(R8396t7070) I(R8396t7024) I(R8396t8039) I(R8396t6871) I(R8396t1998) I(R8397t3273) I(R8397t8214) I(R8397t4492) I(R8397t7629) I(R8397t2242) I(R8398t2704) I(R8398t6287) I(R8398t458) I(R8398t3658) I(R8398t2885) I(R8399t6401) I(R8399t6450) I(R8399t8008) I(R8399t2875) I(R8399t7745) I(R8400t6963) I(R8400t8261) I(R8400t8207) I(R8400t8054) I(R8401t3661) I(R8401t5481) I(R8401t6301) I(R8401t6638) I(R8402t3621) I(R8402t4039) I(R8402t6443) I(R8403t5554) I(R8403t1941) I(R8403t4329) I(R8404t5197) I(R8404t6310) I(R8404t2035) I(R8404t7057) I(R8404t1923) I(R8404t3385) I(R8404t4635) I(R8405t63) I(R8405t6936) I(R8405t1499) I(R8405t1176) I(R8405t2177) I(R8406t917) I(R8406t3673) I(R8406t4581) I(R8406t2329) I(R8406t6659) I(R8407t1678) I(R8407t8278) I(R8407t6248) I(R8407t5640) I(R8407t7913) I(R8407t6722) I(R8408t466) I(R8408t5765) I(R8408t1393) I(R8408t2456) I(R8409t137) I(R8409t6942) I(R8409t4628) I(R8409t7257) I(R8410t1285) I(R8410t6426) I(R8410t7461) I(R8410t8250) I(R8410t3446) I(R8411t2835) I(R8411t2575) I(R8411t4147) I(R8411t3903) I(R8412t3085) I(R8412t2592) I(R8412t953) I(R8412t7076) I(R8412t2259) I(R8413t5928) I(R8413t6438) I(R8413t8034) I(R8413t1999) I(R8413t1214) I(R8414t1871) I(R8414t8138) I(R8414t6261) I(R8414t2452) I(R8414t6919) I(R8414t238) I(R8414t1101) I(R8415t4964) I(R8415t7116) I(R8415t1478) I(R8415t1850) I(R8415t3807) I(R8415t6210) I(R8416t4117) I(R8416t8312) I(R8416t6522) I(R8416t1561) I(R8417t5325) I(R8417t3106) I(R8417t3009) I(R8417t4416) I(R8418t31) I(R8418t3915) I(R8418t2098) I(R8418t271) I(R8418t580) I(R8418t589) I(R8419t2527) I(R8419t3925) I(R8419t1511) I(R8419t4133) I(R8419t2681) I(R8419t5727) I(R8419t5212) I(R8420t6207) I(R8420t5837) I(R8420t5495) I(R8420t4511) I(R8420t1720) I(R8421t1987) I(R8421t6461) I(R8421t2445) I(R8421t940) I(R8421t5799) I(R8421t7993) I(R8422t5169) I(R8422t5756) I(R8422t7215) I(R8422t7156) I(R8422t8223) I(R8422t5106) I(R8422t5410) I(R8423t555) I(R8423t6086) I(R8423t5236) I(R8423t3397) I(R8423t2617) I(R8423t8300) I(R8424t6420) I(R8424t8061) I(R8424t5115) I(R8424t2161) I(R8424t1311) I(R8425t4126) I(R8425t7345) I(R8425t1431) I(R8425t4248) I(R8425t5972) I(R8426t1005) I(R8426t1785) I(R8426t2950) I(R8426t321) I(R8426t319) I(R8427t7662) I(R8427t2063) I(R8427t3638) I(R8427t5455) I(R8427t6368) I(R8427t2395) I(R8428t542) I(R8428t1081) I(R8428t5239) I(R8428t3422) I(R8428t7137) I(R8428t3415) I(R8429t5561) I(R8429t1851) I(R8429t3650) I(R8429t4956) I(R8429t3596) I(R8429t5131) I(R8430t3279) I(R8430t5465) I(R8430t2399) I(R8430t5093) I(R8431t6194) I(R8431t7841) I(R8431t6449) I(R8431t1382) I(R8431t808) I(R8432t2004) I(R8432t8310) I(R8432t3011) I(R8432t471) I(R8432t3162) I(R8433t7950) I(R8433t4442) I(R8433t54) I(R8434t1972) I(R8434t2136) I(R8434t2208) I(R8434t5762) I(R8434t901) I(R8434t3254) I(R8434t3251) I(R8435t2754) I(R8435t3655) I(R8435t5574) I(R8435t7349) I(R8435t2163) I(R8436t2277) I(R8436t6903) I(R8436t7727) I(R8436t893) I(R8436t7209) I(R8436t5313) I(R8437t192) I(R8437t3570) I(R8437t6950) I(R8437t5057) I(R8437t8188) I(R8437t5240) I(R8437t3139) I(R8437t6961) I(R8438t7077) I(R8438t5285) I(R8438t8202) I(R8439t5753) I(R8439t6337) I(R8439t7350) I(R8439t3015) I(R8439t5733) I(R8440t1117) I(R8440t7471) I(R8440t6874) I(R8440t2246) I(R8440t7570) I(R8440t7764) I(R8440t5427) I(R8441t4535) I(R8441t1474) I(R8441t6276) I(R8441t8318) I(R8441t5774) I(R8442t964) I(R8442t1836) I(R8442t3216) I(R8442t7230) I(R8442t5976) I(R8443t6930) I(R8443t760) I(R8443t6900) I(R8443t2695) I(R8443t2317) I(R8443t6962) I(R8443t5797) I(R8443t974) I(R8444t1) I(R8444t6319) I(R8444t7938) I(R8444t5602) I(R8444t3796) I(R8444t1650) I(R8445t5354) I(R8445t218) I(R8445t7247) I(R8446t1547) I(R8446t6671) I(R8446t6262) I(R8447t1016) I(R8447t2725) I(R8447t3489) I(R8447t4549) I(R8447t6299) I(R8448t4724) I(R8448t5995) I(R8448t2173) I(R8449t1632) I(R8449t5949) I(R8449t2769) I(R8449t8094) I(R8449t1009) I(R8449t8161) I(R8450t5650) I(R8450t6858) I(R8450t8392) I(R8450t3779) I(R8450t1580) I(R8451t2680) I(R8451t5669) I(R8451t3373) I(R8451t3036) I(R8451t1158) I(R8451t12) I(R8452t2990) I(R8452t5020) I(R8452t5063) I(R8452t7709) I(R8452t1399) I(R8453t2037) I(R8453t2171) I(R8453t2577) I(R8453t1662) I(R8453t3042) I(R8453t3685) I(R8454t2224) I(R8454t2065) I(R8454t3019) I(R8454t4490) I(R8454t612) I(R8454t6274) I(R8454t2079) I(R8455t812) I(R8455t2332) I(R8455t1693) I(R8455t7585) I(R8455t5621) I(R8456t2939) I(R8456t1256) I(R8456t3376) I(R8456t2945) I(R8457t2411) I(R8457t6576) I(R8457t2746) I(R8457t3662) I(R8457t359) I(R8457t2880) I(R8457t5031) I(R8457t4282) I(R8457t3921) I(R8458t7459) I(R8458t7817) I(R8458t4684) I(R8458t3100) I(R8458t2353) I(R8458t5694) I(R8458t6459) I(R8459t2188) I(R8459t3652) I(R8459t7435) I(R8459t3953) I(R8460t50) I(R8460t4421) I(R8460t4386) I(R8460t7706) I(R8460t5545) I(R8460t757) I(R8461t1215) I(R8461t2896) I(R8461t7557) I(R8461t1272) I(R8462t4269) I(R8462t5927) I(R8462t5937) I(R8462t3469) I(R8462t5012) I(R8462t2911) I(R8462t3555) I(R8462t358) I(R8462t5127) I(R8463t1911) I(R8463t6532) I(R8463t37) I(R8464t2892) I(R8464t3277) I(R8464t7663) I(R8464t5795) I(R8464t2464) I(R8465t5812) I(R8465t8134) I(R8465t4902) I(R8465t7792) I(R8465t1065) I(R8465t1803) I(R8466t95) I(R8466t699) I(R8466t5624) I(R8466t5778) I(R8466t2913) I(R8466t5466) I(R8467t45) I(R8467t2951) I(R8467t2888) I(R8467t4142) I(R8467t3457) I(R8468t2322) I(R8468t6880) I(R8468t7011) I(R8468t364) I(R8468t6005) I(R8469t547) I(R8469t8052) I(R8469t1467) I(R8469t1415) I(R8469t4105) I(R8470t3327) I(R8470t7005) I(R8470t1547) I(R8470t8446) I(R8470t6262) I(R8470t870) I(R8471t2949) I(R8471t6010) I(R8471t7199) I(R8471t4287) I(R8471t1250) I(R8471t1515) I(R8472t6323) I(R8472t6456) I(R8472t430) I(R8472t1448) I(R8472t7890) I(R8473t2336) I(R8473t3309) I(R8473t349) I(R8473t7605) I(R8473t3986) I(R8473t140) I(R8473t6627) I(R8474t4518) I(R8474t7581) I(R8474t8344) I(R8474t2326) I(R8474t2831) I(R8474t7131) I(R8475t2025) I(R8475t5195) I(R8475t691) I(R8475t5233) I(R8475t6619) I(R8475t6354) I(R8475t8261) I(R8476t5256) I(R8476t6136) I(R8476t2029) I(R8477t5699) I(R8477t8085) I(R8477t3224) I(R8478t5208) I(R8478t5745) I(R8478t194) I(R8479t544) I(R8479t4180) I(R8479t1953) I(R8479t5698) I(R8479t4142) I(R8479t2888) I(R8480t1910) I(R8480t7716) I(R8480t2639) I(R8480t1794) I(R8480t7962) I(R8480t535) I(R8481t2606) I(R8481t4139) I(R8481t1040) I(R8481t2435) I(R8481t5755) I(R8481t4842) I(R8482t826) I(R8482t6137) I(R8482t2508) I(R8482t4856) I(R8482t1353) I(R8483t4677) I(R8483t5346) I(R8483t7538) I(R8483t8039) I(R8483t367) I(R8483t6667) I(R8483t3409) I(R8483t7276) I(R8483t5938) I(R8484t4344) I(R8484t6774) I(R8484t6247) I(R8484t5337) I(R8484t1915) I(R8485t883) I(R8485t3535) I(R8485t6806) I(R8485t1815) I(R8485t3256) I(R8486t89) I(R8486t3416) I(R8486t6995) I(R8486t154) I(R8487t1536) I(R8487t5622) I(R8487t4645) I(R8487t7717) I(R8487t4604) I(R8487t7245) I(R8488t2821) I(R8488t3902) I(R8488t3933) I(R8488t5445) I(R8488t2593) I(R8488t1280) I(R8488t6397) I(R8489t929) I(R8489t3141) I(R8489t3861) I(R8489t835) I(R8489t7193) I(R8489t3045) I(R8490t211) I(R8490t808) I(R8490t7841) I(R8490t1868) I(R8490t366) I(R8490t2818) I(R8491t1707) I(R8491t6551) I(R8491t6188) I(R8491t4262) I(R8491t587) I(R8492t3624) I(R8492t5784) I(R8492t4164) I(R8492t2624) I(R8493t2648) I(R8493t6778) I(R8493t3024) I(R8493t6243) I(R8493t6039) I(R8493t5042) I(R8494t2547) I(R8494t3911) I(R8494t2178) I(R8494t5967) I(R8494t3551) I(R8494t3073) I(R8495t1933) I(R8495t6166) I(R8495t6565) I(R8495t5098) I(R8495t1739) I(R8496t6577) I(R8496t8071) I(R8496t7400) I(R8496t5449) I(R8497t5000) I(R8497t6055) I(R8497t6348) I(R8497t1489) I(R8497t6326) I(R8497t7593) I(R8497t6529) I(R8498t4213) I(R8498t4675) I(R8498t6601) I(R8498t1672) I(R8498t3163) I(R8498t2271) I(R8499t5787) I(R8499t1787) I(R8500t5141) I(R8500t2927) I(R8500t510) I(R8500t8006) I(R8500t1767) I(R8500t3043) I(R8501t5046) I(R8501t6757) I(R8501t3149) I(R8501t4469) I(R8502t1679) I(R8502t5805) I(R8502t2367) I(R8502t8369) I(R8503t3193) I(R8503t1422) I(R8504t4552) I(R8504t5237) I(R8504t7129) I(R8505t5745) I(R8505t6480) I(R8505t8478) I(R8505t5208) I(R8505t4030) I(R8505t6245) I(R8505t1244) I(R8505t1606) I(R8506t4948) I(R8506t5961) I(R8506t6259) I(R8506t5098) I(R8506t8495) I(R8506t6565) I(R8506t2403) I(R8507t2523) I(R8507t199) I(R8507t1253) I(R8507t804) I(R8508t3992) I(R8508t4300) I(R8508t1217) I(R8508t3801) I(R8508t7675) I(R8508t4505) I(R8509t5135) I(R8509t5774) I(R8509t558) I(R8509t2291) I(R8509t476) I(R8510t1228) I(R8510t8393) I(R8510t3688) I(R8510t2519) I(R8511t8017) I(R8511t1412) I(R8511t2308) I(R8511t3708) I(R8511t2977) I(R8512t1955) I(R8512t5216) I(R8512t4464) I(R8512t2221) I(R8512t3808) I(R8513t5956) I(R8513t6905) I(R8513t420) I(R8513t2852) I(R8513t7054) I(R8514t4604) I(R8514t571) I(R8514t5676) I(R8514t7380) I(R8515t8476) I(R8515t2029) I(R8515t6726) I(R8515t5626) I(R8516t5532) I(R8516t5720) I(R8516t6375) I(R8516t6604) I(R8517t3234) I(R8517t7267) I(R8517t2835) I(R8517t8411) I(R8517t2575) I(R8517t6304) I(R8518t5535) I(R8518t2455) I(R8518t212) I(R8519t3228) I(R8519t3995) I(R8519t5089) I(R8519t2150) I(R8519t4028) I(R8520t7885) I(R8520t1855) I(R8520t6399) I(R8520t8305) I(R8520t307) I(R8520t7172) I(R8520t3217) I(R8521t180) I(R8521t7281) I(R8521t2341) I(R8521t6346) I(R8521t6320) I(R8521t4027) I(R8521t5347) I(R8522t7566) I(R8522t1556) I(R8523t7138) I(R8523t4362) I(R8523t3342) I(R8524t2419) I(R8524t2699) I(R8524t5529) I(R8524t5045) I(R8524t3590) I(R8525t1385) I(R8525t2599) I(R8525t4303) I(R8525t2041) I(R8525t6053) I(R8525t4281) I(R8525t7385) I(R8526t3298) I(R8526t5454) I(R8526t3222) I(R8526t5168) I(R8526t7482) I(R8526t8111) I(R8526t4881) I(R8527t1566) I(R8527t4129) I(R8527t2372) I(R8527t1359) I(R8527t2730) I(R8528t4198) I(R8528t6113) I(R8528t5804) I(R8528t1906) I(R8528t5114) I(R8528t6818) I(R8528t7854) I(R8528t593) I(R8528t2720) I(R8529t1342) I(R8529t3438) I(R8529t4979) I(R8529t7399) I(R8529t3360) I(R8530t2970) I(R8530t7344) I(R8530t837) I(R8530t1070) I(R8530t537) I(R8530t3098) I(R8531t4347) I(R8531t7308) I(R8531t777) I(R8531t1509) I(R8531t1417) I(R8531t2204) I(R8531t3142) I(R8531t3157) I(R8532t2348) I(R8532t3263) I(R8532t2611) I(R8532t4871) I(R8532t5026) I(R8532t3354) I(R8532t513) I(R8533t735) I(R8533t6486) I(R8533t2916) I(R8533t8253) I(R8533t5414) I(R8533t3974) I(R8533t7418) I(R8534t2051) I(R8534t3269) I(R8534t529) I(R8534t3592) I(R8534t5958) I(R8535t684) I(R8535t5985) I(R8535t6264) I(R8535t7939) I(R8535t2849) I(R8535t6530) I(R8535t7695) I(R8536t3773) I(R8536t7783) I(R8536t5060) I(R8536t5014) I(R8536t8295) I(R8536t5439) I(R8536t6359) I(R8537t686) I(R8537t8089) I(R8537t3747) I(R8537t4971) I(R8537t4477) I(R8538t1895) I(R8538t4683) I(R8538t5819) I(R8538t7008) I(R8538t8016) I(R8538t437) I(R8539t3052) I(R8539t7295) I(R8539t6333) I(R8540t24) I(R8540t4190) I(R8541t5261) I(R8541t5378) I(R8541t4944) I(R8541t6123) I(R8541t1745) I(R8541t4886) I(R8541t8078) I(R8542t152) I(R8542t6851) I(R8542t6060) I(R8542t4841) I(R8542t2365) I(R8542t4579) I(R8542t5516) I(R8543t261) I(R8543t1535) I(R8543t7626) I(R8543t1738) I(R8543t1914) I(R8543t1497) I(R8544t1234) I(R8544t8040) I(R8544t1828) I(R8544t2087) I(R8544t6447) I(R8545t1996) I(R8545t6469) I(R8545t8499) I(R8545t1787) I(R8545t5330) I(R8546t827) I(R8546t3625) I(R8546t6176) I(R8546t3691) I(R8546t6127) I(R8547t3824) I(R8547t4698) I(R8547t3818) I(R8547t5181) I(R8547t4881) I(R8548t8165) I(R8548t2574) I(R8549t5168) I(R8549t8526) I(R8549t3222) I(R8549t1435) I(R8549t3189) I(R8549t4991) I(R8550t3188) I(R8550t5605) I(R8550t4890) I(R8550t8357) I(R8550t4771) I(R8551t950) I(R8551t559) I(R8551t5538) I(R8552t6998) I(R8552t4444) I(R8552t4998) I(R8552t7141) I(R8552t7914) I(R8552t8170) I(R8553t980) I(R8553t1074) I(R8553t3103) I(R8553t3899) I(R8553t993) I(R8554t7176) I(R8554t3366) I(R8554t3455) I(R8555t2425) I(R8555t7944) I(R8555t3999) I(R8555t2119) I(R8555t6237) I(R8555t4769) I(R8556t4205) I(R8556t363) I(R8556t2870) I(R8556t2033) I(R8556t3604) I(R8557t1126) I(R8557t8260) I(R8557t7374) I(R8558t1551) I(R8558t1806) I(R8558t367) I(R8558t7109) I(R8558t2003) I(R8558t4143) I(R8558t3885) I(R8559t4781) I(R8559t7029) I(R8559t5634) I(R8559t5371) I(R8559t6147) I(R8559t1719) I(R8560t4646) I(R8560t5547) I(R8560t2939) I(R8560t8456) I(R8560t1256) I(R8560t4016) I(R8560t1873) I(R8560t6222) I(R8560t6799) I(R8561t3211) I(R8561t4977) I(R8561t6386) I(R8561t3148) I(R8561t1066) I(R8561t1845) I(R8562t854) I(R8562t8202) I(R8562t8215) I(R8562t2959) I(R8563t1946) I(R8563t2270) I(R8563t519) I(R8563t5023) I(R8563t5355) I(R8563t2642) I(R8563t5949) I(R8564t4039) I(R8564t5294) I(R8564t1810) I(R8564t6515) I(R8564t6061) I(R8564t4603) I(R8564t6643) I(R8565t642) I(R8565t5162) I(R8565t1499) I(R8565t8405) I(R8565t1176) I(R8565t881) I(R8565t3082) I(R8566t2891) I(R8566t4882) I(R8566t715) I(R8566t4707) I(R8566t6838) I(R8566t7021) I(R8566t6236) I(R8567t2203) I(R8567t6771) I(R8567t2654) I(R8567t5563) I(R8567t5120) I(R8567t8271) I(R8567t3630) I(R8568t4531) I(R8568t7843) I(R8568t450) I(R8568t2696) I(R8568t7982) I(R8568t7697) I(R8568t2205) I(R8569t2202) I(R8569t7237) I(R8569t1926) I(R8569t651) I(R8569t7229) I(R8570t1398) I(R8570t3541) I(R8570t8192) I(R8570t3374) I(R8570t2779) I(R8570t3559) I(R8571t3381) I(R8571t4672) I(R8571t5986) I(R8571t7489) I(R8571t8298) I(R8572t356) I(R8572t5134) I(R8572t6234) I(R8572t7074) I(R8572t4293) I(R8573t3040) I(R8573t3262) I(R8573t7497) I(R8573t288) I(R8573t1928) I(R8573t5590) I(R8573t337) I(R8573t6657) I(R8573t1306) I(R8573t4035) I(R8574t4397) I(R8574t6159) I(R8574t333) I(R8574t3148) I(R8574t6843) I(R8575t4697) I(R8575t6665) I(R8575t2925) I(R8575t3800) I(R8575t6443) I(R8575t8402) I(R8575t3621) I(R8576t2234) I(R8576t6499) I(R8576t2130) I(R8576t3825) I(R8576t4660) I(R8577t4546) I(R8577t7885) I(R8577t5687) I(R8577t5891) I(R8577t2120) I(R8577t1741) I(R8577t5751) I(R8577t5913) I(R8577t1855) I(R8577t8520) I(R8578t6381) I(R8578t6779) I(R8578t1361) I(R8578t7580) I(R8579t2783) I(R8579t2932) I(R8579t3995) I(R8579t6621) I(R8579t3676) I(R8579t7978) I(R8579t4990) I(R8580t1402) I(R8580t3123) I(R8580t5741) I(R8580t1342) I(R8580t8529) I(R8581t1342) I(R8581t5741) I(R8581t2342) I(R8582t3371) I(R8582t3278) I(R8582t7440) I(R8582t7103) I(R8582t5551) I(R8583t2891) I(R8583t4882) I(R8583t7597) I(R8583t1160) I(R8583t2324) I(R8584t3982) I(R8584t5744) I(R8584t8242) I(R8584t6515) I(R8584t5357) I(R8584t2787) I(R8584t3749) I(R8585t985) I(R8585t6701) I(R8585t2016) I(R8585t1589) I(R8585t4806) I(R8586t392) I(R8586t6536) I(R8586t1365) I(R8587t3329) I(R8587t7351) I(R8587t1087) I(R8587t5488) I(R8587t1134) I(R8587t116) I(R8587t4575) I(R8588t2600) I(R8588t3421) I(R8588t3585) I(R8588t1541) I(R8589t5367) I(R8589t5671) I(R8589t2906) I(R8589t877) I(R8589t5905) I(R8590t2049) I(R8590t7099) I(R8590t1190) I(R8590t7108) I(R8590t6990) I(R8591t4014) I(R8591t7967) I(R8591t6406) I(R8591t7036) I(R8591t1693) I(R8591t1802) I(R8592t6401) I(R8592t8399) I(R8592t7745) I(R8593t463) I(R8593t2004) I(R8593t4929) I(R8593t275) I(R8593t1909) I(R8593t3793) I(R8594t502) I(R8594t2398) I(R8594t1158) I(R8594t2210) I(R8594t4181) I(R8595t3725) I(R8595t7754) I(R8595t926) I(R8595t6182) I(R8595t1790) I(R8596t1729) I(R8596t3373) I(R8596t2210) I(R8596t4181) I(R8597t4475) I(R8597t6577) I(R8597t3326) I(R8597t2565) I(R8597t1468) I(R8598t3588) I(R8598t4949) I(R8598t3864) I(R8598t687) I(R8598t2942) I(R8598t7128) I(R8598t8369) I(R8598t2367) I(R8598t7012) I(R8599t2721) I(R8599t6425) I(R8599t2916) I(R8599t8533) I(R8599t8253) I(R8600t1692) I(R8600t7657) I(R8600t7964) I(R8600t4335) I(R8601t5231) I(R8601t5283) I(R8601t1559) I(R8601t4787) I(R8601t2996) I(R8601t5169) I(R8602t6691) I(R8602t5442) I(R8603t5900) I(R8603t7292) I(R8603t7968) I(R8603t4417) I(R8603t5782) I(R8603t5267) I(R8604t8448) I(R8604t5995) I(R8604t6232) I(R8604t7635) I(R8605t3316) I(R8605t7495) I(R8605t2819) I(R8605t4121) I(R8605t1196) I(R8605t5701) I(R8605t5482) I(R8606t3532) I(R8606t7285) I(R8606t6513) I(R8606t4752) I(R8606t556) I(R8607t7518) I(R8607t8327) I(R8607t2591) I(R8607t4625) I(R8607t1808) I(R8608t405) I(R8608t4017) I(R8608t7792) I(R8608t7689) I(R8608t4726) I(R8609t3115) I(R8609t6697) I(R8609t3700) I(R8609t6615) I(R8609t1801) I(R8609t2183) I(R8610t1167) I(R8610t5194) I(R8610t4303) I(R8610t2467) I(R8611t289) I(R8611t4787) I(R8611t3781) I(R8611t5828) I(R8611t7193) I(R8611t3045) I(R8611t2650) I(R8612t1670) I(R8612t6342) I(R8612t3389) I(R8612t2247) I(R8613t1399) I(R8613t2531) I(R8613t1730) I(R8614t6599) I(R8614t7947) I(R8614t7064) I(R8614t4819) I(R8615t6731) I(R8615t6834) I(R8615t5538) I(R8615t8551) I(R8615t950) I(R8615t6297) I(R8616t2570) I(R8616t8299) I(R8616t5295) I(R8616t3239) I(R8616t573) I(R8616t4792) I(R8617t653) I(R8617t867) I(R8618t3199) I(R8618t6089) I(R8618t4219) I(R8618t4655) I(R8618t4180) I(R8618t4591) I(R8619t2726) I(R8619t7467) I(R8619t6013) I(R8619t352) I(R8619t1476) I(R8619t4791) I(R8619t852) I(R8620t2826) I(R8620t5327) I(R8620t4310) I(R8620t7548) I(R8620t5117) I(R8621t2959) I(R8621t8562) I(R8621t8215) I(R8621t2504) I(R8622t2952) I(R8622t4991) I(R8622t3732) I(R8622t752) I(R8622t1867) I(R8623t6930) I(R8623t8443) I(R8623t760) I(R8623t4097) I(R8623t4605) I(R8623t5829) I(R8624t2317) I(R8624t7781) I(R8624t4695) I(R8624t3721) I(R8625t2885) I(R8625t8398) I(R8625t2558) I(R8625t3658) I(R8626t348) I(R8626t3473) I(R8626t7160) I(R8626t3957) I(R8627t1014) I(R8627t2064) I(R8627t3359) I(R8627t2206) I(R8627t6544) I(R8627t6829) I(R8627t6088) I(R8628t1283) I(R8628t3506) I(R8628t6103) I(R8628t3085) I(R8628t8412) I(R8628t2592) I(R8629t3315) I(R8629t6983) I(R8629t7172) I(R8629t8520) I(R8629t3217) I(R8629t2330) I(R8630t10) I(R8630t4570) I(R8630t4465) I(R8630t5088) I(R8630t8268) I(R8630t6991) I(R8631t2569) I(R8631t4168) I(R8631t354) I(R8631t5875) I(R8631t5700) I(R8632t4135) I(R8632t5292) I(R8632t5633) I(R8632t5419) I(R8632t8393) I(R8632t4747) I(R8632t6589) I(R8633t4046) I(R8633t5822) I(R8633t6212) I(R8633t5016) I(R8633t930) I(R8634t4947) I(R8634t5256) I(R8634t6832) I(R8634t5598) I(R8635t3904) I(R8635t4925) I(R8635t4859) I(R8635t709) I(R8635t2145) I(R8636t3629) I(R8636t5299) I(R8636t5511) I(R8637t2137) I(R8637t6931) I(R8637t4171) I(R8638t4606) I(R8638t850) I(R8638t3960) I(R8639t1398) I(R8639t3541) I(R8639t7170) I(R8639t4225) I(R8639t205) I(R8639t5304) I(R8639t2893) I(R8640t8175) I(R8640t6068) I(R8640t3631) I(R8640t8326) I(R8641t4107) I(R8641t5684) I(R8641t6121) I(R8641t3529) I(R8641t3215) I(R8641t7565) I(R8641t2560) I(R8642t2748) I(R8642t5988) I(R8643t665) I(R8643t8020) I(R8643t6357) I(R8644t305) I(R8644t6651) I(R8644t2472) I(R8644t488) I(R8644t1090) I(R8644t5469) I(R8645t4583) I(R8645t4777) I(R8645t3109) I(R8645t5327) I(R8645t4310) I(R8646t724) I(R8646t595) I(R8646t57) I(R8646t1694) I(R8646t1433) I(R8647t1778) I(R8647t8297) I(R8647t3282) I(R8647t937) I(R8647t8313) I(R8648t1659) I(R8648t4604) I(R8648t8514) I(R8648t7380) I(R8648t7714) I(R8648t3780) I(R8648t6783) I(R8648t6693) I(R8648t4624) I(R8649t3652) I(R8649t7115) I(R8649t5311) I(R8649t1070) I(R8649t837) I(R8650t2580) I(R8650t2815) I(R8650t698) I(R8650t8292) I(R8651t5201) I(R8651t6134) I(R8651t7563) I(R8651t4075) I(R8651t8378) I(R8652t3133) I(R8652t1259) I(R8652t6073) I(R8653t620) I(R8653t7946) I(R8653t6098) I(R8653t2401) I(R8653t266) I(R8654t1008) I(R8654t1895) I(R8654t3165) I(R8654t6197) I(R8654t4154) I(R8654t437) I(R8655t4053) I(R8655t4649) I(R8655t4120) I(R8655t3809) I(R8655t5403) I(R8655t8259) I(R8656t2630) I(R8656t2742) I(R8656t1490) I(R8656t1593) I(R8656t5895) I(R8656t1667) I(R8656t1106) I(R8656t4278) I(R8657t7657) I(R8657t8600) I(R8657t4335) I(R8657t8380) I(R8657t5175) I(R8657t1524) I(R8657t5767) I(R8658t2414) I(R8658t1936) I(R8658t2392) I(R8658t3076) I(R8658t3859) I(R8659t2361) I(R8659t4492) I(R8659t8397) I(R8659t3273) I(R8659t4799) I(R8660t3305) I(R8660t3426) I(R8660t7429) I(R8660t5794) I(R8660t7674) I(R8660t5977) I(R8660t6549) I(R8661t4470) I(R8661t6028) I(R8661t6780) I(R8661t5157) I(R8661t8308) I(R8661t6482) I(R8661t3244) I(R8661t3552) I(R8662t5321) I(R8662t7331) I(R8662t183) I(R8662t2516) I(R8662t7122) I(R8662t6980) I(R8663t2371) I(R8663t4761) I(R8663t1671) I(R8663t7734) I(R8663t6366) I(R8663t2011) I(R8664t83) I(R8664t1451) I(R8664t1567) I(R8664t1056) I(R8664t1218) I(R8665t8403) I(R8665t5554) I(R8665t2228) I(R8665t3955) I(R8665t1111) I(R8666t7155) I(R8666t520) I(R8666t7148) I(R8667t424) I(R8667t6331) I(R8667t5230) I(R8667t4735) I(R8668t4682) I(R8669t2197) I(R8669t6433) I(R8669t5644) I(R8669t2671) I(R8669t3180) I(R8669t7169) I(R8670t3557) I(R8670t8219) I(R8670t2430) I(R8670t5010) I(R8670t3106) I(R8670t3009) I(R8670t3606) I(R8671t352) I(R8671t6013) I(R8671t8338) I(R8671t8018) I(R8671t4987) I(R8672t6280) I(R8672t8348) I(R8672t5943) I(R8672t5796) I(R8672t1487) I(R8672t6391) I(R8673t7667) I(R8673t8110) I(R8673t711) I(R8673t6489) I(R8673t350) I(R8673t2000) I(R8674t3040) I(R8674t5247) I(R8674t4538) I(R8674t2855) I(R8674t4593) I(R8675t6878) I(R8675t7477) I(R8675t2738) I(R8675t3356) I(R8675t106) I(R8675t2292) I(R8676t7883) I(R8676t5904) I(R8676t7010) I(R8676t3961) I(R8677t1946) I(R8677t8366) I(R8677t2640) I(R8677t2769) I(R8677t5949) I(R8678t3020) I(R8678t5341) I(R8678t1113) I(R8678t5174) I(R8678t635) I(R8678t2370) I(R8678t4613) I(R8678t800) I(R8679t4454) I(R8679t6293) I(R8679t8281) I(R8679t4042) I(R8680t1484) I(R8680t6041) I(R8680t1383) I(R8680t7844) I(R8680t6646) I(R8681t2558) I(R8681t8185) I(R8681t2885) I(R8681t8625) I(R8682t3651) I(R8682t4351) I(R8682t4976) I(R8682t1076) I(R8682t4079) I(R8682t2844) I(R8682t3297) I(R8683t970) I(R8683t2237) I(R8683t484) I(R8683t8518) I(R8683t5535) I(R8684t2266) I(R8684t7370) I(R8684t5790) I(R8684t5136) I(R8684t8395) I(R8684t4274) I(R8685t3757) I(R8685t2448) I(R8685t7044) I(R8685t77) I(R8685t584) I(R8686t3143) I(R8686t3330) I(R8686t1428) I(R8686t5384) I(R8686t8088) I(R8686t4260) I(R8687t3723) I(R8687t7528) I(R8687t2038) I(R8687t6713) I(R8687t1408) I(R8688t6170) I(R8688t7162) I(R8688t2410) I(R8688t4013) I(R8688t6867) I(R8688t6931) I(R8688t6822) I(R8688t6747) I(R8689t5018) I(R8689t7731) I(R8689t1193) I(R8689t1120) I(R8690t6289) I(R8690t7413) I(R8690t3266) I(R8690t1867) I(R8690t6417) I(R8691t5468) I(R8691t7854) I(R8691t8528) I(R8691t593) I(R8691t4209) I(R8692t2040) I(R8692t2656) I(R8692t6913) I(R8692t5666) I(R8692t6203) I(R8693t1300) I(R8693t8322) I(R8693t6322) I(R8693t6338) I(R8693t3865) I(R8693t6238) I(R8693t1330) I(R8694t3724) I(R8694t5286) I(R8694t801) I(R8694t2253) I(R8695t2633) I(R8695t8166) I(R8695t4047) I(R8695t5498) I(R8695t4128) I(R8695t1513) I(R8696t1989) I(R8696t6224) I(R8696t2432) I(R8696t2194) I(R8696t3840) I(R8697t5309) I(R8697t4244) I(R8697t3390) I(R8697t5293) I(R8697t6884) I(R8698t982) I(R8698t3364) I(R8698t7144) I(R8698t7527) I(R8698t3953) I(R8698t7435) I(R8699t8277) I(R8699t482) I(R8699t1326) I(R8699t993) I(R8699t3711) I(R8699t2413) I(R8700t1193) I(R8700t8689) I(R8700t8182) I(R8700t5657) I(R8700t3114) I(R8700t5107) I(R8700t6829) I(R8700t8379) I(R8700t1120) I(R8701t4119) I(R8701t6045) I(R8701t5247) I(R8701t4538) I(R8701t1532) I(R8701t2420) I(R8702t1792) I(R8702t5931) I(R8702t1444) I(R8702t2454) I(R8702t4217) I(R8703t413) I(R8703t3691) I(R8703t1573) I(R8703t190) I(R8703t5769) I(R8704t7539) I(R8704t1262) I(R8704t6782) I(R8705t2159) I(R8705t3929) I(R8705t2733) I(R8705t5165) I(R8705t451) I(R8706t3132) I(R8706t5833) I(R8706t38) I(R8707t2260) I(R8707t4535) I(R8707t739) I(R8707t5654) I(R8707t1474) I(R8707t8441) I(R8708t3548) I(R8708t7889) I(R8708t6571) I(R8708t8205) I(R8708t24) I(R8708t8540) I(R8708t4190) I(R8709t2099) I(R8709t5821) I(R8709t6485) I(R8709t5111) I(R8710t885) I(R8710t4280) I(R8710t1923) I(R8710t2012) I(R8711t744) I(R8711t2194) I(R8711t5058) I(R8711t6525) I(R8711t8220) I(R8711t6000) I(R8711t2928) I(R8712t2382) I(R8712t8296) I(R8712t7981) I(R8712t2794) I(R8713t722) I(R8713t5532) I(R8713t8516) I(R8713t6604) I(R8713t4177) I(R8713t2305) I(R8713t8167) I(R8714t2135) I(R8714t7432) I(R8714t8210) I(R8714t2910) I(R8714t8094) I(R8714t1009) I(R8715t4932) I(R8715t6084) I(R8715t5029) I(R8715t4218) I(R8715t5572) I(R8716t58) I(R8716t6669) I(R8716t5497) I(R8716t456) I(R8716t1970) I(R8717t2799) I(R8717t7246) I(R8717t7323) I(R8717t3485) I(R8717t8380) I(R8717t7678) I(R8717t4782) I(R8717t1651) I(R8718t867) I(R8718t54) I(R8718t8433) I(R8718t4442) I(R8718t7161) I(R8718t653) I(R8718t8617) I(R8719t6420) I(R8719t2899) I(R8719t5832) I(R8719t8061) I(R8719t8424) I(R8720t4411) I(R8720t7899) I(R8720t7381) I(R8720t6557) I(R8721t5879) I(R8721t6814) I(R8721t7403) I(R8721t2228) I(R8721t3955) I(R8721t7510) I(R8722t1892) I(R8722t2525) I(R8722t83) I(R8722t8664) I(R8722t1218) I(R8723t992) I(R8723t1018) I(R8723t5556) I(R8723t6970) I(R8723t3178) I(R8723t754) I(R8723t5896) I(R8723t1035) I(R8723t1370) I(R8723t5970) I(R8724t2369) I(R8724t6108) I(R8724t112) I(R8724t5856) I(R8724t6653) I(R8724t2028) I(R8724t3666) I(R8725t4924) I(R8725t3510) I(R8725t591) I(R8725t1867) I(R8725t6417) I(R8726t4255) I(R8726t6369) I(R8726t427) I(R8726t7720) I(R8726t3067) I(R8726t6777) I(R8726t1793) I(R8727t2743) I(R8727t7852) I(R8727t9) I(R8727t7299) I(R8727t7488) I(R8728t175) I(R8728t4606) I(R8728t751) I(R8729t3585) I(R8729t8588) I(R8729t7088) I(R8729t3459) I(R8729t5999) I(R8729t1541) I(R8730t1788) I(R8730t7753) I(R8730t3311) I(R8730t6584) I(R8730t6340) I(R8731t2322) I(R8731t5263) I(R8731t822) I(R8731t6574) I(R8731t3204) I(R8731t227) I(R8732t3379) I(R8732t5394) I(R8732t8164) I(R8733t4934) I(R8733t6513) I(R8733t1966) I(R8733t5711) I(R8734t2776) I(R8734t3680) I(R8735t4234) I(R8735t7693) I(R8735t2661) I(R8735t5817) I(R8736t3632) I(R8736t4768) I(R8736t3022) I(R8737t7077) I(R8737t6886) I(R8737t2533) I(R8737t81) I(R8737t5285) I(R8738t809) I(R8738t1837) I(R8738t4147) I(R8738t3949) I(R8739t968) I(R8739t7901) I(R8739t2865) I(R8739t6831) I(R8739t632) I(R8740t32) I(R8740t2163) I(R8740t3868) I(R8740t3093) I(R8741t4759) I(R8741t5352) I(R8741t3927) I(R8741t895) I(R8741t4628) I(R8741t8409) I(R8741t7257) I(R8741t1763) I(R8741t2792) I(R8742t5112) I(R8742t7967) I(R8743t1406) I(R8743t3391) I(R8743t8368) I(R8743t5773) I(R8743t6042) I(R8743t7339) I(R8744t3083) I(R8744t5830) I(R8744t7236) I(R8744t6891) I(R8744t1242) I(R8744t2808) I(R8745t2776) I(R8745t8734) I(R8745t7871) I(R8745t4026) I(R8746t997) I(R8746t7908) I(R8746t7827) I(R8746t2839) I(R8746t8294) I(R8746t8238) I(R8746t5036) I(R8747t3754) I(R8747t8279) I(R8747t2711) I(R8747t5456) I(R8747t3172) I(R8748t2953) I(R8748t7631) I(R8748t2245) I(R8748t6156) I(R8748t239) I(R8748t3748) I(R8749t650) I(R8749t6172) I(R8749t1705) I(R8749t4476) I(R8749t3839) I(R8750t2955) I(R8750t6467) I(R8750t7483) I(R8750t4076) I(R8750t6441) I(R8750t4497) I(R8750t3109) I(R8751t3810) I(R8751t7992) I(R8751t1548) I(R8751t3894) I(R8751t1211) I(R8751t7980) I(R8751t8169) I(R8752t6018) I(R8752t8239) I(R8752t1284) I(R8752t2428) I(R8752t3338) I(R8753t273) I(R8753t8053) I(R8753t7844) I(R8753t4880) I(R8753t1655) I(R8754t386) I(R8754t3124) I(R8754t2724) I(R8754t4142) I(R8754t5698) I(R8755t5597) I(R8755t5687) I(R8755t7996) I(R8755t8316) I(R8755t5891) I(R8755t8577) I(R8756t6401) I(R8756t8592) I(R8756t3399) I(R8756t3179) I(R8756t6575) I(R8756t7745) I(R8757t431) I(R8757t8247) I(R8757t2716) I(R8757t1250) I(R8757t1515) I(R8757t6010) I(R8757t3554) I(R8757t3015) I(R8758t272) I(R8758t5804) I(R8758t3116) I(R8758t4824) I(R8758t1950) I(R8758t7559) I(R8759t4629) I(R8759t7530) I(R8759t6006) I(R8759t719) I(R8759t2576) I(R8759t2333) I(R8760t617) I(R8760t5623) I(R8760t7973) I(R8760t6400) I(R8761t8214) I(R8761t8397) I(R8761t6017) I(R8761t2242) I(R8762t577) I(R8762t3041) I(R8762t991) I(R8762t4573) I(R8762t3433) I(R8763t908) I(R8763t3616) I(R8763t7842) I(R8763t6195) I(R8763t2930) I(R8764t1007) I(R8764t3619) I(R8764t5013) I(R8764t1449) I(R8764t3807) I(R8764t3813) I(R8765t2315) I(R8765t3720) I(R8765t6570) I(R8765t5611) I(R8765t7483) I(R8765t5187) I(R8766t7327) I(R8766t2968) I(R8766t4565) I(R8767t816) I(R8767t4055) I(R8767t607) I(R8767t3084) I(R8767t4671) I(R8767t8143) I(R8767t8341) I(R8767t659) I(R8768t4316) I(R8768t4933) I(R8768t7896) I(R8768t7687) I(R8768t4242) I(R8769t141) I(R8769t7690) I(R8769t4394) I(R8770t3402) I(R8770t6019) I(R8770t6107) I(R8771t7941) I(R8771t5376) I(R8771t8347) I(R8771t1333) I(R8771t7123) I(R8771t8328) I(R8772t5002) I(R8772t5831) I(R8772t2555) I(R8772t8151) I(R8772t4473) I(R8772t133) I(R8772t445) I(R8772t7767) I(R8772t5717) I(R8772t1858) I(R8773t1090) I(R8773t488) I(R8773t6898) I(R8774t8017) I(R8774t8511) I(R8774t1412) I(R8774t6142) I(R8774t7110) I(R8775t5460) I(R8775t4679) I(R8775t6218) I(R8776t6577) I(R8776t8496) I(R8776t5449) I(R8776t1116) I(R8776t1468) I(R8777t439) I(R8777t1635) I(R8777t8339) I(R8777t2661) I(R8777t4234) I(R8777t1617) I(R8778t728) I(R8778t1563) I(R8778t7298) I(R8778t7975) I(R8778t2152) I(R8778t1493) I(R8779t115) I(R8779t5338) I(R8779t11) I(R8779t4420) I(R8779t1819) I(R8779t2755) I(R8780t449) I(R8780t2436) I(R8780t2285) I(R8780t3816) I(R8780t2482) I(R8780t2715) I(R8781t7327) I(R8781t8766) I(R8781t4565) I(R8781t2393) I(R8781t532) I(R8782t3453) I(R8782t3739) I(R8782t4001) I(R8782t726) I(R8782t2990) I(R8782t7734) I(R8782t1671) I(R8783t3374) I(R8783t8087) I(R8783t5534) I(R8783t5680) I(R8783t6546) I(R8783t3276) I(R8784t4794) I(R8784t4946) I(R8784t4600) I(R8784t7912) I(R8784t6307) I(R8784t5092) I(R8785t734) I(R8785t5770) I(R8785t5833) I(R8785t7306) I(R8785t6182) I(R8786t8000) I(R8786t8003) I(R8786t1151) I(R8786t6040) I(R8786t1928) I(R8786t927) I(R8787t2200) I(R8787t2347) I(R8787t7091) I(R8787t3163) I(R8787t6324) I(R8787t6078) I(R8788t3000) I(R8788t5841) I(R8788t831) I(R8789t73) I(R8789t5814) I(R8789t1475) I(R8789t3481) I(R8789t6053) I(R8790t5736) I(R8790t7653) I(R8790t4952) I(R8790t7690) I(R8790t8769) I(R8790t4394) I(R8791t6090) I(R8791t4385) I(R8791t5396) I(R8791t6345) I(R8792t1678) I(R8792t8278) I(R8792t3979) I(R8792t3235) I(R8792t3814) I(R8793t1972) I(R8793t5725) I(R8793t5181) I(R8794t854) I(R8794t4179) I(R8794t8562) I(R8794t8202) I(R8794t8120) I(R8794t2543) I(R8795t6680) I(R8795t7742) I(R8795t3639) I(R8795t6906) I(R8795t5262) I(R8796t1470) I(R8796t3049) I(R8796t5551) I(R8796t8582) I(R8796t3371) I(R8797t4208) I(R8797t7020) I(R8797t5937) I(R8797t3469) I(R8797t7478) I(R8797t4043) I(R8798t4263) I(R8798t164) I(R8798t2359) I(R8799t1957) I(R8799t4048) I(R8799t3059) I(R8799t6502) I(R8799t4809) I(R8799t4978) I(R8799t2785) I(R8800t3973) I(R8800t4557) I(R8800t4096) I(R8800t2191) I(R8800t6092) I(R8800t8342) I(R8801t1690) I(R8801t1790) I(R8801t2151) I(R8801t2800) I(R8802t2893) I(R8802t5304) I(R8802t6837) I(R8802t7597) I(R8802t3777) I(R8803t5857) I(R8803t7165) I(R8803t182) I(R8803t2822) I(R8803t142) I(R8804t1494) I(R8804t4546) I(R8804t8577) I(R8804t5687) I(R8804t5597) I(R8804t2174) I(R8805t1372) I(R8805t5422) I(R8805t2954) I(R8805t2709) I(R8805t71) I(R8806t235) I(R8806t2104) I(R8806t6207) I(R8806t8420) I(R8806t1720) I(R8807t4456) I(R8807t7548) I(R8807t4284) I(R8807t5117) I(R8808t2649) I(R8808t7663) I(R8808t3277) I(R8808t3481) I(R8808t684) I(R8808t8258) I(R8809t2932) I(R8809t7214) I(R8809t1764) I(R8809t4990) I(R8809t8579) I(R8810t1130) I(R8810t2359) I(R8810t7925) I(R8810t5589) I(R8810t5361) I(R8810t7472) I(R8811t2770) I(R8811t3069) I(R8811t7145) I(R8811t1786) I(R8811t7920) I(R8811t3101) I(R8811t1030) I(R8811t3799) I(R8812t4637) I(R8812t7995) I(R8812t3505) I(R8812t7095) I(R8812t8372) I(R8813t4345) I(R8813t5693) I(R8813t3899) I(R8813t7960) I(R8813t1002) I(R8813t8224) I(R8814t4528) I(R8814t6302) I(R8814t8317) I(R8814t1119) I(R8814t2500) I(R8815t3380) I(R8815t6170) I(R8815t2398) I(R8815t12) I(R8815t3005) I(R8816t1407) I(R8816t3415) I(R8816t3715) I(R8816t1313) I(R8816t7468) I(R8817t1639) I(R8817t7287) I(R8817t3389) I(R8817t2964) I(R8817t3924) I(R8817t4969) I(R8818t836) I(R8818t890) I(R8818t7608) I(R8819t1386) I(R8819t6420) I(R8819t6427) I(R8819t833) I(R8819t2899) I(R8819t8719) I(R8820t3814) I(R8820t5362) I(R8820t8792) I(R8820t3235) I(R8820t741) I(R8821t5693) I(R8821t8813) I(R8821t747) I(R8821t3103) I(R8821t3899) I(R8822t5261) I(R8822t5900) I(R8822t8603) I(R8822t5267) I(R8823t4434) I(R8823t5559) I(R8823t2119) I(R8823t8555) I(R8823t3999) I(R8823t2989) I(R8823t7604) I(R8824t4101) I(R8824t5068) I(R8824t1274) I(R8824t5792) I(R8825t7501) I(R8825t369) I(R8825t1573) I(R8825t190) I(R8825t3379) I(R8825t8732) I(R8825t8164) I(R8826t4539) I(R8826t4233) I(R8826t6388) I(R8827t8775) I(R8827t2376) I(R8827t3335) I(R8827t7355) I(R8827t265) I(R8827t6218) I(R8828t1514) I(R8828t3199) I(R8828t6286) I(R8828t4219) I(R8828t8618) I(R8829t2620) I(R8829t4876) I(R8829t6674) I(R8829t7898) I(R8829t3577) I(R8830t7323) I(R8830t7383) I(R8830t3485) I(R8830t5175) I(R8830t43) I(R8831t8622) I(R8831t4991) I(R8831t8549) I(R8831t5168) I(R8831t7895) I(R8831t6884) I(R8831t3266) I(R8832t314) I(R8832t4611) I(R8832t903) I(R8832t4359) I(R8832t8330) I(R8832t2986) I(R8833t28) I(R8833t6611) I(R8833t8653) I(R8833t266) I(R8834t198) I(R8834t743) I(R8834t3960) I(R8834t8638) I(R8834t850) I(R8834t666) I(R8835t5118) I(R8835t1014) I(R8835t3359) I(R8835t5840) I(R8836t421) I(R8836t5066) I(R8836t616) I(R8836t7498) I(R8836t4405) I(R8836t6532) I(R8837t8173) I(R8837t6409) I(R8837t5360) I(R8837t5402) I(R8837t6872) I(R8837t4051) I(R8838t3375) I(R8838t8263) I(R8838t6218) I(R8838t5145) I(R8838t4500) I(R8838t2984) I(R8838t3259) I(R8839t2057) I(R8839t5387) I(R8839t5713) I(R8839t66) I(R8839t3192) I(R8839t5476) I(R8840t4368) I(R8840t5072) I(R8840t7112) I(R8840t6032) I(R8840t5479) I(R8840t5303) I(R8841t2743) I(R8841t8727) I(R8841t9) I(R8841t7561) I(R8841t1826) I(R8841t2437) I(R8842t5708) I(R8842t6158) I(R8842t327) I(R8843t323) I(R8843t3342) I(R8843t7166) I(R8843t7089) I(R8843t3890) I(R8843t4362) I(R8843t8523) I(R8844t3343) I(R8844t5105) I(R8844t3771) I(R8844t871) I(R8844t5208) I(R8845t4902) I(R8845t7792) I(R8845t3334) I(R8845t6832) I(R8845t2862) I(R8846t1914) I(R8846t3607) I(R8846t3715) I(R8846t5221) I(R8846t1108) I(R8846t1738) I(R8847t8142) I(R8847t8197) I(R8847t6240) I(R8847t4898) I(R8847t7027) I(R8848t167) I(R8848t4547) I(R8848t3579) I(R8848t392) I(R8848t8586) I(R8848t6536) I(R8849t4442) I(R8849t8433) I(R8849t7950) I(R8849t6492) I(R8849t414) I(R8849t5122) I(R8849t7309) I(R8849t7161) I(R8850t5532) I(R8850t8516) I(R8850t5720) I(R8850t2999) I(R8850t7480) I(R8851t598) I(R8851t4328) I(R8851t2270) I(R8851t1946) I(R8851t8366) I(R8851t7784) I(R8852t692) I(R8852t1161) I(R8852t2900) I(R8852t7416) I(R8852t8274) I(R8852t706) I(R8853t3826) I(R8853t8218) I(R8853t7900) I(R8853t4037) I(R8853t4505) I(R8853t3992) I(R8853t7778) I(R8854t4921) I(R8854t1114) I(R8854t7342) I(R8854t7606) I(R8854t3947) I(R8854t2154) I(R8854t7204) I(R8855t6206) I(R8855t4291) I(R8855t815) I(R8855t5460) I(R8856t8285) I(R8856t3385) I(R8856t4280) I(R8856t3909) I(R8856t7296) I(R8857t2004) I(R8857t8432) I(R8857t3011) I(R8857t1475) I(R8857t3793) I(R8857t8593) I(R8858t1276) I(R8858t2601) I(R8858t5880) I(R8858t3295) I(R8858t2716) I(R8858t6911) I(R8859t7642) I(R8859t6141) I(R8859t7612) I(R8859t3176) I(R8859t4789) I(R8860t499) I(R8860t7970) I(R8860t1169) I(R8860t6168) I(R8860t2698) I(R8860t2669) I(R8860t5893) I(R8861t1632) I(R8861t8449) I(R8861t5949) I(R8861t8563) I(R8861t2642) I(R8861t2350) I(R8862t4083) I(R8862t5256) I(R8862t1958) I(R8862t6136) I(R8862t8476) I(R8863t2607) I(R8863t4426) I(R8863t4488) I(R8863t8133) I(R8863t6725) I(R8863t1599) I(R8864t6741) I(R8864t1935) I(R8864t8045) I(R8864t285) I(R8865t3313) I(R8865t6059) I(R8865t662) I(R8865t284) I(R8865t3430) I(R8865t7051) I(R8865t1554) I(R8866t3925) I(R8866t8004) I(R8866t2887) I(R8866t2549) I(R8866t2137) I(R8866t3354) I(R8866t513) I(R8867t5351) I(R8867t6474) I(R8867t7837) I(R8867t1826) I(R8867t7786) I(R8867t4674) I(R8867t3876) I(R8868t6222) I(R8868t8560) I(R8868t2193) I(R8868t4095) I(R8868t6799) I(R8869t5327) I(R8869t5465) I(R8869t3109) I(R8869t4514) I(R8869t2399) I(R8870t2826) I(R8870t8620) I(R8870t814) I(R8870t6576) I(R8870t3921) I(R8870t5117) I(R8871t3251) I(R8871t5725) I(R8871t3390) I(R8871t5293) I(R8871t4324) I(R8871t7040) I(R8871t128) I(R8872t723) I(R8872t2025) I(R8872t8054) I(R8872t8261) I(R8873t2414) I(R8873t8658) I(R8873t5825) I(R8873t1291) I(R8873t3859) I(R8874t1462) I(R8874t7582) I(R8874t3985) I(R8874t7318) I(R8874t4366) I(R8875t4834) I(R8876t7092) I(R8876t8049) I(R8876t8074) I(R8876t8386) I(R8876t3768) I(R8876t8101) I(R8876t6423) I(R8876t3157) I(R8877t2020) I(R8877t3005) I(R8877t8637) I(R8877t6931) I(R8877t6822) I(R8878t588) I(R8878t4667) I(R8878t6235) I(R8878t7818) I(R8878t5343) I(R8879t2118) I(R8879t4958) I(R8879t440) I(R8879t7873) I(R8879t1249) I(R8879t4166) I(R8880t2685) I(R8880t7227) I(R8880t2545) I(R8880t4113) I(R8880t2657) I(R8880t7893) I(R8881t206) I(R8881t2489) I(R8881t2488) I(R8881t5753) I(R8881t1022) I(R8882t2579) I(R8882t6786) I(R8882t4507) I(R8882t8019) I(R8882t526) I(R8883t2390) I(R8883t6458) I(R8883t8026) I(R8883t4058) I(R8884t1717) I(R8884t4230) I(R8884t2207) I(R8884t1347) I(R8884t1319) I(R8885t4637) I(R8885t6896) I(R8885t8372) I(R8885t7152) I(R8885t7403) I(R8885t2228) I(R8885t3077) I(R8885t3701) I(R8886t5112) I(R8886t8742) I(R8886t1496) I(R8886t8082) I(R8886t2039) I(R8887t626) I(R8887t1684) I(R8887t3574) I(R8887t3744) I(R8888t5883) I(R8888t4011) I(R8888t1676) I(R8888t1657) I(R8888t7338) I(R8888t2139) I(R8889t1451) I(R8889t6864) I(R8889t2480) I(R8889t2638) I(R8889t6917) I(R8890t1392) I(R8890t4499) I(R8890t3227) I(R8890t3569) I(R8890t5497) I(R8890t456) I(R8890t2275) I(R8891t1115) I(R8891t1150) I(R8891t2996) I(R8891t5169) I(R8891t5756) I(R8892t1269) I(R8892t2794) I(R8892t8712) I(R8892t7981) I(R8893t5650) I(R8893t8450) I(R8893t1580) I(R8894t5299) I(R8894t256) I(R8894t2412) I(R8895t914) I(R8895t1938) I(R8895t764) I(R8895t671) I(R8895t5660) I(R8895t2528) I(R8896t3968) I(R8896t4451) I(R8896t5544) I(R8896t4804) I(R8897t5369) I(R8897t7293) I(R8897t7283) I(R8897t2250) I(R8897t7489) I(R8897t5986) I(R8897t2351) I(R8898t927) I(R8898t8786) I(R8898t8191) I(R8898t288) I(R8898t1928) I(R8899t6305) I(R8899t8121) I(R8899t2415) I(R8899t6854) I(R8899t5348) I(R8899t4868) I(R8899t2722) I(R8899t2302) I(R8900t585) I(R8900t3312) I(R8900t2752) I(R8900t794) I(R8900t1784) I(R8900t6706) I(R8901t4995) I(R8901t8005) I(R8901t123) I(R8901t1767) I(R8902t6006) I(R8902t1223) I(R8902t478) I(R8902t3386) I(R8902t6055) I(R8902t1517) I(R8903t7066) I(R8903t8099) I(R8903t3518) I(R8903t3515) I(R8903t5034) I(R8903t118) I(R8904t5818) I(R8904t8170) I(R8904t6998) I(R8904t3207) I(R8904t1588) I(R8904t2809) I(R8905t4927) I(R8905t8375) I(R8905t5246) I(R8905t1139) I(R8906t2278) I(R8906t5388) I(R8906t2508) I(R8906t3596) I(R8906t1170) I(R8907t5915) I(R8907t6150) I(R8907t2719) I(R8907t2233) I(R8908t1549) I(R8908t2111) I(R8908t7634) I(R8908t7245) I(R8908t802) I(R8909t1269) I(R8909t3460) I(R8909t6315) I(R8909t214) I(R8909t1556) I(R8910t5118) I(R8910t8835) I(R8910t5840) I(R8910t3512) I(R8910t557) I(R8911t3886) I(R8911t8096) I(R8911t3618) I(R8911t4067) I(R8911t7330) I(R8911t97) I(R8912t695) I(R8912t1372) I(R8912t4067) I(R8912t3827) I(R8912t748) I(R8912t7436) I(R8912t3428) I(R8913t1351) I(R8913t5191) I(R8913t25) I(R8913t6335) I(R8913t4309) I(R8914t3024) I(R8914t7183) I(R8914t2514) I(R8914t2019) I(R8914t4709) I(R8915t6265) I(R8915t8229) I(R8915t8047) I(R8915t1735) I(R8916t260) I(R8916t4236) I(R8916t7257) I(R8916t2471) I(R8916t8196) I(R8917t3057) I(R8917t5730) I(R8917t2680) I(R8917t3373) I(R8917t8596) I(R8917t1729) I(R8918t4479) I(R8918t6099) I(R8918t4508) I(R8918t5551) I(R8918t8582) I(R8918t7103) I(R8919t1706) I(R8919t5057) I(R8919t8437) I(R8919t6950) I(R8920t4186) I(R8920t5018) I(R8920t3994) I(R8920t1029) I(R8920t3844) I(R8920t1925) I(R8920t1776) I(R8920t7430) I(R8920t1120) I(R8921t4827) I(R8921t1706) I(R8921t6802) I(R8921t1769) I(R8921t848) I(R8921t7105) I(R8922t6068) I(R8922t8640) I(R8922t4592) I(R8922t514) I(R8923t3594) I(R8923t544) I(R8923t4591) I(R8923t6089) I(R8923t8328) I(R8924t3862) I(R8924t8329) I(R8924t6719) I(R8924t2026) I(R8924t6477) I(R8924t5145) I(R8924t4500) I(R8925t4880) I(R8925t8753) I(R8925t7844) I(R8925t8680) I(R8926t2775) I(R8926t5849) I(R8926t3576) I(R8926t2482) I(R8926t4509) I(R8926t5955) I(R8927t1071) I(R8927t5141) I(R8927t2927) I(R8927t2967) I(R8927t2477) I(R8928t1803) I(R8928t3920) I(R8928t4265) I(R8928t5146) I(R8928t4025) I(R8928t4920) I(R8928t1065) I(R8929t1067) I(R8929t8311) I(R8929t4140) I(R8929t1918) I(R8929t503) I(R8930t1350) I(R8930t5246) I(R8930t1307) I(R8930t3824) I(R8930t3818) I(R8931t6022) I(R8931t2377) I(R8931t708) I(R8932t899) I(R8932t8213) I(R8932t3140) I(R8932t1888) I(R8932t8088) I(R8933t5665) I(R8933t5706) I(R8933t618) I(R8934t1990) I(R8934t2839) I(R8934t6696) I(R8934t7393) I(R8934t2933) I(R8935t5263) I(R8935t5508) I(R8935t1762) I(R8935t227) I(R8936t1523) I(R8936t5610) I(R8936t7268) I(R8937t290) I(R8937t308) I(R8937t5983) I(R8937t8265) I(R8938t7167) I(R8938t3702) I(R8938t7670) I(R8938t6629) I(R8938t287) I(R8939t2429) I(R8939t4874) I(R8939t7630) I(R8939t6975) I(R8939t3567) I(R8939t296) I(R8940t5558) I(R8940t5791) I(R8940t8100) I(R8940t183) I(R8940t738) I(R8940t1281) I(R8941t4947) I(R8941t8634) I(R8941t5598) I(R8941t5530) I(R8942t4067) I(R8942t8912) I(R8942t8911) I(R8942t7330) I(R8942t381) I(R8942t7300) I(R8942t6244) I(R8942t3827) I(R8943t7501) I(R8943t8825) I(R8943t369) I(R8943t5280) I(R8943t7974) I(R8944t2524) I(R8944t3984) I(R8944t109) I(R8944t4152) I(R8944t8179) I(R8945t2492) I(R8945t6838) I(R8945t8566) I(R8945t4707) I(R8945t7382) I(R8946t7031) I(R8946t6316) I(R8947t202) I(R8947t8330) I(R8947t8832) I(R8947t4359) I(R8947t3646) I(R8947t191) I(R8947t2647) I(R8948t4332) I(R8948t8367) I(R8948t8139) I(R8948t75) I(R8948t4463) I(R8948t3731) I(R8948t3797) I(R8949t276) I(R8949t3992) I(R8949t8508) I(R8949t4300) I(R8950t3591) I(R8950t7342) I(R8950t7626) I(R8950t4943) I(R8950t2186) I(R8950t3714) I(R8950t5546) I(R8951t4263) I(R8951t8798) I(R8951t146) I(R8951t3762) I(R8951t6046) I(R8952t1428) I(R8952t8686) I(R8952t2017) I(R8952t2213) I(R8952t5384) I(R8953t5325) I(R8953t7532) I(R8953t8417) I(R8953t4416) I(R8953t3620) I(R8954t4648) I(R8954t5550) I(R8954t1321) I(R8954t8358) I(R8954t8271) I(R8954t3486) I(R8954t7010) I(R8955t765) I(R8955t1808) I(R8955t8607) I(R8955t4625) I(R8955t4006) I(R8956t5613) I(R8956t7367) I(R8956t5951) I(R8956t2727) I(R8957t7747) I(R8957t5086) I(R8957t3468) I(R8958t966) I(R8958t3290) I(R8958t5780) I(R8958t6327) I(R8958t1731) I(R8959t2318) I(R8959t6788) I(R8959t7598) I(R8959t8311) I(R8959t8929) I(R8959t4140) I(R8960t2361) I(R8960t4972) I(R8960t4532) I(R8960t3133) I(R8961t6435) I(R8961t6532) I(R8961t8463) I(R8961t1911) I(R8961t3468) I(R8961t3660) I(R8962t3463) I(R8962t6883) I(R8962t8356) I(R8962t198) I(R8962t3960) I(R8962t8638) I(R8962t4606) I(R8962t8728) I(R8962t175) I(R8963t1722) I(R8963t3321) I(R8963t4215) I(R8963t6554) I(R8963t5048) I(R8963t3134) I(R8963t7734) I(R8964t376) I(R8964t1464) I(R8964t701) I(R8964t1920) I(R8964t3789) I(R8965t2272) I(R8965t3599) I(R8965t5014) I(R8965t1391) I(R8966t4898) I(R8966t6240) I(R8966t84) I(R8966t5959) I(R8966t5619) I(R8966t1612) I(R8966t573) I(R8966t1818) I(R8967t781) I(R8967t4341) I(R8967t8050) I(R8967t5964) I(R8967t1445) I(R8967t4021) I(R8967t402) I(R8968t2137) I(R8968t8866) I(R8968t2549) I(R8968t3005) I(R8968t8877) I(R8968t8637) I(R8969t1723) I(R8969t6226) I(R8969t6908) I(R8970t649) I(R8970t3545) I(R8970t5848) I(R8970t1171) I(R8971t3027) I(R8971t4085) I(R8971t2289) I(R8971t8557) I(R8971t1126) I(R8972t461) I(R8972t2918) I(R8972t2114) I(R8972t475) I(R8972t3759) I(R8973t2398) I(R8973t4700) I(R8973t6572) I(R8973t4071) I(R8973t3380) I(R8973t8815) I(R8974t2021) I(R8974t4840) I(R8974t6027) I(R8974t5401) I(R8975t5424) I(R8975t6938) I(R8975t3387) I(R8975t5461) I(R8975t2137) I(R8976t2198) I(R8976t6191) I(R8976t278) I(R8976t6966) I(R8976t8187) I(R8976t2095) I(R8977t1642) I(R8977t7117) I(R8977t796) I(R8977t527) I(R8978t1530) I(R8978t7636) I(R8978t137) I(R8978t8409) I(R8978t7257) I(R8978t2471) I(R8978t787) I(R8979t7070) I(R8979t8396) I(R8979t1998) I(R8979t6871) I(R8979t4231) I(R8979t6111) I(R8980t722) I(R8980t2305) I(R8980t4711) I(R8980t4990) I(R8980t2756) I(R8980t4796) I(R8980t5532) I(R8981t4339) I(R8981t7042) I(R8981t424) I(R8981t6331) I(R8981t1752) I(R8982t966) I(R8982t3290) I(R8982t2746) I(R8982t3333) I(R8982t4739) I(R8983t4413) I(R8983t6412) I(R8983t2427) I(R8983t7299) I(R8983t9) I(R8983t7786) I(R8984t554) I(R8984t2426) I(R8984t8123) I(R8984t7007) I(R8984t2822) I(R8985t7328) I(R8985t7554) I(R8985t327) I(R8985t2080) I(R8986t1148) I(R8986t7977) I(R8986t4393) I(R8986t579) I(R8986t7634) I(R8987t3395) I(R8987t6076) I(R8987t4441) I(R8987t1351) I(R8987t8913) I(R8987t4309) I(R8987t2115) I(R8987t5757) I(R8987t5887) I(R8988t5136) I(R8988t8684) I(R8988t8395) I(R8988t6288) I(R8989t1759) I(R8989t4632) I(R8989t1654) I(R8989t4152) I(R8989t6825) I(R8989t2375) I(R8990t5576) I(R8990t7055) I(R8990t6730) I(R8990t8265) I(R8990t8937) I(R8991t1440) I(R8991t3406) I(R8991t2583) I(R8991t516) I(R8991t5226) I(R8991t1013) I(R8991t5160) I(R8991t4116) I(R8992t2782) I(R8992t7594) I(R8992t5362) I(R8992t741) I(R8992t4439) I(R8993t2672) I(R8993t5561) I(R8993t8429) I(R8993t5131) I(R8994t4445) I(R8994t5474) I(R8994t107) I(R8994t2627) I(R8994t2090) I(R8994t7107) I(R8994t6510) I(R8994t7999) I(R8995t4563) I(R8995t6524) I(R8995t2077) I(R8995t3495) I(R8995t5517) I(R8996t5748) I(R8996t508) I(R8997t263) I(R8997t5049) I(R8997t3212) I(R8997t7658) I(R8997t2534) I(R8997t3589) I(R8998t6289) I(R8998t7240) I(R8998t7080) I(R8998t4266) I(R8998t4924) I(R8998t8725) I(R8998t6417) I(R8999t2040) I(R8999t6203) I(R8999t2358) I(R8999t2873) I(R9000t1003) I(R9000t5735) I(R9000t443) I(R9000t49) I(R9000t5667) I(R9000t2665) I(R9001t688) I(R9001t4921) I(R9001t8854) I(R9001t1114) I(R9001t3591) I(R9001t999) I(R9002t306) I(R9002t2026) I(R9002t6477) I(R9002t2979) I(R9002t1807) I(R9002t6555) I(R9003t1540) I(R9003t5704) I(R9003t7843) I(R9003t8568) I(R9003t450) I(R9003t6216) I(R9004t2749) I(R9004t4995) I(R9004t510) I(R9005t4180) I(R9005t8618) I(R9005t4655) I(R9005t979) I(R9005t860) I(R9005t386) I(R9005t5719) I(R9005t1953) I(R9006t622) I(R9006t7478) I(R9006t8797) I(R9006t4043) I(R9006t8012) I(R9006t4653) I(R9006t8186) I(R9006t2349) I(R9007t1220) I(R9007t5453) I(R9007t2080) I(R9007t7701) I(R9008t1875) I(R9008t4597) I(R9008t2907) I(R9008t2767) I(R9008t8187) I(R9008t5951) I(R9009t1452) I(R9009t3629) I(R9009t196) I(R9009t5849) I(R9009t1159) I(R9009t7919) I(R9010t5074) I(R9010t6139) I(R9010t159) I(R9010t601) I(R9010t2564) I(R9010t6033) I(R9011t7157) I(R9011t8011) I(R9011t1370) I(R9011t7696) I(R9011t5896) I(R9011t5761) I(R9012t2327) I(R9012t2495) I(R9012t7375) I(R9012t5113) I(R9012t1582) I(R9012t3934) I(R9012t7631) I(R9012t8748) I(R9012t3748) I(R9013t4232) I(R9013t8225) I(R9013t7481) I(R9013t7660) I(R9013t3883) I(R9013t7035) I(R9013t6982) I(R9013t2213) I(R9013t8141) I(R9014t1560) I(R9014t3072) I(R9014t4019) I(R9014t5024) I(R9015t1447) I(R9015t6365) I(R9015t1521) I(R9015t4146) I(R9016t13) I(R9016t673) I(R9016t4554) I(R9016t652) I(R9016t1109) I(R9017t3672) I(R9017t6472) I(R9017t3837) I(R9017t5110) I(R9017t6595) I(R9017t108) I(R9018t1650) I(R9018t7490) I(R9018t5490) I(R9018t4362) I(R9018t2595) I(R9018t6002) I(R9019t1355) I(R9019t6958) I(R9019t5308) I(R9019t2752) I(R9019t3151) I(R9019t6060) I(R9019t4841) I(R9020t2551) I(R9020t6545) I(R9020t6769) I(R9020t8090) I(R9020t6813) I(R9021t1086) I(R9021t3407) I(R9021t1254) I(R9021t7356) I(R9021t1024) I(R9022t2393) I(R9022t8781) I(R9022t680) I(R9022t3997) I(R9022t5466) I(R9022t532) I(R9023t5652) I(R9023t8073) I(R9023t2673) I(R9023t2958) I(R9023t4740) I(R9024t335) I(R9024t7564) I(R9024t1172) I(R9024t4165) I(R9025t1765) I(R9025t2167) I(R9025t2450) I(R9025t824) I(R9025t1601) I(R9025t4008) I(R9026t716) I(R9026t7387) I(R9026t994) I(R9026t2983) I(R9026t1194) I(R9026t1525) I(R9027t2272) I(R9027t7303) I(R9027t1442) I(R9028t1876) I(R9028t6519) I(R9028t2855) I(R9028t7681) I(R9028t1038) I(R9029t1905) I(R9029t4551) I(R9029t2166) I(R9029t5697) I(R9029t2058) I(R9030t5510) I(R9030t5784) I(R9030t368) I(R9030t2325) I(R9030t2934) I(R9030t134) I(R9030t8355) I(R9031t1778) I(R9031t8297) I(R9031t2493) I(R9031t140) I(R9031t3986) I(R9031t4545) I(R9031t3173) I(R9031t7410) I(R9032t7139) I(R9032t8082) I(R9032t8334) I(R9032t3297) I(R9032t4351) I(R9032t1075) I(R9032t1066) I(R9032t1845) I(R9032t1496) I(R9033t3084) I(R9033t8767) I(R9033t2073) I(R9033t7936) I(R9033t3668) I(R9033t2946) I(R9033t2829) I(R9033t4671) I(R9034t6911) I(R9034t37) I(R9034t6699) I(R9034t4287) I(R9034t1250) I(R9035t8178) I(R9035t7683) I(R9035t6424) I(R9035t3550) I(R9036t2926) I(R9036t7343) I(R9036t5401) I(R9036t2303) I(R9036t3444) I(R9036t6132) I(R9036t6495) I(R9037t1994) I(R9037t4455) I(R9037t7402) I(R9037t6640) I(R9037t4201) I(R9037t4916) I(R9038t4033) I(R9038t8175) I(R9038t8640) I(R9038t8922) I(R9038t514) I(R9038t6850) I(R9038t3665) I(R9039t4423) I(R9039t5614) I(R9039t2567) I(R9039t444) I(R9039t4812) I(R9039t1083) I(R9040t3132) I(R9040t6202) I(R9040t5349) I(R9040t7958) I(R9040t38) I(R9040t8706) I(R9041t5441) I(R9041t6204) I(R9042t230) I(R9042t1415) I(R9042t1421) I(R9042t2840) I(R9042t2947) I(R9042t5000) I(R9043t2574) I(R9043t8548) I(R9043t4089) I(R9043t7616) I(R9043t4689) I(R9044t6154) I(R9044t6984) I(R9044t703) I(R9044t1857) I(R9044t6853) I(R9044t4045) I(R9045t3331) I(R9045t4821) I(R9045t3867) I(R9045t8239) I(R9045t7798) I(R9045t5344) I(R9045t6560) I(R9046t3751) I(R9046t7713) I(R9046t949) I(R9046t8032) I(R9046t7441) I(R9047t3493) I(R9047t4004) I(R9047t4963) I(R9048t6374) I(R9048t8894) I(R9048t2412) I(R9048t5786) I(R9049t663) I(R9049t3201) I(R9049t6190) I(R9049t8826) I(R9049t6388) I(R9049t1135) I(R9050t6723) I(R9050t6768) I(R9050t4414) I(R9050t6706) I(R9050t8900) I(R9050t1784) I(R9051t2318) I(R9051t8959) I(R9051t1245) I(R9051t3857) I(R9051t6788) I(R9052t206) I(R9052t8881) I(R9052t2489) I(R9052t102) I(R9052t5108) I(R9052t842) I(R9053t590) I(R9053t4822) I(R9053t7126) I(R9053t6925) I(R9053t1358) I(R9053t4661) I(R9054t3230) I(R9054t6451) I(R9054t6909) I(R9054t6558) I(R9054t1440) I(R9055t1366) I(R9055t5436) I(R9055t5245) I(R9055t2164) I(R9055t1181) I(R9055t3235) I(R9056t257) I(R9056t6468) I(R9056t1949) I(R9056t3006) I(R9056t8230) I(R9056t761) I(R9057t1063) I(R9057t4356) I(R9057t7095) I(R9057t8372) I(R9057t7152) I(R9058t8393) I(R9058t8510) I(R9058t5419) I(R9058t2857) I(R9058t4491) I(R9058t1809) I(R9058t3688) I(R9059t714) I(R9059t3756) I(R9059t2515) I(R9059t8384) I(R9059t4506) I(R9059t7496) I(R9059t1308) I(R9059t731) I(R9060t701) I(R9060t2739) I(R9060t3831) I(R9061t743) I(R9061t8834) I(R9061t666) I(R9061t6677) I(R9061t7959) I(R9062t8173) I(R9062t8837) I(R9062t4051) I(R9062t3049) I(R9062t5551) I(R9062t4508) I(R9062t615) I(R9063t6110) I(R9063t4205) I(R9063t4470) I(R9063t8661) I(R9063t6780) I(R9063t4911) I(R9064t5979) I(R9064t6350) I(R9064t3679) I(R9064t7469) I(R9064t2238) I(R9064t6625) I(R9064t1423) I(R9064t7093) I(R9065t1363) I(R9065t7947) I(R9065t8614) I(R9065t4819) I(R9066t5805) I(R9066t6600) I(R9066t1619) I(R9066t4150) I(R9067t2242) I(R9067t8761) I(R9067t6017) I(R9067t3774) I(R9067t7091) I(R9068t3674) I(R9068t4220) I(R9068t6797) I(R9068t5289) I(R9068t1337) I(R9069t2182) I(R9069t8144) I(R9069t4835) I(R9069t6470) I(R9069t3542) I(R9069t2123) I(R9069t2584) I(R9070t3652) I(R9070t8649) I(R9070t7452) I(R9070t1305) I(R9070t7694) I(R9070t1569) I(R9070t837) I(R9071t3604) I(R9071t6110) I(R9071t8556) I(R9071t4205) I(R9071t9063) I(R9072t885) I(R9072t5389) I(R9072t3096) I(R9072t6063) I(R9072t3324) I(R9072t7862) I(R9073t2563) I(R9073t5382) I(R9073t8349) I(R9073t7815) I(R9073t5777) I(R9073t1656) I(R9074t5789) I(R9074t6384) I(R9074t2196) I(R9074t6789) I(R9074t4769) I(R9075t7039) I(R9075t7757) I(R9075t7050) I(R9075t5870) I(R9076t5699) I(R9076t8477) I(R9076t3224) I(R9076t1144) I(R9076t6742) I(R9077t1693) I(R9077t8591) I(R9077t3499) I(R9077t8169) I(R9077t1802) I(R9078t384) I(R9078t2330) I(R9078t8629) I(R9079t2758) I(R9079t7867) I(R9079t4409) I(R9079t7704) I(R9079t2925) I(R9079t2304) I(R9080t1552) I(R9080t5345) I(R9080t3325) I(R9080t5291) I(R9080t3847) I(R9080t4890) I(R9080t8357) I(R9081t5435) I(R9081t7361) I(R9081t6691) I(R9081t5393) I(R9082t2215) I(R9082t5413) I(R9082t1756) I(R9082t6688) I(R9082t7723) I(R9083t8109) I(R9083t7766) I(R9083t7244) I(R9083t5301) I(R9084t272) I(R9084t5586) I(R9084t584) I(R9084t8685) I(R9084t3757) I(R9084t787) I(R9084t7851) I(R9085t209) I(R9085t7614) I(R9085t6749) I(R9085t2432) I(R9085t6885) I(R9086t1303) I(R9086t4562) I(R9086t5771) I(R9086t2219) I(R9086t8296) I(R9087t6473) I(R9087t7051) I(R9087t6426) I(R9087t4342) I(R9087t7059) I(R9087t864) I(R9088t3115) I(R9088t5946) I(R9088t5970) I(R9088t3192) I(R9088t8839) I(R9088t66) I(R9089t1695) I(R9089t6241) I(R9089t4072) I(R9089t1041) I(R9089t5366) I(R9090t2388) I(R9090t6149) I(R9090t6472) I(R9090t3837) I(R9090t818) I(R9091t3320) I(R9091t7041) I(R9091t3622) I(R9091t6689) I(R9092t1653) I(R9092t6142) I(R9092t7110) I(R9092t2537) I(R9092t3991) I(R9093t217) I(R9093t2263) I(R9093t1634) I(R9093t7381) I(R9093t8720) I(R9093t1543) I(R9093t2401) I(R9093t6098) I(R9094t779) I(R9094t4217) I(R9094t8702) I(R9094t1792) I(R9095t3821) I(R9095t4308) I(R9095t4396) I(R9095t8264) I(R9095t6782) I(R9095t7768) I(R9095t6957) I(R9095t5655) I(R9096t1686) I(R9096t3392) I(R9096t5989) I(R9096t2031) I(R9096t4211) I(R9096t7916) I(R9096t4513) I(R9096t7800) I(R9097t7624) I(R9097t8146) I(R9097t440) I(R9097t7873) I(R9098t2876) I(R9098t6682) I(R9098t7639) I(R9098t5243) I(R9098t7197) I(R9098t7799) I(R9099t2761) I(R9099t4450) I(R9099t8275) I(R9099t7290) I(R9099t1312) I(R9099t220) I(R9100t4061) I(R9100t6952) I(R9100t7768) I(R9100t4401) I(R9100t4021) I(R9101t8036) I(R9101t1047) I(R9101t3341) I(R9102t5736) I(R9102t7653) I(R9102t7685) I(R9102t8875) I(R9102t5082) I(R9102t3320) I(R9103t568) I(R9103t3060) I(R9103t3616) I(R9103t7907) I(R9103t8059) I(R9104t1475) I(R9104t8789) I(R9104t8857) I(R9104t3793) I(R9104t1909) I(R9104t2892) I(R9104t3277) I(R9104t3481) I(R9105t2361) I(R9105t8960) I(R9105t3133) I(R9105t8652) I(R9105t6073) I(R9105t4799) I(R9105t8659) I(R9106t4003) I(R9106t4167) I(R9106t756) I(R9106t384) I(R9106t9078) I(R9106t2330) I(R9106t5166) I(R9106t8153) I(R9107t3441) I(R9107t6805) I(R9107t4278) I(R9107t8656) I(R9107t2630) I(R9108t3580) I(R9108t7490) I(R9108t1252) I(R9108t5370) I(R9108t2595) I(R9108t6002) I(R9109t375) I(R9109t6133) I(R9109t6803) I(R9109t1055) I(R9109t7399) I(R9110t1058) I(R9110t8301) I(R9110t1329) I(R9110t6992) I(R9110t5050) I(R9111t308) I(R9111t5922) I(R9111t8023) I(R9111t165) I(R9112t3257) I(R9112t6891) I(R9112t1103) I(R9112t7491) I(R9112t1152) I(R9113t1796) I(R9113t3726) I(R9113t7779) I(R9113t6014) I(R9113t2639) I(R9113t6496) I(R9114t4742) I(R9114t7837) I(R9114t5351) I(R9114t6474) I(R9114t6075) I(R9114t479) I(R9115t1302) I(R9115t2405) I(R9115t2836) I(R9115t3791) I(R9115t3131) I(R9116t3391) I(R9116t4374) I(R9116t5773) I(R9116t8368) I(R9117t3159) I(R9117t5510) I(R9117t8193) I(R9117t4058) I(R9117t2390) I(R9117t3047) I(R9117t4164) I(R9117t8492) I(R9117t5784) I(R9118t2043) I(R9118t4009) I(R9118t1270) I(R9118t4798) I(R9118t902) I(R9118t6257) I(R9119t1375) I(R9119t6656) I(R9119t7238) I(R9119t5939) I(R9119t5868) I(R9120t6374) I(R9120t9048) I(R9120t7919) I(R9120t3629) I(R9120t8636) I(R9120t5299) I(R9120t8894) I(R9121t1470) I(R9121t5158) I(R9121t6198) I(R9121t16) I(R9121t3371) I(R9122t4449) I(R9122t7252) I(R9122t3681) I(R9122t1110) I(R9122t4082) I(R9122t4355) I(R9123t360) I(R9123t3164) I(R9123t7785) I(R9123t6567) I(R9123t2529) I(R9123t2681) I(R9124t230) I(R9124t3153) I(R9124t204) I(R9124t3519) I(R9124t1415) I(R9125t4255) I(R9125t5279) I(R9125t2189) I(R9125t2072) I(R9125t6369) I(R9125t8726) I(R9126t3380) I(R9126t6170) I(R9126t7003) I(R9126t7571) I(R9126t4905) I(R9126t2536) I(R9126t7000) I(R9126t253) I(R9126t1410) I(R9127t5016) I(R9127t8633) I(R9127t4365) I(R9127t3882) I(R9127t2833) I(R9127t930) I(R9128t2351) I(R9128t7293) I(R9128t3657) I(R9128t6348) I(R9128t1887) I(R9129t1269) I(R9129t8909) I(R9129t3460) I(R9129t6988) I(R9129t2068) I(R9129t7981) I(R9129t8892) I(R9130t6108) I(R9130t7195) I(R9130t3666) I(R9130t3496) I(R9131t554) I(R9131t7872) I(R9131t182) I(R9131t8803) I(R9131t2822) I(R9132t2498) I(R9132t6103) I(R9132t2169) I(R9132t8129) I(R9132t5104) I(R9132t4988) I(R9133t6377) I(R9133t8216) I(R9133t2806) I(R9133t5021) I(R9133t4279) I(R9133t2380) I(R9133t240) I(R9134t300) I(R9134t4415) I(R9134t3189) I(R9134t6460) I(R9135t4904) I(R9135t7474) I(R9135t2933) I(R9135t6875) I(R9135t7524) I(R9135t7492) I(R9136t650) I(R9136t3839) I(R9136t203) I(R9136t7985) I(R9137t4472) I(R9137t4224) I(R9137t7639) I(R9137t9098) I(R9138t632) I(R9138t4788) I(R9138t508) I(R9138t6831) I(R9139t3471) I(R9139t6100) I(R9139t7650) I(R9139t5659) I(R9139t2312) I(R9140t4431) I(R9140t703) I(R9140t9044) I(R9140t1857) I(R9140t3427) I(R9141t4844) I(R9141t5729) I(R9141t4686) I(R9141t527) I(R9141t8977) I(R9141t1642) I(R9141t6208) I(R9142t8720) I(R9142t9093) I(R9142t1543) I(R9142t7899) I(R9143t1312) I(R9143t2776) I(R9143t3680) I(R9143t8734) I(R9144t2378) I(R9144t2967) I(R9144t3497) I(R9144t6439) I(R9144t3784) I(R9145t3550) I(R9145t6151) I(R9145t9035) I(R9145t8178) I(R9145t7507) I(R9145t2209) I(R9146t4696) I(R9146t5381) I(R9146t1656) I(R9146t5777) I(R9146t6840) I(R9147t2560) I(R9147t7565) I(R9147t1577) I(R9147t5282) I(R9147t4210) I(R9147t8112) I(R9148t577) I(R9148t8762) I(R9148t1989) I(R9148t873) I(R9148t1601) I(R9148t3433) I(R9149t1614) I(R9149t4259) I(R9149t4707) I(R9149t715) I(R9149t2891) I(R9149t7597) I(R9149t8802) I(R9149t6837) I(R9149t2861) I(R9150t7039) I(R9150t9075) I(R9150t6429) I(R9150t6861) I(R9150t1528) I(R9150t7757) I(R9151t7718) I(R9151t7882) I(R9152t2563) I(R9152t6058) I(R9152t3683) I(R9153t5086) I(R9153t8957) I(R9153t4433) I(R9153t7836) I(R9153t6226) I(R9153t8969) I(R9153t6908) I(R9153t3468) I(R9154t4453) I(R9154t7728) I(R9154t5574) I(R9154t7349) I(R9155t4502) I(R9155t5221) I(R9155t2383) I(R9155t999) I(R9155t9001) I(R9155t3591) I(R9156t1615) I(R9156t6809) I(R9156t3877) I(R9156t5499) I(R9156t5718) I(R9156t1869) I(R9156t1472) I(R9157t698) I(R9157t1595) I(R9157t8650) I(R9157t2580) I(R9157t2961) I(R9157t2002) I(R9157t4136) I(R9157t1485) I(R9158t1815) I(R9158t3579) I(R9159t1420) I(R9159t634) I(R9159t3368) I(R9159t2700) I(R9160t1899) I(R9160t5183) I(R9160t4240) I(R9160t5530) I(R9160t4947) I(R9161t1332) I(R9161t3274) I(R9161t3970) I(R9161t5496) I(R9161t3208) I(R9162t3964) I(R9162t2216) I(R9162t7042) I(R9162t6328) I(R9163t1332) I(R9163t3274) I(R9163t1718) I(R9163t7028) I(R9164t303) I(R9164t13) I(R9164t9016) I(R9165t1085) I(R9165t2079) I(R9165t8454) I(R9165t2224) I(R9165t5413) I(R9165t7723) I(R9166t6328) I(R9166t6767) I(R9166t9162) I(R9166t3964) I(R9166t5232) I(R9166t5601) I(R9167t1545) I(R9167t1739) I(R9167t947) I(R9167t6325) I(R9167t6259) I(R9167t8506) I(R9167t5098) I(R9168t1593) I(R9168t3247) I(R9168t668) I(R9168t2052) I(R9169t3298) I(R9169t5560) I(R9169t8526) I(R9169t3222) I(R9170t806) I(R9170t384) I(R9170t9106) I(R9170t756) I(R9170t3931) I(R9171t1718) I(R9171t3751) I(R9171t9163) I(R9171t7028) I(R9171t7332) I(R9172t4935) I(R9172t7290) I(R9172t1312) I(R9172t9143) I(R9172t3680) I(R9173t541) I(R9173t5075) I(R9173t1202) I(R9173t2371) I(R9173t2011) I(R9174t4905) I(R9174t7571) I(R9174t2717) I(R9174t564) I(R9174t6) I(R9174t799) I(R9174t4071) I(R9174t7003) I(R9175t1692) I(R9175t7238) I(R9175t1375) I(R9175t8600) I(R9176t7370) I(R9176t8221) I(R9176t7866) I(R9176t6269) I(R9176t1455) I(R9176t5349) I(R9176t4274) I(R9177t711) I(R9177t7667) I(R9177t2477) I(R9177t8927) I(R9177t2967) I(R9177t3784) I(R9178t2623) I(R9178t4424) I(R9178t4660) I(R9178t994) I(R9178t1736) I(R9178t5629) I(R9178t6540) I(R9178t5171) I(R9179t6444) I(R9179t7072) I(R9179t768) I(R9179t8114) I(R9179t2081) I(R9179t2373) I(R9180t6081) I(R9180t6720) I(R9180t20) I(R9180t7186) I(R9180t2737) I(R9180t5143) I(R9181t1822) I(R9181t3738) I(R9181t7069) I(R9181t2485) I(R9181t3130) I(R9181t1917) I(R9182t2360) I(R9182t3090) I(R9182t2438) I(R9182t2301) I(R9183t1098) I(R9183t3871) I(R9183t7210) I(R9183t391) I(R9184t6096) I(R9184t6740) I(R9184t4448) I(R9184t7917) I(R9185t5700) I(R9185t7267) I(R9185t828) I(R9185t7576) I(R9185t1232) I(R9185t6841) I(R9186t1544) I(R9186t5045) I(R9186t4321) I(R9186t3590) I(R9186t8524) I(R9187t6447) I(R9187t6873) I(R9187t8544) I(R9187t2087) I(R9187t1129) I(R9187t2254) I(R9188t1680) I(R9188t7014) I(R9188t7405) I(R9188t8104) I(R9188t5994) I(R9188t2008) I(R9188t4701) I(R9189t8264) I(R9189t7539) I(R9189t8704) I(R9189t1052) I(R9189t6271) I(R9189t1698) I(R9190t2133) I(R9190t3404) I(R9190t6676) I(R9190t7540) I(R9190t5969) I(R9191t3260) I(R9191t4946) I(R9191t3303) I(R9191t1082) I(R9191t7912) I(R9191t4600) I(R9192t6268) I(R9192t8321) I(R9192t7766) I(R9192t9083) I(R9192t8109) I(R9193t5637) I(R9193t6727) I(R9193t189) I(R9193t7325) I(R9193t8350) I(R9193t6511) I(R9194t2914) I(R9194t5522) I(R9194t6894) I(R9194t5692) I(R9194t5095) I(R9195t64) I(R9195t3072) I(R9195t245) I(R9195t460) I(R9196t46) I(R9196t289) I(R9196t4483) I(R9196t2650) I(R9196t8611) I(R9197t1514) I(R9197t3703) I(R9197t3199) I(R9197t6089) I(R9197t8328) I(R9197t7123) I(R9197t5957) I(R9198t295) I(R9198t4927) I(R9198t5246) I(R9198t1350) I(R9198t872) I(R9199t926) I(R9199t7754) I(R9199t1594) I(R9199t6062) I(R9199t5206) I(R9200t695) I(R9200t5802) I(R9200t3129) I(R9200t5422) I(R9200t1372) I(R9201t4924) I(R9201t5329) I(R9201t8725) I(R9201t3510) I(R9201t1156) I(R9201t7145) I(R9202t413) I(R9202t6176) I(R9202t4485) I(R9202t7829) I(R9202t7732) I(R9202t5769) I(R9202t8703) I(R9203t4586) I(R9203t7307) I(R9203t7877) I(R9203t8045) I(R9203t40) I(R9203t5437) I(R9204t3085) I(R9204t6933) I(R9204t5574) I(R9204t3384) I(R9204t2259) I(R9205t6167) I(R9205t4012) I(R9205t5463) I(R9205t5309) I(R9205t8697) I(R9206t1107) I(R9206t1527) I(R9206t1329) I(R9206t4012) I(R9206t9205) I(R9206t6167) I(R9207t8) I(R9207t3026) I(R9207t6460) I(R9207t3802) I(R9208t5658) I(R9208t7463) I(R9208t1762) I(R9208t7909) I(R9208t7631) I(R9209t6688) I(R9209t8065) I(R9209t8151) I(R9209t3852) I(R9209t6062) I(R9209t469) I(R9209t5689) I(R9209t4615) I(R9210t2707) I(R9210t6130) I(R9210t2297) I(R9210t506) I(R9211t171) I(R9211t4509) I(R9211t2482) I(R9211t8780) I(R9211t2715) I(R9211t7377) I(R9211t1531) I(R9211t7078) I(R9212t7138) I(R9212t8523) I(R9212t4362) I(R9212t1889) I(R9212t42) I(R9213t2714) I(R9213t4464) I(R9213t6485) I(R9213t2099) I(R9213t952) I(R9214t5821) I(R9214t8077) I(R9214t3126) I(R9214t5111) I(R9214t8709) I(R9215t7882) I(R9215t4510) I(R9215t4870) I(R9215t6523) I(R9215t7718) I(R9215t9151) I(R9216t2664) I(R9216t5266) I(R9216t96) I(R9216t4256) I(R9216t1763) I(R9216t7257) I(R9217t2715) I(R9217t6862) I(R9217t151) I(R9217t6164) I(R9217t7450) I(R9217t904) I(R9218t2006) I(R9218t4651) I(R9218t8032) I(R9218t949) I(R9218t4676) I(R9219t4364) I(R9219t6289) I(R9219t6167) I(R9219t9205) I(R9219t8697) I(R9219t6884) I(R9219t7413) I(R9220t1205) I(R9220t4370) I(R9220t4762) I(R9220t2311) I(R9220t7759) I(R9220t512) I(R9220t1833) I(R9221t1089) I(R9221t6551) I(R9221t6188) I(R9221t6237) I(R9221t1286) I(R9221t90) I(R9221t4757) I(R9222t1750) I(R9222t4097) I(R9222t4605) I(R9222t6291) I(R9222t5229) I(R9223t1086) I(R9223t9021) I(R9223t3407) I(R9223t6373) I(R9223t2005) I(R9223t8140) I(R9224t1831) I(R9224t4673) I(R9224t6297) I(R9224t950) I(R9225t5258) I(R9225t7812) I(R9226t491) I(R9226t6173) I(R9226t7043) I(R9226t3795) I(R9226t8019) I(R9226t526) I(R9227t4802) I(R9227t6178) I(R9227t1209) I(R9227t7419) I(R9227t4206) I(R9227t8201) I(R9228t2327) I(R9228t7375) I(R9228t771) I(R9228t5113) I(R9229t2927) I(R9229t2967) I(R9229t510) I(R9229t9004) I(R9229t2749) I(R9229t2378) I(R9230t1447) I(R9230t9015) I(R9230t2158) I(R9230t3873) I(R9230t121) I(R9230t6723) I(R9230t7181) I(R9230t4146) I(R9231t4245) I(R9231t4606) I(R9231t8728) I(R9231t751) I(R9232t7230) I(R9232t8442) I(R9232t6669) I(R9232t1970) I(R9232t3216) I(R9233t16) I(R9233t9121) I(R9233t6198) I(R9233t6399) I(R9233t1855) I(R9233t5913) I(R9234t4492) I(R9234t7263) I(R9234t8659) I(R9234t2361) I(R9235t1805) I(R9235t8015) I(R9235t5205) I(R9235t7031) I(R9235t8946) I(R9235t6316) I(R9236t4717) I(R9236t4930) I(R9236t6823) I(R9236t1846) I(R9236t4875) I(R9237t299) I(R9237t8389) I(R9237t4727) I(R9237t2908) I(R9237t3556) I(R9238t1561) I(R9238t4872) I(R9238t1785) I(R9238t7974) I(R9239t5518) I(R9239t7644) I(R9239t585) I(R9239t3312) I(R9239t4863) I(R9239t4544) I(R9239t5224) I(R9240t2441) I(R9240t2478) I(R9240t2917) I(R9240t7718) I(R9240t9215) I(R9240t6523) I(R9240t6679) I(R9241t2384) I(R9241t5648) I(R9241t2783) I(R9241t7643) I(R9242t3023) I(R9242t4852) I(R9242t2335) I(R9242t8323) I(R9242t2683) I(R9243t813) I(R9243t2687) I(R9243t6694) I(R9243t6273) I(R9243t7737) I(R9244t7083) I(R9244t7764) I(R9244t8046) I(R9244t2905) I(R9244t1788) I(R9245t2923) I(R9245t3411) I(R9245t5987) I(R9245t1900) I(R9245t1608) I(R9246t2419) I(R9246t6695) I(R9246t4440) I(R9246t4961) I(R9246t2699) I(R9246t8524) I(R9247t908) I(R9247t7732) I(R9247t5769) I(R9247t8148) I(R9247t1885) I(R9247t388) I(R9247t3616) I(R9247t8763) I(R9248t5563) I(R9248t8219) I(R9248t3557) I(R9248t4860) I(R9248t5577) I(R9248t2654) I(R9248t8567) I(R9249t4696) I(R9249t5618) I(R9249t7852) I(R9249t1656) I(R9249t9146) I(R9250t3003) I(R9250t6980) I(R9250t1224) I(R9250t7331) I(R9251t1426) I(R9251t6381) I(R9251t6929) I(R9251t2191) I(R9251t8800) I(R9251t6092) I(R9252t6614) I(R9252t3533) I(R9252t237) I(R9252t7879) I(R9253t2274) I(R9253t7970) I(R9253t3775) I(R9253t7142) I(R9253t4406) I(R9253t1138) I(R9253t3746) I(R9254t3621) I(R9254t8402) I(R9254t6718) I(R9254t6643) I(R9254t8564) I(R9254t4039) I(R9255t6182) I(R9255t8595) I(R9255t7306) I(R9255t1594) I(R9255t9199) I(R9255t926) I(R9256t3940) I(R9256t7174) I(R9256t2345) I(R9256t7948) I(R9256t5128) I(R9256t1875) I(R9257t7929) I(R9257t8122) I(R9257t2400) I(R9257t1316) I(R9257t162) I(R9257t2751) I(R9258t3883) I(R9258t4185) I(R9258t4191) I(R9258t2456) I(R9258t8408) I(R9258t466) I(R9259t3921) I(R9259t5117) I(R9259t8870) I(R9260t2758) I(R9260t7867) I(R9260t4892) I(R9260t2819) I(R9260t4121) I(R9260t1196) I(R9261t6004) I(R9261t6415) I(R9261t2364) I(R9261t3018) I(R9262t1167) I(R9262t2467) I(R9262t1854) I(R9262t6596) I(R9262t4056) I(R9262t6547) I(R9262t5573) I(R9263t3276) I(R9263t3374) I(R9263t1664) I(R9263t4709) I(R9263t4516) I(R9264t5464) I(R9264t7462) I(R9264t4113) I(R9264t4155) I(R9265t188) I(R9265t428) I(R9265t856) I(R9265t4598) I(R9265t4640) I(R9265t6692) I(R9265t7202) I(R9266t4543) I(R9266t6321) I(R9266t524) I(R9266t2896) I(R9266t5449) I(R9267t4706) I(R9267t8818) I(R9267t890) I(R9267t5690) I(R9267t260) I(R9267t3684) I(R9268t2337) I(R9268t2774) I(R9268t1498) I(R9268t7962) I(R9268t6836) I(R9268t5689) I(R9269t4039) I(R9269t6443) I(R9269t3872) I(R9269t5294) I(R9270t2886) I(R9270t7277) I(R9270t7320) I(R9270t4611) I(R9270t8078) I(R9270t4886) I(R9271t2390) I(R9271t8883) I(R9271t6458) I(R9271t153) I(R9271t4752) I(R9271t8606) I(R9271t556) I(R9271t8325) I(R9272t1048) I(R9272t7677) I(R9272t3778) I(R9272t6353) I(R9272t4252) I(R9272t6197) I(R9272t6703) I(R9273t4354) I(R9273t6896) I(R9273t3776) I(R9273t7995) I(R9273t4637) I(R9274t4151) I(R9274t5452) I(R9274t2585) I(R9274t5087) I(R9274t965) I(R9274t1533) I(R9274t7879) I(R9274t237) I(R9275t575) I(R9275t6029) I(R9275t4130) I(R9275t2532) I(R9275t7744) I(R9275t977) I(R9276t973) I(R9276t3733) I(R9276t5961) I(R9276t2396) I(R9277t7025) I(R9277t7397) I(R9277t6380) I(R9278t226) I(R9278t1026) I(R9278t3065) I(R9278t1892) I(R9278t8722) I(R9279t3968) I(R9279t4451) I(R9279t3349) I(R9280t2) I(R9280t4784) I(R9280t3086) I(R9280t7407) I(R9281t6090) I(R9281t8791) I(R9281t6345) I(R9281t7351) I(R9281t6445) I(R9282t211) I(R9282t8490) I(R9282t808) I(R9282t4064) I(R9282t7997) I(R9282t1509) I(R9283t2616) I(R9283t7408) I(R9283t3771) I(R9283t5703) I(R9283t4917) I(R9283t1600) I(R9283t7619) I(R9284t2507) I(R9284t2625) I(R9284t1947) I(R9284t2818) I(R9284t3600) I(R9284t1570) I(R9285t8742) I(R9285t8886) I(R9285t2039) I(R9285t3839) I(R9285t9136) I(R9285t203) I(R9285t7967) I(R9286t3583) I(R9286t5881) I(R9286t6410) I(R9286t4937) I(R9286t7519) I(R9286t5244) I(R9287t5850) I(R9287t6893) I(R9287t6267) I(R9287t7449) I(R9287t3302) I(R9287t4249) I(R9287t6685) I(R9287t5603) I(R9287t4765) I(R9287t4823) I(R9288t871) I(R9288t8844) I(R9288t69) I(R9288t3791) I(R9288t194) I(R9288t8478) I(R9288t5208) I(R9289t8501) I(R9289t3149) I(R9289t7329) I(R9289t8036) I(R9289t9101) I(R9289t1047) I(R9290t5450) I(R9290t5542) I(R9290t6607) I(R9290t4914) I(R9291t7263) I(R9291t9234) I(R9291t2361) I(R9291t7859) I(R9291t7708) I(R9291t3958) I(R9291t6817) I(R9291t5625) I(R9292t179) I(R9292t6364) I(R9292t1541) I(R9292t8729) I(R9292t5999) I(R9292t236) I(R9293t4410) I(R9293t7314) I(R9293t7154) I(R9293t7243) I(R9293t5356) I(R9293t3998) I(R9294t8277) I(R9294t8699) I(R9294t6411) I(R9294t7498) I(R9294t616) I(R9294t2413) I(R9295t3427) I(R9295t4431) I(R9295t945) I(R9295t3038) I(R9295t703) I(R9295t9140) I(R9296t1090) I(R9296t8773) I(R9297t6511) I(R9297t8350) I(R9297t6379) I(R9297t7620) I(R9297t550) I(R9297t7305) I(R9298t5565) I(R9298t7057) I(R9298t8404) I(R9298t1923) I(R9298t8710) I(R9298t2012) I(R9298t3464) I(R9298t7284) I(R9299t891) I(R9299t6999) I(R9299t2435) I(R9299t7224) I(R9300t2926) I(R9300t5364) I(R9300t6495) I(R9300t9036) I(R9301t684) I(R9301t8535) I(R9301t5985) I(R9301t553) I(R9301t3481) I(R9301t8808) I(R9302t1679) I(R9302t6976) I(R9302t6995) I(R9302t8486) I(R9302t154) I(R9303t3221) I(R9303t5500) I(R9303t7575) I(R9303t809) I(R9303t5123) I(R9303t2521) I(R9304t51) I(R9304t6667) I(R9304t3409) I(R9304t1463) I(R9304t8130) I(R9304t4825) I(R9305t3997) I(R9305t9022) I(R9305t680) I(R9305t3528) I(R9305t3275) I(R9306t2835) I(R9306t8411) I(R9306t3903) I(R9306t4994) I(R9306t354) I(R9306t8631) I(R9306t5875) I(R9307t6402) I(R9307t6853) I(R9307t3257) I(R9307t8286) I(R9308t197) I(R9308t4154) I(R9308t8654) I(R9308t437) I(R9308t6735) I(R9308t2693) I(R9308t4815) I(R9308t6662) I(R9309t2021) I(R9309t8974) I(R9309t5401) I(R9309t9036) I(R9309t2303) I(R9310t8518) I(R9310t8683) I(R9310t212) I(R9310t7456) I(R9310t3259) I(R9310t4595) I(R9310t484) I(R9311t4293) I(R9311t8578) I(R9311t7580) I(R9311t7074) I(R9311t8572) I(R9312t80) I(R9312t7632) I(R9312t2294) I(R9312t2286) I(R9312t3038) I(R9312t945) I(R9312t5567) I(R9312t4745) I(R9313t3753) I(R9313t6812) I(R9313t8098) I(R9313t6106) I(R9314t491) I(R9314t6173) I(R9314t7670) I(R9314t6629) I(R9314t3106) I(R9314t5010) I(R9314t526) I(R9315t2362) I(R9315t2436) I(R9315t8308) I(R9315t6034) I(R9315t4577) I(R9315t2803) I(R9316t3292) I(R9316t5942) I(R9316t4817) I(R9316t6552) I(R9316t5032) I(R9316t2659) I(R9317t280) I(R9317t1595) I(R9317t7049) I(R9317t2094) I(R9317t5126) I(R9317t3447) I(R9318t2019) I(R9318t3276) I(R9318t6546) I(R9318t7075) I(R9318t5959) I(R9318t5619) I(R9318t6389) I(R9319t4242) I(R9319t7158) I(R9319t8768) I(R9319t7687) I(R9319t6562) I(R9319t1432) I(R9319t4537) I(R9319t1043) I(R9320t2488) I(R9320t8881) I(R9320t2195) I(R9320t4596) I(R9320t3370) I(R9320t5753) I(R9321t2760) I(R9321t3718) I(R9321t7213) I(R9321t330) I(R9321t2215) I(R9321t9082) I(R9321t1756) I(R9321t4615) I(R9322t2394) I(R9322t5429) I(R9322t218) I(R9323t1871) I(R9323t7006) I(R9323t1309) I(R9323t2889) I(R9323t1101) I(R9323t8414) I(R9324t6368) I(R9325t5852) I(R9325t6690) I(R9325t5312) I(R9325t3636) I(R9325t2637) I(R9325t5837) I(R9325t2748) I(R9326t2507) I(R9326t3768) I(R9326t5636) I(R9326t1202) I(R9326t2371) I(R9326t267) I(R9326t2993) I(R9327t4932) I(R9327t1329) I(R9327t5572) I(R9328t1641) I(R9328t1852) I(R9328t2394) I(R9328t8733) I(R9328t5711) I(R9328t5768) I(R9329t1155) I(R9329t4569) I(R9329t2232) I(R9329t4789) I(R9329t7226) I(R9330t2858) I(R9330t3436) I(R9330t7613) I(R9330t935) I(R9331t3115) I(R9331t9088) I(R9331t5970) I(R9331t1370) I(R9331t2183) I(R9332t6590) I(R9332t6614) I(R9332t6969) I(R9332t2288) I(R9332t3533) I(R9332t9252) I(R9333t809) I(R9333t8738) I(R9333t3949) I(R9333t3191) I(R9333t8280) I(R9333t7575) I(R9334t2510) I(R9334t6339) I(R9334t56) I(R9334t975) I(R9335t3914) I(R9335t5215) I(R9336t5215) I(R9336t9335) I(R9336t892) I(R9336t1317) I(R9336t8116) I(R9336t6795) I(R9336t3914) I(R9337t4689) I(R9337t7386) I(R9337t6309) I(R9337t7835) I(R9337t7616) I(R9337t9043) I(R9338t3307) I(R9338t8320) I(R9338t453) I(R9338t4918) I(R9338t8668) I(R9338t4682) I(R9339t6190) I(R9339t9049) I(R9339t248) I(R9339t4233) I(R9339t8826) I(R9340t64) I(R9340t3072) I(R9340t9014) I(R9340t4019) I(R9340t5375) I(R9341t504) I(R9341t792) I(R9341t1867) I(R9341t8725) I(R9341t591) I(R9341t3510) I(R9341t3351) I(R9341t4708) I(R9342t5117) I(R9342t8620) I(R9342t8807) I(R9342t7548) I(R9343t3170) I(R9343t7473) I(R9343t573) I(R9343t8966) I(R9343t1818) I(R9344t2169) I(R9344t8129) I(R9344t505) I(R9344t1753) I(R9344t5739) I(R9344t191) I(R9344t3646) I(R9344t4923) I(R9344t4334) I(R9344t5199) I(R9345t2157) I(R9345t6080) I(R9345t946) I(R9345t954) I(R9345t3016) I(R9345t4706) I(R9345t1137) I(R9346t4138) I(R9346t4344) I(R9346t2523) I(R9346t8507) I(R9346t804) I(R9346t228) I(R9347t1971) I(R9347t9083) I(R9347t7244) I(R9348t3792) I(R9348t6492) I(R9348t414) I(R9348t6388) I(R9348t8826) I(R9348t4539) I(R9348t6491) I(R9349t2020) I(R9349t3005) I(R9349t8815) I(R9349t6170) I(R9349t6747) I(R9350t2901) I(R9350t5405) I(R9350t6649) I(R9350t1195) I(R9351t29) I(R9351t3930) I(R9351t811) I(R9351t3887) I(R9351t5297) I(R9352t2579) I(R9352t7883) I(R9352t8676) I(R9352t5904) I(R9352t7949) I(R9352t6786) I(R9352t8882) I(R9353t5128) I(R9353t7948) I(R9353t4283) I(R9353t4065) I(R9353t1207) I(R9353t5339) I(R9353t4086) I(R9353t7341) I(R9354t2907) I(R9354t9008) I(R9354t1505) I(R9354t4283) I(R9354t5128) I(R9354t9256) I(R9354t1875) I(R9355t8) I(R9355t9207) I(R9355t7775) I(R9355t5324) I(R9355t3026) I(R9356t3279) I(R9356t8430) I(R9356t928) I(R9356t5093) I(R9357t2754) I(R9357t7557) I(R9357t524) I(R9358t364) I(R9358t7011) I(R9358t4549) I(R9358t7652) I(R9358t7065) I(R9359t7374) I(R9359t8557) I(R9359t1126) I(R9360t7395) I(R9360t7860) I(R9360t3229) I(R9360t218) I(R9360t6458) I(R9360t8026) I(R9361t1107) I(R9361t7746) I(R9361t1058) I(R9361t8301) I(R9361t2590) I(R9361t7840) I(R9362t4792) I(R9362t8299) I(R9362t1612) I(R9362t8966) I(R9362t5619) I(R9362t6797) I(R9362t4220) I(R9363t4212) I(R9363t5643) I(R9363t4294) I(R9363t7089) I(R9363t8843) I(R9363t7166) I(R9364t297) I(R9364t1494) I(R9364t6246) I(R9364t6367) I(R9364t5003) I(R9364t4915) I(R9365t5439) I(R9365t6359) I(R9365t5860) I(R9365t4386) I(R9365t1973) I(R9366t4528) I(R9366t8814) I(R9366t2500) I(R9366t3209) I(R9366t460) I(R9367t1870) I(R9367t4135) I(R9367t8293) I(R9367t6228) I(R9367t5292) I(R9367t8632) I(R9368t1602) I(R9368t2855) I(R9368t4957) I(R9368t2101) I(R9368t4728) I(R9369t168) I(R9369t1048) I(R9369t226) I(R9369t9278) I(R9369t8722) I(R9369t1218) I(R9369t746) I(R9370t561) I(R9370t1534) I(R9370t7495) I(R9370t3299) I(R9370t4315) I(R9371t1411) I(R9371t4070) I(R9371t7951) I(R9371t7684) I(R9371t1001) I(R9371t6292) I(R9372t1217) I(R9372t7546) I(R9372t8508) I(R9372t4300) I(R9372t956) I(R9372t6772) I(R9373t4549) I(R9373t6299) I(R9373t7135) I(R9373t797) I(R9373t518) I(R9373t6745) I(R9373t7011) I(R9374t115) I(R9374t4190) I(R9374t2730) I(R9374t8527) I(R9374t1566) I(R9374t7800) I(R9375t3113) I(R9375t4793) I(R9375t5101) I(R9375t1298) I(R9375t7087) I(R9375t249) I(R9376t2465) I(R9376t6510) I(R9376t5391) I(R9376t7107) I(R9376t8994) I(R9377t4834) I(R9377t6898) I(R9377t685) I(R9377t361) I(R9377t1861) I(R9377t7685) I(R9377t9102) I(R9377t8875) I(R9378t4450) I(R9378t9099) I(R9378t8275) I(R9378t4143) I(R9378t5418) I(R9378t834) I(R9379t4932) I(R9379t6084) I(R9379t9327) I(R9379t1329) I(R9379t3677) I(R9379t4088) I(R9379t7033) I(R9380t4732) I(R9380t5965) I(R9380t3782) I(R9380t1255) I(R9380t7096) I(R9380t8156) I(R9381t3544) I(R9381t8142) I(R9381t7812) I(R9381t9225) I(R9381t5258) I(R9382t3530) I(R9382t3594) I(R9382t8923) I(R9382t8328) I(R9382t8771) I(R9382t7941) I(R9382t1804) I(R9383t5426) I(R9383t7182) I(R9383t5257) I(R9383t5888) I(R9383t6487) I(R9384t663) I(R9384t2940) I(R9384t3201) I(R9384t1135) I(R9384t5439) I(R9384t5860) I(R9385t8094) I(R9385t8449) I(R9385t7379) I(R9385t540) I(R9385t2640) I(R9385t2769) I(R9386t2140) I(R9386t2407) I(R9386t3264) I(R9386t2075) I(R9386t210) I(R9386t6345) I(R9386t9281) I(R9386t7351) I(R9387t687) I(R9387t2709) I(R9387t4646) I(R9387t6568) I(R9387t7412) I(R9387t1380) I(R9388t4604) I(R9388t8514) I(R9388t7717) I(R9388t4645) I(R9388t6628) I(R9388t571) I(R9389t2272) I(R9389t8965) I(R9389t1391) I(R9389t9027) I(R9390t448) I(R9390t3523) I(R9390t7268) I(R9390t1916) I(R9390t3939) I(R9390t8021) I(R9391t2553) I(R9391t4375) I(R9391t5993) I(R9391t1260) I(R9391t1249) I(R9392t2671) I(R9392t8669) I(R9392t811) I(R9392t9351) I(R9392t3887) I(R9392t7362) I(R9392t3180) I(R9393t6402) I(R9393t9307) I(R9393t44) I(R9393t6673) I(R9393t8286) I(R9394t3572) I(R9394t7942) I(R9394t5639) I(R9394t7904) I(R9394t1571) I(R9394t7560) I(R9395t5727) I(R9395t8419) I(R9395t5212) I(R9395t1711) I(R9396t1315) I(R9396t7892) I(R9396t1698) I(R9396t9189) I(R9396t8264) I(R9397t7964) I(R9397t8600) I(R9397t9175) I(R9397t1375) I(R9398t2269) I(R9398t3123) I(R9398t1055) I(R9398t3360) I(R9398t8529) I(R9398t8580) I(R9399t982) I(R9399t1568) I(R9399t7435) I(R9399t8459) I(R9399t2188) I(R9399t6663) I(R9399t5032) I(R9399t7001) I(R9400t5172) I(R9400t6670) I(R9400t7770) I(R9400t2678) I(R9401t1844) I(R9401t6419) I(R9401t4755) I(R9401t3412) I(R9401t5012) I(R9402t784) I(R9402t6163) I(R9402t4728) I(R9402t2101) I(R9402t5897) I(R9403t1823) I(R9403t120) I(R9403t4314) I(R9403t3717) I(R9404t2276) I(R9404t6029) I(R9404t4081) I(R9404t611) I(R9404t2460) I(R9404t7094) I(R9404t4130) I(R9405t468) I(R9405t6946) I(R9405t3479) I(R9405t6031) I(R9405t1132) I(R9405t4109) I(R9406t621) I(R9406t7761) I(R9406t7177) I(R9406t6478) I(R9406t6242) I(R9406t4676) I(R9406t4651) I(R9407t1743) I(R9407t7849) I(R9407t1335) I(R9407t1800) I(R9407t5594) I(R9408t1804) I(R9408t7941) I(R9408t3530) I(R9408t3945) I(R9408t3051) I(R9408t8347) I(R9408t5376) I(R9409t5268) I(R9409t7376) I(R9409t4780) I(R9409t7002) I(R9409t4567) I(R9410t1696) I(R9410t7874) I(R9410t1047) I(R9410t9289) I(R9410t8501) I(R9410t5046) I(R9411t1328) I(R9411t7676) I(R9411t6855) I(R9411t2328) I(R9411t2551) I(R9411t163) I(R9412t4325) I(R9412t7852) I(R9412t493) I(R9412t1185) I(R9412t2563) I(R9412t1656) I(R9413t1327) I(R9413t3863) I(R9413t2319) I(R9413t6807) I(R9413t5724) I(R9414t2754) I(R9414t9357) I(R9414t5574) I(R9414t7533) I(R9414t524) I(R9415t1071) I(R9415t5141) I(R9415t2700) I(R9415t3368) I(R9415t3640) I(R9415t2477) I(R9416t4248) I(R9416t7348) I(R9416t4041) I(R9416t1621) I(R9416t4987) I(R9416t1166) I(R9417t4801) I(R9417t6146) I(R9417t2581) I(R9417t1514) I(R9417t5210) I(R9417t1140) I(R9418t2422) I(R9418t6523) I(R9418t7471) I(R9418t1117) I(R9418t5555) I(R9418t4960) I(R9418t3355) I(R9419t494) I(R9419t1390) I(R9419t6732) I(R9419t5133) I(R9419t4722) I(R9419t7026) I(R9420t6173) I(R9420t9226) I(R9420t7043) I(R9420t3702) I(R9421t2178) I(R9421t4590) I(R9421t287) I(R9421t8938) I(R9421t7167) I(R9421t4776) I(R9422t5576) I(R9422t8990) I(R9422t4268) I(R9422t8937) I(R9423t5544) I(R9423t3968) I(R9423t9279) I(R9423t7460) I(R9424t8504) I(R9424t7071) I(R9424t5664) I(R9424t574) I(R9424t1257) I(R9424t7129) I(R9425t517) I(R9425t1497) I(R9426t28) I(R9426t6611) I(R9426t1230) I(R9426t8232) I(R9426t3562) I(R9426t6951) I(R9427t1692) I(R9427t3396) I(R9427t2765) I(R9427t7238) I(R9427t9175) I(R9428t2149) I(R9428t8234) I(R9428t3377) I(R9429t291) I(R9429t3609) I(R9429t5700) I(R9429t8631) I(R9429t2569) I(R9429t6281) I(R9430t3260) I(R9430t6277) I(R9430t2604) I(R9430t3854) I(R9430t1931) I(R9430t47) I(R9431t630) I(R9431t1007) I(R9431t3207) I(R9431t6998) I(R9431t8552) I(R9431t4444) I(R9432t6908) I(R9432t3468) I(R9432t7990) I(R9432t3183) I(R9433t5574) I(R9433t9204) I(R9433t9154) I(R9433t7728) I(R9433t3384) I(R9434t18) I(R9434t1852) I(R9434t7316) I(R9434t218) I(R9434t9322) I(R9434t2394) I(R9434t1641) I(R9435t104) I(R9435t2005) I(R9435t7269) I(R9435t4847) I(R9435t2824) I(R9435t8208) I(R9435t159) I(R9435t1291) I(R9436t4273) I(R9436t5220) I(R9436t4760) I(R9436t1348) I(R9436t4073) I(R9437t6496) I(R9437t7962) I(R9437t1794) I(R9437t8480) I(R9438t4358) I(R9438t7098) I(R9438t6734) I(R9438t2211) I(R9438t2140) I(R9438t7579) I(R9439t4690) I(R9439t6129) I(R9439t1374) I(R9439t68) I(R9440t2453) I(R9440t7842) I(R9440t8763) I(R9440t3616) I(R9440t9103) I(R9440t7907) I(R9441t141) I(R9441t8769) I(R9441t7690) I(R9441t3649) I(R9441t8370) I(R9442t1798) I(R9442t3575) I(R9442t5364) I(R9442t9300) I(R9442t6495) I(R9442t6132) I(R9443t3062) I(R9443t5607) I(R9443t5511) I(R9443t8636) I(R9443t5299) I(R9443t4398) I(R9443t1502) I(R9443t1746) I(R9444t5637) I(R9444t6727) I(R9444t8089) I(R9444t375) I(R9444t6803) I(R9444t5254) I(R9444t7521) I(R9444t7305) I(R9444t9297) I(R9444t6511) I(R9444t9193) I(R9445t3764) I(R9445t5074) I(R9445t159) I(R9445t9435) I(R9445t1291) I(R9445t5270) I(R9445t1737) I(R9446t620) I(R9446t6620) I(R9446t900) I(R9446t6448) I(R9446t5260) I(R9447t2987) I(R9447t8234) I(R9447t9428) I(R9447t769) I(R9447t1683) I(R9447t3465) I(R9448t397) I(R9448t4177) I(R9448t2728) I(R9448t4148) I(R9448t3856) I(R9448t1198) I(R9448t4711) I(R9448t4110) I(R9449t2828) I(R9449t3094) I(R9449t907) I(R9449t5264) I(R9449t1181) I(R9449t2164) I(R9450t1269) I(R9450t7124) I(R9450t8909) I(R9450t1556) I(R9450t8522) I(R9450t805) I(R9450t4704) I(R9450t2757) I(R9450t2636) I(R9451t3269) I(R9451t8534) I(R9451t5958) I(R9451t1669) I(R9451t5241) I(R9451t4212) I(R9452t1052) I(R9452t9189) I(R9452t1378) I(R9452t3155) I(R9452t4176) I(R9452t1262) I(R9452t8704) I(R9453t2543) I(R9453t8794) I(R9453t8120) I(R9453t850) I(R9453t4606) I(R9454t7520) I(R9454t7982) I(R9454t2696) I(R9454t8336) I(R9454t7372) I(R9455t6449) I(R9455t8383) I(R9455t5121) I(R9455t2447) I(R9455t7721) I(R9455t7578) I(R9455t1382) I(R9456t2252) I(R9456t6744) I(R9456t3568) I(R9456t6349) I(R9457t7054) I(R9457t7271) I(R9457t1073) I(R9457t7957) I(R9457t5839) I(R9458t4834) I(R9458t6898) I(R9458t8773) I(R9458t9296) I(R9458t8875) I(R9459t867) I(R9459t8718) I(R9459t54) I(R9459t148) I(R9459t4) I(R9459t4285) I(R9460t2285) I(R9460t3816) I(R9460t3576) I(R9460t5849) I(R9460t196) I(R9460t7640) I(R9461t3437) I(R9461t6012) I(R9461t888) I(R9461t5548) I(R9461t4744) I(R9462t805) I(R9462t9450) I(R9462t495) I(R9462t7566) I(R9462t8522) I(R9463t1364) I(R9463t7530) I(R9463t7293) I(R9463t1517) I(R9463t8902) I(R9463t6006) I(R9464t2277) I(R9464t6355) I(R9464t3817) I(R9464t4939) I(R9464t2112) I(R9465t2848) I(R9465t7208) I(R9465t3717) I(R9465t9403) I(R9465t1823) I(R9466t667) I(R9466t5538) I(R9466t559) I(R9466t8551) I(R9467t622) I(R9467t7478) I(R9467t7740) I(R9467t93) I(R9467t2147) I(R9467t2349) I(R9468t7025) I(R9468t9277) I(R9468t5983) I(R9468t4412) I(R9468t6635) I(R9468t131) I(R9468t6380) I(R9469t784) I(R9469t9402) I(R9469t3078) I(R9469t1301) I(R9469t5897) I(R9470t70) I(R9470t2054) I(R9470t5269) I(R9470t4092) I(R9471t5544) I(R9471t9423) I(R9471t7460) I(R9471t2402) I(R9471t3033) I(R9472t1167) I(R9472t6421) I(R9472t3996) I(R9472t8306) I(R9472t5612) I(R9472t6393) I(R9472t3713) I(R9472t5194) I(R9472t8610) I(R9473t1184) I(R9473t4848) I(R9473t4951) I(R9473t4231) I(R9473t1307) I(R9473t3824) I(R9474t1561) I(R9474t9238) I(R9474t4872) I(R9474t3118) I(R9474t2966) I(R9474t2931) I(R9474t6522) I(R9474t8416) I(R9475t6289) I(R9475t8690) I(R9475t6417) I(R9475t8998) I(R9476t157) I(R9476t5816) I(R9476t5136) I(R9476t2733) I(R9476t5165) I(R9476t451) I(R9476t6767) I(R9477t81) I(R9477t5200) I(R9477t4729) I(R9477t7159) I(R9478t8448) I(R9478t8604) I(R9478t2173) I(R9478t652) I(R9478t9016) I(R9478t1109) I(R9478t4277) I(R9478t7635) I(R9479t3632) I(R9479t8736) I(R9479t874) I(R9479t4977) I(R9479t3211) I(R9479t5594) I(R9479t9407) I(R9479t1743) I(R9479t3022) I(R9480t1372) I(R9480t8912) I(R9480t4067) I(R9480t4989) I(R9480t71) I(R9481t605) I(R9481t3286) I(R9481t4379) I(R9481t2596) I(R9482t1849) I(R9482t7365) I(R9482t2151) I(R9482t8801) I(R9482t1690) I(R9482t7599) I(R9482t2973) I(R9483t620) I(R9483t2042) I(R9483t6611) I(R9483t8833) I(R9483t8653) I(R9484t4050) I(R9484t6235) I(R9484t7818) I(R9484t6910) I(R9484t3937) I(R9484t2146) I(R9484t8067) I(R9485t2952) I(R9485t8622) I(R9485t8831) I(R9485t3266) I(R9486t218) I(R9486t9360) I(R9486t6458) I(R9486t5044) I(R9486t7316) I(R9486t9434) I(R9487t4268) I(R9487t7025) I(R9487t9422) I(R9487t8937) I(R9487t5983) I(R9487t9468) I(R9488t5947) I(R9488t6622) I(R9488t2842) I(R9488t6114) I(R9488t7528) I(R9488t2038) I(R9489t971) I(R9489t5368) I(R9489t4986) I(R9489t4069) I(R9489t2423) I(R9490t1494) I(R9490t8804) I(R9490t4546) I(R9490t7885) I(R9490t8092) I(R9490t465) I(R9491t29) I(R9491t9351) I(R9491t5297) I(R9491t4800) I(R9491t1099) I(R9492t3029) I(R9492t7620) I(R9492t373) I(R9492t550) I(R9492t9297) I(R9493t6792) I(R9493t7596) I(R9493t6204) I(R9493t9041) I(R9493t6457) I(R9493t2530) I(R9494t515) I(R9494t3158) I(R9494t5477) I(R9494t3823) I(R9494t2339) I(R9494t2520) I(R9495t836) I(R9495t3908) I(R9495t8818) I(R9495t9267) I(R9495t4706) I(R9495t8137) I(R9496t8798) I(R9496t8951) I(R9496t6046) I(R9496t3400) I(R9496t2359) I(R9497t2852) I(R9497t8513) I(R9497t7134) I(R9497t419) I(R9497t7054) I(R9498t2370) I(R9498t4613) I(R9498t7379) I(R9498t1832) I(R9499t6738) I(R9499t8238) I(R9499t27) I(R9499t625) I(R9500t329) I(R9500t3474) I(R9500t2284) I(R9500t442) I(R9500t3537) I(R9500t5377) I(R9501t134) I(R9501t7215) I(R9501t8355) I(R9502t5806) I(R9502t6302) I(R9502t8317) I(R9502t2339) I(R9502t3823) I(R9502t8031) I(R9503t1368) I(R9503t2652) I(R9503t1799) I(R9503t3353) I(R9503t7063) I(R9504t4995) I(R9504t8901) I(R9504t9004) I(R9504t510) I(R9504t1767) I(R9505t7617) I(R9505t8176) I(R9505t2944) I(R9505t3717) I(R9505t3661) I(R9505t8401) I(R9505t6301) I(R9506t7141) I(R9506t7914) I(R9506t847) I(R9506t5100) I(R9506t6563) I(R9506t4054) I(R9507t1655) I(R9507t8753) I(R9507t4880) I(R9507t1118) I(R9507t2982) I(R9508t1041) I(R9508t6721) I(R9508t2868) I(R9508t2641) I(R9509t1439) I(R9509t2847) I(R9509t1652) I(R9509t2570) I(R9509t5295) I(R9509t5863) I(R9509t6952) I(R9509t9100) I(R9509t4021) I(R9510t42) I(R9510t4042) I(R9511t1691) I(R9511t2176) I(R9511t322) I(R9511t4329) I(R9511t8403) I(R9511t8665) I(R9511t1111) I(R9512t1841) I(R9512t2649) I(R9512t5502) I(R9512t7353) I(R9512t1853) I(R9512t876) I(R9512t7663) I(R9513t1596) I(R9513t7054) I(R9513t9457) I(R9513t5839) I(R9513t6180) I(R9514t6000) I(R9514t6655) I(R9514t5933) I(R9514t951) I(R9514t1350) I(R9514t8930) I(R9514t1307) I(R9514t6111) I(R9515t2357) I(R9515t5271) I(R9515t8224) I(R9515t1467) I(R9515t1421) I(R9515t8230) I(R9516t4044) I(R9516t4160) I(R9516t4545) I(R9516t7250) I(R9516t252) I(R9516t4739) I(R9517t3188) I(R9517t7200) I(R9517t2121) I(R9517t4861) I(R9517t4404) I(R9517t4771) I(R9517t8550) I(R9518t1992) I(R9518t7934) I(R9518t8045) I(R9518t285) I(R9519t1252) I(R9519t5883) I(R9519t4011) I(R9519t8888) I(R9520t7569) I(R9520t8337) I(R9520t8063) I(R9520t5275) I(R9520t7595) I(R9520t6901) I(R9520t8168) I(R9521t2922) I(R9521t7882) I(R9521t4134) I(R9521t4510) I(R9521t9215) I(R9522t925) I(R9522t6280) I(R9522t8672) I(R9522t8348) I(R9522t2372) I(R9522t4129) I(R9523t2149) I(R9523t9428) I(R9523t9447) I(R9523t769) I(R9523t7214) I(R9523t1764) I(R9524t5526) I(R9524t7445) I(R9524t6340) I(R9524t156) I(R9525t3279) I(R9525t8430) I(R9525t8056) I(R9525t7022) I(R9525t814) I(R9525t2083) I(R9525t5465) I(R9526t2285) I(R9526t9460) I(R9526t7640) I(R9526t4911) I(R9526t6780) I(R9527t1327) I(R9527t3863) I(R9527t2107) I(R9527t639) I(R9527t6637) I(R9527t6267) I(R9527t6893) I(R9528t3694) I(R9528t4382) I(R9528t257) I(R9528t9056) I(R9528t1949) I(R9528t7275) I(R9528t1010) I(R9529t3559) I(R9529t7419) I(R9529t8570) I(R9529t2779) I(R9529t1893) I(R9530t2956) I(R9530t4101) I(R9530t5180) I(R9530t5792) I(R9530t8824) I(R9531t5268) I(R9531t7376) I(R9531t7516) I(R9531t6217) I(R9531t3783) I(R9531t546) I(R9531t3281) I(R9531t4222) I(R9532t1707) I(R9532t8491) I(R9532t3913) I(R9532t4272) I(R9532t377) I(R9532t6551) I(R9533t3331) I(R9533t5848) I(R9533t4936) I(R9533t4922) I(R9533t4430) I(R9534t3389) I(R9534t8817) I(R9534t8612) I(R9534t2247) I(R9534t5531) I(R9534t3819) I(R9534t2964) I(R9535t7293) I(R9535t8897) I(R9535t9128) I(R9535t2351) I(R9536t6180) I(R9536t9513) I(R9536t5839) I(R9536t1976) I(R9536t1400) I(R9536t6660) I(R9537t1749) I(R9537t4471) I(R9537t3834) I(R9537t581) I(R9537t2056) I(R9537t5763) I(R9538t1841) I(R9538t2649) I(R9538t6579) I(R9538t7695) I(R9538t8258) I(R9539t5139) I(R9539t6556) I(R9539t2214) I(R9539t7927) I(R9539t1581) I(R9539t7357) I(R9540t5709) I(R9540t5735) I(R9540t1003) I(R9540t2665) I(R9540t6298) I(R9540t7826) I(R9541t209) I(R9541t8252) I(R9541t8330) I(R9541t202) I(R9541t6683) I(R9541t3586) I(R9541t873) I(R9541t6885) I(R9542t993) I(R9542t8553) I(R9542t1326) I(R9542t3508) I(R9542t1830) I(R9542t3899) I(R9543t2047) I(R9543t4162) I(R9543t1645) I(R9543t7655) I(R9543t7259) I(R9544t9027) I(R9544t9389) I(R9544t1442) I(R9544t7647) I(R9544t7983) I(R9544t1391) I(R9545t2549) I(R9545t5669) I(R9545t8968) I(R9545t3005) I(R9545t12) I(R9545t8451) I(R9546t382) I(R9546t4649) I(R9546t4693) I(R9546t479) I(R9546t9114) I(R9546t4742) I(R9546t5552) I(R9547t6924) I(R9547t8295) I(R9547t8536) I(R9547t5014) I(R9547t7782) I(R9548t5643) I(R9548t7166) I(R9548t5800) I(R9548t2734) I(R9548t79) I(R9548t4893) I(R9549t9439) I(R9549t1374) I(R9549t1311) I(R9549t8424) I(R9549t2161) I(R9550t808) I(R9550t8431) I(R9550t3411) I(R9550t9245) I(R9550t5987) I(R9550t3582) I(R9550t619) I(R9550t1382) I(R9551t1303) I(R9551t7559) I(R9551t4562) I(R9551t1299) I(R9551t378) I(R9552t517) I(R9552t7583) I(R9552t3607) I(R9552t1914) I(R9552t1497) I(R9552t9425) I(R9553t6947) I(R9553t6985) I(R9553t6221) I(R9553t1733) I(R9553t276) I(R9553t8949) I(R9554t2331) I(R9554t3895) I(R9554t964) I(R9554t3401) I(R9555t2567) I(R9555t6610) I(R9555t7165) I(R9555t182) I(R9555t2705) I(R9556t3810) I(R9556t8227) I(R9556t7992) I(R9556t8751) I(R9557t3165) I(R9557t1008) I(R9557t1895) I(R9557t4683) I(R9557t3185) I(R9558t5115) I(R9558t7832) I(R9558t2161) I(R9558t9549) I(R9558t9439) I(R9558t4690) I(R9558t5668) I(R9558t8058) I(R9559t5706) I(R9559t8933) I(R9559t618) I(R9559t3372) I(R9559t2014) I(R9559t3817) I(R9559t4292) I(R9560t6868) I(R9560t7776) I(R9560t3019) I(R9560t766) I(R9560t1579) I(R9560t4529) I(R9561t724) I(R9561t8646) I(R9561t1433) I(R9561t7207) I(R9561t4741) I(R9561t833) I(R9562t2417) I(R9562t5149) I(R9562t4996) I(R9562t8679) I(R9562t8281) I(R9562t7715) I(R9563t2466) I(R9563t3467) I(R9563t3889) I(R9563t4599) I(R9564t5023) I(R9564t5355) I(R9564t6791) I(R9564t751) I(R9564t4993) I(R9565t4533) I(R9565t7493) I(R9565t6805) I(R9565t963) I(R9565t6081) I(R9565t7573) I(R9565t7621) I(R9565t984) I(R9565t5540) I(R9566t8009) I(R9566t8353) I(R9566t4062) I(R9566t2853) I(R9567t1705) I(R9567t8749) I(R9567t6172) I(R9567t5610) I(R9567t8936) I(R9567t1523) I(R9567t3729) I(R9567t4865) I(R9568t5256) I(R9568t8476) I(R9568t5899) I(R9568t5626) I(R9568t8515) I(R9569t7613) I(R9569t9330) I(R9569t4619) I(R9569t4445) I(R9569t2858) I(R9570t242) I(R9570t6626) I(R9570t2711) I(R9570t8279) I(R9570t1162) I(R9571t3128) I(R9571t8038) I(R9571t1051) I(R9571t6883) I(R9571t8356) I(R9572t4027) I(R9572t6320) I(R9572t4163) I(R9572t103) I(R9572t7625) I(R9572t7458) I(R9572t7911) I(R9573t5323) I(R9573t6210) I(R9573t7741) I(R9573t6465) I(R9573t8044) I(R9573t2117) I(R9574t4695) I(R9574t7781) I(R9574t1978) I(R9574t3099) I(R9575t5859) I(R9575t8180) I(R9575t2886) I(R9575t1654) I(R9575t4512) I(R9576t1592) I(R9576t6598) I(R9576t2638) I(R9576t2480) I(R9576t1288) I(R9576t8235) I(R9577t235) I(R9577t5652) I(R9577t6207) I(R9577t2748) I(R9577t8642) I(R9577t5988) I(R9577t5153) I(R9577t2673) I(R9578t3628) I(R9578t8070) I(R9578t1555) I(R9578t3874) I(R9578t1776) I(R9578t2206) I(R9578t3359) I(R9579t2686) I(R9579t6483) I(R9579t3843) I(R9579t4008) I(R9579t9025) I(R9579t1601) I(R9579t873) I(R9580t2526) I(R9580t5920) I(R9580t6719) I(R9580t4125) I(R9580t8057) I(R9580t2736) I(R9580t7621) I(R9581t8219) I(R9581t8670) I(R9581t4261) I(R9581t2268) I(R9581t2430) I(R9582t598) I(R9582t790) I(R9582t8851) I(R9582t4328) I(R9582t7158) I(R9582t4242) I(R9582t4933) I(R9583t5180) I(R9583t9530) I(R9583t6346) I(R9583t8521) I(R9583t2341) I(R9583t2956) I(R9584t515) I(R9584t3158) I(R9584t5477) I(R9584t8193) I(R9584t3180) I(R9584t624) I(R9585t344) I(R9585t6935) I(R9585t1110) I(R9585t5472) I(R9585t89) I(R9585t4124) I(R9585t176) I(R9585t4003) I(R9586t6947) I(R9586t9553) I(R9586t4300) I(R9586t8949) I(R9587t557) I(R9587t8910) I(R9587t7071) I(R9587t9424) I(R9587t8504) I(R9587t4552) I(R9587t3512) I(R9588t8775) I(R9588t8827) I(R9588t2376) I(R9588t5219) I(R9588t6206) I(R9588t8855) I(R9588t5460) I(R9589t351) I(R9589t7273) I(R9589t4833) I(R9589t3232) I(R9589t4772) I(R9589t6609) I(R9589t3478) I(R9589t477) I(R9590t1900) I(R9590t2265) I(R9590t2801) I(R9590t1688) I(R9590t4673) I(R9590t1831) I(R9590t5948) I(R9590t4712) I(R9590t1608) I(R9591t5417) I(R9591t6128) I(R9591t3080) I(R9591t6652) I(R9591t5335) I(R9591t3615) I(R9591t2721) I(R9592t1790) I(R9592t8801) I(R9592t2800) I(R9592t7966) I(R9592t3725) I(R9593t6363) I(R9593t6370) I(R9593t4495) I(R9593t1206) I(R9593t2668) I(R9594t2987) I(R9594t9447) I(R9594t3465) I(R9594t8156) I(R9594t9380) I(R9594t7096) I(R9595t4727) I(R9595t8389) I(R9595t1193) I(R9595t8182) I(R9595t6516) I(R9595t7857) I(R9596t110) I(R9596t5616) I(R9596t7052) I(R9596t4860) I(R9596t3104) I(R9597t3027) I(R9597t5895) I(R9597t4691) I(R9597t4049) I(R9597t5214) I(R9597t7374) I(R9597t9359) I(R9597t1126) I(R9598t1413) I(R9598t7833) I(R9598t48) I(R9598t2892) I(R9598t8464) I(R9598t2464) I(R9598t2660) I(R9599t273) I(R9599t8053) I(R9599t3) I(R9599t6028) I(R9599t4172) I(R9599t6047) I(R9599t1655) I(R9600t1602) I(R9600t2855) I(R9600t9028) I(R9600t6519) I(R9600t3008) I(R9601t6597) I(R9601t8215) I(R9601t7612) I(R9601t6141) I(R9602t6384) I(R9602t9074) I(R9602t4769) I(R9602t6188) I(R9602t4262) I(R9603t6908) I(R9603t9432) I(R9603t8969) I(R9603t1723) I(R9603t3028) I(R9604t806) I(R9604t9170) I(R9604t384) I(R9604t9078) I(R9604t8629) I(R9604t3315) I(R9604t3003) I(R9605t7460) I(R9605t9423) I(R9605t9279) I(R9605t3349) I(R9605t2667) I(R9606t1388) I(R9606t6514) I(R9606t2424) I(R9606t6624) I(R9606t7771) I(R9606t1881) I(R9606t1572) I(R9607t5699) I(R9607t6742) I(R9607t4114) I(R9607t6229) I(R9607t1610) I(R9607t4967) I(R9608t527) I(R9608t6848) I(R9608t4686) I(R9608t7871) I(R9608t4026) I(R9608t6964) I(R9608t4062) I(R9609t8548) I(R9609t9043) I(R9609t4689) I(R9609t8165) I(R9610t3800) I(R9610t6443) I(R9610t7058) I(R9610t5475) I(R9610t3872) I(R9610t9269) I(R9611t3792) I(R9611t7173) I(R9611t7950) I(R9611t8433) I(R9611t54) I(R9611t161) I(R9611t7163) I(R9612t3113) I(R9612t5785) I(R9612t3391) I(R9612t9116) I(R9612t4374) I(R9612t4793) I(R9613t72) I(R9613t7034) I(R9613t1019) I(R9613t7745) I(R9613t6575) I(R9614t5741) I(R9614t8084) I(R9614t8580) I(R9614t1402) I(R9614t3358) I(R9615t2843) I(R9615t8132) I(R9615t7752) I(R9615t7224) I(R9616t886) I(R9616t2820) I(R9616t4710) I(R9616t4047) I(R9616t4907) I(R9616t6588) I(R9617t928) I(R9617t5973) I(R9617t9356) I(R9617t5093) I(R9617t2399) I(R9617t6644) I(R9618t5833) I(R9618t8785) I(R9618t8706) I(R9618t3132) I(R9618t2912) I(R9618t1594) I(R9618t7306) I(R9619t2507) I(R9619t9284) I(R9619t1947) I(R9619t7454) I(R9619t8074) I(R9619t8386) I(R9619t3768) I(R9619t9326) I(R9620t4062) I(R9620t4196) I(R9620t9566) I(R9620t2853) I(R9620t796) I(R9620t8977) I(R9620t527) I(R9621t2651) I(R9621t6948) I(R9621t843) I(R9621t8252) I(R9621t2986) I(R9621t6979) I(R9622t2260) I(R9622t8707) I(R9622t3650) I(R9622t739) I(R9623t3196) I(R9623t3203) I(R9623t2369) I(R9623t8724) I(R9623t112) I(R9623t7862) I(R9624t2665) I(R9624t5667) I(R9624t2189) I(R9624t934) I(R9625t1493) I(R9625t2152) I(R9625t3522) I(R9625t5276) I(R9625t4100) I(R9625t4804) I(R9625t5544) I(R9626t2906) I(R9626t4576) I(R9626t5015) I(R9626t7572) I(R9627t428) I(R9627t2938) I(R9627t4096) I(R9627t1929) I(R9627t856) I(R9627t9265) I(R9628t711) I(R9628t3034) I(R9628t9177) I(R9628t2477) I(R9629t5009) I(R9629t6065) I(R9629t3089) I(R9629t7709) I(R9629t1399) I(R9629t8613) I(R9629t1730) I(R9629t3378) I(R9630t4013) I(R9630t5408) I(R9630t8688) I(R9630t2410) I(R9630t7288) I(R9630t6591) I(R9631t6454) I(R9631t6994) I(R9631t3227) I(R9631t8890) I(R9631t3569) I(R9631t6079) I(R9631t6608) I(R9632t7868) I(R9632t8394) I(R9632t572) I(R9632t749) I(R9632t2723) I(R9632t6709) I(R9632t2355) I(R9633t1699) I(R9633t4467) I(R9633t6116) I(R9633t6653) I(R9633t5856) I(R9634t573) I(R9634t9343) I(R9634t3239) I(R9634t5887) I(R9634t5757) I(R9634t3170) I(R9635t1329) I(R9635t9327) I(R9635t9206) I(R9635t4012) I(R9635t7712) I(R9635t5572) I(R9636t5332) I(R9636t7905) I(R9636t5809) I(R9636t7296) I(R9636t8856) I(R9636t8285) I(R9637t3702) I(R9637t7043) I(R9637t7603) I(R9637t4009) I(R9637t268) I(R9638t6214) I(R9638t7915) I(R9638t6915) I(R9638t4255) I(R9638t1793) I(R9639t7983) I(R9639t9544) I(R9639t7647) I(R9639t1448) I(R9639t7890) I(R9639t8364) I(R9640t551) I(R9640t683) I(R9640t480) I(R9640t82) I(R9640t8177) I(R9640t1840) I(R9640t6018) I(R9641t387) I(R9641t1942) I(R9641t1456) I(R9641t3108) I(R9641t7496) I(R9641t3263) I(R9642t2872) I(R9642t3869) I(R9642t2568) I(R9642t6914) I(R9643t830) I(R9643t6521) I(R9643t7500) I(R9643t7812) I(R9643t9225) I(R9643t5258) I(R9644t3476) I(R9644t7138) I(R9644t4042) I(R9644t9510) I(R9644t42) I(R9644t9212) I(R9645t1176) I(R9645t2176) I(R9645t6102) I(R9645t7251) I(R9645t1691) I(R9646t4635) I(R9646t6256) I(R9646t1165) I(R9647t5254) I(R9647t6774) I(R9647t7922) I(R9647t5646) I(R9648t3638) I(R9648t8427) I(R9648t2738) I(R9648t3356) I(R9648t1727) I(R9648t2063) I(R9649t2282) I(R9649t4959) I(R9649t1972) I(R9649t8793) I(R9649t5181) I(R9649t3818) I(R9649t1139) I(R9650t9432) I(R9650t9603) I(R9650t3028) I(R9650t6752) I(R9650t2317) I(R9650t3183) I(R9651t2463) I(R9651t7701) I(R9651t9007) I(R9651t1220) I(R9651t4633) I(R9651t5512) I(R9652t3061) I(R9652t7897) I(R9652t764) I(R9652t8895) I(R9652t914) I(R9652t7698) I(R9653t1729) I(R9653t8596) I(R9653t4181) I(R9654t7747) I(R9654t8957) I(R9654t5086) I(R9654t3833) I(R9654t2342) I(R9654t8581) I(R9654t5741) I(R9655t665) I(R9655t8643) I(R9655t325) I(R9655t6259) I(R9655t5961) I(R9655t6357) I(R9656t2131) I(R9656t4950) I(R9656t5447) I(R9656t7217) I(R9656t5373) I(R9657t982) I(R9657t7208) I(R9657t1568) I(R9658t3565) I(R9658t4598) I(R9658t5363) I(R9658t1979) I(R9659t3472) I(R9659t4493) I(R9659t7105) I(R9659t8921) I(R9659t4827) I(R9659t4427) I(R9659t2066) I(R9660t2143) I(R9660t7278) I(R9660t423) I(R9660t6291) I(R9660t2404) I(R9660t6708) I(R9660t8125) I(R9661t1109) I(R9661t5710) I(R9661t9016) I(R9661t9164) I(R9661t303) I(R9662t653) I(R9662t6101) I(R9662t4285) I(R9662t9459) I(R9662t867) I(R9662t8617) I(R9663t2786) I(R9663t6463) I(R9663t172) I(R9663t4744) I(R9663t9461) I(R9663t5548) I(R9663t7431) I(R9664t2558) I(R9664t4305) I(R9664t2653) I(R9664t6044) I(R9664t2392) I(R9664t1927) I(R9665t5082) I(R9665t9102) I(R9665t8875) I(R9665t9458) I(R9665t9296) I(R9665t1090) I(R9665t1967) I(R9665t7304) I(R9666t1436) I(R9666t7540) I(R9667t1026) I(R9667t3165) I(R9667t3730) I(R9667t3185) I(R9667t9557) I(R9668t331) I(R9668t582) I(R9668t1016) I(R9668t8447) I(R9668t6299) I(R9668t4610) I(R9668t7758) I(R9669t565) I(R9669t6961) I(R9669t8118) I(R9669t6525) I(R9669t5058) I(R9669t5288) I(R9669t4098) I(R9669t425) I(R9670t2141) I(R9670t3169) I(R9670t7542) I(R9670t7471) I(R9670t9418) I(R9670t2422) I(R9671t4871) I(R9671t6938) I(R9671t4466) I(R9671t2611) I(R9672t8734) I(R9672t8745) I(R9672t3680) I(R9672t6475) I(R9672t7871) I(R9673t3613) I(R9673t3625) I(R9673t827) I(R9673t6897) I(R9673t1521) I(R9673t6365) I(R9673t4122) I(R9673t7487) I(R9673t6127) I(R9674t669) I(R9674t7184) I(R9674t1141) I(R9674t1820) I(R9674t1905) I(R9674t3400) I(R9675t6309) I(R9675t8128) I(R9675t4974) I(R9675t1935) I(R9675t8864) I(R9675t6741) I(R9675t6362) I(R9676t784) I(R9676t5028) I(R9676t8315) I(R9676t3762) I(R9676t3175) I(R9676t3980) I(R9677t2457) I(R9677t4031) I(R9677t5515) I(R9677t2255) I(R9677t4435) I(R9677t4901) I(R9678t4779) I(R9678t7150) I(R9678t8356) I(R9678t3669) I(R9678t3365) I(R9678t7679) I(R9678t2745) I(R9679t3874) I(R9679t4170) I(R9679t9578) I(R9679t1555) I(R9679t5237) I(R9679t670) I(R9679t2125) I(R9679t5721) I(R9680t2154) I(R9680t3947) I(R9680t7625) I(R9680t9572) I(R9680t7458) I(R9680t1620) I(R9681t5116) I(R9681t6434) I(R9681t6835) I(R9681t8293) I(R9681t9367) I(R9681t1870) I(R9681t4169) I(R9682t3385) I(R9682t7905) I(R9682t5332) I(R9682t2854) I(R9682t8183) I(R9682t7519) I(R9682t4937) I(R9683t6532) I(R9683t8463) I(R9683t37) I(R9683t9034) I(R9683t6911) I(R9683t6617) I(R9683t4405) I(R9683t8836) I(R9684t5300) I(R9684t5493) I(R9684t1609) I(R9684t8062) I(R9684t4866) I(R9684t1138) I(R9685t3521) I(R9685t6381) I(R9685t8578) I(R9685t9311) I(R9685t4293) I(R9685t2602) I(R9686t286) I(R9686t6219) I(R9686t1553) I(R9686t3549) I(R9686t8165) I(R9686t8548) I(R9686t2574) I(R9687t4522) I(R9687t4888) I(R9687t5787) I(R9687t5396) I(R9687t210) I(R9688t5638) I(R9688t6517) I(R9688t496) I(R9688t1922) I(R9688t3912) I(R9688t4590) I(R9688t4776) I(R9689t2480) I(R9689t8889) I(R9689t1288) I(R9689t83) I(R9689t1451) I(R9690t4163) I(R9690t6346) I(R9690t3589) I(R9690t2534) I(R9690t8243) I(R9690t103) I(R9691t7987) I(R9691t8043) I(R9691t8117) I(R9691t3326) I(R9691t1425) I(R9692t1183) I(R9692t5073) I(R9692t1703) I(R9692t5758) I(R9692t851) I(R9692t7032) I(R9692t3395) I(R9692t6076) I(R9693t1229) I(R9693t6280) I(R9693t5929) I(R9693t6391) I(d2) I(d3) I(d4) I(d5) I(d6) I(d7) I(d8) I(d9) I(d10) I(d11) I(d12) I(d13) I(d14) I(d15) I(d16) I(d17) I(d18) I(d19) I(d20) I(d21) I(d22) I(d23) I(d24) I(d25) I(d26) I(d27) I(d28) I(d29) I(d30) I(d31) I(d32) I(d33) I(d34) I(d35) I(d36) I(d37) I(d38) I(d39) I(d40) I(d41) I(d42) I(d43) I(d44) I(d45) I(d46) I(d47) I(d48) I(d49) I(d50) I(d51) I(d52) I(d53) I(d54) I(d55) I(d56) I(d57) I(d58) I(d59) I(d60) I(d61) I(d62) I(d63) I(d64) I(d65) I(d66) I(d67) I(d68) I(d69) I(d70) I(d71) I(d72) I(d73) I(d74) I(d75) I(d76) I(d77) I(d78) I(d79) I(d80) I(d81) I(d82) I(d83) I(d84) I(d85) I(d86) I(d87) I(d88) I(d89) I(d90) I(d91) I(d92) I(d93) I(d94) I(d95) I(d96) I(d97) I(d98) I(d99) I(d100) I(d101) I(d102) I(d103) I(d104) I(d105) I(d106) I(d107) I(d108) I(d109) I(d110) I(d111) I(d112) I(d113) I(d114) I(d115) I(d116) I(d117) I(d118) I(d119) I(d120) I(d121) I(d122) I(d123) I(d124) I(d125) I(d126) I(d127) I(d128) I(d129) I(d130) I(d131) I(d132) I(d133) I(d134) I(d135) I(d136) I(d137) I(d138) I(d139) I(d140) I(d141) I(d142) I(d143) I(d144) I(d145) I(d146) I(d147) I(d148) I(d149) I(d150) I(d151) I(d152) I(d153) I(d154) I(d155) I(d156) I(d157) I(d158) I(d159) I(d160) I(d161) I(d162) I(d163) I(d164) I(d165) I(d166) I(d167) I(d168) I(d169) I(d170) I(d171) I(d172) I(d173) I(d174) I(d175) I(d176) I(d177) I(d178) I(d179) I(d180) I(d181) I(d182) I(d183) I(d184) I(d185) I(d186) I(d187) I(d188) I(d189) I(d190) I(d191) I(d192) I(d193) I(d194) I(d195) I(d196) I(d197) I(d198) I(d199) I(d200) I(d201) I(d202) I(d203) I(d204) I(d205) I(d206) I(d207) I(d208) I(d209) I(d210) I(d211) I(d212) I(d213) I(d214) I(d215) I(d216) I(d217) I(d218) I(d219) I(d220) I(d221) I(d222) I(d223) I(d224) I(d225) I(d226) I(d227) I(d228) I(d229) I(d230) I(d231) I(d232) I(d233) I(d234) I(d235) I(d236) I(d237) I(d238) I(d239) I(d240) I(d241) I(d242) I(d243) I(d244) I(d245) I(d246) I(d247) I(d248) I(d249) I(d250) I(d251) I(d252) I(d253) I(d254) I(d255) I(d256) I(d257) I(d258) I(d259) I(d260) I(d261) I(d262) I(d263) I(d264) I(d265) I(d266) I(d267) I(d268) I(d269) I(d270) I(d271) I(d272) I(d273) I(d274) I(d275) I(d276) I(d277) I(d278) I(d279) I(d280) I(d281) I(d282) I(d283) I(d284) I(d285) I(d286) I(d287) I(d288) I(d289) I(d290) I(d291) I(d292) I(d293) I(d294) I(d295) I(d296) I(d297) I(d298) I(d299) I(d300) I(d301) I(d302) I(d303) I(d304) I(d305) I(d306) I(d307) I(d308) I(d309) I(d310) I(d311) I(d312) I(d313) I(d314) I(d315) I(d316) I(d317) I(d318) I(d319) I(d320) I(d321) I(d322) I(d323) I(d324) I(d325) I(d326) I(d327) I(d328) I(d329) I(d330) I(d331) I(d332) I(d333) I(d334) I(d335) I(d336) I(d337) I(d338) I(d339) I(d340) I(d341) I(d342) I(d343) I(d344) I(d345) I(d346) I(d347) I(d348) I(d349) I(d350) I(d351) I(d352) I(d353) I(d354) I(d355) I(d356) I(d357) I(d358) I(d359) I(d360) I(d361) I(d362) I(d363) I(d364) I(d365) I(d366) I(d367) I(d368) I(d369) I(d370) I(d371) I(d372) I(d373) I(d374) I(d375) I(d376) I(d377) I(d378) I(d379) I(d380) I(d381) I(d382) I(d383) I(d384) I(d385) I(d386) I(d387) I(d388) I(d389) I(d390) I(d391) I(d392) I(d393) I(d394) I(d395) I(d396) I(d397) I(d398) I(d399) I(d400) I(d401) I(d402) I(d403) I(d404) I(d405) I(d406) I(d407) I(d408) I(d409) I(d410) I(d411) I(d412) I(d413) I(d414) I(d415) I(d416) I(d417) I(d418) I(d419) I(d420) I(d421) I(d422) I(d423) I(d424) I(d425) I(d426) I(d427) I(d428) I(d429) I(d430) I(d431) I(d432) I(d433) I(d434) I(d435) I(d436) I(d437) I(d438) I(d439) I(d440) I(d441) I(d442) I(d443) I(d444) I(d445) I(d446) I(d447) I(d448) I(d449) I(d450) I(d451) I(d452) I(d453) I(d454) I(d455) I(d456) I(d457) I(d458) I(d459) I(d460) I(d461) I(d462) I(d463) I(d464) I(d465) I(d466) I(d467) I(d468) I(d469) I(d470) I(d471) I(d472) I(d473) I(d474) I(d475) I(d476) I(d477) I(d478) I(d479) I(d480) I(d481) I(d482) I(d483) I(d484) I(d485) I(d486) I(d487) I(d488) I(d489) I(d490) I(d491) I(d492) I(d493) I(d494) I(d495) I(d496) I(d497) I(d498) I(d499) I(d500) I(d501) I(d502) I(d503) I(d504) I(d505) I(d506) I(d507) I(d508) I(d509) I(d510) I(d511) I(d512) I(d513) I(d514) I(d515) I(d516) I(d517) I(d518) I(d519) I(d520) I(d521) I(d522) I(d523) I(d524) I(d525) I(d526) I(d527) I(d528) I(d529) I(d530) I(d531) I(d532) I(d533) I(d534) I(d535) I(d536) I(d537) I(d538) I(d539) I(d540) I(d541) I(d542) I(d543) I(d544) I(d545) I(d546) I(d547) I(d548) I(d549) I(d550) I(d551) I(d552) I(d553) I(d554) I(d555) I(d556) I(d557) I(d558) I(d559) I(d560) I(d561) I(d562) I(d563) I(d564) I(d565) I(d566) I(d567) I(d568) I(d569) I(d570) I(d571) I(d572) I(d573) I(d574) I(d575) I(d576) I(d577) I(d578) I(d579) I(d580) I(d581) I(d582) I(d583) I(d584) I(d585) I(d586) I(d587) I(d588) I(d589) I(d590) I(d591) I(d592) I(d593) I(d594) I(d595) I(d596) I(d597) I(d598) I(d599) I(d600) I(d601) I(d602) I(d603) I(d604) I(d605) I(d606) I(d607) I(d608) I(d609) I(d610) I(d611) I(d612) I(d613) I(d614) I(d615) I(d616) I(d617) I(d618) I(d619) I(d620) I(d621) I(d622) I(d623) I(d624) I(d625) I(d626) I(d627) I(d628) I(d629) I(d630) I(d631) I(d632) I(d633) I(d634) I(d635) I(d636) I(d637) I(d638) I(d639) I(d640) I(d641) I(d642) I(d643) I(d644) I(d645) I(d646) I(d647) I(d648) I(d649) I(d650) I(d651) I(d652) I(d653) I(d654) I(d655) I(d656) I(d657) I(d658) I(d659) I(d660) I(d661) I(d662) I(d663) I(d664) I(d665) I(d666) I(d667) I(d668) I(d669) I(d670) I(d671) I(d672) I(d673) I(d674) I(d675) I(d676) I(d677) I(d678) I(d679) I(d680) I(d681) I(d682) I(d683) I(d684) I(d685) I(d686) I(d687) I(d688) I(d689) I(d690) I(d691) I(d692) I(d693) I(d694) I(d695) I(d696) I(d697) I(d698) I(d699) I(d700) I(d701) I(d702) I(d703) I(d704) I(d705) I(d706) I(d707) I(d708) I(d709) I(d710) I(d711) I(d712) I(d713) I(d714) I(d715) I(d716) I(d717) I(d718) I(d719) I(d720) I(d721) I(d722) I(d723) I(d724) I(d725) I(d726) I(d727) I(d728) I(d729) I(d730) I(d731) I(d732) I(d733) I(d734) I(d735) I(d736) I(d737) I(d738) I(d739) I(d740) I(d741) I(d742) I(d743) I(d744) I(d745) I(d746) I(d747) I(d748) I(d749) I(d750) I(d751) I(d752) I(d753) I(d754) I(d755) I(d756) I(d757) I(d758) I(d759) I(d760) I(d761) I(d762) I(d763) I(d764) I(d765) I(d766) I(d767) I(d768) I(d769) I(d770) I(d771) I(d772) I(d773) I(d774) I(d775) I(d776) I(d777) I(d778) I(d779) I(d780) I(d781) I(d782) I(d783) I(d784) I(d785) I(d786) I(d787) I(d788) I(d789) I(d790) I(d791) I(d792) I(d793) I(d794) I(d795) I(d796) I(d797) I(d798) I(d799) I(d800) I(d801) I(d802) I(d803) I(d804) I(d805) I(d806) I(d807) I(d808) I(d809) I(d810) I(d811) I(d812) I(d813) I(d814) I(d815) I(d816) I(d817) I(d818) I(d819) I(d820) I(d821) I(d822) I(d823) I(d824) I(d825) I(d826) I(d827) I(d828) I(d829) I(d830) I(d831) I(d832) I(d833) I(d834) I(d835) I(d836) I(d837) I(d838) I(d839) I(d840) I(d841) I(d842) I(d843) I(d844) I(d845) I(d846) I(d847) I(d848) I(d849) I(d850) I(d851) I(d852) I(d853) I(d854) I(d855) I(d856) I(d857) I(d858) I(d859) I(d860) I(d861) I(d862) I(d863) I(d864) I(d865) I(d866) I(d867) I(d868) I(d869) I(d870) I(d871) I(d872) I(d873) I(d874) I(d875) I(d876) I(d877) I(d878) I(d879) I(d880) I(d881) I(d882) I(d883) I(d884) I(d885) I(d886) I(d887) I(d888) I(d889) I(d890) I(d891) I(d892) I(d893) I(d894) I(d895) I(d896) I(d897) I(d898) I(d899) I(d900) I(d901) I(d902) I(d903) I(d904) I(d905) I(d906) I(d907) I(d908) I(d909) I(d910) I(d911) I(d912) I(d913) I(d914) I(d915) I(d916) I(d917) I(d918) I(d919) I(d920) I(d921) I(d922) I(d923) I(d924) I(d925) I(d926) I(d927) I(d928) I(d929) I(d930) I(d931) I(d932) I(d933) I(d934) I(d935) I(d936) I(d937) I(d938) I(d939) I(d940) I(d941) I(d942) I(d943) I(d944) I(d945) I(d946) I(d947) I(d948) I(d949) I(d950) I(d951) I(d952) I(d953) I(d954) I(d955) I(d956) I(d957) I(d958) I(d959) I(d960) I(d961) I(d962) I(d963) I(d964) I(d965) I(d966) I(d967) I(d968) I(d969) I(d970) I(d971) I(d972) I(d973) I(d974) I(d975) I(d976) I(d977) I(d978) I(d979) I(d980) I(d981) I(d982) I(d983) I(d984) I(d985) I(d986) I(d987) I(d988) I(d989) I(d990) I(d991) I(d992) I(d993) I(d994) I(d995) I(d996) I(d997) I(d998) I(d999) I(d1000) I(d1001) I(d1002) I(d1003) I(d1004) I(d1005) I(d1006) I(d1007) I(d1008) I(d1009) I(d1010) I(d1011) I(d1012) I(d1013) I(d1014) I(d1015) I(d1016) I(d1017) I(d1018) I(d1019) I(d1020) I(d1021) I(d1022) I(d1023) I(d1024) I(d1025) I(d1026) I(d1027) I(d1028) I(d1029) I(d1030) I(d1031) I(d1032) I(d1033) I(d1034) I(d1035) I(d1036) I(d1037) I(d1038) I(d1039) I(d1040) I(d1041) I(d1042) I(d1043) I(d1044) I(d1045) I(d1046) I(d1047) I(d1048) I(d1049) I(d1050) I(d1051) I(d1052) I(d1053) I(d1054) I(d1055) I(d1056) I(d1057) I(d1058) I(d1059) I(d1060) I(d1061) I(d1062) I(d1063) I(d1064) I(d1065) I(d1066) I(d1067) I(d1068) I(d1069) I(d1070) I(d1071) I(d1072) I(d1073) I(d1074) I(d1075) I(d1076) I(d1077) I(d1078) I(d1079) I(d1080) I(d1081) I(d1082) I(d1083) I(d1084) I(d1085) I(d1086) I(d1087) I(d1088) I(d1089) I(d1090) I(d1091) I(d1092) I(d1093) I(d1094) I(d1095) I(d1096) I(d1097) I(d1098) I(d1099) I(d1100) I(d1101) I(d1102) I(d1103) I(d1104) I(d1105) I(d1106) I(d1107) I(d1108) I(d1109) I(d1110) I(d1111) I(d1112) I(d1113) I(d1114) I(d1115) I(d1116) I(d1117) I(d1118) I(d1119) I(d1120) I(d1121) I(d1122) I(d1123) I(d1124) I(d1125) I(d1126) I(d1127) I(d1128) I(d1129) I(d1130) I(d1131) I(d1132) I(d1133) I(d1134) I(d1135) I(d1136) I(d1137) I(d1138) I(d1139) I(d1140) I(d1141) I(d1142) I(d1143) I(d1144) I(d1145) I(d1146) I(d1147) I(d1148) I(d1149) I(d1150) I(d1151) I(d1152) I(d1153) I(d1154) I(d1155) I(d1156) I(d1157) I(d1158) I(d1159) I(d1160) I(d1161) I(d1162) I(d1163) I(d1164) I(d1165) I(d1166) I(d1167) I(d1168) I(d1169) I(d1170) I(d1171) I(d1172) I(d1173) I(d1174) I(d1175) I(d1176) I(d1177) I(d1178) I(d1179) I(d1180) I(d1181) I(d1182) I(d1183) I(d1184) I(d1185) I(d1186) I(d1187) I(d1188) I(d1189) I(d1190) I(d1191) I(d1192) I(d1193) I(d1194) I(d1195) I(d1196) I(d1197) I(d1198) I(d1199) I(d1200) I(d1201) I(d1202) I(d1203) I(d1204) I(d1205) I(d1206) I(d1207) I(d1208) I(d1209) I(d1210) I(d1211) I(d1212) I(d1213) I(d1214) I(d1215) I(d1216) I(d1217) I(d1218) I(d1219) I(d1220) I(d1221) I(d1222) I(d1223) I(d1224) I(d1225) I(d1226) I(d1227) I(d1228) I(d1229) I(d1230) I(d1231) I(d1232) I(d1233) I(d1234) I(d1235) I(d1236) I(d1237) I(d1238) I(d1239) I(d1240) I(d1241) I(d1242) I(d1243) I(d1244) I(d1245) I(d1246) I(d1247) I(d1248) I(d1249) I(d1250) I(d1251) I(d1252) I(d1253) I(d1254) I(d1255) I(d1256) I(d1257) I(d1258) I(d1259) I(d1260) I(d1261) I(d1262) I(d1263) I(d1264) I(d1265) I(d1266) I(d1267) I(d1268) I(d1269) I(d1270) I(d1271) I(d1272) I(d1273) I(d1274) I(d1275) I(d1276) I(d1277) I(d1278) I(d1279) I(d1280) I(d1281) I(d1282) I(d1283) I(d1284) I(d1285) I(d1286) I(d1287) I(d1288) I(d1289) I(d1290) I(d1291) I(d1292) I(d1293) I(d1294) I(d1295) I(d1296) I(d1297) I(d1298) I(d1299) I(d1300) I(d1301) I(d1302) I(d1303) I(d1304) I(d1305) I(d1306) I(d1307) I(d1308) I(d1309) I(d1310) I(d1311) I(d1312) I(d1313) I(d1314) I(d1315) I(d1316) I(d1317) I(d1318) I(d1319) I(d1320) I(d1321) I(d1322) I(d1323) I(d1324) I(d1325) I(d1326) I(d1327) I(d1328) I(d1329) I(d1330) I(d1331) I(d1332) I(d1333) I(d1334) I(d1335) I(d1336) I(d1337) I(d1338) I(d1339) I(d1340) I(d1341) I(d1342) I(d1343) I(d1344) I(d1345) I(d1346) I(d1347) I(d1348) I(d1349) I(d1350) I(d1351) I(d1352) I(d1353) I(d1354) I(d1355) I(d1356) I(d1357) I(d1358) I(d1359) I(d1360) I(d1361) I(d1362) I(d1363) I(d1364) I(d1365) I(d1366) I(d1367) I(d1368) I(d1369) I(d1370) I(d1371) I(d1372) I(d1373) I(d1374) I(d1375) I(d1376) I(d1377) I(d1378) I(d1379) I(d1380) I(d1381) I(d1382) I(d1383) I(d1384) I(d1385) I(d1386) I(d1387) I(d1388) I(d1389) I(d1390) I(d1391) I(d1392) I(d1393) I(d1394) I(d1395) I(d1396) I(d1397) I(d1398) I(d1399) I(d1400) I(d1401) I(d1402) I(d1403) I(d1404) I(d1405) I(d1406) I(d1407) I(d1408) I(d1409) I(d1410) I(d1411) I(d1412) I(d1413) I(d1414) I(d1415) I(d1416) I(d1417) I(d1418) I(d1419) I(d1420) I(d1421) I(d1422) I(d1423) I(d1424) I(d1425) I(d1426) I(d1427) I(d1428) I(d1429) I(d1430) I(d1431) I(d1432) I(d1433) I(d1434) I(d1435) I(d1436) I(d1437) I(d1438) I(d1439) I(d1440) I(d1441) I(d1442) I(d1443) I(d1444) I(d1445) I(d1446) I(d1447) I(d1448) I(d1449) I(d1450) I(d1451) I(d1452) I(d1453) I(d1454) I(d1455) I(d1456) I(d1457) I(d1458) I(d1459) I(d1460) I(d1461) I(d1462) I(d1463) I(d1464) I(d1465) I(d1466) I(d1467) I(d1468) I(d1469) I(d1470) I(d1471) I(d1472) I(d1473) I(d1474) I(d1475) I(d1476) I(d1477) I(d1478) I(d1479) I(d1480) I(d1481) I(d1482) I(d1483) I(d1484) I(d1485) I(d1486) I(d1487) I(d1488) I(d1489) I(d1490) I(d1491) I(d1492) I(d1493) I(d1494) I(d1495) I(d1496) I(d1497) I(d1498) I(d1499) I(d1500) I(d1501) I(d1502) I(d1503) I(d1504) I(d1505) I(d1506) I(d1507) I(d1508) I(d1509) I(d1510) I(d1511) I(d1512) I(d1513) I(d1514) I(d1515) I(d1516) I(d1517) I(d1518) I(d1519) I(d1520) I(d1521) I(d1522) I(d1523) I(d1524) I(d1525) I(d1526) I(d1527) I(d1528) I(d1529) I(d1530) I(d1531) I(d1532) I(d1533) I(d1534) I(d1535) I(d1536) I(d1537) I(d1538) I(d1539) I(d1540) I(d1541) I(d1542) I(d1543) I(d1544) I(d1545) I(d1546) I(d1547) I(d1548) I(d1549) I(d1550) I(d1551) I(d1552) I(d1553) I(d1554) I(d1555) I(d1556) I(d1557) I(d1558) I(d1559) I(d1560) I(d1561) I(d1562) I(d1563) I(d1564) I(d1565) I(d1566) I(d1567) I(d1568) I(d1569) I(d1570) I(d1571) I(d1572) I(d1573) I(d1574) I(d1575) I(d1576) I(d1577) I(d1578) I(d1579) I(d1580) I(d1581) I(d1582) I(d1583) I(d1584) I(d1585) I(d1586) I(d1587) I(d1588) I(d1589) I(d1590) I(d1591) I(d1592) I(d1593) I(d1594) I(d1595) I(d1596) I(d1597) I(d1598) I(d1599) I(d1600) I(d1601) I(d1602) I(d1603) I(d1604) I(d1605) I(d1606) I(d1607) I(d1608) I(d1609) I(d1610) I(d1611) I(d1612) I(d1613) I(d1614) I(d1615) I(d1616) I(d1617) I(d1618) I(d1619) I(d1620) I(d1621) I(d1622) I(d1623) I(d1624) I(d1625) I(d1626) I(d1627) I(d1628) I(d1629) I(d1630) I(d1631) I(d1632) I(d1633) I(d1634) I(d1635) I(d1636) I(d1637) I(d1638) I(d1639) I(d1640) I(d1641) I(d1642) I(d1643) I(d1644) I(d1645) I(d1646) I(d1647) I(d1648) I(d1649) I(d1650) I(d1651) I(d1652) I(d1653) I(d1654) I(d1655) I(d1656) I(d1657) I(d1658) I(d1659) I(d1660) I(d1661) I(d1662) I(d1663) I(d1664) I(d1665) I(d1666) I(d1667) I(d1668) I(d1669) I(d1670) I(d1671) I(d1672) I(d1673) I(d1674) I(d1675) I(d1676) I(d1677) I(d1678) I(d1679) I(d1680) I(d1681) I(d1682) I(d1683) I(d1684) I(d1685) I(d1686) I(d1687) I(d1688) I(d1689) I(d1690) I(d1691) I(d1692) I(d1693) I(d1694) I(d1695) I(d1696) I(d1697) I(d1698) I(d1699) I(d1700) I(d1701) I(d1702) I(d1703) I(d1704) I(d1705) I(d1706) I(d1707) I(d1708) I(d1709) I(d1710) I(d1711) I(d1712) I(d1713) I(d1714) I(d1715) I(d1716) I(d1717) I(d1718) I(d1719) I(d1720) I(d1721) I(d1722) I(d1723) I(d1724) I(d1725) I(d1726) I(d1727) I(d1728) I(d1729) I(d1730) I(d1731) I(d1732) I(d1733) I(d1734) I(d1735) I(d1736) I(d1737) I(d1738) I(d1739) I(d1740) I(d1741) I(d1742) I(d1743) I(d1744) I(d1745) I(d1746) I(d1747) I(d1748) I(d1749) I(d1750) I(d1751) I(d1752) I(d1753) I(d1754) I(d1755) I(d1756) I(d1757) I(d1758) I(d1759) I(d1760) I(d1761) I(d1762) I(d1763) I(d1764) I(d1765) I(d1766) I(d1767) I(d1768) I(d1769) I(d1770) I(d1771) I(d1772) I(d1773) I(d1774) I(d1775) I(d1776) I(d1777) I(d1778) I(d1779) I(d1780) I(d1781) I(d1782) I(d1783) I(d1784) I(d1785) I(d1786) I(d1787) I(d1788) I(d1789) I(d1790) I(d1791) I(d1792) I(d1793) I(d1794) I(d1795) I(d1796) I(d1797) I(d1798) I(d1799) I(d1800) I(d1801) I(d1802) I(d1803) I(d1804) I(d1805) I(d1806) I(d1807) I(d1808) I(d1809) I(d1810) I(d1811) I(d1812) I(d1813) I(d1814) I(d1815) I(d1816) I(d1817) I(d1818) I(d1819) I(d1820) I(d1821) I(d1822) I(d1823) I(d1824) I(d1825) I(d1826) I(d1827) I(d1828) I(d1829) I(d1830) I(d1831) I(d1832) I(d1833) I(d1834) I(d1835) I(d1836) I(d1837) I(d1838) I(d1839) I(d1840) I(d1841) I(d1842) I(d1843) I(d1844) I(d1845) I(d1846) I(d1847) I(d1848) I(d1849) I(d1850) I(d1851) I(d1852) I(d1853) I(d1854) I(d1855) I(d1856) I(d1857) I(d1858) I(d1859) I(d1860) I(d1861) I(d1862) I(d1863) I(d1864) I(d1865) I(d1866) I(d1867) I(d1868) I(d1869) I(d1870) I(d1871) I(d1872) I(d1873) I(d1874) I(d1875) I(d1876) I(d1877) I(d1878) I(d1879) I(d1880) I(d1881) I(d1882) I(d1883) I(d1884) I(d1885) I(d1886) I(d1887) I(d1888) I(d1889) I(d1890) I(d1891) I(d1892) I(d1893) I(d1894) I(d1895) I(d1896) I(d1897) I(d1898) I(d1899) I(d1900) I(d1901) I(d1902) I(d1903) I(d1904) I(d1905) I(d1906) I(d1907) I(d1908) I(d1909) I(d1910) I(d1911) I(d1912) I(d1913) I(d1914) I(d1915) I(d1916) I(d1917) I(d1918) I(d1919) I(d1920) I(d1921) I(d1922) I(d1923) I(d1924) I(d1925) I(d1926) I(d1927) I(d1928) I(d1929) I(d1930) I(d1931) I(d1932) I(d1933) I(d1934) I(d1935) I(d1936) I(d1937) I(d1938) I(d1939) I(d1940) I(d1941) I(d1942) I(d1943) I(d1944) I(d1945) I(d1946) I(d1947) I(d1948) I(d1949) I(d1950) I(d1951) I(d1952) I(d1953) I(d1954) I(d1955) I(d1956) I(d1957) I(d1958) I(d1959) I(d1960) I(d1961) I(d1962) I(d1963) I(d1964) I(d1965) I(d1966) I(d1967) I(d1968) I(d1969) I(d1970) I(d1971) I(d1972) I(d1973) I(d1974) I(d1975) I(d1976) I(d1977) I(d1978) I(d1979) I(d1980) I(d1981) I(d1982) I(d1983) I(d1984) I(d1985) I(d1986) I(d1987) I(d1988) I(d1989) I(d1990) I(d1991) I(d1992) I(d1993) I(d1994) I(d1995) I(d1996) I(d1997) I(d1998) I(d1999) I(d2000) I(d2001) I(d2002) I(d2003) I(d2004) I(d2005) I(d2006) I(d2007) I(d2008) I(d2009) I(d2010) I(d2011) I(d2012) I(d2013) I(d2014) I(d2015) I(d2016) I(d2017) I(d2018) I(d2019) I(d2020) I(d2021) I(d2022) I(d2023) I(d2024) I(d2025) I(d2026) I(d2027) I(d2028) I(d2029) I(d2030) I(d2031) I(d2032) I(d2033) I(d2034) I(d2035) I(d2036) I(d2037) I(d2038) I(d2039) I(d2040) I(d2041) I(d2042) I(d2043) I(d2044) I(d2045) I(d2046) I(d2047) I(d2048) I(d2049) I(d2050) I(d2051) I(d2052) I(d2053) I(d2054) I(d2055) I(d2056) I(d2057) I(d2058) I(d2059) I(d2060) I(d2061) I(d2062) I(d2063) I(d2064) I(d2065) I(d2066) I(d2067) I(d2068) I(d2069) I(d2070) I(d2071) I(d2072) I(d2073) I(d2074) I(d2075) I(d2076) I(d2077) I(d2078) I(d2079) I(d2080) I(d2081) I(d2082) I(d2083) I(d2084) I(d2085) I(d2086) I(d2087) I(d2088) I(d2089) I(d2090) I(d2091) I(d2092) I(d2093) I(d2094) I(d2095) I(d2096) I(d2097) I(d2098) I(d2099) I(d2100) I(d2101) I(d2102) I(d2103) I(d2104) I(d2105) I(d2106) I(d2107) I(d2108) I(d2109) I(d2110) I(d2111) I(d2112) I(d2113) I(d2114) I(d2115) I(d2116) I(d2117) I(d2118) I(d2119) I(d2120) I(d2121) I(d2122) I(d2123) I(d2124) I(d2125) I(d2126) I(d2127) I(d2128) I(d2129) I(d2130) I(d2131) I(d2132) I(d2133) I(d2134) I(d2135) I(d2136) I(d2137) I(d2138) I(d2139) I(d2140) I(d2141) I(d2142) I(d2143) I(d2144) I(d2145) I(d2146) I(d2147) I(d2148) I(d2149) I(d2150) I(d2151) I(d2152) I(d2153) I(d2154) I(d2155) I(d2156) I(d2157) I(d2158) I(d2159) I(d2160) I(d2161) I(d2162) I(d2163) I(d2164) I(d2165) I(d2166) I(d2167) I(d2168) I(d2169) I(d2170) I(d2171) I(d2172) I(d2173) I(d2174) I(d2175) I(d2176) I(d2177) I(d2178) I(d2179) I(d2180) I(d2181) I(d2182) I(d2183) I(d2184) I(d2185) I(d2186) I(d2187) I(d2188) I(d2189) I(d2190) I(d2191) I(d2192) I(d2193) I(d2194) I(d2195) I(d2196) I(d2197) I(d2198) I(d2199) I(d2200) I(d2201) I(d2202) I(d2203) I(d2204) I(d2205) I(d2206) I(d2207) I(d2208) I(d2209) I(d2210) I(d2211) I(d2212) I(d2213) I(d2214) I(d2215) I(d2216) I(d2217) I(d2218) I(d2219) I(d2220) I(d2221) I(d2222) I(d2223) I(d2224) I(d2225) I(d2226) I(d2227) I(d2228) I(d2229) I(d2230) I(d2231) I(d2232) I(d2233) I(d2234) I(d2235) I(d2236) I(d2237) I(d2238) I(d2239) I(d2240) I(d2241) I(d2242) I(d2243) I(d2244) I(d2245) I(d2246) I(d2247) I(d2248) I(d2249) I(d2250) I(d2251) I(d2252) I(d2253) I(d2254) I(d2255) I(d2256) I(d2257) I(d2258) I(d2259) I(d2260) I(d2261) I(d2262) I(d2263) I(d2264) I(d2265) I(d2266) I(d2267) I(d2268) I(d2269) I(d2270) I(d2271) I(d2272) I(d2273) I(d2274) I(d2275) I(d2276) I(d2277) I(d2278) I(d2279) I(d2280) I(d2281) I(d2282) I(d2283) I(d2284) I(d2285) I(d2286) I(d2287) I(d2288) I(d2289) I(d2290) I(d2291) I(d2292) I(d2293) I(d2294) I(d2295) I(d2296) I(d2297) I(d2298) I(d2299) I(d2300) I(d2301) I(d2302) I(d2303) I(d2304) I(d2305) I(d2306) I(d2307) I(d2308) I(d2309) I(d2310) I(d2311) I(d2312) I(d2313) I(d2314) I(d2315) I(d2316) I(d2317) I(d2318) I(d2319) I(d2320) I(d2321) I(d2322) I(d2323) I(d2324) I(d2325) I(d2326) I(d2327) I(d2328) I(d2329) I(d2330) I(d2331) I(d2332) I(d2333) I(d2334) I(d2335) I(d2336) I(d2337) I(d2338) I(d2339) I(d2340) I(d2341) I(d2342) I(d2343) I(d2344) I(d2345) I(d2346) I(d2347) I(d2348) I(d2349) I(d2350) I(d2351) I(d2352) I(d2353) I(d2354) I(d2355) I(d2356) I(d2357) I(d2358) I(d2359) I(d2360) I(d2361) I(d2362) I(d2363) I(d2364) I(d2365) I(d2366) I(d2367) I(d2368) I(d2369) I(d2370) I(d2371) I(d2372) I(d2373) I(d2374) I(d2375) I(d2376) I(d2377) I(d2378) I(d2379) I(d2380) I(d2381) I(d2382) I(d2383) I(d2384) I(d2385) I(d2386) I(d2387) I(d2388) I(d2389) I(d2390) I(d2391) I(d2392) I(d2393) I(d2394) I(d2395) I(d2396) I(d2397) I(d2398) I(d2399) I(d2400) I(d2401) I(d2402) I(d2403) I(d2404) I(d2405) I(d2406) I(d2407) I(d2408) I(d2409) I(d2410) I(d2411) I(d2412) I(d2413) I(d2414) I(d2415) I(d2416) I(d2417) I(d2418) I(d2419) I(d2420) I(d2421) I(d2422) I(d2423) I(d2424) I(d2425) I(d2426) I(d2427) I(d2428) I(d2429) I(d2430) I(d2431) I(d2432) I(d2433) I(d2434) I(d2435) I(d2436) I(d2437) I(d2438) I(d2439) I(d2440) I(d2441) I(d2442) I(d2443) I(d2444) I(d2445) I(d2446) I(d2447) I(d2448) I(d2449) I(d2450) I(d2451) I(d2452) I(d2453) I(d2454) I(d2455) I(d2456) I(d2457) I(d2458) I(d2459) I(d2460) I(d2461) I(d2462) I(d2463) I(d2464) I(d2465) I(d2466) I(d2467) I(d2468) I(d2469) I(d2470) I(d2471) I(d2472) I(d2473) I(d2474) I(d2475) I(d2476) I(d2477) I(d2478) I(d2479) I(d2480) I(d2481) I(d2482) I(d2483) I(d2484) I(d2485) I(d2486) I(d2487) I(d2488) I(d2489) I(d2490) I(d2491) I(d2492) I(d2493) I(d2494) I(d2495) I(d2496) I(d2497) I(d2498) I(d2499) I(d2500) I(d2501) I(d2502) I(d2503) I(d2504) I(d2505) I(d2506) I(d2507) I(d2508) I(d2509) I(d2510) I(d2511) I(d2512) I(d2513) I(d2514) I(d2515) I(d2516) I(d2517) I(d2518) I(d2519) I(d2520) I(d2521) I(d2522) I(d2523) I(d2524) I(d2525) I(d2526) I(d2527) I(d2528) I(d2529) I(d2530) I(d2531) I(d2532) I(d2533) I(d2534) I(d2535) I(d2536) I(d2537) I(d2538) I(d2539) I(d2540) I(d2541) I(d2542) I(d2543) I(d2544) I(d2545) I(d2546) I(d2547) I(d2548) I(d2549) I(d2550) I(d2551) I(d2552) I(d2553) I(d2554) I(d2555) I(d2556) I(d2557) I(d2558) I(d2559) I(d2560) I(d2561) I(d2562) I(d2563) I(d2564) I(d2565) I(d2566) I(d2567) I(d2568) I(d2569) I(d2570) I(d2571) I(d2572) I(d2573) I(d2574) I(d2575) I(d2576) I(d2577) I(d2578) I(d2579) I(d2580) I(d2581) I(d2582) I(d2583) I(d2584) I(d2585) I(d2586) I(d2587) I(d2588) I(d2589) I(d2590) I(d2591) I(d2592) I(d2593) I(d2594) I(d2595) I(d2596) I(d2597) I(d2598) I(d2599) I(d2600) I(d2601) I(d2602) I(d2603) I(d2604) I(d2605) I(d2606) I(d2607) I(d2608) I(d2609) I(d2610) I(d2611) I(d2612) I(d2613) I(d2614) I(d2615) I(d2616) I(d2617) I(d2618) I(d2619) I(d2620) I(d2621) I(d2622) I(d2623) I(d2624) I(d2625) I(d2626) I(d2627) I(d2628) I(d2629) I(d2630) I(d2631) I(d2632) I(d2633) I(d2634) I(d2635) I(d2636) I(d2637) I(d2638) I(d2639) I(d2640) I(d2641) I(d2642) I(d2643) I(d2644) I(d2645) I(d2646) I(d2647) I(d2648) I(d2649) I(d2650) I(d2651) I(d2652) I(d2653) I(d2654) I(d2655) I(d2656) I(d2657) I(d2658) I(d2659) I(d2660) I(d2661) I(d2662) I(d2663) I(d2664) I(d2665) I(d2666) I(d2667) I(d2668) I(d2669) I(d2670) I(d2671) I(d2672) I(d2673) I(d2674) I(d2675) I(d2676) I(d2677) I(d2678) I(d2679) I(d2680) I(d2681) I(d2682) I(d2683) I(d2684) I(d2685) I(d2686) I(d2687) I(d2688) I(d2689) I(d2690) I(d2691) I(d2692) I(d2693) I(d2694) I(d2695) I(d2696) I(d2697) I(d2698) I(d2699) I(d2700) I(d2701) I(d2702) I(d2703) I(d2704) I(d2705) I(d2706) I(d2707) I(d2708) I(d2709) I(d2710) I(d2711) I(d2712) I(d2713) I(d2714) I(d2715) I(d2716) I(d2717) I(d2718) I(d2719) I(d2720) I(d2721) I(d2722) I(d2723) I(d2724) I(d2725) I(d2726) I(d2727) I(d2728) I(d2729) I(d2730) I(d2731) I(d2732) I(d2733) I(d2734) I(d2735) I(d2736) I(d2737) I(d2738) I(d2739) I(d2740) I(d2741) I(d2742) I(d2743) I(d2744) I(d2745) I(d2746) I(d2747) I(d2748) I(d2749) I(d2750) I(d2751) I(d2752) I(d2753) I(d2754) I(d2755) I(d2756) I(d2757) I(d2758) I(d2759) I(d2760) I(d2761) I(d2762) I(d2763) I(d2764) I(d2765) I(d2766) I(d2767) I(d2768) I(d2769) I(d2770) I(d2771) I(d2772) I(d2773) I(d2774) I(d2775) I(d2776) I(d2777) I(d2778) I(d2779) I(d2780) I(d2781) I(d2782) I(d2783) I(d2784) I(d2785) I(d2786) I(d2787) I(d2788) I(d2789) I(d2790) I(d2791) I(d2792) I(d2793) I(d2794) I(d2795) I(d2796) I(d2797) I(d2798) I(d2799) I(d2800) I(d2801) I(d2802) I(d2803) I(d2804) I(d2805) I(d2806) I(d2807) I(d2808) I(d2809) I(d2810) I(d2811) I(d2812) I(d2813) I(d2814) I(d2815) I(d2816) I(d2817) I(d2818) I(d2819) I(d2820) I(d2821) I(d2822) I(d2823) I(d2824) I(d2825) I(d2826) I(d2827) I(d2828) I(d2829) I(d2830) I(d2831) I(d2832) I(d2833) I(d2834) I(d2835) I(d2836) I(d2837) I(d2838) I(d2839) I(d2840) I(d2841) I(d2842) I(d2843) I(d2844) I(d2845) I(d2846) I(d2847) I(d2848) I(d2849) I(d2850) I(d2851) I(d2852) I(d2853) I(d2854) I(d2855) I(d2856) I(d2857) I(d2858) I(d2859) I(d2860) I(d2861) I(d2862) I(d2863) I(d2864) I(d2865) I(d2866) I(d2867) I(d2868) I(d2869) I(d2870) I(d2871) I(d2872) I(d2873) I(d2874) I(d2875) I(d2876) I(d2877) I(d2878) I(d2879) I(d2880) I(d2881) I(d2882) I(d2883) I(d2884) I(d2885) I(d2886) I(d2887) I(d2888) I(d2889) I(d2890) I(d2891) I(d2892) I(d2893) I(d2894) I(d2895) I(d2896) I(d2897) I(d2898) I(d2899) I(d2900) I(d2901) I(d2902) I(d2903) I(d2904) I(d2905) I(d2906) I(d2907) I(d2908) I(d2909) I(d2910) I(d2911) I(d2912) I(d2913) I(d2914) I(d2915) I(d2916) I(d2917) I(d2918) I(d2919) I(d2920) I(d2921) I(d2922) I(d2923) I(d2924) I(d2925) I(d2926) I(d2927) I(d2928) I(d2929) I(d2930) I(d2931) I(d2932) I(d2933) I(d2934) I(d2935) I(d2936) I(d2937) I(d2938) I(d2939) I(d2940) I(d2941) I(d2942) I(d2943) I(d2944) I(d2945) I(d2946) I(d2947) I(d2948) I(d2949) I(d2950) I(d2951) I(d2952) I(d2953) I(d2954) I(d2955) I(d2956) I(d2957) I(d2958) I(d2959) I(d2960) I(d2961) I(d2962) I(d2963) I(d2964) I(d2965) I(d2966) I(d2967) I(d2968) I(d2969) I(d2970) I(d2971) I(d2972) I(d2973) I(d2974) I(d2975) I(d2976) I(d2977) I(d2978) I(d2979) I(d2980) I(d2981) I(d2982) I(d2983) I(d2984) I(d2985) I(d2986) I(d2987) I(d2988) I(d2989) I(d2990) I(d2991) I(d2992) I(d2993) I(d2994) I(d2995) I(d2996) I(d2997) I(d2998) I(d2999) I(d3000) I(d3001) I(d3002) I(d3003) I(d3004) I(d3005) I(d3006) I(d3007) I(d3008) I(d3009) I(d3010) I(d3011) I(d3012) I(d3013) I(d3014) I(d3015) I(d3016) I(d3017) I(d3018) I(d3019) I(d3020) I(d3021) I(d3022) I(d3023) I(d3024) I(d3025) I(d3026) I(d3027) I(d3028) I(d3029) I(d3030) I(d3031) I(d3032) I(d3033) I(d3034) I(d3035) I(d3036) I(d3037) I(d3038) I(d3039) I(d3040) I(d3041) I(d3042) I(d3043) I(d3044) I(d3045) I(d3046) I(d3047) I(d3048) I(d3049) I(d3050) I(d3051) I(d3052) I(d3053) I(d3054) I(d3055) I(d3056) I(d3057) I(d3058) I(d3059) I(d3060) I(d3061) I(d3062) I(d3063) I(d3064) I(d3065) I(d3066) I(d3067) I(d3068) I(d3069) I(d3070) I(d3071) I(d3072) I(d3073) I(d3074) I(d3075) I(d3076) I(d3077) I(d3078) I(d3079) I(d3080) I(d3081) I(d3082) I(d3083) I(d3084) I(d3085) I(d3086) I(d3087) I(d3088) I(d3089) I(d3090) I(d3091) I(d3092) I(d3093) I(d3094) I(d3095) I(d3096) I(d3097) I(d3098) I(d3099) I(d3100) I(d3101) I(d3102) I(d3103) I(d3104) I(d3105) I(d3106) I(d3107) I(d3108) I(d3109) I(d3110) I(d3111) I(d3112) I(d3113) I(d3114) I(d3115) I(d3116) I(d3117) I(d3118) I(d3119) I(d3120) I(d3121) I(d3122) I(d3123) I(d3124) I(d3125) I(d3126) I(d3127) I(d3128) I(d3129) I(d3130) I(d3131) I(d3132) I(d3133) I(d3134) I(d3135) I(d3136) I(d3137) I(d3138) I(d3139) I(d3140) I(d3141) I(d3142) I(d3143) I(d3144) I(d3145) I(d3146) I(d3147) I(d3148) I(d3149) I(d3150) I(d3151) I(d3152) I(d3153) I(d3154) I(d3155) I(d3156) I(d3157) I(d3158) I(d3159) I(d3160) I(d3161) I(d3162) I(d3163) I(d3164) I(d3165) I(d3166) I(d3167) I(d3168) I(d3169) I(d3170) I(d3171) I(d3172) I(d3173) I(d3174) I(d3175) I(d3176) I(d3177) I(d3178) I(d3179) I(d3180) I(d3181) I(d3182) I(d3183) I(d3184) I(d3185) I(d3186) I(d3187) I(d3188) I(d3189) I(d3190) I(d3191) I(d3192) I(d3193) I(d3194) I(d3195) I(d3196) I(d3197) I(d3198) I(d3199) I(d3200) I(d3201) I(d3202) I(d3203) I(d3204) I(d3205) I(d3206) I(d3207) I(d3208) I(d3209) I(d3210) I(d3211) I(d3212) I(d3213) I(d3214) I(d3215) I(d3216) I(d3217) I(d3218) I(d3219) I(d3220) I(d3221) I(d3222) I(d3223) I(d3224) I(d3225) I(d3226) I(d3227) I(d3228) I(d3229) I(d3230) I(d3231) I(d3232) I(d3233) I(d3234) I(d3235) I(d3236) I(d3237) I(d3238) I(d3239) I(d3240) I(d3241) I(d3242) I(d3243) I(d3244) I(d3245) I(d3246) I(d3247) I(d3248) I(d3249) I(d3250) I(d3251) I(d3252) I(d3253) I(d3254) I(d3255) I(d3256) I(d3257) I(d3258) I(d3259) I(d3260) I(d3261) I(d3262) I(d3263) I(d3264) I(d3265) I(d3266) I(d3267) I(d3268) I(d3269) I(d3270) I(d3271) I(d3272) I(d3273) I(d3274) I(d3275) I(d3276) I(d3277) I(d3278) I(d3279) I(d3280) I(d3281) I(d3282) I(d3283) I(d3284) I(d3285) I(d3286) I(d3287) I(d3288) I(d3289) I(d3290) I(d3291) I(d3292) I(d3293) I(d3294) I(d3295) I(d3296) I(d3297) I(d3298) I(d3299) I(d3300) I(d3301) I(d3302) I(d3303) I(d3304) I(d3305) I(d3306) I(d3307) I(d3308) I(d3309) I(d3310) I(d3311) I(d3312) I(d3313) I(d3314) I(d3315) I(d3316) I(d3317) I(d3318) I(d3319) I(d3320) I(d3321) I(d3322) I(d3323) I(d3324) I(d3325) I(d3326) I(d3327) I(d3328) I(d3329) I(d3330) I(d3331) I(d3332) I(d3333) I(d3334) I(d3335) I(d3336) I(d3337) I(d3338) I(d3339) I(d3340) I(d3341) I(d3342) I(d3343) I(d3344) I(d3345) I(d3346) I(d3347) I(d3348) I(d3349) I(d3350) I(d3351) I(d3352) I(d3353) I(d3354) I(d3355) I(d3356) I(d3357) I(d3358) I(d3359) I(d3360) I(d3361) I(d3362) I(d3363) I(d3364) I(d3365) I(d3366) I(d3367) I(d3368) I(d3369) I(d3370) I(d3371) I(d3372) I(d3373) I(d3374) I(d3375) I(d3376) I(d3377) I(d3378) I(d3379) I(d3380) I(d3381) I(d3382) I(d3383) I(d3384) I(d3385) I(d3386) I(d3387) I(d3388) I(d3389) I(d3390) I(d3391) I(d3392) I(d3393) I(d3394) I(d3395) I(d3396) I(d3397) I(d3398) I(d3399) I(d3400) I(d3401) I(d3402) I(d3403) I(d3404) I(d3405) I(d3406) I(d3407) I(d3408) I(d3409) I(d3410) I(d3411) I(d3412) I(d3413) I(d3414) I(d3415) I(d3416) I(d3417) I(d3418) I(d3419) I(d3420) I(d3421) I(d3422) I(d3423) I(d3424) I(d3425) I(d3426) I(d3427) I(d3428) I(d3429) I(d3430) I(d3431) I(d3432) I(d3433) I(d3434) I(d3435) I(d3436) I(d3437) I(d3438) I(d3439) I(d3440) I(d3441) I(d3442) I(d3443) I(d3444) I(d3445) I(d3446) I(d3447) I(d3448) I(d3449) I(d3450) I(d3451) I(d3452) I(d3453) I(d3454) I(d3455) I(d3456) I(d3457) I(d3458) I(d3459) I(d3460) I(d3461) I(d3462) I(d3463) I(d3464) I(d3465) I(d3466) I(d3467) I(d3468) I(d3469) I(d3470) I(d3471) I(d3472) I(d3473) I(d3474) I(d3475) I(d3476) I(d3477) I(d3478) I(d3479) I(d3480) I(d3481) I(d3482) I(d3483) I(d3484) I(d3485) I(d3486) I(d3487) I(d3488) I(d3489) I(d3490) I(d3491) I(d3492) I(d3493) I(d3494) I(d3495) I(d3496) I(d3497) I(d3498) I(d3499) I(d3500) I(d3501) I(d3502) I(d3503) I(d3504) I(d3505) I(d3506) I(d3507) I(d3508) I(d3509) I(d3510) I(d3511) I(d3512) I(d3513) I(d3514) I(d3515) I(d3516) I(d3517) I(d3518) I(d3519) I(d3520) I(d3521) I(d3522) I(d3523) I(d3524) I(d3525) I(d3526) I(d3527) I(d3528) I(d3529) I(d3530) I(d3531) I(d3532) I(d3533) I(d3534) I(d3535) I(d3536) I(d3537) I(d3538) I(d3539) I(d3540) I(d3541) I(d3542) I(d3543) I(d3544) I(d3545) I(d3546) I(d3547) I(d3548) I(d3549) I(d3550) I(d3551) I(d3552) I(d3553) I(d3554) I(d3555) I(d3556) I(d3557) I(d3558) I(d3559) I(d3560) I(d3561) I(d3562) I(d3563) I(d3564) I(d3565) I(d3566) I(d3567) I(d3568) I(d3569) I(d3570) I(d3571) I(d3572) I(d3573) I(d3574) I(d3575) I(d3576) I(d3577) I(d3578) I(d3579) I(d3580) I(d3581) I(d3582) I(d3583) I(d3584) I(d3585) I(d3586) I(d3587) I(d3588) I(d3589) I(d3590) I(d3591) I(d3592) I(d3593) I(d3594) I(d3595) I(d3596) I(d3597) I(d3598) I(d3599) I(d3600) I(d3601) I(d3602) I(d3603) I(d3604) I(d3605) I(d3606) I(d3607) I(d3608) I(d3609) I(d3610) I(d3611) I(d3612) I(d3613) I(d3614) I(d3615) I(d3616) I(d3617) I(d3618) I(d3619) I(d3620) I(d3621) I(d3622) I(d3623) I(d3624) I(d3625) I(d3626) I(d3627) I(d3628) I(d3629) I(d3630) I(d3631) I(d3632) I(d3633) I(d3634) I(d3635) I(d3636) I(d3637) I(d3638) I(d3639) I(d3640) I(d3641) I(d3642) I(d3643) I(d3644) I(d3645) I(d3646) I(d3647) I(d3648) I(d3649) I(d3650) I(d3651) I(d3652) I(d3653) I(d3654) I(d3655) I(d3656) I(d3657) I(d3658) I(d3659) I(d3660) I(d3661) I(d3662) I(d3663) I(d3664) I(d3665) I(d3666) I(d3667) I(d3668) I(d3669) I(d3670) I(d3671) I(d3672) I(d3673) I(d3674) I(d3675) I(d3676) I(d3677) I(d3678) I(d3679) I(d3680) I(d3681) I(d3682) I(d3683) I(d3684) I(d3685) I(d3686) I(d3687) I(d3688) I(d3689) I(d3690) I(d3691) I(d3692) I(d3693) I(d3694) I(d3695) I(d3696) I(d3697) I(d3698) I(d3699) I(d3700) I(d3701) I(d3702) I(d3703) I(d3704) I(d3705) I(d3706) I(d3707) I(d3708) I(d3709) I(d3710) I(d3711) I(d3712) I(d3713) I(d3714) I(d3715) I(d3716) I(d3717) I(d3718) I(d3719) I(d3720) I(d3721) I(d3722) I(d3723) I(d3724) I(d3725) I(d3726) I(d3727) I(d3728) I(d3729) I(d3730) I(d3731) I(d3732) I(d3733) I(d3734) I(d3735) I(d3736) I(d3737) I(d3738) I(d3739) I(d3740) I(d3741) I(d3742) I(d3743) I(d3744) I(d3745) I(d3746) I(d3747) I(d3748) I(d3749) I(d3750) I(d3751) I(d3752) I(d3753) I(d3754) I(d3755) I(d3756) I(d3757) I(d3758) I(d3759) I(d3760) I(d3761) I(d3762) I(d3763) I(d3764) I(d3765) I(d3766) I(d3767) I(d3768) I(d3769) I(d3770) I(d3771) I(d3772) I(d3773) I(d3774) I(d3775) I(d3776) I(d3777) I(d3778) I(d3779) I(d3780) I(d3781) I(d3782) I(d3783) I(d3784) I(d3785) I(d3786) I(d3787) I(d3788) I(d3789) I(d3790) I(d3791) I(d3792) I(d3793) I(d3794) I(d3795) I(d3796) I(d3797) I(d3798) I(d3799) I(d3800) I(d3801) I(d3802) I(d3803) I(d3804) I(d3805) I(d3806) I(d3807) I(d3808) I(d3809) I(d3810) I(d3811) I(d3812) I(d3813) I(d3814) I(d3815) I(d3816) I(d3817) I(d3818) I(d3819) I(d3820) I(d3821) I(d3822) I(d3823) I(d3824) I(d3825) I(d3826) I(d3827) I(d3828) I(d3829) I(d3830) I(d3831) I(d3832) I(d3833) I(d3834) I(d3835) I(d3836) I(d3837) I(d3838) I(d3839) I(d3840) I(d3841) I(d3842) I(d3843) I(d3844) I(d3845) I(d3846) I(d3847) I(d3848) I(d3849) I(d3850) I(d3851) I(d3852) I(d3853) I(d3854) I(d3855) I(d3856) I(d3857) I(d3858) I(d3859) I(d3860) I(d3861) I(d3862) I(d3863) I(d3864) I(d3865) I(d3866) I(d3867) I(d3868) I(d3869) I(d3870) I(d3871) I(d3872) I(d3873) I(d3874) I(d3875) I(d3876) I(d3877) I(d3878) I(d3879) I(d3880) I(d3881) I(d3882) I(d3883) I(d3884) I(d3885) I(d3886) I(d3887) I(d3888) I(d3889) I(d3890) I(d3891) I(d3892) I(d3893) I(d3894) I(d3895) I(d3896) I(d3897) I(d3898) I(d3899) I(d3900) I(d3901) I(d3902) I(d3903) I(d3904) I(d3905) I(d3906) I(d3907) I(d3908) I(d3909) I(d3910) I(d3911) I(d3912) I(d3913) I(d3914) I(d3915) I(d3916) I(d3917) I(d3918) I(d3919) I(d3920) I(d3921) I(d3922) I(d3923) I(d3924) I(d3925) I(d3926) I(d3927) I(d3928) I(d3929) I(d3930) I(d3931) I(d3932) I(d3933) I(d3934) I(d3935) I(d3936) I(d3937) I(d3938) I(d3939) I(d3940) I(d3941) I(d3942) I(d3943) I(d3944) I(d3945) I(d3946) I(d3947) I(d3948) I(d3949) I(d3950) I(d3951) I(d3952) I(d3953) I(d3954) I(d3955) I(d3956) I(d3957) I(d3958) I(d3959) I(d3960) I(d3961) I(d3962) I(d3963) I(d3964) I(d3965) I(d3966) I(d3967) I(d3968) I(d3969) I(d3970) I(d3971) I(d3972) I(d3973) I(d3974) I(d3975) I(d3976) I(d3977) I(d3978) I(d3979) I(d3980) I(d3981) I(d3982) I(d3983) I(d3984) I(d3985) I(d3986) I(d3987) I(d3988) I(d3989) I(d3990) I(d3991) I(d3992) I(d3993) I(d3994) I(d3995) I(d3996) I(d3997) I(d3998) I(d3999) I(d4000) I(d4001) I(d4002) I(d4003) I(d4004) I(d4005) I(d4006) I(d4007) I(d4008) I(d4009) I(d4010) I(d4011) I(d4012) I(d4013) I(d4014) I(d4015) I(d4016) I(d4017) I(d4018) I(d4019) I(d4020) I(d4021) I(d4022) I(d4023) I(d4024) I(d4025) I(d4026) I(d4027) I(d4028) I(d4029) I(d4030) I(d4031) I(d4032) I(d4033) I(d4034) I(d4035) I(d4036) I(d4037) I(d4038) I(d4039) I(d4040) I(d4041) I(d4042) I(d4043) I(d4044) I(d4045) I(d4046) I(d4047) I(d4048) I(d4049) I(d4050) I(d4051) I(d4052) I(d4053) I(d4054) I(d4055) I(d4056) I(d4057) I(d4058) I(d4059) I(d4060) I(d4061) I(d4062) I(d4063) I(d4064) I(d4065) I(d4066) I(d4067) I(d4068) I(d4069) I(d4070) I(d4071) I(d4072) I(d4073) I(d4074) I(d4075) I(d4076) I(d4077) I(d4078) I(d4079) I(d4080) I(d4081) I(d4082) I(d4083) I(d4084) I(d4085) I(d4086) I(d4087) I(d4088) I(d4089) I(d4090) I(d4091) I(d4092) I(d4093) I(d4094) I(d4095) I(d4096) I(d4097) I(d4098) I(d4099) I(d4100) I(d4101) I(d4102) I(d4103) I(d4104) I(d4105) I(d4106) I(d4107) I(d4108) I(d4109) I(d4110) I(d4111) I(d4112) I(d4113) I(d4114) I(d4115) I(d4116) I(d4117) I(d4118) I(d4119) I(d4120) I(d4121) I(d4122) I(d4123) I(d4124) I(d4125) I(d4126) I(d4127) I(d4128) I(d4129) I(d4130) I(d4131) I(d4132) I(d4133) I(d4134) I(d4135) I(d4136) I(d4137) I(d4138) I(d4139) I(d4140) I(d4141) I(d4142) I(d4143) I(d4144) I(d4145) I(d4146) I(d4147) I(d4148) I(d4149) I(d4150) I(d4151) I(d4152) I(d4153) I(d4154) I(d4155) I(d4156) I(d4157) I(d4158) I(d4159) I(d4160) I(d4161) I(d4162) I(d4163) I(d4164) I(d4165) I(d4166) I(d4167) I(d4168) I(d4169) I(d4170) I(d4171) I(d4172) I(d4173) I(d4174) I(d4175) I(d4176) I(d4177) I(d4178) I(d4179) I(d4180) I(d4181) I(d4182) I(d4183) I(d4184) I(d4185) I(d4186) I(d4187) I(d4188) I(d4189) I(d4190) I(d4191) I(d4192) I(d4193) I(d4194) I(d4195) I(d4196) I(d4197) I(d4198) I(d4199) I(d4200) I(d4201) I(d4202) I(d4203) I(d4204) I(d4205) I(d4206) I(d4207) I(d4208) I(d4209) I(d4210) I(d4211) I(d4212) I(d4213) I(d4214) I(d4215) I(d4216) I(d4217) I(d4218) I(d4219) I(d4220) I(d4221) I(d4222) I(d4223) I(d4224) I(d4225) I(d4226) I(d4227) I(d4228) I(d4229) I(d4230) I(d4231) I(d4232) I(d4233) I(d4234) I(d4235) I(d4236) I(d4237) I(d4238) I(d4239) I(d4240) I(d4241) I(d4242) I(d4243) I(d4244) I(d4245) I(d4246) I(d4247) I(d4248) I(d4249) I(d4250) I(d4251) I(d4252) I(d4253) I(d4254) I(d4255) I(d4256) I(d4257) I(d4258) I(d4259) I(d4260) I(d4261) I(d4262) I(d4263) I(d4264) I(d4265) I(d4266) I(d4267) I(d4268) I(d4269) I(d4270) I(d4271) I(d4272) I(d4273) I(d4274) I(d4275) I(d4276) I(d4277) I(d4278) I(d4279) I(d4280) I(d4281) I(d4282) I(d4283) I(d4284) I(d4285) I(d4286) I(d4287) I(d4288) I(d4289) I(d4290) I(d4291) I(d4292) I(d4293) I(d4294) I(d4295) I(d4296) I(d4297) I(d4298) I(d4299) I(d4300) I(d4301) I(d4302) I(d4303) I(d4304) I(d4305) I(d4306) I(d4307) I(d4308) I(d4309) I(d4310) I(d4311) I(d4312) I(d4313) I(d4314) I(d4315) I(d4316) I(d4317) I(d4318) I(d4319) I(d4320) I(d4321) I(d4322) I(d4323) I(d4324) I(d4325) I(d4326) I(d4327) I(d4328) I(d4329) I(d4330) I(d4331) I(d4332) I(d4333) I(d4334) I(d4335) I(d4336) I(d4337) I(d4338) I(d4339) I(d4340) I(d4341) I(d4342) I(d4343) I(d4344) I(d4345) I(d4346) I(d4347) I(d4348) I(d4349) I(d4350) I(d4351) I(d4352) I(d4353) I(d4354) I(d4355) I(d4356) I(d4357) I(d4358) I(d4359) I(d4360) I(d4361) I(d4362) I(d4363) I(d4364) I(d4365) I(d4366) I(d4367) I(d4368) I(d4369) I(d4370) I(d4371) I(d4372) I(d4373) I(d4374) I(d4375) I(d4376) I(d4377) I(d4378) I(d4379) I(d4380) I(d4381) I(d4382) I(d4383) I(d4384) I(d4385) I(d4386) I(d4387) I(d4388) I(d4389) I(d4390) I(d4391) I(d4392) I(d4393) I(d4394) I(d4395) I(d4396) I(d4397) I(d4398) I(d4399) I(d4400) I(d4401) I(d4402) I(d4403) I(d4404) I(d4405) I(d4406) I(d4407) I(d4408) I(d4409) I(d4410) I(d4411) I(d4412) I(d4413) I(d4414) I(d4415) I(d4416) I(d4417) I(d4418) I(d4419) I(d4420) I(d4421) I(d4422) I(d4423) I(d4424) I(d4425) I(d4426) I(d4427) I(d4428) I(d4429) I(d4430) I(d4431) I(d4432) I(d4433) I(d4434) I(d4435) I(d4436) I(d4437) I(d4438) I(d4439) I(d4440) I(d4441) I(d4442) I(d4443) I(d4444) I(d4445) I(d4446) I(d4447) I(d4448) I(d4449) I(d4450) I(d4451) I(d4452) I(d4453) I(d4454) I(d4455) I(d4456) I(d4457) I(d4458) I(d4459) I(d4460) I(d4461) I(d4462) I(d4463) I(d4464) I(d4465) I(d4466) I(d4467) I(d4468) I(d4469) I(d4470) I(d4471) I(d4472) I(d4473) I(d4474) I(d4475) I(d4476) I(d4477) I(d4478) I(d4479) I(d4480) I(d4481) I(d4482) I(d4483) I(d4484) I(d4485) I(d4486) I(d4487) I(d4488) I(d4489) I(d4490) I(d4491) I(d4492) I(d4493) I(d4494) I(d4495) I(d4496) I(d4497) I(d4498) I(d4499) I(d4500) I(d4501) I(d4502) I(d4503) I(d4504) I(d4505) I(d4506) I(d4507) I(d4508) I(d4509) I(d4510) I(d4511) I(d4512) I(d4513) I(d4514) I(d4515) I(d4516) I(d4517) I(d4518) I(d4519) I(d4520) I(d4521) I(d4522) I(d4523) I(d4524) I(d4525) I(d4526) I(d4527) I(d4528) I(d4529) I(d4530) I(d4531) I(d4532) I(d4533) I(d4534) I(d4535) I(d4536) I(d4537) I(d4538) I(d4539) I(d4540) I(d4541) I(d4542) I(d4543) I(d4544) I(d4545) I(d4546) I(d4547) I(d4548) I(d4549) I(d4550) I(d4551) I(d4552) I(d4553) I(d4554) I(d4555) I(d4556) I(d4557) I(d4558) I(d4559) I(d4560) I(d4561) I(d4562) I(d4563) I(d4564) I(d4565) I(d4566) I(d4567) I(d4568) I(d4569) I(d4570) I(d4571) I(d4572) I(d4573) I(d4574) I(d4575) I(d4576) I(d4577) I(d4578) I(d4579) I(d4580) I(d4581) I(d4582) I(d4583) I(d4584) I(d4585) I(d4586) I(d4587) I(d4588) I(d4589) I(d4590) I(d4591) I(d4592) I(d4593) I(d4594) I(d4595) I(d4596) I(d4597) I(d4598) I(d4599) I(d4600) I(d4601) I(d4602) I(d4603) I(d4604) I(d4605) I(d4606) I(d4607) I(d4608) I(d4609) I(d4610) I(d4611) I(d4612) I(d4613) I(d4614) I(d4615) I(d4616) I(d4617) I(d4618) I(d4619) I(d4620) I(d4621) I(d4622) I(d4623) I(d4624) I(d4625) I(d4626) I(d4627) I(d4628) I(d4629) I(d4630) I(d4631) I(d4632) I(d4633) I(d4634) I(d4635) I(d4636) I(d4637) I(d4638) I(d4639) I(d4640) I(d4641) I(d4642) I(d4643) I(d4644) I(d4645) I(d4646) I(d4647) I(d4648) I(d4649) I(d4650) I(d4651) I(d4652) I(d4653) I(d4654) I(d4655) I(d4656) I(d4657) I(d4658) I(d4659) I(d4660) I(d4661) I(d4662) I(d4663) I(d4664) I(d4665) I(d4666) I(d4667) I(d4668) I(d4669) I(d4670) I(d4671) I(d4672) I(d4673) I(d4674) I(d4675) I(d4676) I(d4677) I(d4678) I(d4679) I(d4680) I(d4681) I(d4682) I(d4683) I(d4684) I(d4685) I(d4686) I(d4687) I(d4688) I(d4689) I(d4690) I(d4691) I(d4692) I(d4693) I(d4694) I(d4695) I(d4696) I(d4697) I(d4698) I(d4699) I(d4700) I(d4701) I(d4702) I(d4703) I(d4704) I(d4705) I(d4706) I(d4707) I(d4708) I(d4709) I(d4710) I(d4711) I(d4712) I(d4713) I(d4714) I(d4715) I(d4716) I(d4717) I(d4718) I(d4719) I(d4720) I(d4721) I(d4722) I(d4723) I(d4724) I(d4725) I(d4726) I(d4727) I(d4728) I(d4729) I(d4730) I(d4731) I(d4732) I(d4733) I(d4734) I(d4735) I(d4736) I(d4737) I(d4738) I(d4739) I(d4740) I(d4741) I(d4742) I(d4743) I(d4744) I(d4745) I(d4746) I(d4747) I(d4748) I(d4749) I(d4750) I(d4751) I(d4752) I(d4753) I(d4754) I(d4755) I(d4756) I(d4757) I(d4758) I(d4759) I(d4760) I(d4761) I(d4762) I(d4763) I(d4764) I(d4765) I(d4766) I(d4767) I(d4768) I(d4769) I(d4770) I(d4771) I(d4772) I(d4773) I(d4774) I(d4775) I(d4776) I(d4777) I(d4778) I(d4779) I(d4780) I(d4781) I(d4782) I(d4783) I(d4784) I(d4785) I(d4786) I(d4787) I(d4788) I(d4789) I(d4790) I(d4791) I(d4792) I(d4793) I(d4794) I(d4795) I(d4796) I(d4797) I(d4798) I(d4799) I(d4800) I(d4801) I(d4802) I(d4803) I(d4804) I(d4805) I(d4806) I(d4807) I(d4808) I(d4809) I(d4810) I(d4811) I(d4812) I(d4813) I(d4814) I(d4815) I(d4816) I(d4817) I(d4818) I(d4819) I(d4820) I(d4821) I(d4822) I(d4823) I(d4824) I(d4825) I(d4826) I(d4827) I(d4828) I(d4829) I(d4830) I(d4831) I(d4832) I(d4833) I(d4834) I(d4835) I(d4836) I(d4837) I(d4838) I(d4839) I(d4840) I(d4841) I(d4842) I(d4843) I(d4844) I(d4845) I(d4846) I(d4847) I(d4848) I(d4849) I(d4850) I(d4851) I(d4852) I(d4853) I(d4854) I(d4855) I(d4856) I(d4857) I(d4858) I(d4859) I(d4860) I(d4861) I(d4862) I(d4863) I(d4864) I(d4865) I(d4866) I(d4867) I(d4868) I(d4869) I(d4870) I(d4871) I(d4872) I(d4873) I(d4874) I(d4875) I(d4876) I(d4877) I(d4878) I(d4879) I(d4880) I(d4881) I(d4882) I(d4883) I(d4884) I(d4885) I(d4886) I(d4887) I(d4888) I(d4889) I(d4890) I(d4891) I(d4892) I(d4893) I(d4894) I(d4895) I(d4896) I(d4897) I(d4898) I(d4899) I(d4900) I(d4901) I(d4902) I(d4903) I(d4904) I(d4905) I(d4906) I(d4907) I(d4908) I(d4909) I(d4910) I(d4911) I(d4912) I(d4913) I(d4914) I(d4915) I(d4916) I(d4917) I(d4918) I(d4919) I(d4920) I(d4921) I(d4922) I(d4923) I(d4924) I(d4925) I(d4926) I(d4927) I(d4928) I(d4929) I(d4930) I(d4931) I(d4932) I(d4933) I(d4934) I(d4935) I(d4936) I(d4937) I(d4938) I(d4939) I(d4940) I(d4941) I(d4942) I(d4943) I(d4944) I(d4945) I(d4946) I(d4947) I(d4948) I(d4949) I(d4950) I(d4951) I(d4952) I(d4953) I(d4954) I(d4955) I(d4956) I(d4957) I(d4958) I(d4959) I(d4960) I(d4961) I(d4962) I(d4963) I(d4964) I(d4965) I(d4966) I(d4967) I(d4968) I(d4969) I(d4970) I(d4971) I(d4972) I(d4973) I(d4974) I(d4975) I(d4976) I(d4977) I(d4978) I(d4979) I(d4980) I(d4981) I(d4982) I(d4983) I(d4984) I(d4985) I(d4986) I(d4987) I(d4988) I(d4989) I(d4990) I(d4991) I(d4992) I(d4993) I(d4994) I(d4995) I(d4996) I(d4997) I(d4998) I(d4999) I(d5000) I(d5001) I(d5002) I(d5003) I(d5004) I(d5005) I(d5006) I(d5007) I(d5008) I(d5009) I(d5010) I(d5011) I(d5012) I(d5013) I(d5014) I(d5015) I(d5016) I(d5017) I(d5018) I(d5019) I(d5020) I(d5021) I(d5022) I(d5023) I(d5024) I(d5025) I(d5026) I(d5027) I(d5028) I(d5029) I(d5030) I(d5031) I(d5032) I(d5033) I(d5034) I(d5035) I(d5036) I(d5037) I(d5038) I(d5039) I(d5040) I(d5041) I(d5042) I(d5043) I(d5044) I(d5045) I(d5046) I(d5047) I(d5048) I(d5049) I(d5050) I(d5051) I(d5052) I(d5053) I(d5054) I(d5055) I(d5056) I(d5057) I(d5058) I(d5059) I(d5060) I(d5061) I(d5062) I(d5063) I(d5064) I(d5065) I(d5066) I(d5067) I(d5068) I(d5069) I(d5070) I(d5071) I(d5072) I(d5073) I(d5074) I(d5075) I(d5076) I(d5077) I(d5078) I(d5079) I(d5080) I(d5081) I(d5082) I(d5083) I(d5084) I(d5085) I(d5086) I(d5087) I(d5088) I(d5089) I(d5090) I(d5091) I(d5092) I(d5093) I(d5094) I(d5095) I(d5096) I(d5097) I(d5098) I(d5099) I(d5100) I(d5101) I(d5102) I(d5103) I(d5104) I(d5105) I(d5106) I(d5107) I(d5108) I(d5109) I(d5110) I(d5111) I(d5112) I(d5113) I(d5114) I(d5115) I(d5116) I(d5117) I(d5118) I(d5119) I(d5120) I(d5121) I(d5122) I(d5123) I(d5124) I(d5125) I(d5126) I(d5127) I(d5128) I(d5129) I(d5130) I(d5131) I(d5132) I(d5133) I(d5134) I(d5135) I(d5136) I(d5137) I(d5138) I(d5139) I(d5140) I(d5141) I(d5142) I(d5143) I(d5144) I(d5145) I(d5146) I(d5147) I(d5148) I(d5149) I(d5150) I(d5151) I(d5152) I(d5153) I(d5154) I(d5155) I(d5156) I(d5157) I(d5158) I(d5159) I(d5160) I(d5161) I(d5162) I(d5163) I(d5164) I(d5165) I(d5166) I(d5167) I(d5168) I(d5169) I(d5170) I(d5171) I(d5172) I(d5173) I(d5174) I(d5175) I(d5176) I(d5177) I(d5178) I(d5179) I(d5180) I(d5181) I(d5182) I(d5183) I(d5184) I(d5185) I(d5186) I(d5187) I(d5188) I(d5189) I(d5190) I(d5191) I(d5192) I(d5193) I(d5194) I(d5195) I(d5196) I(d5197) I(d5198) I(d5199) I(d5200) I(d5201) I(d5202) I(d5203) I(d5204) I(d5205) I(d5206) I(d5207) I(d5208) I(d5209) I(d5210) I(d5211) I(d5212) I(d5213) I(d5214) I(d5215) I(d5216) I(d5217) I(d5218) I(d5219) I(d5220) I(d5221) I(d5222) I(d5223) I(d5224) I(d5225) I(d5226) I(d5227) I(d5228) I(d5229) I(d5230) I(d5231) I(d5232) I(d5233) I(d5234) I(d5235) I(d5236) I(d5237) I(d5238) I(d5239) I(d5240) I(d5241) I(d5242) I(d5243) I(d5244) I(d5245) I(d5246) I(d5247) I(d5248) I(d5249) I(d5250) I(d5251) I(d5252) I(d5253) I(d5254) I(d5255) I(d5256) I(d5257) I(d5258) I(d5259) I(d5260) I(d5261) I(d5262) I(d5263) I(d5264) I(d5265) I(d5266) I(d5267) I(d5268) I(d5269) I(d5270) I(d5271) I(d5272) I(d5273) I(d5274) I(d5275) I(d5276) I(d5277) I(d5278) I(d5279) I(d5280) I(d5281) I(d5282) I(d5283) I(d5284) I(d5285) I(d5286) I(d5287) I(d5288) I(d5289) I(d5290) I(d5291) I(d5292) I(d5293) I(d5294) I(d5295) I(d5296) I(d5297) I(d5298) I(d5299) I(d5300) I(d5301) I(d5302) I(d5303) I(d5304) I(d5305) I(d5306) I(d5307) I(d5308) I(d5309) I(d5310) I(d5311) I(d5312) I(d5313) I(d5314) I(d5315) I(d5316) I(d5317) I(d5318) I(d5319) I(d5320) I(d5321) I(d5322) I(d5323) I(d5324) I(d5325) I(d5326) I(d5327) I(d5328) I(d5329) I(d5330) I(d5331) I(d5332) I(d5333) I(d5334) I(d5335) I(d5336) I(d5337) I(d5338) I(d5339) I(d5340) I(d5341) I(d5342) I(d5343) I(d5344) I(d5345) I(d5346) I(d5347) I(d5348) I(d5349) I(d5350) I(d5351) I(d5352) I(d5353) I(d5354) I(d5355) I(d5356) I(d5357) I(d5358) I(d5359) I(d5360) I(d5361) I(d5362) I(d5363) I(d5364) I(d5365) I(d5366) I(d5367) I(d5368) I(d5369) I(d5370) I(d5371) I(d5372) I(d5373) I(d5374) I(d5375) I(d5376) I(d5377) I(d5378) I(d5379) I(d5380) I(d5381) I(d5382) I(d5383) I(d5384) I(d5385) I(d5386) I(d5387) I(d5388) I(d5389) I(d5390) I(d5391) I(d5392) I(d5393) I(d5394) I(d5395) I(d5396) I(d5397) I(d5398) I(d5399) I(d5400) I(d5401) I(d5402) I(d5403) I(d5404) I(d5405) I(d5406) I(d5407) I(d5408) I(d5409) I(d5410) I(d5411) I(d5412) I(d5413) I(d5414) I(d5415) I(d5416) I(d5417) I(d5418) I(d5419) I(d5420) I(d5421) I(d5422) I(d5423) I(d5424) I(d5425) I(d5426) I(d5427) I(d5428) I(d5429) I(d5430) I(d5431) I(d5432) I(d5433) I(d5434) I(d5435) I(d5436) I(d5437) I(d5438) I(d5439) I(d5440) I(d5441) I(d5442) I(d5443) I(d5444) I(d5445) I(d5446) I(d5447) I(d5448) I(d5449) I(d5450) I(d5451) I(d5452) I(d5453) I(d5454) I(d5455) I(d5456) I(d5457) I(d5458) I(d5459) I(d5460) I(d5461) I(d5462) I(d5463) I(d5464) I(d5465) I(d5466) I(d5467) I(d5468) I(d5469) I(d5470) I(d5471) I(d5472) I(d5473) I(d5474) I(d5475) I(d5476) I(d5477) I(d5478) I(d5479) I(d5480) I(d5481) I(d5482) I(d5483) I(d5484) I(d5485) I(d5486) I(d5487) I(d5488) I(d5489) I(d5490) I(d5491) I(d5492) I(d5493) I(d5494) I(d5495) I(d5496) I(d5497) I(d5498) I(d5499) I(d5500) I(d5501) I(d5502) I(d5503) I(d5504) I(d5505) I(d5506) I(d5507) I(d5508) I(d5509) I(d5510) I(d5511) I(d5512) I(d5513) I(d5514) I(d5515) I(d5516) I(d5517) I(d5518) I(d5519) I(d5520) I(d5521) I(d5522) I(d5523) I(d5524) I(d5525) I(d5526) I(d5527) I(d5528) I(d5529) I(d5530) I(d5531) I(d5532) I(d5533) I(d5534) I(d5535) I(d5536) I(d5537) I(d5538) I(d5539) I(d5540) I(d5541) I(d5542) I(d5543) I(d5544) I(d5545) I(d5546) I(d5547) I(d5548) I(d5549) I(d5550) I(d5551) I(d5552) I(d5553) I(d5554) I(d5555) I(d5556) I(d5557) I(d5558) I(d5559) I(d5560) I(d5561) I(d5562) I(d5563) I(d5564) I(d5565) I(d5566) I(d5567) I(d5568) I(d5569) I(d5570) I(d5571) I(d5572) I(d5573) I(d5574) I(d5575) I(d5576) I(d5577) I(d5578) I(d5579) I(d5580) I(d5581) I(d5582) I(d5583) I(d5584) I(d5585) I(d5586) I(d5587) I(d5588) I(d5589) I(d5590) I(d5591) I(d5592) I(d5593) I(d5594) I(d5595) I(d5596) I(d5597) I(d5598) I(d5599) I(d5600) I(d5601) I(d5602) I(d5603) I(d5604) I(d5605) I(d5606) I(d5607) I(d5608) I(d5609) I(d5610) I(d5611) I(d5612) I(d5613) I(d5614) I(d5615) I(d5616) I(d5617) I(d5618) I(d5619) I(d5620) I(d5621) I(d5622) I(d5623) I(d5624) I(d5625) I(d5626) I(d5627) I(d5628) I(d5629) I(d5630) I(d5631) I(d5632) I(d5633) I(d5634) I(d5635) I(d5636) I(d5637) I(d5638) I(d5639) I(d5640) I(d5641) I(d5642) I(d5643) I(d5644) I(d5645) I(d5646) I(d5647) I(d5648) I(d5649) I(d5650) I(d5651) I(d5652) I(d5653) I(d5654) I(d5655) I(d5656) I(d5657) I(d5658) I(d5659) I(d5660) I(d5661) I(d5662) I(d5663) I(d5664) I(d5665) I(d5666) I(d5667) I(d5668) I(d5669) I(d5670) I(d5671) I(d5672) I(d5673) I(d5674) I(d5675) I(d5676) I(d5677) I(d5678) I(d5679) I(d5680) I(d5681) I(d5682) I(d5683) I(d5684) I(d5685) I(d5686) I(d5687) I(d5688) I(d5689) I(d5690) I(d5691) I(d5692) I(d5693) I(d5694) I(d5695) I(d5696) I(d5697) I(d5698) I(d5699) I(d5700) I(d5701) I(d5702) I(d5703) I(d5704) I(d5705) I(d5706) I(d5707) I(d5708) I(d5709) I(d5710) I(d5711) I(d5712) I(d5713) I(d5714) I(d5715) I(d5716) I(d5717) I(d5718) I(d5719) I(d5720) I(d5721) I(d5722) I(d5723) I(d5724) I(d5725) I(d5726) I(d5727) I(d5728) I(d5729) I(d5730) I(d5731) I(d5732) I(d5733) I(d5734) I(d5735) I(d5736) I(d5737) I(d5738) I(d5739) I(d5740) I(d5741) I(d5742) I(d5743) I(d5744) I(d5745) I(d5746) I(d5747) I(d5748) I(d5749) I(d5750) I(d5751) I(d5752) I(d5753) I(d5754) I(d5755) I(d5756) I(d5757) I(d5758) I(d5759) I(d5760) I(d5761) I(d5762) I(d5763) I(d5764) I(d5765) I(d5766) I(d5767) I(d5768) I(d5769) I(d5770) I(d5771) I(d5772) I(d5773) I(d5774) I(d5775) I(d5776) I(d5777) I(d5778) I(d5779) I(d5780) I(d5781) I(d5782) I(d5783) I(d5784) I(d5785) I(d5786) I(d5787) I(d5788) I(d5789) I(d5790) I(d5791) I(d5792) I(d5793) I(d5794) I(d5795) I(d5796) I(d5797) I(d5798) I(d5799) I(d5800) I(d5801) I(d5802) I(d5803) I(d5804) I(d5805) I(d5806) I(d5807) I(d5808) I(d5809) I(d5810) I(d5811) I(d5812) I(d5813) I(d5814) I(d5815) I(d5816) I(d5817) I(d5818) I(d5819) I(d5820) I(d5821) I(d5822) I(d5823) I(d5824) I(d5825) I(d5826) I(d5827) I(d5828) I(d5829) I(d5830) I(d5831) I(d5832) I(d5833) I(d5834) I(d5835) I(d5836) I(d5837) I(d5838) I(d5839) I(d5840) I(d5841) I(d5842) I(d5843) I(d5844) I(d5845) I(d5846) I(d5847) I(d5848) I(d5849) I(d5850) I(d5851) I(d5852) I(d5853) I(d5854) I(d5855) I(d5856) I(d5857) I(d5858) I(d5859) I(d5860) I(d5861) I(d5862) I(d5863) I(d5864) I(d5865) I(d5866) I(d5867) I(d5868) I(d5869) I(d5870) I(d5871) I(d5872) I(d5873) I(d5874) I(d5875) I(d5876) I(d5877) I(d5878) I(d5879) I(d5880) I(d5881) I(d5882) I(d5883) I(d5884) I(d5885) I(d5886) I(d5887) I(d5888) I(d5889) I(d5890) I(d5891) I(d5892) I(d5893) I(d5894) I(d5895) I(d5896) I(d5897) I(d5898) I(d5899) I(d5900) I(d5901) I(d5902) I(d5903) I(d5904) I(d5905) I(d5906) I(d5907) I(d5908) I(d5909) I(d5910) I(d5911) I(d5912) I(d5913) I(d5914) I(d5915) I(d5916) I(d5917) I(d5918) I(d5919) I(d5920) I(d5921) I(d5922) I(d5923) I(d5924) I(d5925) I(d5926) I(d5927) I(d5928) I(d5929) I(d5930) I(d5931) I(d5932) I(d5933) I(d5934) I(d5935) I(d5936) I(d5937) I(d5938) I(d5939) I(d5940) I(d5941) I(d5942) I(d5943) I(d5944) I(d5945) I(d5946) I(d5947) I(d5948) I(d5949) I(d5950) I(d5951) I(d5952) I(d5953) I(d5954) I(d5955) I(d5956) I(d5957) I(d5958) I(d5959) I(d5960) I(d5961) I(d5962) I(d5963) I(d5964) I(d5965) I(d5966) I(d5967) I(d5968) I(d5969) I(d5970) I(d5971) I(d5972) I(d5973) I(d5974) I(d5975) I(d5976) I(d5977) I(d5978) I(d5979) I(d5980) I(d5981) I(d5982) I(d5983) I(d5984) I(d5985) I(d5986) I(d5987) I(d5988) I(d5989) I(d5990) I(d5991) I(d5992) I(d5993) I(d5994) I(d5995) I(d5996) I(d5997) I(d5998) I(d5999) I(d6000) I(d6001) I(d6002) I(d6003) I(d6004) I(d6005) I(d6006) I(d6007) I(d6008) I(d6009) I(d6010) I(d6011) I(d6012) I(d6013) I(d6014) I(d6015) I(d6016) I(d6017) I(d6018) I(d6019) I(d6020) I(d6021) I(d6022) I(d6023) I(d6024) I(d6025) I(d6026) I(d6027) I(d6028) I(d6029) I(d6030) I(d6031) I(d6032) I(d6033) I(d6034) I(d6035) I(d6036) I(d6037) I(d6038) I(d6039) I(d6040) I(d6041) I(d6042) I(d6043) I(d6044) I(d6045) I(d6046) I(d6047) I(d6048) I(d6049) I(d6050) I(d6051) I(d6052) I(d6053) I(d6054) I(d6055) I(d6056) I(d6057) I(d6058) I(d6059) I(d6060) I(d6061) I(d6062) I(d6063) I(d6064) I(d6065) I(d6066) I(d6067) I(d6068) I(d6069) I(d6070) I(d6071) I(d6072) I(d6073) I(d6074) I(d6075) I(d6076) I(d6077) I(d6078) I(d6079) I(d6080) I(d6081) I(d6082) I(d6083) I(d6084) I(d6085) I(d6086) I(d6087) I(d6088) I(d6089) I(d6090) I(d6091) I(d6092) I(d6093) I(d6094) I(d6095) I(d6096) I(d6097) I(d6098) I(d6099) I(d6100) I(d6101) I(d6102) I(d6103) I(d6104) I(d6105) I(d6106) I(d6107) I(d6108) I(d6109) I(d6110) I(d6111) I(d6112) I(d6113) I(d6114) I(d6115) I(d6116) I(d6117) I(d6118) I(d6119) I(d6120) I(d6121) I(d6122) I(d6123) I(d6124) I(d6125) I(d6126) I(d6127) I(d6128) I(d6129) I(d6130) I(d6131) I(d6132) I(d6133) I(d6134) I(d6135) I(d6136) I(d6137) I(d6138) I(d6139) I(d6140) I(d6141) I(d6142) I(d6143) I(d6144) I(d6145) I(d6146) I(d6147) I(d6148) I(d6149) I(d6150) I(d6151) I(d6152) I(d6153) I(d6154) I(d6155) I(d6156) I(d6157) I(d6158) I(d6159) I(d6160) I(d6161) I(d6162) I(d6163) I(d6164) I(d6165) I(d6166) I(d6167) I(d6168) I(d6169) I(d6170) I(d6171) I(d6172) I(d6173) I(d6174) I(d6175) I(d6176) I(d6177) I(d6178) I(d6179) I(d6180) I(d6181) I(d6182) I(d6183) I(d6184) I(d6185) I(d6186) I(d6187) I(d6188) I(d6189) I(d6190) I(d6191) I(d6192) I(d6193) I(d6194) I(d6195) I(d6196) I(d6197) I(d6198) I(d6199) I(d6200) I(d6201) I(d6202) I(d6203) I(d6204) I(d6205) I(d6206) I(d6207) I(d6208) I(d6209) I(d6210) I(d6211) I(d6212) I(d6213) I(d6214) I(d6215) I(d6216) I(d6217) I(d6218) I(d6219) I(d6220) I(d6221) I(d6222) I(d6223) I(d6224) I(d6225) I(d6226) I(d6227) I(d6228) I(d6229) I(d6230) I(d6231) I(d6232) I(d6233) I(d6234) I(d6235) I(d6236) I(d6237) I(d6238) I(d6239) I(d6240) I(d6241) I(d6242) I(d6243) I(d6244) I(d6245) I(d6246) I(d6247) I(d6248) I(d6249) I(d6250) I(d6251) I(d6252) I(d6253) I(d6254) I(d6255) I(d6256) I(d6257) I(d6258) I(d6259) I(d6260) I(d6261) I(d6262) I(d6263) I(d6264) I(d6265) I(d6266) I(d6267) I(d6268) I(d6269) I(d6270) I(d6271) I(d6272) I(d6273) I(d6274) I(d6275) I(d6276) I(d6277) I(d6278) I(d6279) I(d6280) I(d6281) I(d6282) I(d6283) I(d6284) I(d6285) I(d6286) I(d6287) I(d6288) I(d6289) I(d6290) I(d6291) I(d6292) I(d6293) I(d6294) I(d6295) I(d6296) I(d6297) I(d6298) I(d6299) I(d6300) I(d6301) I(d6302) I(d6303) I(d6304) I(d6305) I(d6306) I(d6307) I(d6308) I(d6309) I(d6310) I(d6311) I(d6312) I(d6313) I(d6314) I(d6315) I(d6316) I(d6317) I(d6318) I(d6319) I(d6320) I(d6321) I(d6322) I(d6323) I(d6324) I(d6325) I(d6326) I(d6327) I(d6328) I(d6329) I(d6330) I(d6331) I(d6332) I(d6333) I(d6334) I(d6335) I(d6336) I(d6337) I(d6338) I(d6339) I(d6340) I(d6341) I(d6342) I(d6343) I(d6344) I(d6345) I(d6346) I(d6347) I(d6348) I(d6349) I(d6350) I(d6351) I(d6352) I(d6353) I(d6354) I(d6355) I(d6356) I(d6357) I(d6358) I(d6359) I(d6360) I(d6361) I(d6362) I(d6363) I(d6364) I(d6365) I(d6366) I(d6367) I(d6368) I(d6369) I(d6370) I(d6371) I(d6372) I(d6373) I(d6374) I(d6375) I(d6376) I(d6377) I(d6378) I(d6379) I(d6380) I(d6381) I(d6382) I(d6383) I(d6384) I(d6385) I(d6386) I(d6387) I(d6388) I(d6389) I(d6390) I(d6391) I(d6392) I(d6393) I(d6394) I(d6395) I(d6396) I(d6397) I(d6398) I(d6399) I(d6400) I(d6401) I(d6402) I(d6403) I(d6404) I(d6405) I(d6406) I(d6407) I(d6408) I(d6409) I(d6410) I(d6411) I(d6412) I(d6413) I(d6414) I(d6415) I(d6416) I(d6417) I(d6418) I(d6419) I(d6420) I(d6421) I(d6422) I(d6423) I(d6424) I(d6425) I(d6426) I(d6427) I(d6428) I(d6429) I(d6430) I(d6431) I(d6432) I(d6433) I(d6434) I(d6435) I(d6436) I(d6437) I(d6438) I(d6439) I(d6440) I(d6441) I(d6442) I(d6443) I(d6444) I(d6445) I(d6446) I(d6447) I(d6448) I(d6449) I(d6450) I(d6451) I(d6452) I(d6453) I(d6454) I(d6455) I(d6456) I(d6457) I(d6458) I(d6459) I(d6460) I(d6461) I(d6462) I(d6463) I(d6464) I(d6465) I(d6466) I(d6467) I(d6468) I(d6469) I(d6470) I(d6471) I(d6472) I(d6473) I(d6474) I(d6475) I(d6476) I(d6477) I(d6478) I(d6479) I(d6480) I(d6481) I(d6482) I(d6483) I(d6484) I(d6485) I(d6486) I(d6487) I(d6488) I(d6489) I(d6490) I(d6491) I(d6492) I(d6493) I(d6494) I(d6495) I(d6496) I(d6497) I(d6498) I(d6499) I(d6500) I(d6501) I(d6502) I(d6503) I(d6504) I(d6505) I(d6506) I(d6507) I(d6508) I(d6509) I(d6510) I(d6511) I(d6512) I(d6513) I(d6514) I(d6515) I(d6516) I(d6517) I(d6518) I(d6519) I(d6520) I(d6521) I(d6522) I(d6523) I(d6524) I(d6525) I(d6526) I(d6527) I(d6528) I(d6529) I(d6530) I(d6531) I(d6532) I(d6533) I(d6534) I(d6535) I(d6536) I(d6537) I(d6538) I(d6539) I(d6540) I(d6541) I(d6542) I(d6543) I(d6544) I(d6545) I(d6546) I(d6547) I(d6548) I(d6549) I(d6550) I(d6551) I(d6552) I(d6553) I(d6554) I(d6555) I(d6556) I(d6557) I(d6558) I(d6559) I(d6560) I(d6561) I(d6562) I(d6563) I(d6564) I(d6565) I(d6566) I(d6567) I(d6568) I(d6569) I(d6570) I(d6571) I(d6572) I(d6573) I(d6574) I(d6575) I(d6576) I(d6577) I(d6578) I(d6579) I(d6580) I(d6581) I(d6582) I(d6583) I(d6584) I(d6585) I(d6586) I(d6587) I(d6588) I(d6589) I(d6590) I(d6591) I(d6592) I(d6593) I(d6594) I(d6595) I(d6596) I(d6597) I(d6598) I(d6599) I(d6600) I(d6601) I(d6602) I(d6603) I(d6604) I(d6605) I(d6606) I(d6607) I(d6608) I(d6609) I(d6610) I(d6611) I(d6612) I(d6613) I(d6614) I(d6615) I(d6616) I(d6617) I(d6618) I(d6619) I(d6620) I(d6621) I(d6622) I(d6623) I(d6624) I(d6625) I(d6626) I(d6627) I(d6628) I(d6629) I(d6630) I(d6631) I(d6632) I(d6633) I(d6634) I(d6635) I(d6636) I(d6637) I(d6638) I(d6639) I(d6640) I(d6641) I(d6642) I(d6643) I(d6644) I(d6645) I(d6646) I(d6647) I(d6648) I(d6649) I(d6650) I(d6651) I(d6652) I(d6653) I(d6654) I(d6655) I(d6656) I(d6657) I(d6658) I(d6659) I(d6660) I(d6661) I(d6662) I(d6663) I(d6664) I(d6665) I(d6666) I(d6667) I(d6668) I(d6669) I(d6670) I(d6671) I(d6672) I(d6673) I(d6674) I(d6675) I(d6676) I(d6677) I(d6678) I(d6679) I(d6680) I(d6681) I(d6682) I(d6683) I(d6684) I(d6685) I(d6686) I(d6687) I(d6688) I(d6689) I(d6690) I(d6691) I(d6692) I(d6693) I(d6694) I(d6695) I(d6696) I(d6697) I(d6698) I(d6699) I(d6700) I(d6701) I(d6702) I(d6703) I(d6704) I(d6705) I(d6706) I(d6707) I(d6708) I(d6709) I(d6710) I(d6711) I(d6712) I(d6713) I(d6714) I(d6715) I(d6716) I(d6717) I(d6718) I(d6719) I(d6720) I(d6721) I(d6722) I(d6723) I(d6724) I(d6725) I(d6726) I(d6727) I(d6728) I(d6729) I(d6730) I(d6731) I(d6732) I(d6733) I(d6734) I(d6735) I(d6736) I(d6737) I(d6738) I(d6739) I(d6740) I(d6741) I(d6742) I(d6743) I(d6744) I(d6745) I(d6746) I(d6747) I(d6748) I(d6749) I(d6750) I(d6751) I(d6752) I(d6753) I(d6754) I(d6755) I(d6756) I(d6757) I(d6758) I(d6759) I(d6760) I(d6761) I(d6762) I(d6763) I(d6764) I(d6765) I(d6766) I(d6767) I(d6768) I(d6769) I(d6770) I(d6771) I(d6772) I(d6773) I(d6774) I(d6775) I(d6776) I(d6777) I(d6778) I(d6779) I(d6780) I(d6781) I(d6782) I(d6783) I(d6784) I(d6785) I(d6786) I(d6787) I(d6788) I(d6789) I(d6790) I(d6791) I(d6792) I(d6793) I(d6794) I(d6795) I(d6796) I(d6797) I(d6798) I(d6799) I(d6800) I(d6801) I(d6802) I(d6803) I(d6804) I(d6805) I(d6806) I(d6807) I(d6808) I(d6809) I(d6810) I(d6811) I(d6812) I(d6813) I(d6814) I(d6815) I(d6816) I(d6817) I(d6818) I(d6819) I(d6820) I(d6821) I(d6822) I(d6823) I(d6824) I(d6825) I(d6826) I(d6827) I(d6828) I(d6829) I(d6830) I(d6831) I(d6832) I(d6833) I(d6834) I(d6835) I(d6836) I(d6837) I(d6838) I(d6839) I(d6840) I(d6841) I(d6842) I(d6843) I(d6844) I(d6845) I(d6846) I(d6847) I(d6848) I(d6849) I(d6850) I(d6851) I(d6852) I(d6853) I(d6854) I(d6855) I(d6856) I(d6857) I(d6858) I(d6859) I(d6860) I(d6861) I(d6862) I(d6863) I(d6864) I(d6865) I(d6866) I(d6867) I(d6868) I(d6869) I(d6870) I(d6871) I(d6872) I(d6873) I(d6874) I(d6875) I(d6876) I(d6877) I(d6878) I(d6879) I(d6880) I(d6881) I(d6882) I(d6883) I(d6884) I(d6885) I(d6886) I(d6887) I(d6888) I(d6889) I(d6890) I(d6891) I(d6892) I(d6893) I(d6894) I(d6895) I(d6896) I(d6897) I(d6898) I(d6899) I(d6900) I(d6901) I(d6902) I(d6903) I(d6904) I(d6905) I(d6906) I(d6907) I(d6908) I(d6909) I(d6910) I(d6911) I(d6912) I(d6913) I(d6914) I(d6915) I(d6916) I(d6917) I(d6918) I(d6919) I(d6920) I(d6921) I(d6922) I(d6923) I(d6924) I(d6925) I(d6926) I(d6927) I(d6928) I(d6929) I(d6930) I(d6931) I(d6932) I(d6933) I(d6934) I(d6935) I(d6936) I(d6937) I(d6938) I(d6939) I(d6940) I(d6941) I(d6942) I(d6943) I(d6944) I(d6945) I(d6946) I(d6947) I(d6948) I(d6949) I(d6950) I(d6951) I(d6952) I(d6953) I(d6954) I(d6955) I(d6956) I(d6957) I(d6958) I(d6959) I(d6960) I(d6961) I(d6962) I(d6963) I(d6964) I(d6965) I(d6966) I(d6967) I(d6968) I(d6969) I(d6970) I(d6971) I(d6972) I(d6973) I(d6974) I(d6975) I(d6976) I(d6977) I(d6978) I(d6979) I(d6980) I(d6981) I(d6982) I(d6983) I(d6984) I(d6985) I(d6986) I(d6987) I(d6988) I(d6989) I(d6990) I(d6991) I(d6992) I(d6993) I(d6994) I(d6995) I(d6996) I(d6997) I(d6998) I(d6999) I(d7000) I(d7001) I(d7002) I(d7003) I(d7004) I(d7005) I(d7006) I(d7007) I(d7008) I(d7009) I(d7010) I(d7011) I(d7012) I(d7013) I(d7014) I(d7015) I(d7016) I(d7017) I(d7018) I(d7019) I(d7020) I(d7021) I(d7022) I(d7023) I(d7024) I(d7025) I(d7026) I(d7027) I(d7028) I(d7029) I(d7030) I(d7031) I(d7032) I(d7033) I(d7034) I(d7035) I(d7036) I(d7037) I(d7038) I(d7039) I(d7040) I(d7041) I(d7042) I(d7043) I(d7044) I(d7045) I(d7046) I(d7047) I(d7048) I(d7049) I(d7050) I(d7051) I(d7052) I(d7053) I(d7054) I(d7055) I(d7056) I(d7057) I(d7058) I(d7059) I(d7060) I(d7061) I(d7062) I(d7063) I(d7064) I(d7065) I(d7066) I(d7067) I(d7068) I(d7069) I(d7070) I(d7071) I(d7072) I(d7073) I(d7074) I(d7075) I(d7076) I(d7077) I(d7078) I(d7079) I(d7080) I(d7081) I(d7082) I(d7083) I(d7084) I(d7085) I(d7086) I(d7087) I(d7088) I(d7089) I(d7090) I(d7091) I(d7092) I(d7093) I(d7094) I(d7095) I(d7096) I(d7097) I(d7098) I(d7099) I(d7100) I(d7101) I(d7102) I(d7103) I(d7104) I(d7105) I(d7106) I(d7107) I(d7108) I(d7109) I(d7110) I(d7111) I(d7112) I(d7113) I(d7114) I(d7115) I(d7116) I(d7117) I(d7118) I(d7119) I(d7120) I(d7121) I(d7122) I(d7123) I(d7124) I(d7125) I(d7126) I(d7127) I(d7128) I(d7129) I(d7130) I(d7131) I(d7132) I(d7133) I(d7134) I(d7135) I(d7136) I(d7137) I(d7138) I(d7139) I(d7140) I(d7141) I(d7142) I(d7143) I(d7144) I(d7145) I(d7146) I(d7147) I(d7148) I(d7149) I(d7150) I(d7151) I(d7152) I(d7153) I(d7154) I(d7155) I(d7156) I(d7157) I(d7158) I(d7159) I(d7160) I(d7161) I(d7162) I(d7163) I(d7164) I(d7165) I(d7166) I(d7167) I(d7168) I(d7169) I(d7170) I(d7171) I(d7172) I(d7173) I(d7174) I(d7175) I(d7176) I(d7177) I(d7178) I(d7179) I(d7180) I(d7181) I(d7182) I(d7183) I(d7184) I(d7185) I(d7186) I(d7187) I(d7188) I(d7189) I(d7190) I(d7191) I(d7192) I(d7193) I(d7194) I(d7195) I(d7196) I(d7197) I(d7198) I(d7199) I(d7200) I(d7201) I(d7202) I(d7203) I(d7204) I(d7205) I(d7206) I(d7207) I(d7208) I(d7209) I(d7210) I(d7211) I(d7212) I(d7213) I(d7214) I(d7215) I(d7216) I(d7217) I(d7218) I(d7219) I(d7220) I(d7221) I(d7222) I(d7223) I(d7224) I(d7225) I(d7226) I(d7227) I(d7228) I(d7229) I(d7230) I(d7231) I(d7232) I(d7233) I(d7234) I(d7235) I(d7236) I(d7237) I(d7238) I(d7239) I(d7240) I(d7241) I(d7242) I(d7243) I(d7244) I(d7245) I(d7246) I(d7247) I(d7248) I(d7249) I(d7250) I(d7251) I(d7252) I(d7253) I(d7254) I(d7255) I(d7256) I(d7257) I(d7258) I(d7259) I(d7260) I(d7261) I(d7262) I(d7263) I(d7264) I(d7265) I(d7266) I(d7267) I(d7268) I(d7269) I(d7270) I(d7271) I(d7272) I(d7273) I(d7274) I(d7275) I(d7276) I(d7277) I(d7278) I(d7279) I(d7280) I(d7281) I(d7282) I(d7283) I(d7284) I(d7285) I(d7286) I(d7287) I(d7288) I(d7289) I(d7290) I(d7291) I(d7292) I(d7293) I(d7294) I(d7295) I(d7296) I(d7297) I(d7298) I(d7299) I(d7300) I(d7301) I(d7302) I(d7303) I(d7304) I(d7305) I(d7306) I(d7307) I(d7308) I(d7309) I(d7310) I(d7311) I(d7312) I(d7313) I(d7314) I(d7315) I(d7316) I(d7317) I(d7318) I(d7319) I(d7320) I(d7321) I(d7322) I(d7323) I(d7324) I(d7325) I(d7326) I(d7327) I(d7328) I(d7329) I(d7330) I(d7331) I(d7332) I(d7333) I(d7334) I(d7335) I(d7336) I(d7337) I(d7338) I(d7339) I(d7340) I(d7341) I(d7342) I(d7343) I(d7344) I(d7345) I(d7346) I(d7347) I(d7348) I(d7349) I(d7350) I(d7351) I(d7352) I(d7353) I(d7354) I(d7355) I(d7356) I(d7357) I(d7358) I(d7359) I(d7360) I(d7361) I(d7362) I(d7363) I(d7364) I(d7365) I(d7366) I(d7367) I(d7368) I(d7369) I(d7370) I(d7371) I(d7372) I(d7373) I(d7374) I(d7375) I(d7376) I(d7377) I(d7378) I(d7379) I(d7380) I(d7381) I(d7382) I(d7383) I(d7384) I(d7385) I(d7386) I(d7387) I(d7388) I(d7389) I(d7390) I(d7391) I(d7392) I(d7393) I(d7394) I(d7395) I(d7396) I(d7397) I(d7398) I(d7399) I(d7400) I(d7401) I(d7402) I(d7403) I(d7404) I(d7405) I(d7406) I(d7407) I(d7408) I(d7409) I(d7410) I(d7411) I(d7412) I(d7413) I(d7414) I(d7415) I(d7416) I(d7417) I(d7418) I(d7419) I(d7420) I(d7421) I(d7422) I(d7423) I(d7424) I(d7425) I(d7426) I(d7427) I(d7428) I(d7429) I(d7430) I(d7431) I(d7432) I(d7433) I(d7434) I(d7435) I(d7436) I(d7437) I(d7438) I(d7439) I(d7440) I(d7441) I(d7442) I(d7443) I(d7444) I(d7445) I(d7446) I(d7447) I(d7448) I(d7449) I(d7450) I(d7451) I(d7452) I(d7453) I(d7454) I(d7455) I(d7456) I(d7457) I(d7458) I(d7459) I(d7460) I(d7461) I(d7462) I(d7463) I(d7464) I(d7465) I(d7466) I(d7467) I(d7468) I(d7469) I(d7470) I(d7471) I(d7472) I(d7473) I(d7474) I(d7475) I(d7476) I(d7477) I(d7478) I(d7479) I(d7480) I(d7481) I(d7482) I(d7483) I(d7484) I(d7485) I(d7486) I(d7487) I(d7488) I(d7489) I(d7490) I(d7491) I(d7492) I(d7493) I(d7494) I(d7495) I(d7496) I(d7497) I(d7498) I(d7499) I(d7500) I(d7501) I(d7502) I(d7503) I(d7504) I(d7505) I(d7506) I(d7507) I(d7508) I(d7509) I(d7510) I(d7511) I(d7512) I(d7513) I(d7514) I(d7515) I(d7516) I(d7517) I(d7518) I(d7519) I(d7520) I(d7521) I(d7522) I(d7523) I(d7524) I(d7525) I(d7526) I(d7527) I(d7528) I(d7529) I(d7530) I(d7531) I(d7532) I(d7533) I(d7534) I(d7535) I(d7536) I(d7537) I(d7538) I(d7539) I(d7540) I(d7541) I(d7542) I(d7543) I(d7544) I(d7545) I(d7546) I(d7547) I(d7548) I(d7549) I(d7550) I(d7551) I(d7552) I(d7553) I(d7554) I(d7555) I(d7556) I(d7557) I(d7558) I(d7559) I(d7560) I(d7561) I(d7562) I(d7563) I(d7564) I(d7565) I(d7566) I(d7567) I(d7568) I(d7569) I(d7570) I(d7571) I(d7572) I(d7573) I(d7574) I(d7575) I(d7576) I(d7577) I(d7578) I(d7579) I(d7580) I(d7581) I(d7582) I(d7583) I(d7584) I(d7585) I(d7586) I(d7587) I(d7588) I(d7589) I(d7590) I(d7591) I(d7592) I(d7593) I(d7594) I(d7595) I(d7596) I(d7597) I(d7598) I(d7599) I(d7600) I(d7601) I(d7602) I(d7603) I(d7604) I(d7605) I(d7606) I(d7607) I(d7608) I(d7609) I(d7610) I(d7611) I(d7612) I(d7613) I(d7614) I(d7615) I(d7616) I(d7617) I(d7618) I(d7619) I(d7620) I(d7621) I(d7622) I(d7623) I(d7624) I(d7625) I(d7626) I(d7627) I(d7628) I(d7629) I(d7630) I(d7631) I(d7632) I(d7633) I(d7634) I(d7635) I(d7636) I(d7637) I(d7638) I(d7639) I(d7640) I(d7641) I(d7642) I(d7643) I(d7644) I(d7645) I(d7646) I(d7647) I(d7648) I(d7649) I(d7650) I(d7651) I(d7652) I(d7653) I(d7654) I(d7655) I(d7656) I(d7657) I(d7658) I(d7659) I(d7660) I(d7661) I(d7662) I(d7663) I(d7664) I(d7665) I(d7666) I(d7667) I(d7668) I(d7669) I(d7670) I(d7671) I(d7672) I(d7673) I(d7674) I(d7675) I(d7676) I(d7677) I(d7678) I(d7679) I(d7680) I(d7681) I(d7682) I(d7683) I(d7684) I(d7685) I(d7686) I(d7687) I(d7688) I(d7689) I(d7690) I(d7691) I(d7692) I(d7693) I(d7694) I(d7695) I(d7696) I(d7697) I(d7698) I(d7699) I(d7700) I(d7701) I(d7702) I(d7703) I(d7704) I(d7705) I(d7706) I(d7707) I(d7708) I(d7709) I(d7710) I(d7711) I(d7712) I(d7713) I(d7714) I(d7715) I(d7716) I(d7717) I(d7718) I(d7719) I(d7720) I(d7721) I(d7722) I(d7723) I(d7724) I(d7725) I(d7726) I(d7727) I(d7728) I(d7729) I(d7730) I(d7731) I(d7732) I(d7733) I(d7734) I(d7735) I(d7736) I(d7737) I(d7738) I(d7739) I(d7740) I(d7741) I(d7742) I(d7743) I(d7744) I(d7745) I(d7746) I(d7747) I(d7748) I(d7749) I(d7750) I(d7751) I(d7752) I(d7753) I(d7754) I(d7755) I(d7756) I(d7757) I(d7758) I(d7759) I(d7760) I(d7761) I(d7762) I(d7763) I(d7764) I(d7765) I(d7766) I(d7767) I(d7768) I(d7769) I(d7770) I(d7771) I(d7772) I(d7773) I(d7774) I(d7775) I(d7776) I(d7777) I(d7778) I(d7779) I(d7780) I(d7781) I(d7782) I(d7783) I(d7784) I(d7785) I(d7786) I(d7787) I(d7788) I(d7789) I(d7790) I(d7791) I(d7792) I(d7793) I(d7794) I(d7795) I(d7796) I(d7797) I(d7798) I(d7799) I(d7800) I(d7801) I(d7802) I(d7803) I(d7804) I(d7805) I(d7806) I(d7807) I(d7808) I(d7809) I(d7810) I(d7811) I(d7812) I(d7813) I(d7814) I(d7815) I(d7816) I(d7817) I(d7818) I(d7819) I(d7820) I(d7821) I(d7822) I(d7823) I(d7824) I(d7825) I(d7826) I(d7827) I(d7828) I(d7829) I(d7830) I(d7831) I(d7832) I(d7833) I(d7834) I(d7835) I(d7836) I(d7837) I(d7838) I(d7839) I(d7840) I(d7841) I(d7842) I(d7843) I(d7844) I(d7845) I(d7846) I(d7847) I(d7848) I(d7849) I(d7850) I(d7851) I(d7852) I(d7853) I(d7854) I(d7855) I(d7856) I(d7857) I(d7858) I(d7859) I(d7860) I(d7861) I(d7862) I(d7863) I(d7864) I(d7865) I(d7866) I(d7867) I(d7868) I(d7869) I(d7870) I(d7871) I(d7872) I(d7873) I(d7874) I(d7875) I(d7876) I(d7877) I(d7878) I(d7879) I(d7880) I(d7881) I(d7882) I(d7883) I(d7884) I(d7885) I(d7886) I(d7887) I(d7888) I(d7889) I(d7890) I(d7891) I(d7892) I(d7893) I(d7894) I(d7895) I(d7896) I(d7897) I(d7898) I(d7899) I(d7900) I(d7901) I(d7902) I(d7903) I(d7904) I(d7905) I(d7906) I(d7907) I(d7908) I(d7909) I(d7910) I(d7911) I(d7912) I(d7913) I(d7914) I(d7915) I(d7916) I(d7917) I(d7918) I(d7919) I(d7920) I(d7921) I(d7922) I(d7923) I(d7924) I(d7925) I(d7926) I(d7927) I(d7928) I(d7929) I(d7930) I(d7931) I(d7932) I(d7933) I(d7934) I(d7935) I(d7936) I(d7937) I(d7938) I(d7939) I(d7940) I(d7941) I(d7942) I(d7943) I(d7944) I(d7945) I(d7946) I(d7947) I(d7948) I(d7949) I(d7950) I(d7951) I(d7952) I(d7953) I(d7954) I(d7955) I(d7956) I(d7957) I(d7958) I(d7959) I(d7960) I(d7961) I(d7962) I(d7963) I(d7964) I(d7965) I(d7966) I(d7967) I(d7968) I(d7969) I(d7970) I(d7971) I(d7972) I(d7973) I(d7974) I(d7975) I(d7976) I(d7977) I(d7978) I(d7979) I(d7980) I(d7981) I(d7982) I(d7983) I(d7984) I(d7985) I(d7986) I(d7987) I(d7988) I(d7989) I(d7990) I(d7991) I(d7992) I(d7993) I(d7994) I(d7995) I(d7996) I(d7997) I(d7998) I(d7999) I(d8000) I(d8001) I(d8002) I(d8003) I(d8004) I(d8005) I(d8006) I(d8007) I(d8008) I(d8009) I(d8010) I(d8011) I(d8012) I(d8013) I(d8014) I(d8015) I(d8016) I(d8017) I(d8018) I(d8019) I(d8020) I(d8021) I(d8022) I(d8023) I(d8024) I(d8025) I(d8026) I(d8027) I(d8028) I(d8029) I(d8030) I(d8031) I(d8032) I(d8033) I(d8034) I(d8035) I(d8036) I(d8037) I(d8038) I(d8039) I(d8040) I(d8041) I(d8042) I(d8043) I(d8044) I(d8045) I(d8046) I(d8047) I(d8048) I(d8049) I(d8050) I(d8051) I(d8052) I(d8053) I(d8054) I(d8055) I(d8056) I(d8057) I(d8058) I(d8059) I(d8060) I(d8061) I(d8062) I(d8063) I(d8064) I(d8065) I(d8066) I(d8067) I(d8068) I(d8069) I(d8070) I(d8071) I(d8072) I(d8073) I(d8074) I(d8075) I(d8076) I(d8077) I(d8078) I(d8079) I(d8080) I(d8081) I(d8082) I(d8083) I(d8084) I(d8085) I(d8086) I(d8087) I(d8088) I(d8089) I(d8090) I(d8091) I(d8092) I(d8093) I(d8094) I(d8095) I(d8096) I(d8097) I(d8098) I(d8099) I(d8100) I(d8101) I(d8102) I(d8103) I(d8104) I(d8105) I(d8106) I(d8107) I(d8108) I(d8109) I(d8110) I(d8111) I(d8112) I(d8113) I(d8114) I(d8115) I(d8116) I(d8117) I(d8118) I(d8119) I(d8120) I(d8121) I(d8122) I(d8123) I(d8124) I(d8125) I(d8126) I(d8127) I(d8128) I(d8129) I(d8130) I(d8131) I(d8132) I(d8133) I(d8134) I(d8135) I(d8136) I(d8137) I(d8138) I(d8139) I(d8140) I(d8141) I(d8142) I(d8143) I(d8144) I(d8145) I(d8146) I(d8147) I(d8148) I(d8149) I(d8150) I(d8151) I(d8152) I(d8153) I(d8154) I(d8155) I(d8156) I(d8157) I(d8158) I(d8159) I(d8160) I(d8161) I(d8162) I(d8163) I(d8164) I(d8165) I(d8166) I(d8167) I(d8168) I(d8169) I(d8170) I(d8171) I(d8172) I(d8173) I(d8174) I(d8175) I(d8176) I(d8177) I(d8178) I(d8179) I(d8180) I(d8181) I(d8182) I(d8183) I(d8184) I(d8185) I(d8186) I(d8187) I(d8188) I(d8189) I(d8190) I(d8191) I(d8192) I(d8193) I(d8194) I(d8195) I(d8196) I(d8197) I(d8198) I(d8199) I(d8200) I(d8201) I(d8202) I(d8203) I(d8204) I(d8205) I(d8206) I(d8207) I(d8208) I(d8209) I(d8210) I(d8211) I(d8212) I(d8213) I(d8214) I(d8215) I(d8216) I(d8217) I(d8218) I(d8219) I(d8220) I(d8221) I(d8222) I(d8223) I(d8224) I(d8225) I(d8226) I(d8227) I(d8228) I(d8229) I(d8230) I(d8231) I(d8232) I(d8233) I(d8234) I(d8235) I(d8236) I(d8237) I(d8238) I(d8239) I(d8240) I(d8241) I(d8242) I(d8243) I(d8244) I(d8245) I(d8246) I(d8247) I(d8248) I(d8249) I(d8250) I(d8251) I(d8252) I(d8253) I(d8254) I(d8255) I(d8256) I(d8257) I(d8258) I(d8259) I(d8260) I(d8261) I(d8262) I(d8263) I(d8264) I(d8265) I(d8266) I(d8267) I(d8268) I(d8269) I(d8270) I(d8271) I(d8272) I(d8273) I(d8274) I(d8275) I(d8276) I(d8277) I(d8278) I(d8279) I(d8280) I(d8281) I(d8282) I(d8283) I(d8284) I(d8285) I(d8286) I(d8287) I(d8288) I(d8289) I(d8290) I(d8291) I(d8292) I(d8293) I(d8294) I(d8295) I(d8296) I(d8297) I(d8298) I(d8299) I(d8300) I(d8301) I(d8302) I(d8303) I(d8304) I(d8305) I(d8306) I(d8307) I(d8308) I(d8309) I(d8310) I(d8311) I(d8312) I(d8313) I(d8314) I(d8315) I(d8316) I(d8317) I(d8318) I(d8319) I(d8320) I(d8321) I(d8322) I(d8323) I(d8324) I(d8325) I(d8326) I(d8327) I(d8328) I(d8329) I(d8330) I(d8331) I(d8332) I(d8333) I(d8334) I(d8335) I(d8336) I(d8337) I(d8338) I(d8339) I(d8340) I(d8341) I(d8342) I(d8343) I(d8344) I(d8345) I(d8346) I(d8347) I(d8348) I(d8349) I(d8350) I(d8351) I(d8352) I(d8353) I(d8354) I(d8355) I(d8356) I(d8357) I(d8358) I(d8359) I(d8360) I(d8361) I(d8362) I(d8363) I(d8364) I(d8365) I(d8366) I(d8367) I(d8368) I(d8369) I(d8370) I(d8371) I(d8372) I(d8373) I(d8374) I(d8375) I(d8376) I(d8377) I(d8378) I(d8379) I(d8380) I(d8381) I(d8382) I(d8383) I(d8384) I(d8385) I(d8386) I(d8387) I(d8388) I(d8389) I(d8390) I(d8391) I(d8392) I(d8393) I(d8394) I(d8395) I(d8396) I(d8397) I(d8398) I(d8399) I(d8400) I(d8401) I(d8402) I(d8403) I(d8404) I(d8405) I(d8406) I(d8407) I(d8408) I(d8409) I(d8410) I(d8411) I(d8412) I(d8413) I(d8414) I(d8415) I(d8416) I(d8417) I(d8418) I(d8419) I(d8420) I(d8421) I(d8422) I(d8423) I(d8424) I(d8425) I(d8426) I(d8427) I(d8428) I(d8429) I(d8430) I(d8431) I(d8432) I(d8433) I(d8434) I(d8435) I(d8436) I(d8437) I(d8438) I(d8439) I(d8440) I(d8441) I(d8442) I(d8443) I(d8444) I(d8445) I(d8446) I(d8447) I(d8448) I(d8449) I(d8450) I(d8451) I(d8452) I(d8453) I(d8454) I(d8455) I(d8456) I(d8457) I(d8458) I(d8459) I(d8460) I(d8461) I(d8462) I(d8463) I(d8464) I(d8465) I(d8466) I(d8467) I(d8468) I(d8469) I(d8470) I(d8471) I(d8472) I(d8473) I(d8474) I(d8475) I(d8476) I(d8477) I(d8478) I(d8479) I(d8480) I(d8481) I(d8482) I(d8483) I(d8484) I(d8485) I(d8486) I(d8487) I(d8488) I(d8489) I(d8490) I(d8491) I(d8492) I(d8493) I(d8494) I(d8495) I(d8496) I(d8497) I(d8498) I(d8499) I(d8500) I(d8501) I(d8502) I(d8503) I(d8504) I(d8505) I(d8506) I(d8507) I(d8508) I(d8509) I(d8510) I(d8511) I(d8512) I(d8513) I(d8514) I(d8515) I(d8516) I(d8517) I(d8518) I(d8519) I(d8520) I(d8521) I(d8522) I(d8523) I(d8524) I(d8525) I(d8526) I(d8527) I(d8528) I(d8529) I(d8530) I(d8531) I(d8532) I(d8533) I(d8534) I(d8535) I(d8536) I(d8537) I(d8538) I(d8539) I(d8540) I(d8541) I(d8542) I(d8543) I(d8544) I(d8545) I(d8546) I(d8547) I(d8548) I(d8549) I(d8550) I(d8551) I(d8552) I(d8553) I(d8554) I(d8555) I(d8556) I(d8557) I(d8558) I(d8559) I(d8560) I(d8561) I(d8562) I(d8563) I(d8564) I(d8565) I(d8566) I(d8567) I(d8568) I(d8569) I(d8570) I(d8571) I(d8572) I(d8573) I(d8574) I(d8575) I(d8576) I(d8577) I(d8578) I(d8579) I(d8580) I(d8581) I(d8582) I(d8583) I(d8584) I(d8585) I(d8586) I(d8587) I(d8588) I(d8589) I(d8590) I(d8591) I(d8592) I(d8593) I(d8594) I(d8595) I(d8596) I(d8597) I(d8598) I(d8599) I(d8600) I(d8601) I(d8602) I(d8603) I(d8604) I(d8605) I(d8606) I(d8607) I(d8608) I(d8609) I(d8610) I(d8611) I(d8612) I(d8613) I(d8614) I(d8615) I(d8616) I(d8617) I(d8618) I(d8619) I(d8620) I(d8621) I(d8622) I(d8623) I(d8624) I(d8625) I(d8626) I(d8627) I(d8628) I(d8629) I(d8630) I(d8631) I(d8632) I(d8633) I(d8634) I(d8635) I(d8636) I(d8637) I(d8638) I(d8639) I(d8640) I(d8641) I(d8642) I(d8643) I(d8644) I(d8645) I(d8646) I(d8647) I(d8648) I(d8649) I(d8650) I(d8651) I(d8652) I(d8653) I(d8654) I(d8655) I(d8656) I(d8657) I(d8658) I(d8659) I(d8660) I(d8661) I(d8662) I(d8663) I(d8664) I(d8665) I(d8666) I(d8667) I(d8668) I(d8669) I(d8670) I(d8671) I(d8672) I(d8673) I(d8674) I(d8675) I(d8676) I(d8677) I(d8678) I(d8679) I(d8680) I(d8681) I(d8682) I(d8683) I(d8684) I(d8685) I(d8686) I(d8687) I(d8688) I(d8689) I(d8690) I(d8691) I(d8692) I(d8693) I(d8694) I(d8695) I(d8696) I(d8697) I(d8698) I(d8699) I(d8700) I(d8701) I(d8702) I(d8703) I(d8704) I(d8705) I(d8706) I(d8707) I(d8708) I(d8709) I(d8710) I(d8711) I(d8712) I(d8713) I(d8714) I(d8715) I(d8716) I(d8717) I(d8718) I(d8719) I(d8720) I(d8721) I(d8722) I(d8723) I(d8724) I(d8725) I(d8726) I(d8727) I(d8728) I(d8729) I(d8730) I(d8731) I(d8732) I(d8733) I(d8734) I(d8735) I(d8736) I(d8737) I(d8738) I(d8739) I(d8740) I(d8741) I(d8742) I(d8743) I(d8744) I(d8745) I(d8746) I(d8747) I(d8748) I(d8749) I(d8750) I(d8751) I(d8752) I(d8753) I(d8754) I(d8755) I(d8756) I(d8757) I(d8758) I(d8759) I(d8760) I(d8761) I(d8762) I(d8763) I(d8764) I(d8765) I(d8766) I(d8767) I(d8768) I(d8769) I(d8770) I(d8771) I(d8772) I(d8773) I(d8774) I(d8775) I(d8776) I(d8777) I(d8778) I(d8779) I(d8780) I(d8781) I(d8782) I(d8783) I(d8784) I(d8785) I(d8786) I(d8787) I(d8788) I(d8789) I(d8790) I(d8791) I(d8792) I(d8793) I(d8794) I(d8795) I(d8796) I(d8797) I(d8798) I(d8799) I(d8800) I(d8801) I(d8802) I(d8803) I(d8804) I(d8805) I(d8806) I(d8807) I(d8808) I(d8809) I(d8810) I(d8811) I(d8812) I(d8813) I(d8814) I(d8815) I(d8816) I(d8817) I(d8818) I(d8819) I(d8820) I(d8821) I(d8822) I(d8823) I(d8824) I(d8825) I(d8826) I(d8827) I(d8828) I(d8829) I(d8830) I(d8831) I(d8832) I(d8833) I(d8834) I(d8835) I(d8836) I(d8837) I(d8838) I(d8839) I(d8840) I(d8841) I(d8842) I(d8843) I(d8844) I(d8845) I(d8846) I(d8847) I(d8848) I(d8849) I(d8850) I(d8851) I(d8852) I(d8853) I(d8854) I(d8855) I(d8856) I(d8857) I(d8858) I(d8859) I(d8860) I(d8861) I(d8862) I(d8863) I(d8864) I(d8865) I(d8866) I(d8867) I(d8868) I(d8869) I(d8870) I(d8871) I(d8872) I(d8873) I(d8874) I(d8875) I(d8876) I(d8877) I(d8878) I(d8879) I(d8880) I(d8881) I(d8882) I(d8883) I(d8884) I(d8885) I(d8886) I(d8887) I(d8888) I(d8889) I(d8890) I(d8891) I(d8892) I(d8893) I(d8894) I(d8895) I(d8896) I(d8897) I(d8898) I(d8899) I(d8900) I(d8901) I(d8902) I(d8903) I(d8904) I(d8905) I(d8906) I(d8907) I(d8908) I(d8909) I(d8910) I(d8911) I(d8912) I(d8913) I(d8914) I(d8915) I(d8916) I(d8917) I(d8918) I(d8919) I(d8920) I(d8921) I(d8922) I(d8923) I(d8924) I(d8925) I(d8926) I(d8927) I(d8928) I(d8929) I(d8930) I(d8931) I(d8932) I(d8933) I(d8934) I(d8935) I(d8936) I(d8937) I(d8938) I(d8939) I(d8940) I(d8941) I(d8942) I(d8943) I(d8944) I(d8945) I(d8946) I(d8947) I(d8948) I(d8949) I(d8950) I(d8951) I(d8952) I(d8953) I(d8954) I(d8955) I(d8956) I(d8957) I(d8958) I(d8959) I(d8960) I(d8961) I(d8962) I(d8963) I(d8964) I(d8965) I(d8966) I(d8967) I(d8968) I(d8969) I(d8970) I(d8971) I(d8972) I(d8973) I(d8974) I(d8975) I(d8976) I(d8977) I(d8978) I(d8979) I(d8980) I(d8981) I(d8982) I(d8983) I(d8984) I(d8985) I(d8986) I(d8987) I(d8988) I(d8989) I(d8990) I(d8991) I(d8992) I(d8993) I(d8994) I(d8995) I(d8996) I(d8997) I(d8998) I(d8999) I(d9000) I(d9001) I(d9002) I(d9003) I(d9004) I(d9005) I(d9006) I(d9007) I(d9008) I(d9009) I(d9010) I(d9011) I(d9012) I(d9013) I(d9014) I(d9015) I(d9016) I(d9017) I(d9018) I(d9019) I(d9020) I(d9021) I(d9022) I(d9023) I(d9024) I(d9025) I(d9026) I(d9027) I(d9028) I(d9029) I(d9030) I(d9031) I(d9032) I(d9033) I(d9034) I(d9035) I(d9036) I(d9037) I(d9038) I(d9039) I(d9040) I(d9041) I(d9042) I(d9043) I(d9044) I(d9045) I(d9046) I(d9047) I(d9048) I(d9049) I(d9050) I(d9051) I(d9052) I(d9053) I(d9054) I(d9055) I(d9056) I(d9057) I(d9058) I(d9059) I(d9060) I(d9061) I(d9062) I(d9063) I(d9064) I(d9065) I(d9066) I(d9067) I(d9068) I(d9069) I(d9070) I(d9071) I(d9072) I(d9073) I(d9074) I(d9075) I(d9076) I(d9077) I(d9078) I(d9079) I(d9080) I(d9081) I(d9082) I(d9083) I(d9084) I(d9085) I(d9086) I(d9087) I(d9088) I(d9089) I(d9090) I(d9091) I(d9092) I(d9093) I(d9094) I(d9095) I(d9096) I(d9097) I(d9098) I(d9099) I(d9100) I(d9101) I(d9102) I(d9103) I(d9104) I(d9105) I(d9106) I(d9107) I(d9108) I(d9109) I(d9110) I(d9111) I(d9112) I(d9113) I(d9114) I(d9115) I(d9116) I(d9117) I(d9118) I(d9119) I(d9120) I(d9121) I(d9122) I(d9123) I(d9124) I(d9125) I(d9126) I(d9127) I(d9128) I(d9129) I(d9130) I(d9131) I(d9132) I(d9133) I(d9134) I(d9135) I(d9136) I(d9137) I(d9138) I(d9139) I(d9140) I(d9141) I(d9142) I(d9143) I(d9144) I(d9145) I(d9146) I(d9147) I(d9148) I(d9149) I(d9150) I(d9151) I(d9152) I(d9153) I(d9154) I(d9155) I(d9156) I(d9157) I(d9158) I(d9159) I(d9160) I(d9161) I(d9162) I(d9163) I(d9164) I(d9165) I(d9166) I(d9167) I(d9168) I(d9169) I(d9170) I(d9171) I(d9172) I(d9173) I(d9174) I(d9175) I(d9176) I(d9177) I(d9178) I(d9179) I(d9180) I(d9181) I(d9182) I(d9183) I(d9184) I(d9185) I(d9186) I(d9187) I(d9188) I(d9189) I(d9190) I(d9191) I(d9192) I(d9193) I(d9194) I(d9195) I(d9196) I(d9197) I(d9198) I(d9199) I(d9200) I(d9201) I(d9202) I(d9203) I(d9204) I(d9205) I(d9206) I(d9207) I(d9208) I(d9209) I(d9210) I(d9211) I(d9212) I(d9213) I(d9214) I(d9215) I(d9216) I(d9217) I(d9218) I(d9219) I(d9220) I(d9221) I(d9222) I(d9223) I(d9224) I(d9225) I(d9226) I(d9227) I(d9228) I(d9229) I(d9230) I(d9231) I(d9232) I(d9233) I(d9234) I(d9235) I(d9236) I(d9237) I(d9238) I(d9239) I(d9240) I(d9241) I(d9242) I(d9243) I(d9244) I(d9245) I(d9246) I(d9247) I(d9248) I(d9249) I(d9250) I(d9251) I(d9252) I(d9253) I(d9254) I(d9255) I(d9256) I(d9257) I(d9258) I(d9259) I(d9260) I(d9261) I(d9262) I(d9263) I(d9264) I(d9265) I(d9266) I(d9267) I(d9268) I(d9269) I(d9270) I(d9271) I(d9272) I(d9273) I(d9274) I(d9275) I(d9276) I(d9277) I(d9278) I(d9279) I(d9280) I(d9281) I(d9282) I(d9283) I(d9284) I(d9285) I(d9286) I(d9287) I(d9288) I(d9289) I(d9290) I(d9291) I(d9292) I(d9293) I(d9294) I(d9295) I(d9296) I(d9297) I(d9298) I(d9299) I(d9300) I(d9301) I(d9302) I(d9303) I(d9304) I(d9305) I(d9306) I(d9307) I(d9308) I(d9309) I(d9310) I(d9311) I(d9312) I(d9313) I(d9314) I(d9315) I(d9316) I(d9317) I(d9318) I(d9319) I(d9320) I(d9321) I(d9322) I(d9323) I(d9324) I(d9325) I(d9326) I(d9327) I(d9328) I(d9329) I(d9330) I(d9331) I(d9332) I(d9333) I(d9334) I(d9335) I(d9336) I(d9337) I(d9338) I(d9339) I(d9340) I(d9341) I(d9342) I(d9343) I(d9344) I(d9345) I(d9346) I(d9347) I(d9348) I(d9349) I(d9350) I(d9351) I(d9352) I(d9353) I(d9354) I(d9355) I(d9356) I(d9357) I(d9358) I(d9359) I(d9360) I(d9361) I(d9362) I(d9363) I(d9364) I(d9365) I(d9366) I(d9367) I(d9368) I(d9369) I(d9370) I(d9371) I(d9372) I(d9373) I(d9374) I(d9375) I(d9376) I(d9377) I(d9378) I(d9379) I(d9380) I(d9381) I(d9382) I(d9383) I(d9384) I(d9385) I(d9386) I(d9387) I(d9388) I(d9389) I(d9390) I(d9391) I(d9392) I(d9393) I(d9394) I(d9395) I(d9396) I(d9397) I(d9398) I(d9399) I(d9400) I(d9401) I(d9402) I(d9403) I(d9404) I(d9405) I(d9406) I(d9407) I(d9408) I(d9409) I(d9410) I(d9411) I(d9412) I(d9413) I(d9414) I(d9415) I(d9416) I(d9417) I(d9418) I(d9419) I(d9420) I(d9421) I(d9422) I(d9423) I(d9424) I(d9425) I(d9426) I(d9427) I(d9428) I(d9429) I(d9430) I(d9431) I(d9432) I(d9433) I(d9434) I(d9435) I(d9436) I(d9437) I(d9438) I(d9439) I(d9440) I(d9441) I(d9442) I(d9443) I(d9444) I(d9445) I(d9446) I(d9447) I(d9448) I(d9449) I(d9450) I(d9451) I(d9452) I(d9453) I(d9454) I(d9455) I(d9456) I(d9457) I(d9458) I(d9459) I(d9460) I(d9461) I(d9462) I(d9463) I(d9464) I(d9465) I(d9466) I(d9467) I(d9468) I(d9469) I(d9470) I(d9471) I(d9472) I(d9473) I(d9474) I(d9475) I(d9476) I(d9477) I(d9478) I(d9479) I(d9480) I(d9481) I(d9482) I(d9483) I(d9484) I(d9485) I(d9486) I(d9487) I(d9488) I(d9489) I(d9490) I(d9491) I(d9492) I(d9493) I(d9494) I(d9495) I(d9496) I(d9497) I(d9498) I(d9499) I(d9500) I(d9501) I(d9502) I(d9503) I(d9504) I(d9505) I(d9506) I(d9507) I(d9508) I(d9509) I(d9510) I(d9511) I(d9512) I(d9513) I(d9514) I(d9515) I(d9516) I(d9517) I(d9518) I(d9519) I(d9520) I(d9521) I(d9522) I(d9523) I(d9524) I(d9525) I(d9526) I(d9527) I(d9528) I(d9529) I(d9530) I(d9531) I(d9532) I(d9533) I(d9534) I(d9535) I(d9536) I(d9537) I(d9538) I(d9539) I(d9540) I(d9541) I(d9542) I(d9543) I(d9544) I(d9545) I(d9546) I(d9547) I(d9548) I(d9549) I(d9550) I(d9551) I(d9552) I(d9553) I(d9554) I(d9555) I(d9556) I(d9557) I(d9558) I(d9559) I(d9560) I(d9561) I(d9562) I(d9563) I(d9564) I(d9565) I(d9566) I(d9567) I(d9568) I(d9569) I(d9570) I(d9571) I(d9572) I(d9573) I(d9574) I(d9575) I(d9576) I(d9577) I(d9578) I(d9579) I(d9580) I(d9581) I(d9582) I(d9583) I(d9584) I(d9585) I(d9586) I(d9587) I(d9588) I(d9589) I(d9590) I(d9591) I(d9592) I(d9593) I(d9594) I(d9595) I(d9596) I(d9597) I(d9598) I(d9599) I(d9600) I(d9601) I(d9602) I(d9603) I(d9604) I(d9605) I(d9606) I(d9607) I(d9608) I(d9609) I(d9610) I(d9611) I(d9612) I(d9613) I(d9614) I(d9615) I(d9616) I(d9617) I(d9618) I(d9619) I(d9620) I(d9621) I(d9622) I(d9623) I(d9624) I(d9625) I(d9626) I(d9627) I(d9628) I(d9629) I(d9630) I(d9631) I(d9632) I(d9633) I(d9634) I(d9635) I(d9636) I(d9637) I(d9638) I(d9639) I(d9640) I(d9641) I(d9642) I(d9643) I(d9644) I(d9645) I(d9646) I(d9647) I(d9648) I(d9649) I(d9650) I(d9651) I(d9652) I(d9653) I(d9654) I(d9655) I(d9656) I(d9657) I(d9658) I(d9659) I(d9660) I(d9661) I(d9662) I(d9663) I(d9664) I(d9665) I(d9666) I(d9667) I(d9668) I(d9669) I(d9670) I(d9671) I(d9672) I(d9673) I(d9674) I(d9675) I(d9676) I(d9677) I(d9678) I(d9679) I(d9680) I(d9681) I(d9682) I(d9683) I(d9684) I(d9685) I(d9686) I(d9687) I(d9688) I(d9689) I(d9690) I(d9691) I(d9692) I(d9693)


*** END 
.end 

