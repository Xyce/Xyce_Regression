*******************************************************************************
* This netlist is equivalent to Step 0 for the Off_TimeTest.cir netlist.
* It has VS1:VA=1
*
*******************************************************************************
*
* a few sources of different types
VS  1  0  SIN(0 1 1KHz 0 0)
VP  2  0  PULSE( 0 100 0.2ms 0.2ms 0.2ms 1ms 2ms )

R1  1  0  100
R2  2  0  100

* Use MEASFAIL to test the reset of the default calculation value
.OPTIONS MEASURE MEASFAIL=0

.TRAN 0  250ms
.PRINT TRAN FORMAT=NOINDEX V(1) V(2)

.measure tran off1KHz OFF_TIME V(1) OFF=.25
.measure tran offTop OFF_TIME V(2) OFF=25

* add TO-FROM modifiers
.measure tran sineHalfInterval off_time V(1) OFF=0.25 FROM=0 TO=0.5

* mix in TDs before and after FROM value.
.measure tran sineTDbetween off_time V(1) OFF=0.25 FROM=0 TO=0.25 TD=0.01
.measure tran sineTDbefore off_time V(1) OFF=0.25 FROM=0.01 TO=0.25 TD=0.005

* this test should return -1 
.measure tran returnNegOne off_time V(1) OFF=0.25 FROM=0.2e-3 TO=0.25e-3 TD=0.5e-3 default_val=-1

*this test should return 0
.measure tran returnZero off_time V(1) OFF=-2.0

.END

