* Test SNDR measure type for .MEASURE FFT for a .TRAN
* analysis.  Test covers voltage-difference operators,
* lead currents and expressions.
*
* See SON Bugs 1280 and 1327 for more details.
******************************************************

.TRAN 0 1
.OPTIONS FFT FFT_ACCURATE=1 FFTOUT=1

V1 1 0 1
R1 1 2 1
R2 2 0 1

V3 3 0 SIN(0 1 1)
R3 3 0 1

* This will be used to test with FREQ=2 on the .FFT line
V4 4 0 1
R4 4 0 1

* Test with multiple .FFT lines. The second .FFT V(1)
* line should get used by .MEASURE FFT.
.FFT V(1) NP=8 WINDOW=BART
.FFT V(1) NP=8 WINDOW=HANN
.FFT V(1,2) NP=8 WINDOW=HARRIS
.FFT V(3) NP=8 WINDOW=HARRIS
.FFT {I(V3)} NP=8 WINDOW=HANN
.FFT I(R3) NP=8 WINDOW=HARRIS
.FFT V(4) NP=16 WINDOW=HANN FREQ=2

.MEASURE FFT SNDRV1 SNDR V(1)

* Test with voltage difference syntax
.MEASURE FFT SNDRV12 SNDR V(1,2)

* Test expression and lead current
.MEASURE FFT SNDREXP SNDR {I(V3)}
.MEASURE FFT SNDRIR3 SNDR I(R3)

* Test that TRAN and FFT measure modes
* work in the same netlist
.MEASURE TRAN MAXV3 MAX V(3)

* Test with FFT-mode measure values in EQN measures
.MEASURE FFT EQN1 EQN SNDRV1
.MEASURE FFT EQN2 EQN SNDRV1
.MEASURE FFT PARAM1 PARAM {SNDREXP}

* Test that .MEASURE FFT line uses the FREQ value
* specified on the associated .FFT line.
.MEASURE FFT SNDRV4 SNDR V(4)

.PRINT TRAN V(1) V(2) V(3) I(V3) I(R3) V(4)
.END
