Test for OCT capability in DC sweeps. baseline
*
VT1 4 0 0V
R1  4 5 10
R2  5 0 5

.DC OCT VT1  0.125 66 3
.print DC V(4) V(5)

.END

