* This circuit tests a set of 1000 nested .funcs.

.param arg1=0.5
.param arg2=0.25
.param a=1
.param b=a

.func f0(x0) {x0+b}
.func f1(x1) { f0(x1)+b}
.func f2(x2) { f1(x2)+b}
.func f3(x3) { f2(x3)+b}
.func f4(x4) { f3(x4)+b}
.func f5(x5) { f4(x5)+b}
.func f6(x6) { f5(x6)+b}
.func f7(x7) { f6(x7)+b}
.func f8(x8) { f7(x8)+b}
.func f9(x9) { f8(x9)+b}
.func f10(x10) { f9(x10)+b}
.func f11(x11) { f10(x11)+b}
.func f12(x12) { f11(x12)+b}
.func f13(x13) { f12(x13)+b}
.func f14(x14) { f13(x14)+b}
.func f15(x15) { f14(x15)+b}
.func f16(x16) { f15(x16)+b}
.func f17(x17) { f16(x17)+b}
.func f18(x18) { f17(x18)+b}
.func f19(x19) { f18(x19)+b}
.func f20(x20) { f19(x20)+b}
.func f21(x21) { f20(x21)+b}
.func f22(x22) { f21(x22)+b}
.func f23(x23) { f22(x23)+b}
.func f24(x24) { f23(x24)+b}
.func f25(x25) { f24(x25)+b}
.func f26(x26) { f25(x26)+b}
.func f27(x27) { f26(x27)+b}
.func f28(x28) { f27(x28)+b}
.func f29(x29) { f28(x29)+b}
.func f30(x30) { f29(x30)+b}
.func f31(x31) { f30(x31)+b}
.func f32(x32) { f31(x32)+b}
.func f33(x33) { f32(x33)+b}
.func f34(x34) { f33(x34)+b}
.func f35(x35) { f34(x35)+b}
.func f36(x36) { f35(x36)+b}
.func f37(x37) { f36(x37)+b}
.func f38(x38) { f37(x38)+b}
.func f39(x39) { f38(x39)+b}
.func f40(x40) { f39(x40)+b}
.func f41(x41) { f40(x41)+b}
.func f42(x42) { f41(x42)+b}
.func f43(x43) { f42(x43)+b}
.func f44(x44) { f43(x44)+b}
.func f45(x45) { f44(x45)+b}
.func f46(x46) { f45(x46)+b}
.func f47(x47) { f46(x47)+b}
.func f48(x48) { f47(x48)+b}
.func f49(x49) { f48(x49)+b}
.func f50(x50) { f49(x50)+b}
.func f51(x51) { f50(x51)+b}
.func f52(x52) { f51(x52)+b}
.func f53(x53) { f52(x53)+b}
.func f54(x54) { f53(x54)+b}
.func f55(x55) { f54(x55)+b}
.func f56(x56) { f55(x56)+b}
.func f57(x57) { f56(x57)+b}
.func f58(x58) { f57(x58)+b}
.func f59(x59) { f58(x59)+b}
.func f60(x60) { f59(x60)+b}
.func f61(x61) { f60(x61)+b}
.func f62(x62) { f61(x62)+b}
.func f63(x63) { f62(x63)+b}
.func f64(x64) { f63(x64)+b}
.func f65(x65) { f64(x65)+b}
.func f66(x66) { f65(x66)+b}
.func f67(x67) { f66(x67)+b}
.func f68(x68) { f67(x68)+b}
.func f69(x69) { f68(x69)+b}
.func f70(x70) { f69(x70)+b}
.func f71(x71) { f70(x71)+b}
.func f72(x72) { f71(x72)+b}
.func f73(x73) { f72(x73)+b}
.func f74(x74) { f73(x74)+b}
.func f75(x75) { f74(x75)+b}
.func f76(x76) { f75(x76)+b}
.func f77(x77) { f76(x77)+b}
.func f78(x78) { f77(x78)+b}
.func f79(x79) { f78(x79)+b}
.func f80(x80) { f79(x80)+b}
.func f81(x81) { f80(x81)+b}
.func f82(x82) { f81(x82)+b}
.func f83(x83) { f82(x83)+b}
.func f84(x84) { f83(x84)+b}
.func f85(x85) { f84(x85)+b}
.func f86(x86) { f85(x86)+b}
.func f87(x87) { f86(x87)+b}
.func f88(x88) { f87(x88)+b}
.func f89(x89) { f88(x89)+b}
.func f90(x90) { f89(x90)+b}
.func f91(x91) { f90(x91)+b}
.func f92(x92) { f91(x92)+b}
.func f93(x93) { f92(x93)+b}
.func f94(x94) { f93(x94)+b}
.func f95(x95) { f94(x95)+b}
.func f96(x96) { f95(x96)+b}
.func f97(x97) { f96(x97)+b}
.func f98(x98) { f97(x98)+b}
.func f99(x99) { f98(x99)+b}
.func f100(x100) { f99(x100)+b}
.func f101(x101) { f100(x101)+b}
.func f102(x102) { f101(x102)+b}
.func f103(x103) { f102(x103)+b}
.func f104(x104) { f103(x104)+b}
.func f105(x105) { f104(x105)+b}
.func f106(x106) { f105(x106)+b}
.func f107(x107) { f106(x107)+b}
.func f108(x108) { f107(x108)+b}
.func f109(x109) { f108(x109)+b}
.func f110(x110) { f109(x110)+b}
.func f111(x111) { f110(x111)+b}
.func f112(x112) { f111(x112)+b}
.func f113(x113) { f112(x113)+b}
.func f114(x114) { f113(x114)+b}
.func f115(x115) { f114(x115)+b}
.func f116(x116) { f115(x116)+b}
.func f117(x117) { f116(x117)+b}
.func f118(x118) { f117(x118)+b}
.func f119(x119) { f118(x119)+b}
.func f120(x120) { f119(x120)+b}
.func f121(x121) { f120(x121)+b}
.func f122(x122) { f121(x122)+b}
.func f123(x123) { f122(x123)+b}
.func f124(x124) { f123(x124)+b}
.func f125(x125) { f124(x125)+b}
.func f126(x126) { f125(x126)+b}
.func f127(x127) { f126(x127)+b}
.func f128(x128) { f127(x128)+b}
.func f129(x129) { f128(x129)+b}
.func f130(x130) { f129(x130)+b}
.func f131(x131) { f130(x131)+b}
.func f132(x132) { f131(x132)+b}
.func f133(x133) { f132(x133)+b}
.func f134(x134) { f133(x134)+b}
.func f135(x135) { f134(x135)+b}
.func f136(x136) { f135(x136)+b}
.func f137(x137) { f136(x137)+b}
.func f138(x138) { f137(x138)+b}
.func f139(x139) { f138(x139)+b}
.func f140(x140) { f139(x140)+b}
.func f141(x141) { f140(x141)+b}
.func f142(x142) { f141(x142)+b}
.func f143(x143) { f142(x143)+b}
.func f144(x144) { f143(x144)+b}
.func f145(x145) { f144(x145)+b}
.func f146(x146) { f145(x146)+b}
.func f147(x147) { f146(x147)+b}
.func f148(x148) { f147(x148)+b}
.func f149(x149) { f148(x149)+b}
.func f150(x150) { f149(x150)+b}
.func f151(x151) { f150(x151)+b}
.func f152(x152) { f151(x152)+b}
.func f153(x153) { f152(x153)+b}
.func f154(x154) { f153(x154)+b}
.func f155(x155) { f154(x155)+b}
.func f156(x156) { f155(x156)+b}
.func f157(x157) { f156(x157)+b}
.func f158(x158) { f157(x158)+b}
.func f159(x159) { f158(x159)+b}
.func f160(x160) { f159(x160)+b}
.func f161(x161) { f160(x161)+b}
.func f162(x162) { f161(x162)+b}
.func f163(x163) { f162(x163)+b}
.func f164(x164) { f163(x164)+b}
.func f165(x165) { f164(x165)+b}
.func f166(x166) { f165(x166)+b}
.func f167(x167) { f166(x167)+b}
.func f168(x168) { f167(x168)+b}
.func f169(x169) { f168(x169)+b}
.func f170(x170) { f169(x170)+b}
.func f171(x171) { f170(x171)+b}
.func f172(x172) { f171(x172)+b}
.func f173(x173) { f172(x173)+b}
.func f174(x174) { f173(x174)+b}
.func f175(x175) { f174(x175)+b}
.func f176(x176) { f175(x176)+b}
.func f177(x177) { f176(x177)+b}
.func f178(x178) { f177(x178)+b}
.func f179(x179) { f178(x179)+b}
.func f180(x180) { f179(x180)+b}
.func f181(x181) { f180(x181)+b}
.func f182(x182) { f181(x182)+b}
.func f183(x183) { f182(x183)+b}
.func f184(x184) { f183(x184)+b}
.func f185(x185) { f184(x185)+b}
.func f186(x186) { f185(x186)+b}
.func f187(x187) { f186(x187)+b}
.func f188(x188) { f187(x188)+b}
.func f189(x189) { f188(x189)+b}
.func f190(x190) { f189(x190)+b}
.func f191(x191) { f190(x191)+b}
.func f192(x192) { f191(x192)+b}
.func f193(x193) { f192(x193)+b}
.func f194(x194) { f193(x194)+b}
.func f195(x195) { f194(x195)+b}
.func f196(x196) { f195(x196)+b}
.func f197(x197) { f196(x197)+b}
.func f198(x198) { f197(x198)+b}
.func f199(x199) { f198(x199)+b}
.func f200(x200) { f199(x200)+b}
.func f201(x201) { f200(x201)+b}
.func f202(x202) { f201(x202)+b}
.func f203(x203) { f202(x203)+b}
.func f204(x204) { f203(x204)+b}
.func f205(x205) { f204(x205)+b}
.func f206(x206) { f205(x206)+b}
.func f207(x207) { f206(x207)+b}
.func f208(x208) { f207(x208)+b}
.func f209(x209) { f208(x209)+b}
.func f210(x210) { f209(x210)+b}
.func f211(x211) { f210(x211)+b}
.func f212(x212) { f211(x212)+b}
.func f213(x213) { f212(x213)+b}
.func f214(x214) { f213(x214)+b}
.func f215(x215) { f214(x215)+b}
.func f216(x216) { f215(x216)+b}
.func f217(x217) { f216(x217)+b}
.func f218(x218) { f217(x218)+b}
.func f219(x219) { f218(x219)+b}
.func f220(x220) { f219(x220)+b}
.func f221(x221) { f220(x221)+b}
.func f222(x222) { f221(x222)+b}
.func f223(x223) { f222(x223)+b}
.func f224(x224) { f223(x224)+b}
.func f225(x225) { f224(x225)+b}
.func f226(x226) { f225(x226)+b}
.func f227(x227) { f226(x227)+b}
.func f228(x228) { f227(x228)+b}
.func f229(x229) { f228(x229)+b}
.func f230(x230) { f229(x230)+b}
.func f231(x231) { f230(x231)+b}
.func f232(x232) { f231(x232)+b}
.func f233(x233) { f232(x233)+b}
.func f234(x234) { f233(x234)+b}
.func f235(x235) { f234(x235)+b}
.func f236(x236) { f235(x236)+b}
.func f237(x237) { f236(x237)+b}
.func f238(x238) { f237(x238)+b}
.func f239(x239) { f238(x239)+b}
.func f240(x240) { f239(x240)+b}
.func f241(x241) { f240(x241)+b}
.func f242(x242) { f241(x242)+b}
.func f243(x243) { f242(x243)+b}
.func f244(x244) { f243(x244)+b}
.func f245(x245) { f244(x245)+b}
.func f246(x246) { f245(x246)+b}
.func f247(x247) { f246(x247)+b}
.func f248(x248) { f247(x248)+b}
.func f249(x249) { f248(x249)+b}
.func f250(x250) { f249(x250)+b}
.func f251(x251) { f250(x251)+b}
.func f252(x252) { f251(x252)+b}
.func f253(x253) { f252(x253)+b}
.func f254(x254) { f253(x254)+b}
.func f255(x255) { f254(x255)+b}
.func f256(x256) { f255(x256)+b}
.func f257(x257) { f256(x257)+b}
.func f258(x258) { f257(x258)+b}
.func f259(x259) { f258(x259)+b}
.func f260(x260) { f259(x260)+b}
.func f261(x261) { f260(x261)+b}
.func f262(x262) { f261(x262)+b}
.func f263(x263) { f262(x263)+b}
.func f264(x264) { f263(x264)+b}
.func f265(x265) { f264(x265)+b}
.func f266(x266) { f265(x266)+b}
.func f267(x267) { f266(x267)+b}
.func f268(x268) { f267(x268)+b}
.func f269(x269) { f268(x269)+b}
.func f270(x270) { f269(x270)+b}
.func f271(x271) { f270(x271)+b}
.func f272(x272) { f271(x272)+b}
.func f273(x273) { f272(x273)+b}
.func f274(x274) { f273(x274)+b}
.func f275(x275) { f274(x275)+b}
.func f276(x276) { f275(x276)+b}
.func f277(x277) { f276(x277)+b}
.func f278(x278) { f277(x278)+b}
.func f279(x279) { f278(x279)+b}
.func f280(x280) { f279(x280)+b}
.func f281(x281) { f280(x281)+b}
.func f282(x282) { f281(x282)+b}
.func f283(x283) { f282(x283)+b}
.func f284(x284) { f283(x284)+b}
.func f285(x285) { f284(x285)+b}
.func f286(x286) { f285(x286)+b}
.func f287(x287) { f286(x287)+b}
.func f288(x288) { f287(x288)+b}
.func f289(x289) { f288(x289)+b}
.func f290(x290) { f289(x290)+b}
.func f291(x291) { f290(x291)+b}
.func f292(x292) { f291(x292)+b}
.func f293(x293) { f292(x293)+b}
.func f294(x294) { f293(x294)+b}
.func f295(x295) { f294(x295)+b}
.func f296(x296) { f295(x296)+b}
.func f297(x297) { f296(x297)+b}
.func f298(x298) { f297(x298)+b}
.func f299(x299) { f298(x299)+b}
.func f300(x300) { f299(x300)+b}
.func f301(x301) { f300(x301)+b}
.func f302(x302) { f301(x302)+b}
.func f303(x303) { f302(x303)+b}
.func f304(x304) { f303(x304)+b}
.func f305(x305) { f304(x305)+b}
.func f306(x306) { f305(x306)+b}
.func f307(x307) { f306(x307)+b}
.func f308(x308) { f307(x308)+b}
.func f309(x309) { f308(x309)+b}
.func f310(x310) { f309(x310)+b}
.func f311(x311) { f310(x311)+b}
.func f312(x312) { f311(x312)+b}
.func f313(x313) { f312(x313)+b}
.func f314(x314) { f313(x314)+b}
.func f315(x315) { f314(x315)+b}
.func f316(x316) { f315(x316)+b}
.func f317(x317) { f316(x317)+b}
.func f318(x318) { f317(x318)+b}
.func f319(x319) { f318(x319)+b}
.func f320(x320) { f319(x320)+b}
.func f321(x321) { f320(x321)+b}
.func f322(x322) { f321(x322)+b}
.func f323(x323) { f322(x323)+b}
.func f324(x324) { f323(x324)+b}
.func f325(x325) { f324(x325)+b}
.func f326(x326) { f325(x326)+b}
.func f327(x327) { f326(x327)+b}
.func f328(x328) { f327(x328)+b}
.func f329(x329) { f328(x329)+b}
.func f330(x330) { f329(x330)+b}
.func f331(x331) { f330(x331)+b}
.func f332(x332) { f331(x332)+b}
.func f333(x333) { f332(x333)+b}
.func f334(x334) { f333(x334)+b}
.func f335(x335) { f334(x335)+b}
.func f336(x336) { f335(x336)+b}
.func f337(x337) { f336(x337)+b}
.func f338(x338) { f337(x338)+b}
.func f339(x339) { f338(x339)+b}
.func f340(x340) { f339(x340)+b}
.func f341(x341) { f340(x341)+b}
.func f342(x342) { f341(x342)+b}
.func f343(x343) { f342(x343)+b}
.func f344(x344) { f343(x344)+b}
.func f345(x345) { f344(x345)+b}
.func f346(x346) { f345(x346)+b}
.func f347(x347) { f346(x347)+b}
.func f348(x348) { f347(x348)+b}
.func f349(x349) { f348(x349)+b}
.func f350(x350) { f349(x350)+b}
.func f351(x351) { f350(x351)+b}
.func f352(x352) { f351(x352)+b}
.func f353(x353) { f352(x353)+b}
.func f354(x354) { f353(x354)+b}
.func f355(x355) { f354(x355)+b}
.func f356(x356) { f355(x356)+b}
.func f357(x357) { f356(x357)+b}
.func f358(x358) { f357(x358)+b}
.func f359(x359) { f358(x359)+b}
.func f360(x360) { f359(x360)+b}
.func f361(x361) { f360(x361)+b}
.func f362(x362) { f361(x362)+b}
.func f363(x363) { f362(x363)+b}
.func f364(x364) { f363(x364)+b}
.func f365(x365) { f364(x365)+b}
.func f366(x366) { f365(x366)+b}
.func f367(x367) { f366(x367)+b}
.func f368(x368) { f367(x368)+b}
.func f369(x369) { f368(x369)+b}
.func f370(x370) { f369(x370)+b}
.func f371(x371) { f370(x371)+b}
.func f372(x372) { f371(x372)+b}
.func f373(x373) { f372(x373)+b}
.func f374(x374) { f373(x374)+b}
.func f375(x375) { f374(x375)+b}
.func f376(x376) { f375(x376)+b}
.func f377(x377) { f376(x377)+b}
.func f378(x378) { f377(x378)+b}
.func f379(x379) { f378(x379)+b}
.func f380(x380) { f379(x380)+b}
.func f381(x381) { f380(x381)+b}
.func f382(x382) { f381(x382)+b}
.func f383(x383) { f382(x383)+b}
.func f384(x384) { f383(x384)+b}
.func f385(x385) { f384(x385)+b}
.func f386(x386) { f385(x386)+b}
.func f387(x387) { f386(x387)+b}
.func f388(x388) { f387(x388)+b}
.func f389(x389) { f388(x389)+b}
.func f390(x390) { f389(x390)+b}
.func f391(x391) { f390(x391)+b}
.func f392(x392) { f391(x392)+b}
.func f393(x393) { f392(x393)+b}
.func f394(x394) { f393(x394)+b}
.func f395(x395) { f394(x395)+b}
.func f396(x396) { f395(x396)+b}
.func f397(x397) { f396(x397)+b}
.func f398(x398) { f397(x398)+b}
.func f399(x399) { f398(x399)+b}
.func f400(x400) { f399(x400)+b}
.func f401(x401) { f400(x401)+b}
.func f402(x402) { f401(x402)+b}
.func f403(x403) { f402(x403)+b}
.func f404(x404) { f403(x404)+b}
.func f405(x405) { f404(x405)+b}
.func f406(x406) { f405(x406)+b}
.func f407(x407) { f406(x407)+b}
.func f408(x408) { f407(x408)+b}
.func f409(x409) { f408(x409)+b}
.func f410(x410) { f409(x410)+b}
.func f411(x411) { f410(x411)+b}
.func f412(x412) { f411(x412)+b}
.func f413(x413) { f412(x413)+b}
.func f414(x414) { f413(x414)+b}
.func f415(x415) { f414(x415)+b}
.func f416(x416) { f415(x416)+b}
.func f417(x417) { f416(x417)+b}
.func f418(x418) { f417(x418)+b}
.func f419(x419) { f418(x419)+b}
.func f420(x420) { f419(x420)+b}
.func f421(x421) { f420(x421)+b}
.func f422(x422) { f421(x422)+b}
.func f423(x423) { f422(x423)+b}
.func f424(x424) { f423(x424)+b}
.func f425(x425) { f424(x425)+b}
.func f426(x426) { f425(x426)+b}
.func f427(x427) { f426(x427)+b}
.func f428(x428) { f427(x428)+b}
.func f429(x429) { f428(x429)+b}
.func f430(x430) { f429(x430)+b}
.func f431(x431) { f430(x431)+b}
.func f432(x432) { f431(x432)+b}
.func f433(x433) { f432(x433)+b}
.func f434(x434) { f433(x434)+b}
.func f435(x435) { f434(x435)+b}
.func f436(x436) { f435(x436)+b}
.func f437(x437) { f436(x437)+b}
.func f438(x438) { f437(x438)+b}
.func f439(x439) { f438(x439)+b}
.func f440(x440) { f439(x440)+b}
.func f441(x441) { f440(x441)+b}
.func f442(x442) { f441(x442)+b}
.func f443(x443) { f442(x443)+b}
.func f444(x444) { f443(x444)+b}
.func f445(x445) { f444(x445)+b}
.func f446(x446) { f445(x446)+b}
.func f447(x447) { f446(x447)+b}
.func f448(x448) { f447(x448)+b}
.func f449(x449) { f448(x449)+b}
.func f450(x450) { f449(x450)+b}
.func f451(x451) { f450(x451)+b}
.func f452(x452) { f451(x452)+b}
.func f453(x453) { f452(x453)+b}
.func f454(x454) { f453(x454)+b}
.func f455(x455) { f454(x455)+b}
.func f456(x456) { f455(x456)+b}
.func f457(x457) { f456(x457)+b}
.func f458(x458) { f457(x458)+b}
.func f459(x459) { f458(x459)+b}
.func f460(x460) { f459(x460)+b}
.func f461(x461) { f460(x461)+b}
.func f462(x462) { f461(x462)+b}
.func f463(x463) { f462(x463)+b}
.func f464(x464) { f463(x464)+b}
.func f465(x465) { f464(x465)+b}
.func f466(x466) { f465(x466)+b}
.func f467(x467) { f466(x467)+b}
.func f468(x468) { f467(x468)+b}
.func f469(x469) { f468(x469)+b}
.func f470(x470) { f469(x470)+b}
.func f471(x471) { f470(x471)+b}
.func f472(x472) { f471(x472)+b}
.func f473(x473) { f472(x473)+b}
.func f474(x474) { f473(x474)+b}
.func f475(x475) { f474(x475)+b}
.func f476(x476) { f475(x476)+b}
.func f477(x477) { f476(x477)+b}
.func f478(x478) { f477(x478)+b}
.func f479(x479) { f478(x479)+b}
.func f480(x480) { f479(x480)+b}
.func f481(x481) { f480(x481)+b}
.func f482(x482) { f481(x482)+b}
.func f483(x483) { f482(x483)+b}
.func f484(x484) { f483(x484)+b}
.func f485(x485) { f484(x485)+b}
.func f486(x486) { f485(x486)+b}
.func f487(x487) { f486(x487)+b}
.func f488(x488) { f487(x488)+b}
.func f489(x489) { f488(x489)+b}
.func f490(x490) { f489(x490)+b}
.func f491(x491) { f490(x491)+b}
.func f492(x492) { f491(x492)+b}
.func f493(x493) { f492(x493)+b}
.func f494(x494) { f493(x494)+b}
.func f495(x495) { f494(x495)+b}
.func f496(x496) { f495(x496)+b}
.func f497(x497) { f496(x497)+b}
.func f498(x498) { f497(x498)+b}
.func f499(x499) { f498(x499)+b}
.func f500(x500) { f499(x500)+b}
.func f501(x501) { f500(x501)+b}
.func f502(x502) { f501(x502)+b}
.func f503(x503) { f502(x503)+b}
.func f504(x504) { f503(x504)+b}
.func f505(x505) { f504(x505)+b}
.func f506(x506) { f505(x506)+b}
.func f507(x507) { f506(x507)+b}
.func f508(x508) { f507(x508)+b}
.func f509(x509) { f508(x509)+b}
.func f510(x510) { f509(x510)+b}
.func f511(x511) { f510(x511)+b}
.func f512(x512) { f511(x512)+b}
.func f513(x513) { f512(x513)+b}
.func f514(x514) { f513(x514)+b}
.func f515(x515) { f514(x515)+b}
.func f516(x516) { f515(x516)+b}
.func f517(x517) { f516(x517)+b}
.func f518(x518) { f517(x518)+b}
.func f519(x519) { f518(x519)+b}
.func f520(x520) { f519(x520)+b}
.func f521(x521) { f520(x521)+b}
.func f522(x522) { f521(x522)+b}
.func f523(x523) { f522(x523)+b}
.func f524(x524) { f523(x524)+b}
.func f525(x525) { f524(x525)+b}
.func f526(x526) { f525(x526)+b}
.func f527(x527) { f526(x527)+b}
.func f528(x528) { f527(x528)+b}
.func f529(x529) { f528(x529)+b}
.func f530(x530) { f529(x530)+b}
.func f531(x531) { f530(x531)+b}
.func f532(x532) { f531(x532)+b}
.func f533(x533) { f532(x533)+b}
.func f534(x534) { f533(x534)+b}
.func f535(x535) { f534(x535)+b}
.func f536(x536) { f535(x536)+b}
.func f537(x537) { f536(x537)+b}
.func f538(x538) { f537(x538)+b}
.func f539(x539) { f538(x539)+b}
.func f540(x540) { f539(x540)+b}
.func f541(x541) { f540(x541)+b}
.func f542(x542) { f541(x542)+b}
.func f543(x543) { f542(x543)+b}
.func f544(x544) { f543(x544)+b}
.func f545(x545) { f544(x545)+b}
.func f546(x546) { f545(x546)+b}
.func f547(x547) { f546(x547)+b}
.func f548(x548) { f547(x548)+b}
.func f549(x549) { f548(x549)+b}
.func f550(x550) { f549(x550)+b}
.func f551(x551) { f550(x551)+b}
.func f552(x552) { f551(x552)+b}
.func f553(x553) { f552(x553)+b}
.func f554(x554) { f553(x554)+b}
.func f555(x555) { f554(x555)+b}
.func f556(x556) { f555(x556)+b}
.func f557(x557) { f556(x557)+b}
.func f558(x558) { f557(x558)+b}
.func f559(x559) { f558(x559)+b}
.func f560(x560) { f559(x560)+b}
.func f561(x561) { f560(x561)+b}
.func f562(x562) { f561(x562)+b}
.func f563(x563) { f562(x563)+b}
.func f564(x564) { f563(x564)+b}
.func f565(x565) { f564(x565)+b}
.func f566(x566) { f565(x566)+b}
.func f567(x567) { f566(x567)+b}
.func f568(x568) { f567(x568)+b}
.func f569(x569) { f568(x569)+b}
.func f570(x570) { f569(x570)+b}
.func f571(x571) { f570(x571)+b}
.func f572(x572) { f571(x572)+b}
.func f573(x573) { f572(x573)+b}
.func f574(x574) { f573(x574)+b}
.func f575(x575) { f574(x575)+b}
.func f576(x576) { f575(x576)+b}
.func f577(x577) { f576(x577)+b}
.func f578(x578) { f577(x578)+b}
.func f579(x579) { f578(x579)+b}
.func f580(x580) { f579(x580)+b}
.func f581(x581) { f580(x581)+b}
.func f582(x582) { f581(x582)+b}
.func f583(x583) { f582(x583)+b}
.func f584(x584) { f583(x584)+b}
.func f585(x585) { f584(x585)+b}
.func f586(x586) { f585(x586)+b}
.func f587(x587) { f586(x587)+b}
.func f588(x588) { f587(x588)+b}
.func f589(x589) { f588(x589)+b}
.func f590(x590) { f589(x590)+b}
.func f591(x591) { f590(x591)+b}
.func f592(x592) { f591(x592)+b}
.func f593(x593) { f592(x593)+b}
.func f594(x594) { f593(x594)+b}
.func f595(x595) { f594(x595)+b}
.func f596(x596) { f595(x596)+b}
.func f597(x597) { f596(x597)+b}
.func f598(x598) { f597(x598)+b}
.func f599(x599) { f598(x599)+b}
.func f600(x600) { f599(x600)+b}
.func f601(x601) { f600(x601)+b}
.func f602(x602) { f601(x602)+b}
.func f603(x603) { f602(x603)+b}
.func f604(x604) { f603(x604)+b}
.func f605(x605) { f604(x605)+b}
.func f606(x606) { f605(x606)+b}
.func f607(x607) { f606(x607)+b}
.func f608(x608) { f607(x608)+b}
.func f609(x609) { f608(x609)+b}
.func f610(x610) { f609(x610)+b}
.func f611(x611) { f610(x611)+b}
.func f612(x612) { f611(x612)+b}
.func f613(x613) { f612(x613)+b}
.func f614(x614) { f613(x614)+b}
.func f615(x615) { f614(x615)+b}
.func f616(x616) { f615(x616)+b}
.func f617(x617) { f616(x617)+b}
.func f618(x618) { f617(x618)+b}
.func f619(x619) { f618(x619)+b}
.func f620(x620) { f619(x620)+b}
.func f621(x621) { f620(x621)+b}
.func f622(x622) { f621(x622)+b}
.func f623(x623) { f622(x623)+b}
.func f624(x624) { f623(x624)+b}
.func f625(x625) { f624(x625)+b}
.func f626(x626) { f625(x626)+b}
.func f627(x627) { f626(x627)+b}
.func f628(x628) { f627(x628)+b}
.func f629(x629) { f628(x629)+b}
.func f630(x630) { f629(x630)+b}
.func f631(x631) { f630(x631)+b}
.func f632(x632) { f631(x632)+b}
.func f633(x633) { f632(x633)+b}
.func f634(x634) { f633(x634)+b}
.func f635(x635) { f634(x635)+b}
.func f636(x636) { f635(x636)+b}
.func f637(x637) { f636(x637)+b}
.func f638(x638) { f637(x638)+b}
.func f639(x639) { f638(x639)+b}
.func f640(x640) { f639(x640)+b}
.func f641(x641) { f640(x641)+b}
.func f642(x642) { f641(x642)+b}
.func f643(x643) { f642(x643)+b}
.func f644(x644) { f643(x644)+b}
.func f645(x645) { f644(x645)+b}
.func f646(x646) { f645(x646)+b}
.func f647(x647) { f646(x647)+b}
.func f648(x648) { f647(x648)+b}
.func f649(x649) { f648(x649)+b}
.func f650(x650) { f649(x650)+b}
.func f651(x651) { f650(x651)+b}
.func f652(x652) { f651(x652)+b}
.func f653(x653) { f652(x653)+b}
.func f654(x654) { f653(x654)+b}
.func f655(x655) { f654(x655)+b}
.func f656(x656) { f655(x656)+b}
.func f657(x657) { f656(x657)+b}
.func f658(x658) { f657(x658)+b}
.func f659(x659) { f658(x659)+b}
.func f660(x660) { f659(x660)+b}
.func f661(x661) { f660(x661)+b}
.func f662(x662) { f661(x662)+b}
.func f663(x663) { f662(x663)+b}
.func f664(x664) { f663(x664)+b}
.func f665(x665) { f664(x665)+b}
.func f666(x666) { f665(x666)+b}
.func f667(x667) { f666(x667)+b}
.func f668(x668) { f667(x668)+b}
.func f669(x669) { f668(x669)+b}
.func f670(x670) { f669(x670)+b}
.func f671(x671) { f670(x671)+b}
.func f672(x672) { f671(x672)+b}
.func f673(x673) { f672(x673)+b}
.func f674(x674) { f673(x674)+b}
.func f675(x675) { f674(x675)+b}
.func f676(x676) { f675(x676)+b}
.func f677(x677) { f676(x677)+b}
.func f678(x678) { f677(x678)+b}
.func f679(x679) { f678(x679)+b}
.func f680(x680) { f679(x680)+b}
.func f681(x681) { f680(x681)+b}
.func f682(x682) { f681(x682)+b}
.func f683(x683) { f682(x683)+b}
.func f684(x684) { f683(x684)+b}
.func f685(x685) { f684(x685)+b}
.func f686(x686) { f685(x686)+b}
.func f687(x687) { f686(x687)+b}
.func f688(x688) { f687(x688)+b}
.func f689(x689) { f688(x689)+b}
.func f690(x690) { f689(x690)+b}
.func f691(x691) { f690(x691)+b}
.func f692(x692) { f691(x692)+b}
.func f693(x693) { f692(x693)+b}
.func f694(x694) { f693(x694)+b}
.func f695(x695) { f694(x695)+b}
.func f696(x696) { f695(x696)+b}
.func f697(x697) { f696(x697)+b}
.func f698(x698) { f697(x698)+b}
.func f699(x699) { f698(x699)+b}
.func f700(x700) { f699(x700)+b}
.func f701(x701) { f700(x701)+b}
.func f702(x702) { f701(x702)+b}
.func f703(x703) { f702(x703)+b}
.func f704(x704) { f703(x704)+b}
.func f705(x705) { f704(x705)+b}
.func f706(x706) { f705(x706)+b}
.func f707(x707) { f706(x707)+b}
.func f708(x708) { f707(x708)+b}
.func f709(x709) { f708(x709)+b}
.func f710(x710) { f709(x710)+b}
.func f711(x711) { f710(x711)+b}
.func f712(x712) { f711(x712)+b}
.func f713(x713) { f712(x713)+b}
.func f714(x714) { f713(x714)+b}
.func f715(x715) { f714(x715)+b}
.func f716(x716) { f715(x716)+b}
.func f717(x717) { f716(x717)+b}
.func f718(x718) { f717(x718)+b}
.func f719(x719) { f718(x719)+b}
.func f720(x720) { f719(x720)+b}
.func f721(x721) { f720(x721)+b}
.func f722(x722) { f721(x722)+b}
.func f723(x723) { f722(x723)+b}
.func f724(x724) { f723(x724)+b}
.func f725(x725) { f724(x725)+b}
.func f726(x726) { f725(x726)+b}
.func f727(x727) { f726(x727)+b}
.func f728(x728) { f727(x728)+b}
.func f729(x729) { f728(x729)+b}
.func f730(x730) { f729(x730)+b}
.func f731(x731) { f730(x731)+b}
.func f732(x732) { f731(x732)+b}
.func f733(x733) { f732(x733)+b}
.func f734(x734) { f733(x734)+b}
.func f735(x735) { f734(x735)+b}
.func f736(x736) { f735(x736)+b}
.func f737(x737) { f736(x737)+b}
.func f738(x738) { f737(x738)+b}
.func f739(x739) { f738(x739)+b}
.func f740(x740) { f739(x740)+b}
.func f741(x741) { f740(x741)+b}
.func f742(x742) { f741(x742)+b}
.func f743(x743) { f742(x743)+b}
.func f744(x744) { f743(x744)+b}
.func f745(x745) { f744(x745)+b}
.func f746(x746) { f745(x746)+b}
.func f747(x747) { f746(x747)+b}
.func f748(x748) { f747(x748)+b}
.func f749(x749) { f748(x749)+b}
.func f750(x750) { f749(x750)+b}
.func f751(x751) { f750(x751)+b}
.func f752(x752) { f751(x752)+b}
.func f753(x753) { f752(x753)+b}
.func f754(x754) { f753(x754)+b}
.func f755(x755) { f754(x755)+b}
.func f756(x756) { f755(x756)+b}
.func f757(x757) { f756(x757)+b}
.func f758(x758) { f757(x758)+b}
.func f759(x759) { f758(x759)+b}
.func f760(x760) { f759(x760)+b}
.func f761(x761) { f760(x761)+b}
.func f762(x762) { f761(x762)+b}
.func f763(x763) { f762(x763)+b}
.func f764(x764) { f763(x764)+b}
.func f765(x765) { f764(x765)+b}
.func f766(x766) { f765(x766)+b}
.func f767(x767) { f766(x767)+b}
.func f768(x768) { f767(x768)+b}
.func f769(x769) { f768(x769)+b}
.func f770(x770) { f769(x770)+b}
.func f771(x771) { f770(x771)+b}
.func f772(x772) { f771(x772)+b}
.func f773(x773) { f772(x773)+b}
.func f774(x774) { f773(x774)+b}
.func f775(x775) { f774(x775)+b}
.func f776(x776) { f775(x776)+b}
.func f777(x777) { f776(x777)+b}
.func f778(x778) { f777(x778)+b}
.func f779(x779) { f778(x779)+b}
.func f780(x780) { f779(x780)+b}
.func f781(x781) { f780(x781)+b}
.func f782(x782) { f781(x782)+b}
.func f783(x783) { f782(x783)+b}
.func f784(x784) { f783(x784)+b}
.func f785(x785) { f784(x785)+b}
.func f786(x786) { f785(x786)+b}
.func f787(x787) { f786(x787)+b}
.func f788(x788) { f787(x788)+b}
.func f789(x789) { f788(x789)+b}
.func f790(x790) { f789(x790)+b}
.func f791(x791) { f790(x791)+b}
.func f792(x792) { f791(x792)+b}
.func f793(x793) { f792(x793)+b}
.func f794(x794) { f793(x794)+b}
.func f795(x795) { f794(x795)+b}
.func f796(x796) { f795(x796)+b}
.func f797(x797) { f796(x797)+b}
.func f798(x798) { f797(x798)+b}
.func f799(x799) { f798(x799)+b}
.func f800(x800) { f799(x800)+b}
.func f801(x801) { f800(x801)+b}
.func f802(x802) { f801(x802)+b}
.func f803(x803) { f802(x803)+b}
.func f804(x804) { f803(x804)+b}
.func f805(x805) { f804(x805)+b}
.func f806(x806) { f805(x806)+b}
.func f807(x807) { f806(x807)+b}
.func f808(x808) { f807(x808)+b}
.func f809(x809) { f808(x809)+b}
.func f810(x810) { f809(x810)+b}
.func f811(x811) { f810(x811)+b}
.func f812(x812) { f811(x812)+b}
.func f813(x813) { f812(x813)+b}
.func f814(x814) { f813(x814)+b}
.func f815(x815) { f814(x815)+b}
.func f816(x816) { f815(x816)+b}
.func f817(x817) { f816(x817)+b}
.func f818(x818) { f817(x818)+b}
.func f819(x819) { f818(x819)+b}
.func f820(x820) { f819(x820)+b}
.func f821(x821) { f820(x821)+b}
.func f822(x822) { f821(x822)+b}
.func f823(x823) { f822(x823)+b}
.func f824(x824) { f823(x824)+b}
.func f825(x825) { f824(x825)+b}
.func f826(x826) { f825(x826)+b}
.func f827(x827) { f826(x827)+b}
.func f828(x828) { f827(x828)+b}
.func f829(x829) { f828(x829)+b}
.func f830(x830) { f829(x830)+b}
.func f831(x831) { f830(x831)+b}
.func f832(x832) { f831(x832)+b}
.func f833(x833) { f832(x833)+b}
.func f834(x834) { f833(x834)+b}
.func f835(x835) { f834(x835)+b}
.func f836(x836) { f835(x836)+b}
.func f837(x837) { f836(x837)+b}
.func f838(x838) { f837(x838)+b}
.func f839(x839) { f838(x839)+b}
.func f840(x840) { f839(x840)+b}
.func f841(x841) { f840(x841)+b}
.func f842(x842) { f841(x842)+b}
.func f843(x843) { f842(x843)+b}
.func f844(x844) { f843(x844)+b}
.func f845(x845) { f844(x845)+b}
.func f846(x846) { f845(x846)+b}
.func f847(x847) { f846(x847)+b}
.func f848(x848) { f847(x848)+b}
.func f849(x849) { f848(x849)+b}
.func f850(x850) { f849(x850)+b}
.func f851(x851) { f850(x851)+b}
.func f852(x852) { f851(x852)+b}
.func f853(x853) { f852(x853)+b}
.func f854(x854) { f853(x854)+b}
.func f855(x855) { f854(x855)+b}
.func f856(x856) { f855(x856)+b}
.func f857(x857) { f856(x857)+b}
.func f858(x858) { f857(x858)+b}
.func f859(x859) { f858(x859)+b}
.func f860(x860) { f859(x860)+b}
.func f861(x861) { f860(x861)+b}
.func f862(x862) { f861(x862)+b}
.func f863(x863) { f862(x863)+b}
.func f864(x864) { f863(x864)+b}
.func f865(x865) { f864(x865)+b}
.func f866(x866) { f865(x866)+b}
.func f867(x867) { f866(x867)+b}
.func f868(x868) { f867(x868)+b}
.func f869(x869) { f868(x869)+b}
.func f870(x870) { f869(x870)+b}
.func f871(x871) { f870(x871)+b}
.func f872(x872) { f871(x872)+b}
.func f873(x873) { f872(x873)+b}
.func f874(x874) { f873(x874)+b}
.func f875(x875) { f874(x875)+b}
.func f876(x876) { f875(x876)+b}
.func f877(x877) { f876(x877)+b}
.func f878(x878) { f877(x878)+b}
.func f879(x879) { f878(x879)+b}
.func f880(x880) { f879(x880)+b}
.func f881(x881) { f880(x881)+b}
.func f882(x882) { f881(x882)+b}
.func f883(x883) { f882(x883)+b}
.func f884(x884) { f883(x884)+b}
.func f885(x885) { f884(x885)+b}
.func f886(x886) { f885(x886)+b}
.func f887(x887) { f886(x887)+b}
.func f888(x888) { f887(x888)+b}
.func f889(x889) { f888(x889)+b}
.func f890(x890) { f889(x890)+b}
.func f891(x891) { f890(x891)+b}
.func f892(x892) { f891(x892)+b}
.func f893(x893) { f892(x893)+b}
.func f894(x894) { f893(x894)+b}
.func f895(x895) { f894(x895)+b}
.func f896(x896) { f895(x896)+b}
.func f897(x897) { f896(x897)+b}
.func f898(x898) { f897(x898)+b}
.func f899(x899) { f898(x899)+b}
.func f900(x900) { f899(x900)+b}
.func f901(x901) { f900(x901)+b}
.func f902(x902) { f901(x902)+b}
.func f903(x903) { f902(x903)+b}
.func f904(x904) { f903(x904)+b}
.func f905(x905) { f904(x905)+b}
.func f906(x906) { f905(x906)+b}
.func f907(x907) { f906(x907)+b}
.func f908(x908) { f907(x908)+b}
.func f909(x909) { f908(x909)+b}
.func f910(x910) { f909(x910)+b}
.func f911(x911) { f910(x911)+b}
.func f912(x912) { f911(x912)+b}
.func f913(x913) { f912(x913)+b}
.func f914(x914) { f913(x914)+b}
.func f915(x915) { f914(x915)+b}
.func f916(x916) { f915(x916)+b}
.func f917(x917) { f916(x917)+b}
.func f918(x918) { f917(x918)+b}
.func f919(x919) { f918(x919)+b}
.func f920(x920) { f919(x920)+b}
.func f921(x921) { f920(x921)+b}
.func f922(x922) { f921(x922)+b}
.func f923(x923) { f922(x923)+b}
.func f924(x924) { f923(x924)+b}
.func f925(x925) { f924(x925)+b}
.func f926(x926) { f925(x926)+b}
.func f927(x927) { f926(x927)+b}
.func f928(x928) { f927(x928)+b}
.func f929(x929) { f928(x929)+b}
.func f930(x930) { f929(x930)+b}
.func f931(x931) { f930(x931)+b}
.func f932(x932) { f931(x932)+b}
.func f933(x933) { f932(x933)+b}
.func f934(x934) { f933(x934)+b}
.func f935(x935) { f934(x935)+b}
.func f936(x936) { f935(x936)+b}
.func f937(x937) { f936(x937)+b}
.func f938(x938) { f937(x938)+b}
.func f939(x939) { f938(x939)+b}
.func f940(x940) { f939(x940)+b}
.func f941(x941) { f940(x941)+b}
.func f942(x942) { f941(x942)+b}
.func f943(x943) { f942(x943)+b}
.func f944(x944) { f943(x944)+b}
.func f945(x945) { f944(x945)+b}
.func f946(x946) { f945(x946)+b}
.func f947(x947) { f946(x947)+b}
.func f948(x948) { f947(x948)+b}
.func f949(x949) { f948(x949)+b}
.func f950(x950) { f949(x950)+b}
.func f951(x951) { f950(x951)+b}
.func f952(x952) { f951(x952)+b}
.func f953(x953) { f952(x953)+b}
.func f954(x954) { f953(x954)+b}
.func f955(x955) { f954(x955)+b}
.func f956(x956) { f955(x956)+b}
.func f957(x957) { f956(x957)+b}
.func f958(x958) { f957(x958)+b}
.func f959(x959) { f958(x959)+b}
.func f960(x960) { f959(x960)+b}
.func f961(x961) { f960(x961)+b}
.func f962(x962) { f961(x962)+b}
.func f963(x963) { f962(x963)+b}
.func f964(x964) { f963(x964)+b}
.func f965(x965) { f964(x965)+b}
.func f966(x966) { f965(x966)+b}
.func f967(x967) { f966(x967)+b}
.func f968(x968) { f967(x968)+b}
.func f969(x969) { f968(x969)+b}
.func f970(x970) { f969(x970)+b}
.func f971(x971) { f970(x971)+b}
.func f972(x972) { f971(x972)+b}
.func f973(x973) { f972(x973)+b}
.func f974(x974) { f973(x974)+b}
.func f975(x975) { f974(x975)+b}
.func f976(x976) { f975(x976)+b}
.func f977(x977) { f976(x977)+b}
.func f978(x978) { f977(x978)+b}
.func f979(x979) { f978(x979)+b}
.func f980(x980) { f979(x980)+b}
.func f981(x981) { f980(x981)+b}
.func f982(x982) { f981(x982)+b}
.func f983(x983) { f982(x983)+b}
.func f984(x984) { f983(x984)+b}
.func f985(x985) { f984(x985)+b}
.func f986(x986) { f985(x986)+b}
.func f987(x987) { f986(x987)+b}
.func f988(x988) { f987(x988)+b}
.func f989(x989) { f988(x989)+b}
.func f990(x990) { f989(x990)+b}
.func f991(x991) { f990(x991)+b}
.func f992(x992) { f991(x992)+b}
.func f993(x993) { f992(x993)+b}
.func f994(x994) { f993(x994)+b}
.func f995(x995) { f994(x995)+b}
.func f996(x996) { f995(x996)+b}
.func f997(x997) { f996(x997)+b}
.func f998(x998) { f997(x998)+b}
.func f999(x999) { f998(x999)+b}
.global_param test1 = { f999(arg1) + f999(arg2) }

.DC V1 1.0 1.0 1.0
R1 1 0 {test1}
V1 1 0 1.0

.print dc v(1) {R1:R} 

