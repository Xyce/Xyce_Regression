CMOS INVERTER
*
M1 2 1 0 0 NMOS W = 20U L = 5U
M2 2 1 3 3 PMOS W = 40U L = 5U
VDD 3 0 5
VIN 1 0 SIN 2.5 2.5 20MEG
.MODEL NMOS NMOS LEVEL = 3 CGDO = .2N CGSO = .2N CGBO = 2N
.MODEL PMOS PMOS LEVEL = 3 CGDO = .2N CGSO = .2N CGBO = 2N
*.OP
.TRAN 1N 100N
.FOUR 20MEG ID(M1) IG(M1) IS(M1) IB(M1)
.PRINT TRAN ID(M1) IG(M1) IS(M1) IB(M1)
.END
