Noise example adapted from the LTSpice educational examples directory.  
* The original name of the file was noise.asc.
*
Q5 N001 N006 N007 0 2N3904
Q7 N001 N007 OUT 0 2N2219A
Q8 OUT N013 N014 0 2N2219A
Q6 N013 N012 OUT 0 2N3906
V1 N001 0 10
V2 N014 0 -10
R11 N012 N014 5K
R14 OUT 0 8
R9 N006 N008 2K
R10 N008 N012 1K
Q4 N006 N008 N012 0 2N3904
Q1 N002 N009 N011 0 2N3904
Q2 N001 N010 N011 0 2N3904
R2 N001 N002 200
R3 N011 N014 1K
Q3 N006 N005 N004 0 2N3906
R6 N010 0 5K
R7 OUT N010 50K
V3 IN 0 AC 1
R1 N009 IN 5K
R8 N001 N004 100
R4 N003 N002 9K
C2 N006 N005 100p
C1 N003 N002 10p
R13 N013 N014 1K
R12 N007 OUT 1K
C3 N006 N012 .001u
R5 N005 N003 1K
*.model NPN NPN
*.model PNP PNP

.model 2N3904 NPN(IS=1E-14 VAF=100
+  Bf=300 IKF=0.4 XTB=1.5 BR=4
+  CJC=4E-12  CJE=8E-12 RB=20 RC=0.1 RE=0.1
+  TR=250E-9  TF=350E-12 ITF=1 VTF=2 XTF=3 
*+ Vceo=40 Icrating=200m mfg=Philips
+)

.model 2N3906 PNP(IS=1E-14 VAF=100
+  BF=200 IKF=0.4 XTB=1.5 BR=4
+  CJC=4.5E-12 CJE=10E-12 RB=20 RC=0.1 RE=0.1
+  TR=250E-9   TF=350E-12 ITF=1 VTF=2 XTF=3 
*+ Vceo=40  Icrating=200m mfg=Philips
+ )

.model 2N2219A  NPN(Is=14.34f Xti=3 Eg=1.11 Vaf=74.03 Bf=255.9 Ne=1.307 
+ Ise=14.34f Ikf=.2847 Xtb=1.5 Br=6.092 Nc=2 Isc=0 Ikr=0 Rc=1 Cjc=7.306p
+ Mjc=.3416 Vjc=.75 Fc=.5 Cje=22.01p Mje=.377 Vje=.75 Tr=46.91n Tf=411.1p 
+ Itf=.6 Vtf=1.7 Xtf=3 Rb=10 
*+ Vceo=40 Icrating=800m mfg=Philips
+ )

.noise V(out) V3 oct 100 1 20K

.options device debuglevel=-100

.end
