*Xyce netlist for testing E-sources syntaxes

.TRAN 0 1000ns
.PRINT TRAN FORMAT=PROBE V(N382405) V(N382063) V(N381794)
+ V(N386932) V(N395297) V(N395329)
+ V(N384791) V($G_CLK) V(2) V(3) V(4)

E_E1         N382063 0 VALUE 2*V(N382405,0)
E_E2         N381794 0 N380960 0 1.5
V_V2         N381000 0  1
R_R3         N381794 0  1 
R_R2         N382063 0  1 
R_R1         N382405 0  1 
V_V1         N382405 0  SIN(0V 1V 1e6 0 0 0)
V_V3         N380960 0  1

*test the E-Source POLY Syntax
E_E4         N386932 0 POLY(1) N380960 0 0.0 2
R_R7         N386932 0  1

*test the TABLE syntax
R_R21         N395329 0 1 
V_V13         N395297 0 SIN(0V 1V 1e6 0 0 0)
E_E5          N395329 0 TABLE V(N395297, 0) = (-1,-3) (1,3)

* test NOT (~) syntax in E-Source definition.
E_E3         N384791 0 VALUE IF( ~(V(N380960) >= 0) , 0, 1)
R_R4         N384791 0  1 

*Test of E-Source syntaxes with Global Node
RG1 $G_CLK 0 1
VG1 $G_CLK 0  SIN(0V 1V 1e6 0 0 0)

RG2  2 0 1
EG2  2 0 VALUE 2*V($G_CLK) 

RG3  3 0 1
EG3  3 0 VALUE 3*V($G_CLK) 

RG4  4 0 1
EG4  4 0 VALUE IF(((V($G_CLK) >= 0.8)&(V($G_CLK) >= 0.8)),3.5, 3.5)

.END