* Test AC mode support for the EQN measure.
* To be conservative, there are subtests for each
* valid operator (V, VR, VI, VP, VM and VDB) for
* each measure type.
*
* See SON Bug 1140 for more details
*****************************************************

* Trivial high-pass filter (V-C-R) circuit
R1 b 0 2
C1 a b 1u
V1 a 0 DC 0V AC 1

.print AC vr(b) vi(b) vm(b) vp(b) vdb(b)
.ac dec 5 100Hz 1e6
.STEP R1 0.5 2 1.5

* EQN
.MEASURE AC eqnvb eqn {1+v(b)}
.MEASURE AC eqnvmb eqn {1+vm(b)}
.MEASURE AC eqnvrb eqn {1+vr(b)}
.MEASURE AC eqnvib eqn {1+vi(b)}
.MEASURE AC eqnvpb eqn {1+vp(b)}
.MEASURE AC eqnvdbb eqn {1+vdb(b)}

* add FROM-TO
.MEASURE AC eqnvmbFromTo eqn {1+vm(b)} FROM=1e3 TO=1e5

* Tests should return -1 or -100, since the FROM-T0 window 
* has various problems
.measure ac eqnReturnNegOne eqn v(b) FROM=1e7 TO=1e8
.measure ac maxReturnNeg100 max vr(b) FROM=1e6 TO=1e2 DEFAULT_VAL=-100

* Signifies end of test. .sh file looks for a measure named lastMeasure.  
* This is needed for compatibility for testing with a verbose build, which 
* is often used by the Xyce developers.
.measure ac lastMeasure eqn {1+vm(b)} 

.end

