*Id-Vd Characteristics for NMOS 

.include "nmos_b3soi.mod"
.options device temp=25

* --- Voltage Sources ---
vd drain  0 dc 0
vg gate  0 dc 1
vs source 0 dc 0
ve substrate 0 0
 
* --- Transistor ---
m1 drain gate source substrate  nmos1 W=1e-5 L=1e-6  

* --- DC Analysis ---
.dc vd 0 1.2 0.01 vg 0.2 1.2 0.1

.step TEMP list 15 25 35

.print dc v(drain) v(gate) id(m1)
.end
