********************************************************
* Test that .PRINT PCE output in an unsupported format
* (RAW, PROBE, TOUCHSTONE and TOUCHSTONE2) defaults
* to STD format (.prn file with an Index column).  This
* tests with .OP rather than with .DC
*
* See SON Bug 1231 for more details.
********************************************************

.global_param R1value={1000.0}
.global_param R2value={1000.0}
.global_param Vvalue={5.0}

R2 1 0 {R2value}
R1 1 2 {R1value}
Von 2 0 {Vvalue}

.op

.print dc format=tecplot v(1)
.PRINT PCE PRECISION=6 FILE=pce-formats-default-to-prn.cir.PCE.raw FORMAT=RAW
.PRINT PCE PRECISION=6 FILE=pce-formats-default-to-prn.cir.PCE.probe FORMAT=PROBE
.PRINT PCE PRECISION=6 FILE=pce-formats-default-to-prn.cir.PCE.ts1 FORMAT=TOUCHSTONE
.PRINT PCE PRECISION=6 FILE=pce-formats-default-to-prn.cir.PCE.ts2 FORMAT=TOUCHSTONE2

.PCE
+ param=R1value
+ type=normal
+ means=1000.0
+ std_deviations=200.0

.options PCES
+ order=2
+ outputs={v(1)}

.options nonlin nox=0

.end
