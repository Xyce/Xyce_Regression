* Test error handling in the function extractSourceData().
* The instance lines for V1 and I2 are missing a value after
* the DC keyword.  The instance lines for V3 and I4 do not
* have a valid numeric value after the DC keyword. See SON 
* Bug 1087 for details.
V1 1 0 DC
R1 1 0 1

I2 2 0 DC
R2 2 0 1

V3 3 0 DC V
R3 3 0 1

I4 4 0 DC A
I4 4 0 1

.DC V1 1 5 1
.PRINT DC V(1) V(2) V(3) V(4)
.END

