* In this netlist, the multi-character wildcards should be silently
* ignored.  The V(a*) and I(V*) wildcards should work though.
*
* See SON Bug 1211 for more details.
*
* Trivial low-pass filter (V-L-R) circuits.
*

R1 b1 0 2
L1 a1 b1 1u
V1 a1 0 DC 0V AC 1

R2 b2 0 2
L2 a2 b2 1u
V2 a2 0 DC 0V AC 1

.print AC V(a*) VR(a*) VDB(a*) I(V*) IR(V*) IDB(V*)
.ac dec 5 100Hz 10e6

.end
