Lead current test for vdmos
*
VD 0 3 -0.5
VG 0 4 10 pulse(0 -10 300ns 50ns 50ns 400ns 1000ns)
VS 0 2 0
VB 0 1 0
M1 3 4 2 1 IRF130 W=0.386 L=2.5u
*
VDp 0 3p 0.5
VGp 0 4p 10 pulse(0 10 300ns 50ns 50ns 400ns 1000ns)
VSp 0 2p 0
VBp 0 1p 0
M1p 3p 4p 2p 1p IRF130p W=0.386 L=2.5u
*
.MODEL IRF130 NMOS LEVEL=18
+ CV=1
+ CVE=1
+ VTO=3.5
+ RD= 0
+ RS= 0.005
+ LAMBDA=0
+ M=3
+ SIGMA0=0
+ UO=230
+ VMAX=4e4
+ DELTA=5
+ TOX=50nm
*
.MODEL IRF130p PMOS LEVEL=18
+ CV=1
+ CVE=1
+ VTO=-3.5
+ RD= 0
+ RS= 0.005
+ LAMBDA=0
+ M=3
+ SIGMA0=0
+ UO=230
+ VMAX=4e4
+ DELTA=5
+ TOX=50nm
*
.TRAN 0.5n 1u 0u 2n
*COMP {I(VD)-ID(M1)} abstol=2.0e-6 zerotol=1.0e-7
*COMP {I(VG)-IG(M1)} abstol=2.0e-6 zerotol=1.0e-7
*COMP {I(VS)-IS(M1)} abstol=2.0e-6 zerotol=1.0e-7
*COMP {I(VB)-IB(M1)} abstol=2.0e-6 zerotol=1.0e-7
*COMP {I(VDp)-ID(M1p)} abstol=2.0e-6 zerotol=1.0e-7
*COMP {I(VGp)-IG(M1p)} abstol=2.0e-6 zerotol=1.0e-7
*COMP {I(VSp)-IS(M1p)} abstol=2.0e-6 zerotol=1.0e-7
*COMP {I(VBp)-IB(M1p)} abstol=2.0e-6 zerotol=1.0e-7

.PRINT TRAN {I(VD)-ID(M1)} {I(VG)-IG(M1)} {I(VS)-IS(M1)} {I(VB)-IB(M1)}
+ {I(VDp)-ID(M1p)} {I(VGp)-IG(M1p)} {I(VSp)-IS(M1p)} {I(VBp)-IB(M1p)}
.options timeint method=trap newbpstepping=0
.options nonlin-tran rhstol=1.0e-7
.END

