smult20.sp SPICE FILE
.model nenh nmos
+ level = 2
+   vto = 0.688434   kp = 4.769e-05   gamma = 0.399818
+   phi = 0.85
+
+   cgso = 3.54e-10   cgdo = 3.54e-10
+   rsh = 70   cj = 0.000363
+   mj = 0.916   cjsw = 1.83e-10   mjsw = 0.195
+   tox = 2.15e-08   nsub = 1.79246e+16
+   nss = 3e+10   nfs = 10   tpg = 1
+   xj = 9e-07   ld = -8.3e-08   uo = 683.594
+   ucrit = 200   uexp = 0.0177713
+   vmax = 81459.2   neff = 2.18502
+
+   delta = 2.72869
.model penh pmos
+ level = 2
+   vto = -0.635779   kp = 1.91591e-05   gamma = 0.335224
+   phi = 0.85
+
+   cgso = 4.01e-10   cgdo = 4.01e-10
+   rsh = 164   cj = 0.000442
+   mj = 0.3285   cjsw = 2.34e-10   mjsw = 0.307
+   tox = 2.15e-08   nsub = 6e+17
+   nss = 3e+10   nfs = 85.3597   tpg = -1
+   xj = 1e-09   ld = -2.3e-08   uo = 41.2542
+   ucrit = 50408.2   uexp = 0.0976377
+   vmax = 42755.1   neff = 0.0107262
+
+   delta = 4.72482
m0 3 5 4 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m1 1 6 3 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m2 7 8 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m3 1 8 7 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m4 8 5 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m5 1 9 8 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m6 6 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m7 10 5 11 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m8 1 12 10 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m9 13 14 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m10 1 14 13 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m11 14 5 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m12 1 15 14 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m13 12 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m14 4 5 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m15 0 6 4 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m16 7 4 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m17 0 4 7 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m18 16 5 8 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m19 0 9 16 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m20 6 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m21 1 17 5 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m22 18 5 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m23 17 19 18 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m24 11 5 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m25 0 12 11 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m26 13 11 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m27 0 11 13 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m28 20 5 14 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m29 0 15 20 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m30 12 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m31 1 22 21 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m32 23 21 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m33 24 25 23 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m34 22 26 24 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m35 27 28 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m36 1 28 27 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m37 29 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m38 28 31 29 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m39 32 33 28 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m40 1 34 32 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m41 34 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m42 0 17 5 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m43 21 19 17 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m44 0 22 21 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m45 35 21 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m46 22 19 35 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m47 18 5 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m48 22 25 36 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=1.098e-11 ps=8.66e-06 pd=1.33e-05 
+ nrs=0.6 nrd=0.85 
m49 27 26 22 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m50 0 37 22 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m51 27 28 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m52 0 28 27 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m53 38 34 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m54 28 31 38 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m55 39 33 28 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m56 0 30 39 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m57 34 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m58 40 42 41 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m59 1 43 40 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m60 44 45 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m61 1 45 44 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m62 45 42 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m63 1 9 45 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m64 43 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m65 46 42 47 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m66 1 48 46 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m67 49 50 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m68 1 50 49 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m69 50 42 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m70 1 15 50 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m71 48 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m72 41 42 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m73 0 43 41 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m74 44 41 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m75 0 41 44 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m76 51 42 45 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m77 0 9 51 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m78 43 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m79 1 52 42 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m80 53 42 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m81 52 19 53 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m82 47 42 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m83 0 48 47 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m84 49 47 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m85 0 47 49 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m86 54 42 50 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m87 0 15 54 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m88 48 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m89 1 56 55 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m90 57 55 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m91 58 25 57 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m92 56 26 58 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m93 59 60 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m94 1 60 59 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m95 61 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m96 60 62 61 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m97 63 64 60 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m98 1 65 63 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m99 65 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m100 0 52 42 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m101 55 19 52 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m102 0 56 55 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m103 66 55 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m104 56 19 66 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m105 53 42 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m106 56 25 5 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m107 59 26 56 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m108 0 37 56 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m109 59 60 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m110 0 60 59 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m111 67 65 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m112 60 62 67 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m113 68 64 60 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m114 0 30 68 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m115 65 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m116 69 71 70 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m117 1 72 69 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m118 73 74 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m119 1 74 73 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m120 74 71 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m121 1 9 74 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m122 72 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m123 75 71 76 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m124 1 77 75 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m125 78 79 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m126 1 79 78 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m127 79 71 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m128 1 15 79 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m129 77 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m130 70 71 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m131 0 72 70 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m132 73 70 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m133 0 70 73 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m134 80 71 74 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m135 0 9 80 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m136 72 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m137 1 81 71 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m138 82 71 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m139 81 19 82 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m140 76 71 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m141 0 77 76 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m142 78 76 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m143 0 76 78 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m144 83 71 79 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m145 0 15 83 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m146 77 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m147 1 85 84 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m148 86 84 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m149 87 25 86 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m150 85 26 87 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m151 88 89 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m152 1 89 88 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m153 90 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m154 89 91 90 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m155 92 93 89 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m156 1 94 92 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m157 94 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m158 0 81 71 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m159 84 19 81 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m160 0 85 84 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m161 95 84 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m162 85 19 95 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m163 82 71 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m164 85 25 42 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m165 88 26 85 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m166 0 37 85 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m167 88 89 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m168 0 89 88 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m169 96 94 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m170 89 91 96 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m171 97 93 89 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m172 0 30 97 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m173 94 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m174 98 100 99 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m175 1 101 98 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m176 102 103 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m177 1 103 102 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m178 103 100 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m179 1 9 103 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m180 101 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m181 104 100 105 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m182 1 106 104 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m183 107 108 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m184 1 108 107 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m185 108 100 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m186 1 15 108 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m187 106 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m188 99 100 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m189 0 101 99 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m190 102 99 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m191 0 99 102 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m192 109 100 103 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m193 0 9 109 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m194 101 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m195 1 110 100 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m196 111 100 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m197 110 19 111 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m198 105 100 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m199 0 106 105 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m200 107 105 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m201 0 105 107 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m202 112 100 108 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m203 0 15 112 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m204 106 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m205 1 114 113 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m206 115 113 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m207 116 25 115 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m208 114 26 116 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m209 117 118 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m210 1 118 117 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m211 119 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m212 118 120 119 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m213 121 122 118 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m214 1 123 121 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m215 123 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m216 0 110 100 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m217 113 19 110 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m218 0 114 113 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m219 124 113 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m220 114 19 124 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m221 111 100 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m222 114 25 71 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m223 117 26 114 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m224 0 37 114 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m225 117 118 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m226 0 118 117 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m227 125 123 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m228 118 120 125 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m229 126 122 118 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m230 0 30 126 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m231 123 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m232 127 129 128 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m233 1 130 127 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m234 131 132 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m235 1 132 131 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m236 132 129 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m237 1 9 132 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m238 130 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m239 133 129 134 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m240 1 135 133 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m241 136 137 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m242 1 137 136 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m243 137 129 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m244 1 15 137 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m245 135 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m246 128 129 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m247 0 130 128 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m248 131 128 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m249 0 128 131 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m250 138 129 132 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m251 0 9 138 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m252 130 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m253 1 139 129 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m254 140 129 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m255 139 19 140 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m256 134 129 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m257 0 135 134 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m258 136 134 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m259 0 134 136 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m260 141 129 137 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m261 0 15 141 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m262 135 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m263 1 143 142 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m264 144 142 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m265 145 25 144 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m266 143 26 145 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m267 146 147 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m268 1 147 146 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m269 148 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m270 147 149 148 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m271 150 151 147 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m272 1 152 150 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m273 152 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m274 0 139 129 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m275 142 19 139 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m276 0 143 142 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m277 153 142 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m278 143 19 153 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m279 140 129 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m280 143 25 100 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m281 146 26 143 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m282 0 37 143 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m283 146 147 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m284 0 147 146 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m285 154 152 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m286 147 149 154 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m287 155 151 147 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m288 0 30 155 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m289 152 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m290 156 158 157 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m291 1 159 156 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m292 160 161 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m293 1 161 160 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m294 161 158 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m295 1 9 161 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m296 159 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m297 162 158 163 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m298 1 164 162 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m299 165 166 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m300 1 166 165 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m301 166 158 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m302 1 15 166 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m303 164 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m304 157 158 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m305 0 159 157 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m306 160 157 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m307 0 157 160 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m308 167 158 161 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m309 0 9 167 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m310 159 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m311 1 168 158 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m312 169 158 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m313 168 19 169 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m314 163 158 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m315 0 164 163 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m316 165 163 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m317 0 163 165 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m318 170 158 166 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m319 0 15 170 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m320 164 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m321 1 172 171 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m322 173 171 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m323 174 25 173 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m324 172 26 174 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m325 175 176 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m326 1 176 175 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m327 177 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m328 176 178 177 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m329 179 180 176 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m330 1 181 179 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m331 181 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m332 0 168 158 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m333 171 19 168 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m334 0 172 171 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m335 182 171 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m336 172 19 182 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m337 169 158 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m338 172 25 129 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m339 175 26 172 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m340 0 37 172 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m341 175 176 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m342 0 176 175 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m343 183 181 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m344 176 178 183 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m345 184 180 176 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m346 0 30 184 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m347 181 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m348 185 187 186 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m349 1 188 185 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m350 189 190 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m351 1 190 189 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m352 190 187 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m353 1 9 190 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m354 188 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m355 191 187 192 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m356 1 193 191 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m357 194 195 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m358 1 195 194 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m359 195 187 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m360 1 15 195 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m361 193 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m362 186 187 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m363 0 188 186 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m364 189 186 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m365 0 186 189 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m366 196 187 190 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m367 0 9 196 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m368 188 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m369 1 197 187 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m370 198 187 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m371 197 19 198 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m372 192 187 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m373 0 193 192 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m374 194 192 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m375 0 192 194 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m376 199 187 195 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m377 0 15 199 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m378 193 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m379 1 201 200 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m380 202 200 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m381 203 25 202 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m382 201 26 203 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m383 204 205 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m384 1 205 204 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m385 206 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m386 205 207 206 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m387 208 209 205 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m388 1 210 208 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m389 210 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m390 0 197 187 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m391 200 19 197 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m392 0 201 200 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m393 211 200 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m394 201 19 211 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m395 198 187 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m396 201 25 158 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m397 204 26 201 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m398 0 37 201 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m399 204 205 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m400 0 205 204 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m401 212 210 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m402 205 207 212 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m403 213 209 205 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m404 0 30 213 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m405 210 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m406 214 216 215 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m407 1 217 214 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m408 218 219 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m409 1 219 218 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m410 219 216 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m411 1 9 219 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m412 217 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m413 220 216 221 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m414 1 222 220 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m415 223 224 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m416 1 224 223 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m417 224 216 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m418 1 15 224 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m419 222 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m420 215 216 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m421 0 217 215 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m422 218 215 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m423 0 215 218 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m424 225 216 219 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m425 0 9 225 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m426 217 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m427 1 226 216 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m428 227 216 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m429 226 19 227 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m430 221 216 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m431 0 222 221 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m432 223 221 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m433 0 221 223 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m434 228 216 224 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m435 0 15 228 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m436 222 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m437 1 230 229 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m438 231 229 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m439 232 25 231 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m440 230 26 232 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m441 233 234 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m442 1 234 233 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m443 235 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m444 234 236 235 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m445 237 238 234 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m446 1 239 237 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m447 239 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m448 0 226 216 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m449 229 19 226 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m450 0 230 229 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m451 240 229 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m452 230 19 240 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m453 227 216 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m454 230 25 187 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m455 233 26 230 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m456 0 37 230 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m457 233 234 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m458 0 234 233 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m459 241 239 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m460 234 236 241 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m461 242 238 234 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m462 0 30 242 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m463 239 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m464 243 245 244 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m465 1 246 243 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m466 247 248 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m467 1 248 247 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m468 248 245 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m469 1 9 248 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m470 246 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m471 249 245 250 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m472 1 251 249 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m473 252 253 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m474 1 253 252 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m475 253 245 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m476 1 15 253 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m477 251 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m478 244 245 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m479 0 246 244 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m480 247 244 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m481 0 244 247 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m482 254 245 248 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m483 0 9 254 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m484 246 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m485 1 255 245 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m486 256 245 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m487 255 19 256 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m488 250 245 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m489 0 251 250 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m490 252 250 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m491 0 250 252 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m492 257 245 253 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m493 0 15 257 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m494 251 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m495 1 259 258 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m496 260 258 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m497 261 25 260 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m498 259 26 261 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m499 262 263 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m500 1 263 262 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m501 264 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m502 263 265 264 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m503 266 267 263 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m504 1 268 266 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m505 268 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m506 0 255 245 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m507 258 19 255 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m508 0 259 258 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m509 269 258 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m510 259 19 269 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m511 256 245 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m512 259 25 216 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m513 262 26 259 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m514 0 37 259 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m515 262 263 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m516 0 263 262 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m517 270 268 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m518 263 265 270 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m519 271 267 263 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m520 0 30 271 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m521 268 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m522 272 274 273 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m523 1 275 272 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m524 276 277 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m525 1 277 276 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m526 277 274 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m527 1 9 277 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m528 275 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m529 278 274 279 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m530 1 280 278 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m531 281 282 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m532 1 282 281 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m533 282 274 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m534 1 15 282 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m535 280 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m536 273 274 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m537 0 275 273 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m538 276 273 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m539 0 273 276 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m540 283 274 277 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m541 0 9 283 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m542 275 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m543 1 284 274 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m544 285 274 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m545 284 19 285 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m546 279 274 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m547 0 280 279 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m548 281 279 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m549 0 279 281 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m550 286 274 282 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m551 0 15 286 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m552 280 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m553 1 288 287 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m554 289 287 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m555 290 25 289 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m556 288 26 290 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m557 291 292 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m558 1 292 291 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m559 293 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m560 292 294 293 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m561 295 296 292 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m562 1 297 295 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m563 297 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m564 0 284 274 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m565 287 19 284 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m566 0 288 287 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m567 298 287 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m568 288 19 298 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m569 285 274 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m570 288 25 245 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m571 291 26 288 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m572 0 37 288 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m573 291 292 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m574 0 292 291 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m575 299 297 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m576 292 294 299 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m577 300 296 292 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m578 0 30 300 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m579 297 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m580 301 303 302 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m581 1 304 301 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m582 305 306 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m583 1 306 305 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m584 306 303 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m585 1 9 306 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m586 304 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m587 307 303 308 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m588 1 309 307 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m589 310 311 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m590 1 311 310 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m591 311 303 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m592 1 15 311 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m593 309 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m594 302 303 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m595 0 304 302 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m596 305 302 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m597 0 302 305 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m598 312 303 306 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m599 0 9 312 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m600 304 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m601 1 313 303 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m602 314 303 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m603 313 19 314 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m604 308 303 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m605 0 309 308 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m606 310 308 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m607 0 308 310 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m608 315 303 311 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m609 0 15 315 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m610 309 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m611 1 317 316 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m612 318 316 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m613 319 25 318 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m614 317 26 319 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m615 320 321 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m616 1 321 320 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m617 322 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m618 321 323 322 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m619 324 325 321 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m620 1 326 324 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m621 326 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m622 0 313 303 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m623 316 19 313 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m624 0 317 316 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m625 327 316 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m626 317 19 327 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m627 314 303 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m628 317 25 274 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m629 320 26 317 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m630 0 37 317 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m631 320 321 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m632 0 321 320 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m633 328 326 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m634 321 323 328 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m635 329 325 321 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m636 0 30 329 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m637 326 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m638 330 332 331 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m639 1 333 330 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m640 334 335 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m641 1 335 334 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m642 335 332 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m643 1 9 335 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m644 333 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m645 336 332 337 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m646 1 338 336 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m647 339 340 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m648 1 340 339 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m649 340 332 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m650 1 15 340 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m651 338 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m652 331 332 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m653 0 333 331 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m654 334 331 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m655 0 331 334 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m656 341 332 335 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m657 0 9 341 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m658 333 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m659 1 342 332 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m660 343 332 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m661 342 19 343 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m662 337 332 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m663 0 338 337 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m664 339 337 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m665 0 337 339 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m666 344 332 340 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m667 0 15 344 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m668 338 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m669 1 346 345 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m670 347 345 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m671 348 25 347 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m672 346 26 348 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m673 349 350 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m674 1 350 349 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m675 351 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m676 350 352 351 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m677 353 354 350 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m678 1 355 353 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m679 355 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m680 0 342 332 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m681 345 19 342 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m682 0 346 345 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m683 356 345 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m684 346 19 356 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m685 343 332 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m686 346 25 303 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m687 349 26 346 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m688 0 37 346 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m689 349 350 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m690 0 350 349 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m691 357 355 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m692 350 352 357 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m693 358 354 350 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m694 0 30 358 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m695 355 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m696 359 361 360 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m697 1 362 359 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m698 363 364 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m699 1 364 363 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m700 364 361 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m701 1 9 364 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m702 362 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m703 365 361 366 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m704 1 367 365 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m705 368 369 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m706 1 369 368 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m707 369 361 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m708 1 15 369 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m709 367 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m710 360 361 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m711 0 362 360 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m712 363 360 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m713 0 360 363 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m714 370 361 364 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m715 0 9 370 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m716 362 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m717 1 371 361 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m718 372 361 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m719 371 19 372 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m720 366 361 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m721 0 367 366 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m722 368 366 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m723 0 366 368 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m724 373 361 369 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m725 0 15 373 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m726 367 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m727 1 375 374 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m728 376 374 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m729 377 25 376 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m730 375 26 377 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m731 378 379 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m732 1 379 378 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m733 380 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m734 379 381 380 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m735 382 383 379 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m736 1 384 382 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m737 384 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m738 0 371 361 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m739 374 19 371 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m740 0 375 374 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m741 385 374 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m742 375 19 385 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m743 372 361 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m744 375 25 332 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m745 378 26 375 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m746 0 37 375 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m747 378 379 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m748 0 379 378 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m749 386 384 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m750 379 381 386 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m751 387 383 379 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m752 0 30 387 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m753 384 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m754 388 390 389 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m755 1 391 388 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m756 392 393 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m757 1 393 392 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m758 393 390 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m759 1 9 393 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m760 391 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m761 394 390 395 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m762 1 396 394 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m763 397 398 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m764 1 398 397 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m765 398 390 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m766 1 15 398 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m767 396 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m768 389 390 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m769 0 391 389 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m770 392 389 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m771 0 389 392 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m772 399 390 393 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m773 0 9 399 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m774 391 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m775 1 400 390 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m776 401 390 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m777 400 19 401 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m778 395 390 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m779 0 396 395 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m780 397 395 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m781 0 395 397 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m782 402 390 398 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m783 0 15 402 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m784 396 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m785 1 404 403 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m786 405 403 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m787 406 25 405 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m788 404 26 406 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m789 407 408 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m790 1 408 407 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m791 409 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m792 408 410 409 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m793 411 412 408 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m794 1 413 411 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m795 413 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m796 0 400 390 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m797 403 19 400 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m798 0 404 403 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m799 414 403 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m800 404 19 414 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m801 401 390 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m802 404 25 361 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m803 407 26 404 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m804 0 37 404 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m805 407 408 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m806 0 408 407 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m807 415 413 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m808 408 410 415 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m809 416 412 408 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m810 0 30 416 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m811 413 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m812 417 419 418 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m813 1 420 417 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m814 421 422 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m815 1 422 421 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m816 422 419 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m817 1 9 422 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m818 420 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m819 423 419 424 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m820 1 425 423 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m821 426 427 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m822 1 427 426 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m823 427 419 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m824 1 15 427 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m825 425 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m826 418 419 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m827 0 420 418 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m828 421 418 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m829 0 418 421 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m830 428 419 422 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m831 0 9 428 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m832 420 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m833 1 429 419 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m834 430 419 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m835 429 19 430 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m836 424 419 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m837 0 425 424 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m838 426 424 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m839 0 424 426 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m840 431 419 427 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m841 0 15 431 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m842 425 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m843 1 433 432 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m844 434 432 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m845 435 25 434 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m846 433 26 435 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m847 436 437 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m848 1 437 436 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m849 438 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m850 437 439 438 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m851 440 441 437 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m852 1 442 440 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m853 442 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m854 0 429 419 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m855 432 19 429 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m856 0 433 432 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m857 443 432 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m858 433 19 443 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m859 430 419 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m860 433 25 390 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m861 436 26 433 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m862 0 37 433 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m863 436 437 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m864 0 437 436 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m865 444 442 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m866 437 439 444 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m867 445 441 437 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m868 0 30 445 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m869 442 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m870 446 448 447 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m871 1 449 446 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m872 450 451 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m873 1 451 450 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m874 451 448 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m875 1 9 451 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m876 449 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m877 452 448 453 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m878 1 454 452 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m879 455 456 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m880 1 456 455 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m881 456 448 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m882 1 15 456 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m883 454 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m884 447 448 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m885 0 449 447 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m886 450 447 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m887 0 447 450 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m888 457 448 451 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m889 0 9 457 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m890 449 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m891 1 458 448 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m892 459 448 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m893 458 19 459 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m894 453 448 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m895 0 454 453 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m896 455 453 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m897 0 453 455 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m898 460 448 456 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m899 0 15 460 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m900 454 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m901 1 462 461 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m902 463 461 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m903 464 25 463 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m904 462 26 464 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m905 465 466 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m906 1 466 465 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m907 467 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m908 466 468 467 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m909 469 470 466 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m910 1 471 469 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m911 471 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m912 0 458 448 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m913 461 19 458 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m914 0 462 461 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m915 472 461 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m916 462 19 472 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m917 459 448 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m918 462 25 419 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m919 465 26 462 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m920 0 37 462 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m921 465 466 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m922 0 466 465 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m923 473 471 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m924 466 468 473 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m925 474 470 466 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m926 0 30 474 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m927 471 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m928 475 477 476 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m929 1 478 475 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m930 479 480 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m931 1 480 479 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m932 480 477 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m933 1 9 480 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m934 478 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m935 481 477 482 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m936 1 483 481 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m937 484 485 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m938 1 485 484 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m939 485 477 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m940 1 15 485 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m941 483 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m942 476 477 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m943 0 478 476 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m944 479 476 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m945 0 476 479 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m946 486 477 480 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m947 0 9 486 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m948 478 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m949 1 487 477 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m950 488 477 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m951 487 19 488 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m952 482 477 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m953 0 483 482 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m954 484 482 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m955 0 482 484 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m956 489 477 485 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m957 0 15 489 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m958 483 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m959 1 491 490 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m960 492 490 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m961 493 25 492 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m962 491 26 493 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m963 494 495 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m964 1 495 494 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m965 496 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m966 495 497 496 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m967 498 499 495 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m968 1 500 498 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m969 500 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m970 0 487 477 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m971 490 19 487 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m972 0 491 490 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m973 501 490 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m974 491 19 501 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m975 488 477 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m976 491 25 448 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m977 494 26 491 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m978 0 37 491 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m979 494 495 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m980 0 495 494 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m981 502 500 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m982 495 497 502 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m983 503 499 495 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m984 0 30 503 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m985 500 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m986 504 506 505 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m987 1 507 504 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m988 508 509 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m989 1 509 508 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m990 509 506 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m991 1 9 509 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m992 507 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m993 510 506 511 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m994 1 512 510 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m995 513 514 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m996 1 514 513 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m997 514 506 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m998 1 15 514 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m999 512 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m1000 505 506 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m1001 0 507 505 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m1002 508 505 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m1003 0 505 508 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m1004 515 506 509 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m1005 0 9 515 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m1006 507 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m1007 1 516 506 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m1008 517 506 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m1009 516 19 517 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m1010 511 506 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m1011 0 512 511 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m1012 513 511 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m1013 0 511 513 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m1014 518 506 514 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m1015 0 15 518 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m1016 512 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m1017 1 520 519 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1018 521 519 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m1019 522 25 521 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1020 520 26 522 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m1021 523 524 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m1022 1 524 523 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m1023 525 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m1024 524 526 525 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m1025 527 528 524 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m1026 1 529 527 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m1027 529 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m1028 0 516 506 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m1029 519 19 516 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m1030 0 520 519 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m1031 530 519 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m1032 520 19 530 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m1033 517 506 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m1034 520 25 477 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m1035 523 26 520 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m1036 0 37 520 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m1037 523 524 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m1038 0 524 523 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m1039 531 529 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m1040 524 526 531 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m1041 532 528 524 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m1042 0 30 532 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m1043 529 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m1044 533 535 534 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m1045 1 536 533 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m1046 537 538 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m1047 1 538 537 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m1048 538 535 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m1049 1 9 538 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m1050 536 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m1051 539 535 540 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m1052 1 541 539 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m1053 542 543 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m1054 1 543 542 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m1055 543 535 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m1056 1 15 543 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m1057 541 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m1058 534 535 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m1059 0 536 534 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m1060 537 534 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m1061 0 534 537 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m1062 544 535 538 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m1063 0 9 544 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m1064 536 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m1065 1 545 535 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m1066 546 535 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m1067 545 19 546 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m1068 540 535 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m1069 0 541 540 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m1070 542 540 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m1071 0 540 542 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m1072 547 535 543 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m1073 0 15 547 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m1074 541 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m1075 1 549 548 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1076 550 548 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m1077 551 25 550 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1078 549 26 551 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m1079 552 553 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m1080 1 553 552 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m1081 554 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m1082 553 33 554 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m1083 555 556 553 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m1084 1 557 555 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m1085 557 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m1086 0 545 535 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m1087 548 19 545 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m1088 0 549 548 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m1089 558 548 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m1090 549 19 558 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m1091 546 535 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m1092 549 25 506 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m1093 552 26 549 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m1094 0 37 549 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m1095 552 553 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m1096 0 553 552 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m1097 559 557 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m1098 553 33 559 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m1099 560 556 553 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m1100 0 30 560 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m1101 557 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m1102 561 563 562 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.744e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.22 
m1103 1 564 561 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m1104 565 566 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m1105 1 566 565 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m1106 566 563 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m1107 1 9 566 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m1108 564 9 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m1109 567 563 568 1 penh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=2.52e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.2 
m1110 1 569 567 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=9.52e-12 ps=2.114e-05 pd=1.29e-05 
+ nrs=0.2 nrd=0.08 
m1111 570 571 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m1112 1 571 570 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m1113 571 563 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m1114 1 15 571 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m1115 569 15 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m1116 562 563 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m1117 0 564 562 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m1118 565 562 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m1119 0 562 565 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m1120 572 563 566 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m1121 0 9 572 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m1122 564 9 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m1123 1 573 563 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=2.572e-11 ps=2.265e-05 pd=2.69e-05 
+ nrs=0.19 nrd=0.18 
m1124 574 563 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=2.587e-11 ad=3.295e-11 ps=2.908e-05 pd=2.794e-05 
+ nrs=0.12 nrd=0.15 
m1125 573 19 574 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.19e-12 ps=1.25e-05 pd=4.72e-06 
+ nrs=1.63 nrd=0.73 
m1126 568 563 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m1127 0 569 568 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m1128 570 568 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.378e-11 ps=1.45e-05 pd=2.249e-05 
+ nrs=0.1 nrd=0.17 
m1129 0 568 570 0 nenh l=1.1e-06 w=1.2e-05 
+ as=2.378e-11 ad=1.452e-11 ps=2.249e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.1 
m1130 575 563 571 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=2.928e-11 ps=1.13e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.32 
m1131 0 15 575 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=8.16e-12 ps=1.799e-05 pd=1.13e-05 
+ nrs=0.21 nrd=0.09 
m1132 569 15 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m1133 1 577 576 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1134 578 576 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m1135 579 25 578 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1136 577 26 579 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m1137 580 581 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.386e-11 ad=2.583e-11 ps=1.41e-05 pd=2.19e-05 
+ nrs=0.1 nrd=0.19 
m1138 1 581 580 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=1.386e-11 ps=2.19e-05 pd=1.41e-05 
+ nrs=0.19 nrd=0.1 
m1139 582 30 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.059e-11 ad=2.405e-11 ps=1.381e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m1140 581 64 582 1 penh l=1.1e-06 w=1e-05 
+ as=1.25e-11 ad=9.81e-12 ps=1.25e-05 pd=1.279e-05 
+ nrs=0.13 nrd=0.1 
m1141 583 584 581 1 penh l=1.1e-06 w=1e-05 
+ as=9.81e-12 ad=1.25e-11 ps=1.279e-05 pd=1.25e-05 
+ nrs=0.1 nrd=0.13 
m1142 1 585 583 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.059e-11 ps=2.039e-05 pd=1.381e-05 
+ nrs=0.21 nrd=0.09 
m1143 585 30 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m1144 0 573 563 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.744e-11 ps=2.099e-05 pd=2.85e-05 
+ nrs=0.18 nrd=0.22 
m1145 576 19 573 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.6e-12 ad=1.098e-11 ps=7.28e-06 pd=1.33e-05 
+ nrs=0.59 nrd=0.85 
m1146 0 577 576 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.182e-11 ps=1.05e-05 pd=1.132e-05 
+ nrs=0.35 nrd=0.38 
m1147 586 576 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m1148 577 19 586 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m1149 574 563 0 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.624e-11 ad=2.537e-11 ps=2.85e-05 pd=2.399e-05 
+ nrs=0.16 nrd=0.15 
m1150 577 25 535 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m1151 580 26 577 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m1152 0 37 577 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m1153 580 581 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=1.11e-11 ps=1.207e-05 pd=1.05e-05 
+ nrs=0.37 nrd=0.35 
m1154 0 581 580 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.169e-11 ps=1.05e-05 pd=1.207e-05 
+ nrs=0.35 nrd=0.37 
m1155 587 585 0 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.007e-11 ad=2.22e-11 ps=1.605e-05 pd=2.099e-05 
+ nrs=0.08 nrd=0.18 
m1156 581 64 587 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.122e-11 ad=6.11e-12 ps=1.01e-05 pd=9.75e-06 
+ nrs=0.24 nrd=0.13 
m1157 588 584 581 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.11e-12 ad=1.122e-11 ps=9.75e-06 pd=1.01e-05 
+ nrs=0.13 nrd=0.24 
m1158 0 30 588 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=1.007e-11 ps=2.099e-05 pd=1.605e-05 
+ nrs=0.18 nrd=0.08 
m1159 585 30 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m1160 1 590 589 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1161 591 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1162 593 589 591 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1163 594 595 593 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1164 1 596 594 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1165 597 26 598 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1166 599 25 597 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1167 1 600 599 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1168 600 598 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1169 598 25 601 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1170 1 602 595 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1171 603 19 595 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1172 602 603 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1173 604 19 598 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1174 0 600 604 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1175 0 590 589 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1176 605 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1177 593 589 605 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1178 606 595 593 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1179 0 592 606 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1180 598 26 593 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1181 600 598 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1182 603 19 600 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1183 0 37 598 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1184 0 602 595 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=4.976e-11 ps=3.374e-05 pd=6.197e-05 
+ nrs=0.11 nrd=0.15 
m1185 602 603 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.455e-11 ad=3.726e-11 ps=6.627e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1186 1 608 607 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1187 609 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1188 610 607 609 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1189 611 612 610 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1190 1 596 611 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1191 613 26 614 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1192 615 25 613 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1193 1 616 615 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1194 616 614 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1195 614 25 617 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1196 1 601 612 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1197 618 19 612 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1198 601 618 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1199 619 19 614 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1200 0 616 619 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1201 0 608 607 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1202 620 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1203 610 607 620 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1204 621 612 610 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1205 0 592 621 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1206 614 26 610 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1207 616 614 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1208 618 19 616 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1209 0 37 614 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1210 0 601 612 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1211 601 618 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1212 1 623 622 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1213 624 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1214 625 622 624 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1215 626 627 625 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1216 1 596 626 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1217 628 26 629 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1218 630 25 628 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1219 1 631 630 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1220 631 629 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1221 629 25 632 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1222 1 617 627 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1223 633 19 627 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1224 617 633 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1225 634 19 629 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1226 0 631 634 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1227 0 623 622 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1228 635 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1229 625 622 635 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1230 636 627 625 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1231 0 592 636 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1232 629 26 625 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1233 631 629 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1234 633 19 631 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1235 0 37 629 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1236 0 617 627 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1237 617 633 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1238 1 638 637 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1239 639 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1240 640 637 639 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1241 641 642 640 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1242 1 596 641 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1243 643 26 644 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1244 645 25 643 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1245 1 646 645 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1246 646 644 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1247 644 25 647 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1248 1 632 642 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1249 648 19 642 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1250 632 648 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1251 649 19 644 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1252 0 646 649 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1253 0 638 637 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1254 650 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1255 640 637 650 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1256 651 642 640 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1257 0 592 651 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1258 644 26 640 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1259 646 644 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1260 648 19 646 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1261 0 37 644 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1262 0 632 642 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1263 632 648 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1264 1 653 652 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1265 654 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1266 655 652 654 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1267 656 657 655 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1268 1 596 656 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1269 658 26 659 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1270 660 25 658 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1271 1 661 660 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1272 661 659 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1273 659 25 662 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1274 1 647 657 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1275 663 19 657 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1276 647 663 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1277 664 19 659 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1278 0 661 664 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1279 0 653 652 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1280 665 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1281 655 652 665 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1282 666 657 655 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1283 0 592 666 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1284 659 26 655 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1285 661 659 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1286 663 19 661 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1287 0 37 659 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1288 0 647 657 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1289 647 663 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1290 1 668 667 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1291 669 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1292 670 667 669 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1293 671 672 670 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1294 1 596 671 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1295 673 26 674 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1296 675 25 673 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1297 1 676 675 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1298 676 674 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1299 674 25 677 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1300 1 662 672 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1301 678 19 672 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1302 662 678 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1303 679 19 674 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1304 0 676 679 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1305 0 668 667 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1306 680 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1307 670 667 680 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1308 681 672 670 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1309 0 592 681 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1310 674 26 670 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1311 676 674 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1312 678 19 676 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1313 0 37 674 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1314 0 662 672 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1315 662 678 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1316 1 683 682 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1317 684 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1318 685 682 684 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1319 686 687 685 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1320 1 596 686 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1321 688 26 689 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1322 690 25 688 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1323 1 691 690 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1324 691 689 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1325 689 25 692 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1326 1 677 687 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1327 693 19 687 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1328 677 693 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1329 694 19 689 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1330 0 691 694 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1331 0 683 682 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1332 695 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1333 685 682 695 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1334 696 687 685 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1335 0 592 696 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1336 689 26 685 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1337 691 689 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1338 693 19 691 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1339 0 37 689 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1340 0 677 687 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1341 677 693 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1342 1 698 697 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1343 699 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1344 700 697 699 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1345 701 702 700 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1346 1 596 701 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1347 703 26 704 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1348 705 25 703 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1349 1 706 705 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1350 706 704 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1351 704 25 707 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1352 1 692 702 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1353 708 19 702 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1354 692 708 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1355 709 19 704 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1356 0 706 709 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1357 0 698 697 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1358 710 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1359 700 697 710 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1360 711 702 700 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1361 0 592 711 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1362 704 26 700 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1363 706 704 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1364 708 19 706 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1365 0 37 704 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1366 0 692 702 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1367 692 708 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1368 1 713 712 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1369 714 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1370 715 712 714 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1371 716 717 715 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1372 1 596 716 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1373 718 26 719 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1374 720 25 718 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1375 1 721 720 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1376 721 719 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1377 719 25 722 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1378 1 707 717 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1379 723 19 717 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1380 707 723 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1381 724 19 719 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1382 0 721 724 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1383 0 713 712 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1384 725 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1385 715 712 725 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1386 726 717 715 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1387 0 592 726 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1388 719 26 715 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1389 721 719 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1390 723 19 721 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1391 0 37 719 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1392 0 707 717 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1393 707 723 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1394 1 728 727 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1395 729 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1396 730 727 729 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1397 731 732 730 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1398 1 596 731 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1399 733 26 734 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1400 735 25 733 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1401 1 736 735 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1402 736 734 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1403 734 25 737 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1404 1 722 732 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1405 738 19 732 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1406 722 738 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1407 739 19 734 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1408 0 736 739 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1409 0 728 727 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1410 740 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1411 730 727 740 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1412 741 732 730 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1413 0 592 741 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1414 734 26 730 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1415 736 734 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1416 738 19 736 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1417 0 37 734 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1418 0 722 732 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1419 722 738 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1420 1 743 742 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1421 744 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1422 745 742 744 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1423 746 747 745 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1424 1 596 746 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1425 748 26 749 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1426 750 25 748 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1427 1 751 750 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1428 751 749 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1429 749 25 752 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1430 1 737 747 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1431 753 19 747 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1432 737 753 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1433 754 19 749 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1434 0 751 754 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1435 0 743 742 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1436 755 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1437 745 742 755 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1438 756 747 745 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1439 0 592 756 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1440 749 26 745 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1441 751 749 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1442 753 19 751 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1443 0 37 749 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1444 0 737 747 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1445 737 753 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1446 1 758 757 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1447 759 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1448 760 757 759 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1449 761 762 760 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1450 1 596 761 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1451 763 26 764 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1452 765 25 763 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1453 1 766 765 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1454 766 764 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1455 764 25 767 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1456 1 752 762 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1457 768 19 762 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1458 752 768 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1459 769 19 764 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1460 0 766 769 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1461 0 758 757 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1462 770 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1463 760 757 770 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1464 771 762 760 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1465 0 592 771 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1466 764 26 760 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1467 766 764 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1468 768 19 766 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1469 0 37 764 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1470 0 752 762 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1471 752 768 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1472 1 773 772 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1473 774 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1474 775 772 774 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1475 776 777 775 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1476 1 596 776 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1477 778 26 779 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1478 780 25 778 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1479 1 781 780 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1480 781 779 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1481 779 25 782 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1482 1 767 777 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1483 783 19 777 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1484 767 783 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1485 784 19 779 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1486 0 781 784 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1487 0 773 772 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1488 785 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1489 775 772 785 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1490 786 777 775 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1491 0 592 786 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1492 779 26 775 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1493 781 779 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1494 783 19 781 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1495 0 37 779 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1496 0 767 777 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1497 767 783 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1498 1 788 787 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1499 789 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1500 790 787 789 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1501 791 792 790 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1502 1 596 791 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1503 793 26 794 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1504 795 25 793 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1505 1 796 795 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1506 796 794 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1507 794 25 797 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1508 1 782 792 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1509 798 19 792 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1510 782 798 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1511 799 19 794 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1512 0 796 799 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1513 0 788 787 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1514 800 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1515 790 787 800 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1516 801 792 790 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1517 0 592 801 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1518 794 26 790 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1519 796 794 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1520 798 19 796 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1521 0 37 794 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1522 0 782 792 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1523 782 798 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1524 1 803 802 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1525 804 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1526 805 802 804 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1527 806 807 805 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1528 1 596 806 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1529 808 26 809 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1530 810 25 808 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1531 1 811 810 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1532 811 809 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1533 809 25 812 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1534 1 797 807 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1535 813 19 807 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1536 797 813 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1537 814 19 809 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1538 0 811 814 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1539 0 803 802 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1540 815 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1541 805 802 815 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1542 816 807 805 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1543 0 592 816 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1544 809 26 805 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1545 811 809 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1546 813 19 811 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1547 0 37 809 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1548 0 797 807 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1549 797 813 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1550 1 818 817 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1551 819 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1552 820 817 819 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1553 821 822 820 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1554 1 596 821 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1555 823 26 824 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1556 825 25 823 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1557 1 826 825 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1558 826 824 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1559 824 25 827 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1560 1 812 822 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1561 828 19 822 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1562 812 828 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1563 829 19 824 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1564 0 826 829 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1565 0 818 817 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1566 830 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1567 820 817 830 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1568 831 822 820 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1569 0 592 831 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1570 824 26 820 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1571 826 824 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1572 828 19 826 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1573 0 37 824 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1574 0 812 822 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1575 812 828 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1576 1 833 832 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1577 834 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1578 835 832 834 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1579 836 837 835 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1580 1 596 836 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1581 838 26 839 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1582 840 25 838 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1583 1 841 840 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1584 841 839 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1585 839 25 842 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.32e-12 ps=1.146e-05 pd=1.093e-05 
+ nrs=1.26 nrd=0.91 
m1586 1 827 837 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1587 843 19 837 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1588 827 843 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1589 844 19 839 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1590 0 841 844 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1591 0 833 832 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1592 845 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1593 835 832 845 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1594 846 837 835 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1595 0 592 846 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1596 839 26 835 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1597 841 839 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1598 843 19 841 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1599 0 37 839 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1600 0 827 837 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1601 827 843 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1602 1 848 847 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1603 849 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1604 850 847 849 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1605 851 852 850 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1606 1 596 851 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1607 853 26 854 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1608 855 25 853 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1609 1 856 855 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1610 856 854 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1611 854 25 857 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=8.27e-12 ps=1.146e-05 pd=9.11e-06 
+ nrs=1.26 nrd=0.81 
m1612 1 858 852 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1613 859 19 852 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1614 858 859 1 1 penh l=1.1e-06 w=1.84e-05 
+ as=2.332e-11 ad=4.097e-11 ps=3.89e-05 pd=3.474e-05 
+ nrs=0.07 nrd=0.12 
m1615 860 19 854 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1616 0 856 860 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1617 0 848 847 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1618 861 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1619 850 847 861 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1620 862 852 850 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1621 0 592 862 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1622 854 26 850 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1623 856 854 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1624 859 19 856 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1625 0 37 854 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1626 0 858 852 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1627 858 859 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=4.602e-11 ad=3.171e-11 ps=5.54e-05 pd=2.999e-05 
+ nrs=0.18 nrd=0.12 
m1628 1 864 863 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1629 865 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1630 866 863 865 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1631 867 868 866 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1632 1 596 867 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1633 869 26 870 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1634 871 25 869 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1635 1 872 871 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1636 872 870 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1637 870 25 858 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.2e-12 ps=1.146e-05 pd=1.108e-05 
+ nrs=1.26 nrd=0.9 
m1638 1 842 868 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1639 873 19 868 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1640 842 873 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.786e-11 ad=4.72e-11 ps=4.45e-05 pd=4.002e-05 
+ nrs=0.06 nrd=0.11 
m1641 874 19 870 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1642 0 872 874 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1643 0 864 863 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1644 875 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1645 866 863 875 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1646 876 868 866 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1647 0 592 876 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1648 870 26 866 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1649 872 870 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1650 873 19 872 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1651 0 37 870 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1652 0 842 868 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.013e-11 ps=3.374e-05 pd=6.012e-05 
+ nrs=0.11 nrd=0.15 
m1653 842 873 0 0 nenh l=1.1e-06 w=1.88e-05 
+ as=5.474e-11 ad=3.726e-11 ps=6.424e-05 pd=3.524e-05 
+ nrs=0.15 nrd=0.11 
m1654 0 878 877 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.427e-11 ad=1.876e-11 ps=1.35e-05 pd=2.05e-05 
+ nrs=0.28 nrd=0.36 
m1655 878 879 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m1656 0 881 880 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.22e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.76 
m1657 881 882 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.22e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.76 nrd=0.5 
m1658 883 884 0 0 nenh l=1.1e-06 w=4.4e-06 
+ as=7.26e-12 ad=8.72e-12 ps=7.7e-06 pd=8.25e-06 
+ nrs=0.37 nrd=0.45 
m1659 0 884 883 0 nenh l=1.1e-06 w=4.4e-06 
+ as=8.72e-12 ad=7.26e-12 ps=8.25e-06 pd=7.7e-06 
+ nrs=0.45 nrd=0.37 
m1660 885 886 884 0 nenh l=1.1e-06 w=8.8e-06 
+ as=7.66e-12 ad=1.964e-11 ps=1.122e-05 pd=2.37e-05 
+ nrs=0.1 nrd=0.25 
m1661 887 888 885 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.4e-12 ps=1.25e-05 pd=1.378e-05 
+ nrs=0.08 nrd=0.08 
m1662 0 889 887 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m1663 890 886 0 0 nenh l=1.1e-06 w=8.8e-06 
+ as=9.24e-12 ad=1.744e-11 ps=1.13e-05 pd=1.65e-05 
+ nrs=0.12 nrd=0.23 
m1664 0 891 890 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.744e-11 ad=9.24e-12 ps=1.65e-05 pd=1.13e-05 
+ nrs=0.23 nrd=0.12 
m1665 892 893 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=1.665e-11 ps=1.01e-05 pd=1.575e-05 
+ nrs=0.1 nrd=0.24 
m1666 894 895 892 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.89e-11 ad=7.14e-12 ps=2.29e-05 pd=1.01e-05 
+ nrs=0.27 nrd=0.1 
m1667 1 878 877 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=2.346e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.23 
m1668 878 879 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m1669 1 881 880 1 penh l=1.1e-06 w=9.6e-06 
+ as=2.137e-11 ad=2.256e-11 ps=1.812e-05 pd=2.29e-05 
+ nrs=0.23 nrd=0.24 
m1670 881 882 1 1 penh l=1.1e-06 w=9.6e-06 
+ as=2.256e-11 ad=2.137e-11 ps=2.29e-05 pd=1.812e-05 
+ nrs=0.24 nrd=0.23 
m1671 896 888 895 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.27e-12 ad=2.112e-11 ps=1.176e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.23 
m1672 897 889 896 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.31e-12 ps=1.25e-05 pd=1.324e-05 
+ nrs=0.08 nrd=0.08 
m1673 0 898 897 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m1674 899 886 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m1675 900 901 899 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.31e-12 ad=9.18e-12 ps=1.324e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m1676 893 902 900 0 nenh l=1.1e-06 w=9.6e-06 
+ as=2.112e-11 ad=8.27e-12 ps=2.53e-05 pd=1.176e-05 
+ nrs=0.23 nrd=0.09 
m1677 883 884 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.352e-11 ad=2.494e-11 ps=1.37e-05 pd=2.114e-05 
+ nrs=0.11 nrd=0.2 
m1678 1 884 883 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.352e-11 ps=2.114e-05 pd=1.37e-05 
+ nrs=0.2 nrd=0.11 
m1679 1 886 884 1 penh l=1.1e-06 w=9.6e-06 
+ as=2.137e-11 ad=1.315e-11 ps=1.812e-05 pd=1.587e-05 
+ nrs=0.23 nrd=0.14 
m1680 884 888 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.26e-11 ad=2.048e-11 ps=1.521e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m1681 1 889 884 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.26e-11 ps=1.737e-05 pd=1.521e-05 
+ nrs=0.24 nrd=0.15 
m1682 903 886 1 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.122e-11 ad=2.939e-11 ps=1.49e-05 pd=2.492e-05 
+ nrs=0.06 nrd=0.17 
m1683 890 891 903 1 penh l=1.1e-06 w=1.32e-05 
+ as=2.586e-11 ad=1.122e-11 ps=3.01e-05 pd=1.49e-05 
+ nrs=0.15 nrd=0.06 
m1684 894 893 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.466e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.07 nrd=0.15 
m1685 1 895 894 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.466e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.07 
m1686 1 888 895 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.297e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m1687 895 889 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.297e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m1688 1 898 895 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.297e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m1689 893 886 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m1690 1 901 893 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m1691 893 902 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m1692 882 904 1 1 penh l=1.1e-06 w=1e-05 
+ as=2.698e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.27 nrd=0.22 
m1693 904 905 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m1694 906 891 907 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.059e-11 ad=2.892e-11 ps=1.558e-05 pd=3.01e-05 
+ nrs=0.07 nrd=0.2 
m1695 1 898 906 1 penh l=1.1e-06 w=1.28e-05 
+ as=2.85e-11 ad=1.129e-11 ps=2.416e-05 pd=1.662e-05 
+ nrs=0.17 nrd=0.07 
m1696 908 902 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m1697 1 901 908 1 penh l=1.1e-06 w=8e-06 
+ as=1.781e-11 ad=1.075e-11 ps=1.51e-05 pd=1.383e-05 
+ nrs=0.28 nrd=0.17 
m1698 908 898 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m1699 909 908 1 1 penh l=1.1e-06 w=1e-05 
+ as=1.058e-11 ad=2.227e-11 ps=1.25e-05 pd=1.888e-05 
+ nrs=0.11 nrd=0.22 
m1700 1 908 909 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=1.058e-11 ps=1.888e-05 pd=1.25e-05 
+ nrs=0.22 nrd=0.11 
m1701 879 894 1 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=8.54e-12 ps=7.22e-06 pd=1.094e-05 
+ nrs=0.69 nrd=1.09 
m1702 879 883 910 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.88e-12 ps=7.22e-06 pd=1.048e-05 
+ nrs=0.69 nrd=1 
m1703 911 909 879 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m1704 879 890 911 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.91e-12 ps=7.22e-06 pd=1.05e-05 
+ nrs=0.69 nrd=1.01 
m1705 910 907 879 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m1706 0 894 905 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m1707 0 904 882 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.952e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.48 
m1708 0 905 904 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.26e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.4 
m1709 905 909 595 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=9.95e-12 ps=8.18e-06 pd=1.239e-05 
+ nrs=0.54 nrd=0.77 
m1710 602 883 905 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.045e-11 ad=6.95e-12 ps=1.269e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m1711 905 890 910 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.013e-11 ps=8.18e-06 pd=1.347e-05 
+ nrs=0.54 nrd=0.78 
m1712 911 907 905 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.016e-11 ad=6.95e-12 ps=1.35e-05 pd=8.18e-06 
+ nrs=0.78 nrd=0.54 
m1713 912 901 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=2.405e-11 ps=1.41e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m1714 891 902 912 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.046e-11 ad=1.014e-11 ps=1.25e-05 pd=1.41e-05 
+ nrs=0.09 nrd=0.09 
m1715 913 889 891 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=1.046e-11 ps=1.41e-05 pd=1.25e-05 
+ nrs=0.09 nrd=0.09 
m1716 1 888 913 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.014e-11 ps=2.039e-05 pd=1.41e-05 
+ nrs=0.21 nrd=0.09 
m1717 907 891 0 0 nenh l=1.1e-06 w=8e-06 
+ as=8.95e-12 ad=1.586e-11 ps=1.063e-05 pd=1.5e-05 
+ nrs=0.14 nrd=0.25 
m1718 0 898 907 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=9.39e-12 ps=1.575e-05 pd=1.117e-05 
+ nrs=0.24 nrd=0.13 
m1719 914 902 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m1720 915 901 914 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.4e-12 ad=9.18e-12 ps=1.378e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m1721 908 898 915 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.964e-11 ad=7.66e-12 ps=2.37e-05 pd=1.122e-05 
+ nrs=0.25 nrd=0.1 
m1722 909 908 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m1723 0 908 909 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m1724 916 901 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=1.024e-11 ad=2.141e-11 ps=1.384e-05 pd=2.024e-05 
+ nrs=0.09 nrd=0.18 
m1725 891 889 916 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.062e-11 ps=1.29e-05 pd=1.436e-05 
+ nrs=0.09 nrd=0.08 
m1726 917 902 891 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.062e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.08 nrd=0.09 
m1727 0 888 917 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.024e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m1728 918 919 1 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=8.54e-12 ps=6.1e-06 pd=1.094e-05 
+ nrs=0.59 nrd=1.09 
m1729 911 920 918 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=4.62e-12 ps=1.05e-05 pd=6.1e-06 
+ nrs=1.01 nrd=0.59 
m1730 918 921 911 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=7.91e-12 ps=6.1e-06 pd=1.05e-05 
+ nrs=0.59 nrd=1.01 
m1731 910 922 918 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=4.62e-12 ps=1.048e-05 pd=6.1e-06 
+ nrs=1 nrd=0.59 
m1732 0 924 923 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m1733 0 925 924 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m1734 925 919 0 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.46e-12 ad=7.14e-12 ps=1.01e-05 pd=6.75e-06 
+ nrs=0.65 nrd=0.55 
m1735 1 924 923 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=2.186e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.22 
m1736 925 920 595 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.46e-12 ad=9.95e-12 ps=1.01e-05 pd=1.239e-05 
+ nrs=0.65 nrd=0.77 
m1737 925 921 910 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.46e-12 ad=1.013e-11 ps=1.01e-05 pd=1.347e-05 
+ nrs=0.65 nrd=0.78 
m1738 911 922 925 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.016e-11 ad=8.46e-12 ps=1.35e-05 pd=1.01e-05 
+ nrs=0.78 nrd=0.65 
m1739 921 926 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=1.268e-11 ps=8.9e-06 pd=1.2e-05 
+ nrs=0.18 nrd=0.31 
m1740 0 926 921 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=7.2e-12 ps=1.2e-05 pd=8.9e-06 
+ nrs=0.31 nrd=0.18 
m1741 922 927 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=1.268e-11 ps=8.9e-06 pd=1.2e-05 
+ nrs=0.18 nrd=0.31 
m1742 0 927 922 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=7.2e-12 ps=1.2e-05 pd=8.9e-06 
+ nrs=0.31 nrd=0.18 
m1743 928 929 927 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.334e-11 ps=1.25e-05 pd=2.77e-05 
+ nrs=0.08 nrd=0.2 
m1744 0 902 928 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m1745 930 929 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m1746 926 889 930 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.67e-11 ad=9.18e-12 ps=2.77e-05 pd=1.25e-05 
+ nrs=0.23 nrd=0.08 
m1747 1 925 924 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.82e-11 ps=1.057e-05 pd=1.81e-05 
+ nrs=0.4 nrd=0.58 
m1748 921 926 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=9.9e-12 ad=2.048e-11 ps=1.17e-05 pd=1.737e-05 
+ nrs=0.12 nrd=0.24 
m1749 1 926 921 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=9.9e-12 ps=1.737e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.12 
m1750 922 927 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.452e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m1751 1 927 922 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.452e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m1752 927 929 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=9.58e-12 ad=2.048e-11 ps=1.17e-05 pd=1.737e-05 
+ nrs=0.11 nrd=0.24 
m1753 1 902 927 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=9.58e-12 ps=1.737e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.11 
m1754 926 929 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=9.58e-12 ad=2.048e-11 ps=1.17e-05 pd=1.737e-05 
+ nrs=0.11 nrd=0.24 
m1755 1 889 926 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=9.58e-12 ps=1.737e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.11 
m1756 1 932 931 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=2.522e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.25 
m1757 1 934 933 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1758 935 592 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m1759 936 933 935 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m1760 937 910 936 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m1761 1 596 937 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m1762 938 26 939 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.148e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.37 
m1763 940 25 938 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m1764 1 941 940 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m1765 941 939 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.37 nrd=0.4 
m1766 932 918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m1767 0 932 931 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.427e-11 ad=2.196e-11 ps=1.35e-05 pd=2.05e-05 
+ nrs=0.28 nrd=0.42 
m1768 932 918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m1769 939 25 602 0 nenh l=1.1e-06 w=3.2e-06 
+ as=1.294e-11 ad=9.28e-12 ps=1.146e-05 pd=1.128e-05 
+ nrs=1.26 nrd=0.91 
m1770 1 911 910 1 penh l=1.1e-06 w=2.2e-05 
+ as=4.898e-11 ad=5.176e-11 ps=4.153e-05 pd=4.391e-05 
+ nrs=0.1 nrd=0.11 
m1771 920 942 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=9.58e-12 ad=2.048e-11 ps=1.17e-05 pd=1.737e-05 
+ nrs=0.11 nrd=0.24 
m1772 1 942 920 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=9.58e-12 ps=1.737e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.11 
m1773 942 889 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=9.58e-12 ad=2.048e-11 ps=1.17e-05 pd=1.737e-05 
+ nrs=0.11 nrd=0.24 
m1774 1 943 942 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=9.58e-12 ps=1.737e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.11 
m1775 919 944 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=9.58e-12 ad=2.048e-11 ps=1.17e-05 pd=1.737e-05 
+ nrs=0.11 nrd=0.24 
m1776 1 944 919 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=9.58e-12 ps=1.737e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.11 
m1777 944 902 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=9.58e-12 ad=2.048e-11 ps=1.17e-05 pd=1.737e-05 
+ nrs=0.11 nrd=0.24 
m1778 1 943 944 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=9.58e-12 ps=1.737e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.11 
m1779 945 19 910 1 penh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=6.59e-12 ps=1.17e-05 pd=5.59e-06 
+ nrs=1.09 nrd=0.84 
m1780 911 945 1 1 penh l=1.1e-06 w=1.84e-05 
+ as=2.332e-11 ad=4.097e-11 ps=3.89e-05 pd=3.474e-05 
+ nrs=0.07 nrd=0.12 
m1781 946 19 939 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=1.132e-11 ps=4.5e-06 pd=1.003e-05 
+ nrs=0.3 nrd=1.44 
m1782 0 941 946 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m1783 0 934 933 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m1784 947 596 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1785 936 933 947 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m1786 948 910 936 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m1787 0 592 948 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1788 939 26 936 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.456e-11 ad=7.52e-12 ps=1.289e-05 pd=7.76e-06 
+ nrs=1.12 nrd=0.58 
m1789 941 939 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.12e-12 ad=1.11e-11 ps=9.23e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1790 945 19 941 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=8.46e-12 ps=1.65e-05 pd=8.57e-06 
+ nrs=0.41 nrd=0.31 
m1791 0 37 939 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.132e-11 ps=5.25e-06 pd=1.003e-05 
+ nrs=0.71 nrd=1.44 
m1792 920 942 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=1.11e-11 ps=8.9e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1793 0 942 920 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=9.24e-12 ps=1.05e-05 pd=8.9e-06 
+ nrs=0.35 nrd=0.29 
m1794 949 889 942 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.708e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.54 
m1795 0 943 949 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m1796 919 944 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=1.11e-11 ps=8.9e-06 pd=1.05e-05 
+ nrs=0.29 nrd=0.35 
m1797 0 944 919 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=9.24e-12 ps=1.05e-05 pd=8.9e-06 
+ nrs=0.35 nrd=0.29 
m1798 950 902 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m1799 944 943 950 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m1800 0 911 910 0 nenh l=1.1e-06 w=1.8e-05 
+ as=3.568e-11 ad=5.064e-11 ps=3.374e-05 pd=6.734e-05 
+ nrs=0.11 nrd=0.16 
m1801 911 945 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=4.517e-11 ad=3.171e-11 ps=6.002e-05 pd=2.999e-05 
+ nrs=0.18 nrd=0.12 
m1802 951 953 952 0 nenh l=1.1e-06 w=5.2e-06 
+ as=4.42e-12 ad=1.586e-11 ps=6.9e-06 pd=1.65e-05 
+ nrs=0.16 nrd=0.59 
m1803 0 954 951 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.031e-11 ad=4.42e-12 ps=9.75e-06 pd=6.9e-06 
+ nrs=0.38 nrd=0.16 
m1804 0 955 954 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m1805 956 953 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m1806 957 955 956 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m1807 958 954 957 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m1808 0 931 958 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m1809 953 931 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m1810 952 953 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.036e-11 ad=1.247e-11 ps=9.3e-06 pd=1.057e-05 
+ nrs=0.33 nrd=0.4 
m1811 1 954 952 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.036e-11 ps=1.057e-05 pd=9.3e-06 
+ nrs=0.4 nrd=0.33 
m1812 1 955 954 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.622e-11 ps=1.435e-05 pd=2.21e-05 
+ nrs=0.29 nrd=0.45 
m1813 959 953 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.362e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.09 nrd=0.19 
m1814 957 954 959 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.408e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.09 
m1815 960 955 957 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m1816 1 931 960 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m1817 953 931 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.55e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.27 nrd=0.29 
m1818 955 961 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.3e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.3 nrd=0.25 
m1819 961 962 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.26e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.4 nrd=0.4 
m1820 0 894 962 0 nenh l=1.1e-06 w=3.2e-06 
+ as=6.34e-12 ad=6.09e-12 ps=6e-06 pd=7.29e-06 
+ nrs=0.62 nrd=0.6 
m1821 0 961 955 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.952e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.48 
m1822 0 962 961 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.446e-11 ps=1.125e-05 pd=1.81e-05 
+ nrs=0.33 nrd=0.4 
m1823 962 909 612 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.003e-11 ps=8.2e-06 pd=1.202e-05 
+ nrs=0.53 nrd=0.77 
m1824 601 883 962 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.86e-12 ps=1.23e-05 pd=8.2e-06 
+ nrs=0.81 nrd=0.53 
m1825 962 907 602 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.045e-11 ps=8.2e-06 pd=1.269e-05 
+ nrs=0.53 nrd=0.81 
m1826 595 890 962 0 nenh l=1.1e-06 w=3.6e-06 
+ as=9.95e-12 ad=6.86e-12 ps=1.239e-05 pd=8.2e-06 
+ nrs=0.77 nrd=0.53 
m1827 963 964 0 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.298e-11 ad=1.031e-11 ps=1.65e-05 pd=9.75e-06 
+ nrs=0.48 nrd=0.38 
m1828 0 965 964 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.574e-11 ps=1.125e-05 pd=1.81e-05 
+ nrs=0.33 nrd=0.44 
m1829 965 919 0 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.46e-12 ad=7.14e-12 ps=1.01e-05 pd=6.75e-06 
+ nrs=0.65 nrd=0.55 
m1830 1 964 963 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m1831 965 920 612 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.46e-12 ad=1.003e-11 ps=1.01e-05 pd=1.202e-05 
+ nrs=0.65 nrd=0.77 
m1832 965 922 602 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.46e-12 ad=1.045e-11 ps=1.01e-05 pd=1.269e-05 
+ nrs=0.65 nrd=0.81 
m1833 595 921 965 0 nenh l=1.1e-06 w=3.6e-06 
+ as=9.95e-12 ad=8.46e-12 ps=1.239e-05 pd=1.01e-05 
+ nrs=0.77 nrd=0.65 
m1834 1 965 964 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1835 966 967 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m1836 0 968 966 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m1837 0 969 968 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m1838 970 967 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m1839 971 968 970 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m1840 972 969 971 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m1841 0 923 972 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m1842 967 923 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m1843 973 967 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m1844 966 968 973 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m1845 1 969 968 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m1846 974 967 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m1847 971 969 974 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m1848 975 968 971 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m1849 1 923 975 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m1850 967 923 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m1851 969 976 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m1852 976 977 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m1853 0 894 977 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m1854 0 976 969 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m1855 0 977 976 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m1856 977 909 627 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m1857 617 883 977 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m1858 977 907 601 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m1859 612 890 977 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m1860 978 979 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m1861 0 980 979 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m1862 980 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m1863 980 920 627 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m1864 980 922 601 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m1865 612 921 980 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m1866 1 979 978 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m1867 1 980 979 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1868 981 982 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m1869 0 983 981 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m1870 0 984 983 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m1871 985 982 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m1872 986 983 985 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m1873 987 984 986 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m1874 0 963 987 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m1875 982 963 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m1876 988 982 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m1877 981 983 988 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m1878 1 984 983 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m1879 989 982 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m1880 986 984 989 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m1881 990 983 986 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m1882 1 963 990 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m1883 982 963 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m1884 984 991 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m1885 991 992 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m1886 0 894 992 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m1887 0 991 984 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m1888 0 992 991 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m1889 992 909 642 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m1890 632 883 992 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m1891 992 907 617 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m1892 627 890 992 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m1893 993 994 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m1894 0 995 994 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m1895 995 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m1896 995 920 642 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m1897 995 922 617 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m1898 627 921 995 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m1899 1 994 993 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m1900 1 995 994 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1901 996 997 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m1902 0 998 996 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m1903 0 999 998 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m1904 1000 997 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m1905 1001 998 1000 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m1906 1002 999 1001 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m1907 0 978 1002 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m1908 997 978 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m1909 1003 997 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m1910 996 998 1003 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m1911 1 999 998 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m1912 1004 997 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m1913 1001 999 1004 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m1914 1005 998 1001 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m1915 1 978 1005 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m1916 997 978 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m1917 999 1006 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m1918 1006 1007 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m1919 0 894 1007 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m1920 0 1006 999 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m1921 0 1007 1006 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m1922 1007 909 657 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m1923 647 883 1007 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m1924 1007 907 632 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m1925 642 890 1007 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m1926 1008 1009 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m1927 0 1010 1009 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m1928 1010 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m1929 1010 920 657 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m1930 1010 922 632 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m1931 642 921 1010 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m1932 1 1009 1008 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m1933 1 1010 1009 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1934 1011 1012 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m1935 0 1013 1011 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m1936 0 1014 1013 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m1937 1015 1012 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m1938 1016 1013 1015 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m1939 1017 1014 1016 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m1940 0 993 1017 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m1941 1012 993 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m1942 1018 1012 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m1943 1011 1013 1018 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m1944 1 1014 1013 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m1945 1019 1012 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m1946 1016 1014 1019 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m1947 1020 1013 1016 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m1948 1 993 1020 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m1949 1012 993 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m1950 1014 1021 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m1951 1021 1022 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m1952 0 894 1022 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m1953 0 1021 1014 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m1954 0 1022 1021 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m1955 1022 909 672 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m1956 662 883 1022 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m1957 1022 907 647 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m1958 657 890 1022 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m1959 1023 1024 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m1960 0 1025 1024 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m1961 1025 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m1962 1025 920 672 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m1963 1025 922 647 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m1964 657 921 1025 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m1965 1 1024 1023 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m1966 1 1025 1024 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m1967 1026 1027 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m1968 0 1028 1026 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m1969 0 1029 1028 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m1970 1030 1027 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m1971 1031 1028 1030 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m1972 1032 1029 1031 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m1973 0 1008 1032 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m1974 1027 1008 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m1975 1033 1027 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m1976 1026 1028 1033 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m1977 1 1029 1028 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m1978 1034 1027 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m1979 1031 1029 1034 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m1980 1035 1028 1031 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m1981 1 1008 1035 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m1982 1027 1008 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m1983 1029 1036 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m1984 1036 1037 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m1985 0 894 1037 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m1986 0 1036 1029 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m1987 0 1037 1036 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m1988 1037 909 687 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m1989 677 883 1037 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m1990 1037 907 662 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m1991 672 890 1037 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m1992 1038 1039 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m1993 0 1040 1039 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m1994 1040 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m1995 1040 920 687 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m1996 1040 922 662 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m1997 672 921 1040 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m1998 1 1039 1038 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m1999 1 1040 1039 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2000 1041 1042 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m2001 0 1043 1041 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m2002 0 1044 1043 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m2003 1045 1042 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m2004 1046 1043 1045 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m2005 1047 1044 1046 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m2006 0 1023 1047 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m2007 1042 1023 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m2008 1048 1042 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2009 1041 1043 1048 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m2010 1 1044 1043 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m2011 1049 1042 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m2012 1046 1044 1049 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m2013 1050 1043 1046 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m2014 1 1023 1050 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m2015 1042 1023 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m2016 1044 1051 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2017 1051 1052 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2018 0 894 1052 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m2019 0 1051 1044 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m2020 0 1052 1051 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2021 1052 909 702 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m2022 692 883 1052 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m2023 1052 907 677 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m2024 687 890 1052 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m2025 1053 1054 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m2026 0 1055 1054 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m2027 1055 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m2028 1055 920 702 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m2029 1055 922 677 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m2030 687 921 1055 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m2031 1 1054 1053 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m2032 1 1055 1054 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2033 1056 1057 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m2034 0 1058 1056 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m2035 0 1059 1058 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m2036 1060 1057 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m2037 1061 1058 1060 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m2038 1062 1059 1061 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m2039 0 1038 1062 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m2040 1057 1038 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m2041 1063 1057 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2042 1056 1058 1063 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m2043 1 1059 1058 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m2044 1064 1057 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m2045 1061 1059 1064 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m2046 1065 1058 1061 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m2047 1 1038 1065 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m2048 1057 1038 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m2049 1059 1066 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2050 1066 1067 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2051 0 894 1067 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m2052 0 1066 1059 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m2053 0 1067 1066 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2054 1067 909 717 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m2055 707 883 1067 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m2056 1067 907 692 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m2057 702 890 1067 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m2058 1068 1069 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m2059 0 1070 1069 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m2060 1070 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m2061 1070 920 717 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m2062 1070 922 692 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m2063 702 921 1070 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m2064 1 1069 1068 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m2065 1 1070 1069 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2066 1071 1072 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m2067 0 1073 1071 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m2068 0 1074 1073 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m2069 1075 1072 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m2070 1076 1073 1075 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m2071 1077 1074 1076 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m2072 0 1053 1077 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m2073 1072 1053 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m2074 1078 1072 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2075 1071 1073 1078 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m2076 1 1074 1073 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m2077 1079 1072 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m2078 1076 1074 1079 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m2079 1080 1073 1076 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m2080 1 1053 1080 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m2081 1072 1053 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m2082 1074 1081 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2083 1081 1082 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2084 0 894 1082 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m2085 0 1081 1074 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m2086 0 1082 1081 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2087 1082 909 732 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m2088 722 883 1082 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m2089 1082 907 707 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m2090 717 890 1082 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m2091 1083 1084 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m2092 0 1085 1084 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m2093 1085 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m2094 1085 920 732 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m2095 1085 922 707 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m2096 717 921 1085 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m2097 1 1084 1083 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m2098 1 1085 1084 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2099 1086 1087 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m2100 0 1088 1086 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m2101 0 1089 1088 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m2102 1090 1087 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m2103 1091 1088 1090 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m2104 1092 1089 1091 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m2105 0 1068 1092 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m2106 1087 1068 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m2107 1093 1087 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2108 1086 1088 1093 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m2109 1 1089 1088 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m2110 1094 1087 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m2111 1091 1089 1094 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m2112 1095 1088 1091 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m2113 1 1068 1095 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m2114 1087 1068 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m2115 1089 1096 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2116 1096 1097 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2117 0 894 1097 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m2118 0 1096 1089 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m2119 0 1097 1096 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2120 1097 909 747 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m2121 737 883 1097 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m2122 1097 907 722 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m2123 732 890 1097 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m2124 1098 1099 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m2125 0 1100 1099 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m2126 1100 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m2127 1100 920 747 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m2128 1100 922 722 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m2129 732 921 1100 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m2130 1 1099 1098 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m2131 1 1100 1099 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2132 1101 1102 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m2133 0 1103 1101 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m2134 0 1104 1103 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m2135 1105 1102 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m2136 1106 1103 1105 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m2137 1107 1104 1106 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m2138 0 1083 1107 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m2139 1102 1083 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m2140 1108 1102 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2141 1101 1103 1108 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m2142 1 1104 1103 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m2143 1109 1102 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m2144 1106 1104 1109 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m2145 1110 1103 1106 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m2146 1 1083 1110 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m2147 1102 1083 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m2148 1104 1111 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2149 1111 1112 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2150 0 894 1112 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m2151 0 1111 1104 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m2152 0 1112 1111 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2153 1112 909 762 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m2154 752 883 1112 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m2155 1112 907 737 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m2156 747 890 1112 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m2157 1113 1114 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m2158 0 1115 1114 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m2159 1115 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m2160 1115 920 762 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m2161 1115 922 737 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m2162 747 921 1115 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m2163 1 1114 1113 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m2164 1 1115 1114 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2165 1116 1117 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m2166 0 1118 1116 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m2167 0 1119 1118 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m2168 1120 1117 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m2169 1121 1118 1120 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m2170 1122 1119 1121 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m2171 0 1098 1122 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m2172 1117 1098 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m2173 1123 1117 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2174 1116 1118 1123 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m2175 1 1119 1118 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m2176 1124 1117 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m2177 1121 1119 1124 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m2178 1125 1118 1121 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m2179 1 1098 1125 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m2180 1117 1098 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m2181 1119 1126 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2182 1126 1127 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2183 0 894 1127 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m2184 0 1126 1119 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m2185 0 1127 1126 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2186 1127 909 777 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m2187 767 883 1127 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m2188 1127 907 752 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m2189 762 890 1127 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m2190 1128 1129 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m2191 0 1130 1129 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m2192 1130 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m2193 1130 920 777 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m2194 1130 922 752 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m2195 762 921 1130 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m2196 1 1129 1128 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m2197 1 1130 1129 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2198 1131 1132 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m2199 0 1133 1131 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m2200 0 1134 1133 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m2201 1135 1132 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m2202 1136 1133 1135 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m2203 1137 1134 1136 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m2204 0 1113 1137 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m2205 1132 1113 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m2206 1138 1132 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2207 1131 1133 1138 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m2208 1 1134 1133 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m2209 1139 1132 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m2210 1136 1134 1139 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m2211 1140 1133 1136 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m2212 1 1113 1140 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m2213 1132 1113 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m2214 1134 1141 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2215 1141 1142 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2216 0 894 1142 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m2217 0 1141 1134 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m2218 0 1142 1141 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2219 1142 909 792 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m2220 782 883 1142 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m2221 1142 907 767 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m2222 777 890 1142 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m2223 1143 1144 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m2224 0 1145 1144 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m2225 1145 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m2226 1145 920 792 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m2227 1145 922 767 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m2228 777 921 1145 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m2229 1 1144 1143 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m2230 1 1145 1144 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2231 1146 1147 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m2232 0 1148 1146 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m2233 0 1149 1148 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m2234 1150 1147 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m2235 1151 1148 1150 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m2236 1152 1149 1151 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m2237 0 1128 1152 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m2238 1147 1128 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m2239 1153 1147 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2240 1146 1148 1153 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m2241 1 1149 1148 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m2242 1154 1147 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m2243 1151 1149 1154 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m2244 1155 1148 1151 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m2245 1 1128 1155 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m2246 1147 1128 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m2247 1149 1156 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2248 1156 1157 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2249 0 894 1157 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m2250 0 1156 1149 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m2251 0 1157 1156 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2252 1157 909 807 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m2253 797 883 1157 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m2254 1157 907 782 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m2255 792 890 1157 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m2256 1158 1159 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m2257 0 1160 1159 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m2258 1160 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m2259 1160 920 807 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m2260 1160 922 782 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m2261 792 921 1160 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m2262 1 1159 1158 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m2263 1 1160 1159 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2264 1161 1162 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m2265 0 1163 1161 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m2266 0 1164 1163 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m2267 1165 1162 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m2268 1166 1163 1165 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m2269 1167 1164 1166 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m2270 0 1143 1167 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m2271 1162 1143 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m2272 1168 1162 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2273 1161 1163 1168 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m2274 1 1164 1163 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m2275 1169 1162 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m2276 1166 1164 1169 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m2277 1170 1163 1166 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m2278 1 1143 1170 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m2279 1162 1143 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m2280 1164 1171 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2281 1171 1172 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2282 0 894 1172 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m2283 0 1171 1164 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m2284 0 1172 1171 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2285 1172 909 822 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m2286 812 883 1172 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m2287 1172 907 797 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m2288 807 890 1172 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m2289 1173 1174 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m2290 0 1175 1174 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m2291 1175 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m2292 1175 920 822 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m2293 1175 922 797 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m2294 807 921 1175 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m2295 1 1174 1173 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m2296 1 1175 1174 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2297 1176 1177 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m2298 0 1178 1176 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m2299 0 1179 1178 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m2300 1180 1177 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m2301 1181 1178 1180 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m2302 1182 1179 1181 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m2303 0 1158 1182 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m2304 1177 1158 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m2305 1183 1177 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2306 1176 1178 1183 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m2307 1 1179 1178 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m2308 1184 1177 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m2309 1181 1179 1184 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m2310 1185 1178 1181 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m2311 1 1158 1185 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m2312 1177 1158 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m2313 1179 1186 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2314 1186 1187 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2315 0 894 1187 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m2316 0 1186 1179 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m2317 0 1187 1186 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2318 1187 909 837 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m2319 827 883 1187 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m2320 1187 907 812 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m2321 822 890 1187 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m2322 1188 1189 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m2323 0 1190 1189 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m2324 1190 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m2325 1190 920 837 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m2326 1190 922 812 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m2327 822 921 1190 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m2328 1 1189 1188 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m2329 1 1190 1189 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2330 1191 1192 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m2331 0 1193 1191 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m2332 0 1194 1193 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m2333 1195 1192 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m2334 1196 1193 1195 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m2335 1197 1194 1196 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m2336 0 1173 1197 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m2337 1192 1173 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m2338 1198 1192 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2339 1191 1193 1198 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m2340 1 1194 1193 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m2341 1199 1192 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m2342 1196 1194 1199 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m2343 1200 1193 1196 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m2344 1 1173 1200 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m2345 1192 1173 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m2346 1194 1201 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2347 1201 1202 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2348 0 894 1202 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m2349 0 1201 1194 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m2350 0 1202 1201 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2351 1202 909 868 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m2352 842 883 1202 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.76e-12 ps=1.23e-05 pd=8.23e-06 
+ nrs=0.81 nrd=0.52 
m2353 1202 907 827 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m2354 837 890 1202 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m2355 1203 1204 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m2356 0 1205 1204 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m2357 1205 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m2358 1205 920 868 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m2359 1205 922 827 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m2360 837 921 1205 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m2361 1 1204 1203 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m2362 1 1205 1204 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2363 1206 1207 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m2364 0 1208 1206 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m2365 0 1209 1208 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m2366 1210 1207 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m2367 1211 1208 1210 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m2368 1212 1209 1211 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m2369 0 1188 1212 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m2370 1207 1188 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m2371 1213 1207 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2372 1206 1208 1213 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m2373 1 1209 1208 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=2.158e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.37 
m2374 1214 1207 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.173e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.08 nrd=0.19 
m2375 1211 1209 1214 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.213e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.08 
m2376 1215 1208 1211 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m2377 1 1188 1215 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m2378 1207 1188 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.742e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.3 nrd=0.29 
m2379 1209 1216 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2380 1216 1217 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2381 0 894 1217 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m2382 0 1216 1209 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m2383 0 1217 1216 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2384 1217 909 852 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.003e-11 ps=8.23e-06 pd=1.202e-05 
+ nrs=0.52 nrd=0.77 
m2385 858 883 1217 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.036e-11 ad=6.76e-12 ps=1.246e-05 pd=8.23e-06 
+ nrs=0.8 nrd=0.52 
m2386 1217 907 842 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.048e-11 ps=8.23e-06 pd=1.23e-05 
+ nrs=0.52 nrd=0.81 
m2387 868 890 1217 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m2388 1218 1219 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m2389 0 1220 1219 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.664e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.41 
m2390 1220 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m2391 1220 920 852 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.003e-11 ps=1.027e-05 pd=1.202e-05 
+ nrs=0.64 nrd=0.77 
m2392 1220 922 842 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.048e-11 ps=1.027e-05 pd=1.23e-05 
+ nrs=0.64 nrd=0.81 
m2393 868 921 1220 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m2394 1 1219 1218 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.3e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.3 
m2395 1 1220 1219 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2396 1221 1222 0 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=1.189e-11 ps=8.5e-06 pd=1.125e-05 
+ nrs=0.19 nrd=0.33 
m2397 0 1223 1221 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=6.86e-12 ps=1.125e-05 pd=8.5e-06 
+ nrs=0.33 nrd=0.19 
m2398 0 1224 1223 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.076e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.67 
m2399 1225 1222 0 0 nenh l=1.1e-06 w=1.2e-05 
+ as=1.243e-11 ad=2.378e-11 ps=1.583e-05 pd=2.249e-05 
+ nrs=0.09 nrd=0.17 
m2400 1226 1223 1225 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.161e-11 ps=1.29e-05 pd=1.477e-05 
+ nrs=0.09 nrd=0.09 
m2401 1227 1224 1226 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.111e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.09 nrd=0.09 
m2402 0 1203 1227 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.071e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m2403 1222 1203 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.076e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.67 nrd=0.5 
m2404 1228 1222 1221 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.708e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.54 
m2405 1 1223 1228 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m2406 1 1224 1223 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=1.998e-11 ps=1.435e-05 pd=2.13e-05 
+ nrs=0.29 nrd=0.35 
m2407 1229 1222 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.362e-11 ad=2.672e-11 ps=1.505e-05 pd=2.265e-05 
+ nrs=0.09 nrd=0.19 
m2408 1226 1224 1229 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.182e-11 ad=1.408e-11 ps=1.41e-05 pd=1.555e-05 
+ nrs=0.08 nrd=0.09 
m2409 1230 1223 1226 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.208e-11 ad=1.182e-11 ps=1.507e-05 pd=1.41e-05 
+ nrs=0.08 nrd=0.08 
m2410 1 1203 1230 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.052e-11 ps=2.039e-05 pd=1.313e-05 
+ nrs=0.21 nrd=0.09 
m2411 1222 1203 1 1 penh l=1.1e-06 w=7.6e-06 
+ as=2.078e-11 ad=1.692e-11 ps=2.13e-05 pd=1.435e-05 
+ nrs=0.36 nrd=0.29 
m2412 1 1232 1231 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2413 1233 909 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2414 1232 890 1233 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.148e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m2415 1 1234 1224 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=2.444e-11 ps=1.661e-05 pd=2.37e-05 
+ nrs=0.25 nrd=0.32 
m2416 1234 1235 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.202e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.44 nrd=0.43 
m2417 0 1232 1231 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m2418 1232 909 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=5.55e-12 ps=6.1e-06 pd=5.25e-06 
+ nrs=0.59 nrd=0.71 
m2419 0 890 1232 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=4.62e-12 ps=5.25e-06 pd=6.1e-06 
+ nrs=0.71 nrd=0.59 
m2420 0 894 1235 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.26e-12 ps=5.25e-06 pd=6.4e-06 
+ nrs=0.71 nrd=0.67 
m2421 0 1234 1224 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.792e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.44 
m2422 0 1235 1234 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.446e-11 ps=1.125e-05 pd=1.81e-05 
+ nrs=0.33 nrd=0.4 
m2423 1235 909 1 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.098e-11 ps=8.23e-06 pd=1.406e-05 
+ nrs=0.52 nrd=0.85 
m2424 0 883 1235 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.76e-12 ps=6.75e-06 pd=8.23e-06 
+ nrs=0.55 nrd=0.52 
m2425 1235 907 858 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.76e-12 ad=1.036e-11 ps=8.23e-06 pd=1.246e-05 
+ nrs=0.52 nrd=0.8 
m2426 852 890 1235 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.76e-12 ps=1.202e-05 pd=8.23e-06 
+ nrs=0.77 nrd=0.52 
m2427 1236 1237 0 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.952e-11 ad=1.268e-11 ps=1.89e-05 pd=1.2e-05 
+ nrs=0.48 nrd=0.31 
m2428 0 1238 1237 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.574e-11 ps=1.125e-05 pd=1.81e-05 
+ nrs=0.33 nrd=0.44 
m2429 1238 919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.46e-12 ad=5.55e-12 ps=7.99e-06 pd=5.25e-06 
+ nrs=0.82 nrd=0.71 
m2430 1238 920 1 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.098e-11 ps=1.027e-05 pd=1.406e-05 
+ nrs=0.64 nrd=0.85 
m2431 1238 922 858 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.31e-12 ad=1.036e-11 ps=1.027e-05 pd=1.246e-05 
+ nrs=0.64 nrd=0.8 
m2432 852 921 1238 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=8.31e-12 ps=1.202e-05 pd=1.027e-05 
+ nrs=0.77 nrd=0.64 
m2433 0 1240 1239 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=1.078e-11 ps=5.25e-06 pd=1.33e-05 
+ nrs=0.71 nrd=1.38 
m2434 1240 920 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=5.55e-12 ps=6.1e-06 pd=5.25e-06 
+ nrs=0.59 nrd=0.71 
m2435 0 921 1240 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=4.62e-12 ps=5.25e-06 pd=6.1e-06 
+ nrs=0.71 nrd=0.59 
m2436 1 1240 1239 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2437 1241 920 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2438 1240 921 1241 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.372e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.44 nrd=0.15 
m2439 1 1237 1236 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=1.914e-11 ps=1.284e-05 pd=1.97e-05 
+ nrs=0.33 nrd=0.41 
m2440 1237 1238 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.106e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.41 nrd=0.43 
m2441 0 1243 1242 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m2442 1244 1245 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m2443 1246 1242 1244 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m2444 1247 1243 1246 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m2445 0 1248 1247 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m2446 1245 1248 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m2447 0 1246 120 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m2448 1 1246 120 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.562e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m2449 1249 1251 1250 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.57e-11 ps=1.429e-05 pd=2.04e-05 
+ nrs=0.11 nrd=0.12 
m2450 1252 1253 1249 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m2451 1250 1254 1252 0 nenh l=1.1e-06 w=1e-05 
+ as=1.354e-11 ad=8.5e-12 ps=1.759e-05 pd=1.17e-05 
+ nrs=0.14 nrd=0.08 
m2452 0 1254 1250 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m2453 1250 1253 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m2454 0 1253 1255 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m2455 1255 1254 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m2456 1256 1254 1255 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.354e-11 ps=1.17e-05 pd=1.759e-05 
+ nrs=0.08 nrd=0.14 
m2457 1257 1253 1256 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m2458 0 1211 1254 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2459 1258 1254 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m2460 1248 1253 1258 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m2461 1259 1221 1248 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m2462 0 1211 1259 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m2463 1253 1221 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.372e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.44 nrd=0.35 
m2464 1255 1243 1257 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=1.416e-11 ps=2.04e-05 pd=1.429e-05 
+ nrs=0.12 nrd=0.11 
m2465 1 1243 1242 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m2466 1260 1245 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m2467 1246 1243 1260 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m2468 1261 1242 1246 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m2469 1 1248 1261 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m2470 1245 1248 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m2471 1249 1251 1262 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m2472 1263 1253 1249 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m2473 1 1254 1263 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m2474 1262 1254 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m2475 1 1253 1262 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m2476 1264 1253 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m2477 1 1254 1264 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m2478 1265 1254 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m2479 1257 1253 1265 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m2480 1264 1243 1257 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m2481 1 1211 1254 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=2.186e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.22 
m2482 1266 1254 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.45e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m2483 1248 1221 1266 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.033e-11 ad=7.53e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.11 
m2484 1267 1253 1248 1 penh l=1.1e-06 w=7.6e-06 
+ as=6.58e-12 ad=9.35e-12 ps=9.55e-06 pd=9.97e-06 
+ nrs=0.11 nrd=0.16 
m2485 1 1211 1267 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.24e-12 ps=1.359e-05 pd=9.05e-06 
+ nrs=0.31 nrd=0.12 
m2486 1253 1221 1 1 penh l=1.1e-06 w=1e-05 
+ as=2.522e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.25 nrd=0.22 
m2487 1 1268 91 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.562e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m2488 1 1270 1269 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m2489 1271 1272 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m2490 1273 1270 1271 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m2491 1274 1269 1273 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m2492 1 1275 1274 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m2493 1272 1275 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m2494 1268 1273 1 1 penh l=1.1e-06 w=8.4e-06 
+ as=2.562e-11 ad=1.87e-11 ps=2.29e-05 pd=1.586e-05 
+ nrs=0.36 nrd=0.27 
m2495 0 1268 91 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m2496 1268 1273 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m2497 1 1226 1276 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=2.334e-11 ps=2.039e-05 pd=2.77e-05 
+ nrs=0.21 nrd=0.2 
m2498 1277 1278 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=7.69e-12 ad=1.959e-11 ps=1.17e-05 pd=1.661e-05 
+ nrs=0.1 nrd=0.25 
m2499 1275 1226 1277 1 penh l=1.1e-06 w=7.6e-06 
+ as=9.65e-12 ad=6.65e-12 ps=9.97e-06 pd=1.01e-05 
+ nrs=0.17 nrd=0.12 
m2500 1279 1276 1275 1 penh l=1.1e-06 w=8.4e-06 
+ as=7.41e-12 ad=1.067e-11 ps=1.143e-05 pd=1.103e-05 
+ nrs=0.11 nrd=0.15 
m2501 1 1231 1279 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=7.77e-12 ps=1.661e-05 pd=1.197e-05 
+ nrs=0.25 nrd=0.1 
m2502 1278 1231 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.334e-11 ad=2.405e-11 ps=2.77e-05 pd=2.039e-05 
+ nrs=0.2 nrd=0.21 
m2503 1280 1281 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.55e-11 ad=2.672e-11 ps=1.478e-05 pd=2.265e-05 
+ nrs=0.11 nrd=0.19 
m2504 1251 1226 1280 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.151e-11 ad=1.498e-11 ps=1.394e-05 pd=1.428e-05 
+ nrs=0.09 nrd=0.11 
m2505 1280 1231 1251 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.705e-11 ad=1.309e-11 ps=1.625e-05 pd=1.586e-05 
+ nrs=0.1 nrd=0.08 
m2506 1282 1231 1280 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.498e-11 ps=1.33e-05 pd=1.428e-05 
+ nrs=0.07 nrd=0.11 
m2507 1 1226 1282 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m2508 1283 1226 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m2509 1284 1231 1283 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=9.86e-12 ps=1.428e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m2510 1243 1231 1284 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.309e-11 ad=1.705e-11 ps=1.586e-05 pd=1.625e-05 
+ nrs=0.08 nrd=0.1 
m2511 1284 1226 1243 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=1.151e-11 ps=1.428e-05 pd=1.394e-05 
+ nrs=0.11 nrd=0.09 
m2512 1 1270 1284 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.55e-11 ps=2.265e-05 pd=1.478e-05 
+ nrs=0.19 nrd=0.11 
m2513 0 1270 1269 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m2514 1285 1272 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m2515 1273 1269 1285 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m2516 1286 1270 1273 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m2517 0 1275 1286 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m2518 1272 1275 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m2519 0 1226 1276 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2520 1287 1278 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m2521 1275 1276 1287 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m2522 1288 1226 1275 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m2523 0 1231 1288 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m2524 1278 1231 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.372e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.44 nrd=0.35 
m2525 1251 1281 1289 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.175e-11 ad=1.755e-11 ps=1.429e-05 pd=1.841e-05 
+ nrs=0.09 nrd=0.13 
m2526 1290 1226 1251 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.013e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.1 
m2527 0 1231 1290 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=8.5e-12 ps=1.874e-05 pd=1.17e-05 
+ nrs=0.2 nrd=0.08 
m2528 1289 1231 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=2.299e-11 ps=1.841e-05 pd=2.174e-05 
+ nrs=0.13 nrd=0.17 
m2529 0 1226 1289 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=1.513e-11 ps=1.874e-05 pd=1.587e-05 
+ nrs=0.2 nrd=0.15 
m2530 1291 1226 0 0 nenh l=1.1e-06 w=1e-05 
+ as=1.513e-11 ad=1.982e-11 ps=1.587e-05 pd=1.874e-05 
+ nrs=0.15 nrd=0.2 
m2531 0 1231 1291 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.755e-11 ps=2.174e-05 pd=1.841e-05 
+ nrs=0.17 nrd=0.13 
m2532 1292 1231 0 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.982e-11 ps=1.17e-05 pd=1.874e-05 
+ nrs=0.08 nrd=0.2 
m2533 1243 1226 1292 0 nenh l=1.1e-06 w=1e-05 
+ as=1.013e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.1 nrd=0.08 
m2534 1291 1270 1243 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=1.175e-11 ps=1.841e-05 pd=1.429e-05 
+ nrs=0.13 nrd=0.09 
m2535 0 1293 62 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m2536 0 1295 1294 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m2537 1296 1297 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m2538 1293 1294 1296 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m2539 1298 1295 1293 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m2540 0 1218 1298 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m2541 1297 1218 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m2542 1281 1299 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=5.55e-12 ps=6.1e-06 pd=5.25e-06 
+ nrs=0.59 nrd=0.71 
m2543 0 1300 1281 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=4.62e-12 ps=5.25e-06 pd=6.1e-06 
+ nrs=0.71 nrd=0.59 
m2544 1270 1300 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=5.55e-12 ps=6.1e-06 pd=5.25e-06 
+ nrs=0.59 nrd=0.71 
m2545 0 1295 1270 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=4.62e-12 ps=5.25e-06 pd=6.1e-06 
+ nrs=0.71 nrd=0.59 
m2546 1300 1218 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m2547 1 1293 62 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2548 1 1295 1294 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2549 1301 1297 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m2550 1293 1295 1301 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m2551 1302 1294 1293 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m2552 1 1218 1302 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m2553 1297 1218 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2554 1303 1299 1281 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.708e-11 ps=7.3e-06 pd=1.73e-05 
+ nrs=0.15 nrd=0.54 
m2555 1 1300 1303 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.76e-12 ps=1.057e-05 pd=7.3e-06 
+ nrs=0.4 nrd=0.15 
m2556 1304 1300 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m2557 1270 1295 1304 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m2558 1 1218 1300 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2559 1 1305 31 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2560 1305 1306 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2561 1 1236 1307 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m2562 1308 1309 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m2563 1306 1236 1308 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m2564 1310 1307 1306 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m2565 1 1239 1310 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m2566 1309 1239 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2567 1311 1236 1299 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.122e-11 ad=3.114e-11 ps=1.49e-05 pd=3.25e-05 
+ nrs=0.06 nrd=0.18 
m2568 1 1239 1311 1 penh l=1.1e-06 w=1.32e-05 
+ as=2.939e-11 ad=1.122e-11 ps=2.492e-05 pd=1.49e-05 
+ nrs=0.17 nrd=0.06 
m2569 1295 1239 1 1 penh l=1.1e-06 w=1.28e-05 
+ as=1.488e-11 ad=2.85e-11 ps=1.53e-05 pd=2.416e-05 
+ nrs=0.09 nrd=0.17 
m2570 1 1236 1295 1 penh l=1.1e-06 w=1.28e-05 
+ as=2.85e-11 ad=1.488e-11 ps=2.416e-05 pd=1.53e-05 
+ nrs=0.17 nrd=0.09 
m2571 0 1305 31 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m2572 1305 1306 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m2573 0 1236 1307 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m2574 1312 1309 0 0 nenh l=1.1e-06 w=7.2e-06 
+ as=7.02e-12 ad=1.427e-11 ps=1.001e-05 pd=1.35e-05 
+ nrs=0.14 nrd=0.28 
m2575 1306 1307 1312 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=5.46e-12 ps=8.9e-06 pd=7.79e-06 
+ nrs=0.29 nrd=0.17 
m2576 1313 1236 1306 0 nenh l=1.1e-06 w=5.6e-06 
+ as=5.18e-12 ad=9.24e-12 ps=7.79e-06 pd=8.9e-06 
+ nrs=0.17 nrd=0.29 
m2577 0 1239 1313 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.427e-11 ad=6.66e-12 ps=1.35e-05 pd=1.001e-05 
+ nrs=0.28 nrd=0.13 
m2578 1309 1239 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m2579 592 596 1 1 penh l=1.1e-06 w=2.12e-05 
+ as=2.378e-11 ad=4.72e-11 ps=2.29e-05 pd=4.002e-05 
+ nrs=0.05 nrd=0.11 
m2580 1 596 592 1 penh l=1.1e-06 w=2.12e-05 
+ as=4.72e-11 ad=2.378e-11 ps=4.002e-05 pd=2.29e-05 
+ nrs=0.11 nrd=0.05 
m2581 1299 1236 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=1.284e-11 ad=2.061e-11 ps=1.29e-05 pd=1.949e-05 
+ nrs=0.12 nrd=0.19 
m2582 0 1239 1299 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.061e-11 ad=1.284e-11 ps=1.949e-05 pd=1.29e-05 
+ nrs=0.19 nrd=0.12 
m2583 1314 1239 1295 0 nenh l=1.1e-06 w=1.24e-05 
+ as=1.054e-11 ad=3.302e-11 ps=1.41e-05 pd=3.09e-05 
+ nrs=0.07 nrd=0.21 
m2584 0 1236 1314 0 nenh l=1.1e-06 w=1.24e-05 
+ as=2.458e-11 ad=1.054e-11 ps=2.324e-05 pd=1.41e-05 
+ nrs=0.16 nrd=0.07 
m2585 592 596 0 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.806e-11 ad=3.092e-11 ps=1.73e-05 pd=2.924e-05 
+ nrs=0.07 nrd=0.13 
m2586 0 596 592 0 nenh l=1.1e-06 w=1.56e-05 
+ as=3.092e-11 ad=1.806e-11 ps=2.924e-05 pd=1.73e-05 
+ nrs=0.13 nrd=0.07 
m2587 0 1316 1315 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.427e-11 ad=2.196e-11 ps=1.35e-05 pd=2.05e-05 
+ nrs=0.28 nrd=0.42 
m2588 1316 1317 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m2589 0 1319 1318 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.22e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.76 
m2590 1319 1320 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.22e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.76 nrd=0.5 
m2591 1 1316 1315 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m2592 1316 1317 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2593 1321 1322 0 0 nenh l=1.1e-06 w=4e-06 
+ as=6.6e-12 ad=7.93e-12 ps=7.3e-06 pd=7.5e-06 
+ nrs=0.41 nrd=0.5 
m2594 0 1322 1321 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=6.6e-12 ps=7.5e-06 pd=7.3e-06 
+ nrs=0.5 nrd=0.41 
m2595 1323 1324 1322 0 nenh l=1.1e-06 w=8.8e-06 
+ as=7.66e-12 ad=1.964e-11 ps=1.122e-05 pd=2.37e-05 
+ nrs=0.1 nrd=0.25 
m2596 1325 1326 1323 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.4e-12 ps=1.25e-05 pd=1.378e-05 
+ nrs=0.08 nrd=0.08 
m2597 0 898 1325 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m2598 1327 1324 0 0 nenh l=1.1e-06 w=8.8e-06 
+ as=9.24e-12 ad=1.744e-11 ps=1.13e-05 pd=1.65e-05 
+ nrs=0.12 nrd=0.23 
m2599 0 1328 1327 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.744e-11 ad=9.24e-12 ps=1.65e-05 pd=1.13e-05 
+ nrs=0.23 nrd=0.12 
m2600 1329 1330 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=1.665e-11 ps=1.01e-05 pd=1.575e-05 
+ nrs=0.1 nrd=0.24 
m2601 1331 1332 1329 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.89e-11 ad=7.14e-12 ps=2.29e-05 pd=1.01e-05 
+ nrs=0.27 nrd=0.1 
m2602 1 1319 1318 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=2.358e-11 ps=1.737e-05 pd=2.29e-05 
+ nrs=0.24 nrd=0.28 
m2603 1319 1320 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.358e-11 ad=2.048e-11 ps=2.29e-05 pd=1.737e-05 
+ nrs=0.28 nrd=0.24 
m2604 1321 1322 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.128e-11 ad=2.494e-11 ps=1.37e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m2605 1 1322 1321 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.128e-11 ps=2.114e-05 pd=1.37e-05 
+ nrs=0.2 nrd=0.09 
m2606 1333 1326 1332 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.27e-12 ad=2.16e-11 ps=1.176e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.23 
m2607 1334 898 1333 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.31e-12 ps=1.25e-05 pd=1.324e-05 
+ nrs=0.08 nrd=0.08 
m2608 0 1335 1334 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m2609 1336 1324 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m2610 1337 1338 1336 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.31e-12 ad=9.18e-12 ps=1.324e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m2611 1330 886 1337 0 nenh l=1.1e-06 w=9.6e-06 
+ as=2.16e-11 ad=8.27e-12 ps=2.53e-05 pd=1.176e-05 
+ nrs=0.23 nrd=0.09 
m2612 1 1324 1322 1 penh l=1.1e-06 w=9.6e-06 
+ as=2.137e-11 ad=1.315e-11 ps=1.812e-05 pd=1.587e-05 
+ nrs=0.23 nrd=0.14 
m2613 1322 1326 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.26e-11 ad=2.048e-11 ps=1.521e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m2614 1 898 1322 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.26e-11 ps=1.737e-05 pd=1.521e-05 
+ nrs=0.24 nrd=0.15 
m2615 1339 1324 1 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.194e-11 ad=2.939e-11 ps=1.49e-05 pd=2.492e-05 
+ nrs=0.07 nrd=0.17 
m2616 1327 1328 1339 1 penh l=1.1e-06 w=1.32e-05 
+ as=2.586e-11 ad=1.194e-11 ps=3.01e-05 pd=1.49e-05 
+ nrs=0.15 nrd=0.07 
m2617 1331 1330 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.466e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.07 nrd=0.15 
m2618 1 1332 1331 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.466e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.07 
m2619 1 1326 1332 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m2620 1332 898 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m2621 1 1335 1332 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m2622 1330 1324 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m2623 1 1338 1330 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m2624 1330 886 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m2625 1320 1340 1 1 penh l=1.1e-06 w=1e-05 
+ as=2.346e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.23 nrd=0.22 
m2626 1340 1341 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2627 1317 1331 1 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=8.54e-12 ps=7.22e-06 pd=1.094e-05 
+ nrs=0.69 nrd=1.09 
m2628 910 1321 1317 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m2629 1342 1328 1343 1 penh l=1.1e-06 w=1.04e-05 
+ as=8.84e-12 ad=2.596e-11 ps=1.21e-05 pd=2.69e-05 
+ nrs=0.08 nrd=0.24 
m2630 1 1335 1342 1 penh l=1.1e-06 w=1.04e-05 
+ as=2.316e-11 ad=8.84e-12 ps=1.963e-05 pd=1.21e-05 
+ nrs=0.21 nrd=0.08 
m2631 1344 886 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m2632 1 1338 1344 1 penh l=1.1e-06 w=8e-06 
+ as=1.781e-11 ad=1.075e-11 ps=1.51e-05 pd=1.383e-05 
+ nrs=0.28 nrd=0.17 
m2633 1344 1335 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m2634 1345 1344 1 1 penh l=1.1e-06 w=1e-05 
+ as=1.058e-11 ad=2.227e-11 ps=1.25e-05 pd=1.888e-05 
+ nrs=0.11 nrd=0.22 
m2635 1 1344 1345 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=1.058e-11 ps=1.888e-05 pd=1.25e-05 
+ nrs=0.22 nrd=0.11 
m2636 1341 1345 595 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.74e-12 ps=7.22e-06 pd=9.64e-06 
+ nrs=0.69 nrd=0.99 
m2637 602 1321 1341 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=5.4e-12 ps=9.87e-06 pd=7.22e-06 
+ nrs=1.04 nrd=0.69 
m2638 1341 1327 910 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.88e-12 ps=7.22e-06 pd=1.048e-05 
+ nrs=0.69 nrd=1 
m2639 911 1343 1341 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m2640 0 1331 1341 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.4e-12 ps=5.25e-06 pd=7.22e-06 
+ nrs=0.71 nrd=0.69 
m2641 1346 1338 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=2.405e-11 ps=1.41e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m2642 1328 886 1346 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.046e-11 ad=1.014e-11 ps=1.25e-05 pd=1.41e-05 
+ nrs=0.09 nrd=0.09 
m2643 1347 898 1328 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=1.046e-11 ps=1.41e-05 pd=1.25e-05 
+ nrs=0.09 nrd=0.09 
m2644 1 1326 1347 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.014e-11 ps=2.039e-05 pd=1.41e-05 
+ nrs=0.21 nrd=0.09 
m2645 911 1345 1317 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m2646 1317 1327 911 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.91e-12 ps=7.22e-06 pd=1.05e-05 
+ nrs=0.69 nrd=1.01 
m2647 910 1343 1317 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m2648 0 1340 1320 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m2649 0 1341 1340 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m2650 1343 1328 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m2651 0 1335 1343 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m2652 1348 886 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m2653 1349 1338 1348 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.4e-12 ad=9.18e-12 ps=1.378e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m2654 1344 1335 1349 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.964e-11 ad=7.66e-12 ps=2.37e-05 pd=1.122e-05 
+ nrs=0.25 nrd=0.1 
m2655 1345 1344 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m2656 0 1344 1345 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m2657 1350 1338 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=9.84e-12 ad=2.061e-11 ps=1.319e-05 pd=1.949e-05 
+ nrs=0.09 nrd=0.19 
m2658 1328 898 1350 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.06e-11 ps=1.29e-05 pd=1.421e-05 
+ nrs=0.09 nrd=0.08 
m2659 1351 886 1328 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.062e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.08 nrd=0.09 
m2660 0 1326 1351 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.024e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m2661 0 1353 1352 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m2662 1354 1355 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m2663 0 877 1354 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m2664 1356 1355 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m2665 1353 877 1356 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m2666 1354 880 1353 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m2667 1357 880 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m2668 1358 1353 1357 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m2669 1 1353 1352 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m2670 1359 877 1358 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m2671 1360 880 1359 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m2672 0 1355 1360 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m2673 1357 877 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m2674 0 1355 1357 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m2675 1361 1355 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m2676 1362 877 1361 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m2677 1353 1355 1362 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m2678 1362 877 1353 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m2679 1363 1358 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m2680 1 880 1362 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m2681 1358 1353 1364 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m2682 1365 877 1358 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m2683 1366 880 1365 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m2684 1355 1367 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2685 1367 1368 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2686 1364 1355 1366 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m2687 1 877 1364 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m2688 1364 1355 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m2689 1 880 1364 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m2690 1363 1358 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m2691 0 1367 1355 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m2692 0 1368 1367 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m2693 0 1331 1368 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m2694 1368 1345 612 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m2695 601 1321 1368 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m2696 1368 1343 602 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.045e-11 ps=8.18e-06 pd=1.269e-05 
+ nrs=0.54 nrd=0.81 
m2697 595 1327 1368 0 nenh l=1.1e-06 w=3.6e-06 
+ as=9.95e-12 ad=6.95e-12 ps=1.239e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m2698 0 1370 1369 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m2699 1371 1372 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m2700 0 881 1371 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m2701 1373 1372 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m2702 1370 881 1373 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m2703 1371 952 1370 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m2704 1374 952 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m2705 1375 1370 1374 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m2706 1 1370 1369 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m2707 1376 881 1375 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m2708 1377 952 1376 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m2709 0 1372 1377 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m2710 1374 881 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m2711 0 1372 1374 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m2712 1378 1372 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m2713 1379 881 1378 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m2714 1370 1372 1379 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m2715 1379 881 1370 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m2716 1380 1375 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m2717 1 952 1379 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m2718 1375 1370 1381 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m2719 1382 881 1375 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m2720 1383 952 1382 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m2721 1372 1384 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2722 1384 1385 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2723 1381 1372 1383 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m2724 1 881 1381 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m2725 1381 1372 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m2726 1 952 1381 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m2727 1380 1375 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m2728 0 1384 1372 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m2729 0 1385 1384 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m2730 0 1331 1385 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m2731 1385 1345 627 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m2732 617 1321 1385 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m2733 1385 1343 601 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m2734 612 1327 1385 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m2735 0 1387 1386 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m2736 1388 1389 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m2737 0 957 1388 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m2738 1390 1389 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m2739 1387 957 1390 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m2740 1388 966 1387 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m2741 1391 966 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m2742 1392 1387 1391 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m2743 1 1387 1386 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m2744 1393 957 1392 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m2745 1394 966 1393 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m2746 0 1389 1394 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m2747 1391 957 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m2748 0 1389 1391 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m2749 1395 1389 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m2750 1396 957 1395 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m2751 1387 1389 1396 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m2752 1396 957 1387 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m2753 1397 1392 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m2754 1 966 1396 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m2755 1392 1387 1398 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m2756 1399 957 1392 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m2757 1400 966 1399 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m2758 1389 1401 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2759 1401 1402 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2760 1398 1389 1400 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m2761 1 957 1398 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m2762 1398 1389 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m2763 1 966 1398 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m2764 1397 1392 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m2765 0 1401 1389 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m2766 0 1402 1401 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m2767 0 1331 1402 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m2768 1402 1345 642 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m2769 632 1321 1402 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m2770 1402 1343 617 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m2771 627 1327 1402 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m2772 0 1404 1403 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m2773 1405 1406 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m2774 0 971 1405 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m2775 1407 1406 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m2776 1404 971 1407 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m2777 1405 981 1404 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m2778 1408 981 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m2779 1409 1404 1408 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m2780 1 1404 1403 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m2781 1410 971 1409 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m2782 1411 981 1410 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m2783 0 1406 1411 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m2784 1408 971 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m2785 0 1406 1408 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m2786 1412 1406 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m2787 1413 971 1412 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m2788 1404 1406 1413 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m2789 1413 971 1404 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m2790 1414 1409 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m2791 1 981 1413 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m2792 1409 1404 1415 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m2793 1416 971 1409 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m2794 1417 981 1416 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m2795 1406 1418 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2796 1418 1419 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2797 1415 1406 1417 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m2798 1 971 1415 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m2799 1415 1406 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m2800 1 981 1415 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m2801 1414 1409 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m2802 0 1418 1406 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m2803 0 1419 1418 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m2804 0 1331 1419 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m2805 1419 1345 657 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m2806 647 1321 1419 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m2807 1419 1343 632 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m2808 642 1327 1419 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m2809 0 1421 1420 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m2810 1422 1423 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m2811 0 986 1422 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m2812 1424 1423 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m2813 1421 986 1424 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m2814 1422 996 1421 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m2815 1425 996 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m2816 1426 1421 1425 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m2817 1 1421 1420 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m2818 1427 986 1426 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m2819 1428 996 1427 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m2820 0 1423 1428 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m2821 1425 986 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m2822 0 1423 1425 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m2823 1429 1423 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m2824 1430 986 1429 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m2825 1421 1423 1430 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m2826 1430 986 1421 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m2827 1431 1426 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m2828 1 996 1430 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m2829 1426 1421 1432 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m2830 1433 986 1426 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m2831 1434 996 1433 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m2832 1423 1435 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2833 1435 1436 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2834 1432 1423 1434 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m2835 1 986 1432 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m2836 1432 1423 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m2837 1 996 1432 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m2838 1431 1426 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m2839 0 1435 1423 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m2840 0 1436 1435 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m2841 0 1331 1436 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m2842 1436 1345 672 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m2843 662 1321 1436 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m2844 1436 1343 647 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m2845 657 1327 1436 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m2846 0 1438 1437 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m2847 1439 1440 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m2848 0 1001 1439 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m2849 1441 1440 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m2850 1438 1001 1441 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m2851 1439 1011 1438 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m2852 1442 1011 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m2853 1443 1438 1442 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m2854 1 1438 1437 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m2855 1444 1001 1443 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m2856 1445 1011 1444 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m2857 0 1440 1445 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m2858 1442 1001 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m2859 0 1440 1442 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m2860 1446 1440 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m2861 1447 1001 1446 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m2862 1438 1440 1447 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m2863 1447 1001 1438 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m2864 1448 1443 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m2865 1 1011 1447 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m2866 1443 1438 1449 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m2867 1450 1001 1443 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m2868 1451 1011 1450 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m2869 1440 1452 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2870 1452 1453 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2871 1449 1440 1451 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m2872 1 1001 1449 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m2873 1449 1440 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m2874 1 1011 1449 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m2875 1448 1443 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m2876 0 1452 1440 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m2877 0 1453 1452 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m2878 0 1331 1453 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m2879 1453 1345 687 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m2880 677 1321 1453 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m2881 1453 1343 662 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m2882 672 1327 1453 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m2883 0 1455 1454 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m2884 1456 1457 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m2885 0 1016 1456 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m2886 1458 1457 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m2887 1455 1016 1458 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m2888 1456 1026 1455 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m2889 1459 1026 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m2890 1460 1455 1459 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m2891 1 1455 1454 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m2892 1461 1016 1460 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m2893 1462 1026 1461 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m2894 0 1457 1462 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m2895 1459 1016 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m2896 0 1457 1459 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m2897 1463 1457 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m2898 1464 1016 1463 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m2899 1455 1457 1464 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m2900 1464 1016 1455 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m2901 1465 1460 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m2902 1 1026 1464 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m2903 1460 1455 1466 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m2904 1467 1016 1460 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m2905 1468 1026 1467 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m2906 1457 1469 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2907 1469 1470 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2908 1466 1457 1468 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m2909 1 1016 1466 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m2910 1466 1457 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m2911 1 1026 1466 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m2912 1465 1460 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m2913 0 1469 1457 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m2914 0 1470 1469 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m2915 0 1331 1470 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m2916 1470 1345 702 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m2917 692 1321 1470 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m2918 1470 1343 677 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m2919 687 1327 1470 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m2920 0 1472 1471 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m2921 1473 1474 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m2922 0 1031 1473 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m2923 1475 1474 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m2924 1472 1031 1475 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m2925 1473 1041 1472 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m2926 1476 1041 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m2927 1477 1472 1476 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m2928 1 1472 1471 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m2929 1478 1031 1477 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m2930 1479 1041 1478 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m2931 0 1474 1479 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m2932 1476 1031 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m2933 0 1474 1476 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m2934 1480 1474 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m2935 1481 1031 1480 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m2936 1472 1474 1481 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m2937 1481 1031 1472 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m2938 1482 1477 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m2939 1 1041 1481 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m2940 1477 1472 1483 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m2941 1484 1031 1477 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m2942 1485 1041 1484 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m2943 1474 1486 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2944 1486 1487 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2945 1483 1474 1485 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m2946 1 1031 1483 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m2947 1483 1474 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m2948 1 1041 1483 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m2949 1482 1477 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m2950 0 1486 1474 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m2951 0 1487 1486 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m2952 0 1331 1487 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m2953 1487 1345 717 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m2954 707 1321 1487 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m2955 1487 1343 692 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m2956 702 1327 1487 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m2957 0 1489 1488 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m2958 1490 1491 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m2959 0 1046 1490 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m2960 1492 1491 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m2961 1489 1046 1492 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m2962 1490 1056 1489 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m2963 1493 1056 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m2964 1494 1489 1493 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m2965 1 1489 1488 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m2966 1495 1046 1494 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m2967 1496 1056 1495 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m2968 0 1491 1496 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m2969 1493 1046 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m2970 0 1491 1493 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m2971 1497 1491 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m2972 1498 1046 1497 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m2973 1489 1491 1498 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m2974 1498 1046 1489 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m2975 1499 1494 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m2976 1 1056 1498 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m2977 1494 1489 1500 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m2978 1501 1046 1494 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m2979 1502 1056 1501 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m2980 1491 1503 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m2981 1503 1504 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m2982 1500 1491 1502 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m2983 1 1046 1500 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m2984 1500 1491 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m2985 1 1056 1500 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m2986 1499 1494 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m2987 0 1503 1491 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m2988 0 1504 1503 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m2989 0 1331 1504 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m2990 1504 1345 732 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m2991 722 1321 1504 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m2992 1504 1343 707 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m2993 717 1327 1504 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m2994 0 1506 1505 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m2995 1507 1508 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m2996 0 1061 1507 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m2997 1509 1508 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m2998 1506 1061 1509 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m2999 1507 1071 1506 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3000 1510 1071 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3001 1511 1506 1510 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3002 1 1506 1505 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3003 1512 1061 1511 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3004 1513 1071 1512 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3005 0 1508 1513 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3006 1510 1061 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3007 0 1508 1510 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3008 1514 1508 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3009 1515 1061 1514 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3010 1506 1508 1515 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3011 1515 1061 1506 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3012 1516 1511 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3013 1 1071 1515 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3014 1511 1506 1517 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3015 1518 1061 1511 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3016 1519 1071 1518 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3017 1508 1520 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3018 1520 1521 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3019 1517 1508 1519 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3020 1 1061 1517 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3021 1517 1508 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3022 1 1071 1517 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3023 1516 1511 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3024 0 1520 1508 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3025 0 1521 1520 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3026 0 1331 1521 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3027 1521 1345 747 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3028 737 1321 1521 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3029 1521 1343 722 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3030 732 1327 1521 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3031 0 1523 1522 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3032 1524 1525 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3033 0 1076 1524 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3034 1526 1525 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3035 1523 1076 1526 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3036 1524 1086 1523 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3037 1527 1086 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3038 1528 1523 1527 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3039 1 1523 1522 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3040 1529 1076 1528 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3041 1530 1086 1529 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3042 0 1525 1530 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3043 1527 1076 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3044 0 1525 1527 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3045 1531 1525 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3046 1532 1076 1531 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3047 1523 1525 1532 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3048 1532 1076 1523 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3049 1533 1528 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3050 1 1086 1532 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3051 1528 1523 1534 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3052 1535 1076 1528 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3053 1536 1086 1535 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3054 1525 1537 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3055 1537 1538 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3056 1534 1525 1536 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3057 1 1076 1534 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3058 1534 1525 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3059 1 1086 1534 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3060 1533 1528 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3061 0 1537 1525 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3062 0 1538 1537 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3063 0 1331 1538 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3064 1538 1345 762 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3065 752 1321 1538 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3066 1538 1343 737 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3067 747 1327 1538 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3068 0 1540 1539 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3069 1541 1542 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3070 0 1091 1541 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3071 1543 1542 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3072 1540 1091 1543 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3073 1541 1101 1540 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3074 1544 1101 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3075 1545 1540 1544 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3076 1 1540 1539 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3077 1546 1091 1545 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3078 1547 1101 1546 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3079 0 1542 1547 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3080 1544 1091 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3081 0 1542 1544 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3082 1548 1542 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3083 1549 1091 1548 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3084 1540 1542 1549 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3085 1549 1091 1540 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3086 1550 1545 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3087 1 1101 1549 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3088 1545 1540 1551 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3089 1552 1091 1545 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3090 1553 1101 1552 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3091 1542 1554 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3092 1554 1555 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3093 1551 1542 1553 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3094 1 1091 1551 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3095 1551 1542 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3096 1 1101 1551 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3097 1550 1545 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3098 0 1554 1542 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3099 0 1555 1554 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3100 0 1331 1555 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3101 1555 1345 777 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3102 767 1321 1555 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3103 1555 1343 752 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3104 762 1327 1555 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3105 0 1557 1556 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3106 1558 1559 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3107 0 1106 1558 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3108 1560 1559 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3109 1557 1106 1560 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3110 1558 1116 1557 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3111 1561 1116 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3112 1562 1557 1561 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3113 1 1557 1556 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3114 1563 1106 1562 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3115 1564 1116 1563 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3116 0 1559 1564 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3117 1561 1106 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3118 0 1559 1561 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3119 1565 1559 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3120 1566 1106 1565 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3121 1557 1559 1566 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3122 1566 1106 1557 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3123 1567 1562 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3124 1 1116 1566 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3125 1562 1557 1568 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3126 1569 1106 1562 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3127 1570 1116 1569 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3128 1559 1571 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3129 1571 1572 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3130 1568 1559 1570 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3131 1 1106 1568 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3132 1568 1559 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3133 1 1116 1568 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3134 1567 1562 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3135 0 1571 1559 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3136 0 1572 1571 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3137 0 1331 1572 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3138 1572 1345 792 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3139 782 1321 1572 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3140 1572 1343 767 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3141 777 1327 1572 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3142 0 1574 1573 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3143 1575 1576 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3144 0 1121 1575 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3145 1577 1576 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3146 1574 1121 1577 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3147 1575 1131 1574 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3148 1578 1131 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3149 1579 1574 1578 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3150 1 1574 1573 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3151 1580 1121 1579 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3152 1581 1131 1580 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3153 0 1576 1581 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3154 1578 1121 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3155 0 1576 1578 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3156 1582 1576 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3157 1583 1121 1582 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3158 1574 1576 1583 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3159 1583 1121 1574 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3160 1584 1579 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3161 1 1131 1583 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3162 1579 1574 1585 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3163 1586 1121 1579 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3164 1587 1131 1586 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3165 1576 1588 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3166 1588 1589 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3167 1585 1576 1587 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3168 1 1121 1585 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3169 1585 1576 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3170 1 1131 1585 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3171 1584 1579 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3172 0 1588 1576 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3173 0 1589 1588 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3174 0 1331 1589 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3175 1589 1345 807 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3176 797 1321 1589 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3177 1589 1343 782 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3178 792 1327 1589 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3179 0 1591 1590 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3180 1592 1593 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3181 0 1136 1592 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3182 1594 1593 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3183 1591 1136 1594 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3184 1592 1146 1591 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3185 1595 1146 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3186 1596 1591 1595 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3187 1 1591 1590 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3188 1597 1136 1596 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3189 1598 1146 1597 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3190 0 1593 1598 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3191 1595 1136 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3192 0 1593 1595 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3193 1599 1593 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3194 1600 1136 1599 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3195 1591 1593 1600 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3196 1600 1136 1591 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3197 1601 1596 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3198 1 1146 1600 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3199 1596 1591 1602 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3200 1603 1136 1596 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3201 1604 1146 1603 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3202 1593 1605 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3203 1605 1606 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3204 1602 1593 1604 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3205 1 1136 1602 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3206 1602 1593 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3207 1 1146 1602 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3208 1601 1596 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3209 0 1605 1593 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3210 0 1606 1605 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3211 0 1331 1606 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3212 1606 1345 822 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3213 812 1321 1606 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3214 1606 1343 797 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3215 807 1327 1606 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3216 0 1608 1607 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3217 1609 1610 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3218 0 1151 1609 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3219 1611 1610 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3220 1608 1151 1611 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3221 1609 1161 1608 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3222 1612 1161 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3223 1613 1608 1612 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3224 1 1608 1607 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3225 1614 1151 1613 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3226 1615 1161 1614 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3227 0 1610 1615 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3228 1612 1151 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3229 0 1610 1612 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3230 1616 1610 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3231 1617 1151 1616 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3232 1608 1610 1617 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3233 1617 1151 1608 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3234 1618 1613 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3235 1 1161 1617 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3236 1613 1608 1619 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3237 1620 1151 1613 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3238 1621 1161 1620 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3239 1610 1622 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3240 1622 1623 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3241 1619 1610 1621 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3242 1 1151 1619 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3243 1619 1610 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3244 1 1161 1619 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3245 1618 1613 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3246 0 1622 1610 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3247 0 1623 1622 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3248 0 1331 1623 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3249 1623 1345 837 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3250 827 1321 1623 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3251 1623 1343 812 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3252 822 1327 1623 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3253 0 1625 1624 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3254 1626 1627 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3255 0 1166 1626 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3256 1628 1627 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3257 1625 1166 1628 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3258 1626 1176 1625 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3259 1629 1176 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3260 1630 1625 1629 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3261 1 1625 1624 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3262 1631 1166 1630 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3263 1632 1176 1631 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3264 0 1627 1632 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3265 1629 1166 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3266 0 1627 1629 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3267 1633 1627 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3268 1634 1166 1633 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3269 1625 1627 1634 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3270 1634 1166 1625 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3271 1635 1630 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3272 1 1176 1634 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3273 1630 1625 1636 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3274 1637 1166 1630 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3275 1638 1176 1637 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3276 1627 1639 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3277 1639 1640 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3278 1636 1627 1638 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3279 1 1166 1636 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3280 1636 1627 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3281 1 1176 1636 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3282 1635 1630 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3283 0 1639 1627 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3284 0 1640 1639 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3285 0 1331 1640 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3286 1640 1345 868 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3287 842 1321 1640 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3288 1640 1343 827 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3289 837 1327 1640 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3290 0 1642 1641 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3291 1643 1644 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3292 0 1181 1643 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3293 1645 1644 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3294 1642 1181 1645 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3295 1643 1191 1642 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3296 1646 1191 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3297 1647 1642 1646 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3298 1 1642 1641 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3299 1648 1181 1647 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3300 1649 1191 1648 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3301 0 1644 1649 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3302 1646 1181 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3303 0 1644 1646 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3304 1650 1644 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3305 1651 1181 1650 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3306 1642 1644 1651 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3307 1651 1181 1642 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3308 1652 1647 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3309 1 1191 1651 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3310 1647 1642 1653 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3311 1654 1181 1647 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3312 1655 1191 1654 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3313 1644 1656 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3314 1656 1657 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3315 1653 1644 1655 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3316 1 1181 1653 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3317 1653 1644 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3318 1 1191 1653 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3319 1652 1647 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3320 0 1656 1644 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3321 0 1657 1656 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3322 0 1331 1657 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3323 1657 1345 852 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3324 858 1321 1657 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.036e-11 ad=6.95e-12 ps=1.246e-05 pd=8.18e-06 
+ nrs=0.8 nrd=0.54 
m3325 1657 1343 842 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3326 868 1327 1657 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3327 0 1659 1658 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=3.144e-11 ps=2.699e-05 pd=3.25e-05 
+ nrs=0.14 nrd=0.15 
m3328 1660 1661 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.083e-11 ad=3.013e-11 ps=2.27e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m3329 0 1196 1660 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.083e-11 ps=2.849e-05 pd=2.27e-05 
+ nrs=0.13 nrd=0.09 
m3330 1662 1661 0 0 nenh l=1.1e-06 w=1.68e-05 
+ as=1.454e-11 ad=3.33e-11 ps=1.992e-05 pd=3.149e-05 
+ nrs=0.05 nrd=0.12 
m3331 1659 1196 1662 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.246e-11 ps=1.795e-05 pd=1.708e-05 
+ nrs=0.07 nrd=0.06 
m3332 1660 1206 1659 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.919e-11 ad=1.383e-11 ps=2.091e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m3333 1663 1206 0 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.352e-11 ad=2.854e-11 ps=1.61e-05 pd=2.699e-05 
+ nrs=0.07 nrd=0.14 
m3334 1664 1659 1663 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.449e-11 ad=1.352e-11 ps=1.785e-05 pd=1.61e-05 
+ nrs=0.07 nrd=0.07 
m3335 1665 1196 1664 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.489e-11 ps=1.701e-05 pd=1.835e-05 
+ nrs=0.06 nrd=0.07 
m3336 1666 1206 1665 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3337 0 1661 1666 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3338 1663 1196 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.502e-11 ad=3.171e-11 ps=1.789e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3339 0 1661 1663 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.202e-11 ps=2.399e-05 pd=1.431e-05 
+ nrs=0.15 nrd=0.07 
m3340 1 1659 1658 1 penh l=1.1e-06 w=1.8e-05 
+ as=4.008e-11 ad=3.314e-11 ps=3.398e-05 pd=3.89e-05 
+ nrs=0.12 nrd=0.1 
m3341 1667 1664 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3342 1668 1661 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m3343 1669 1196 1668 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m3344 1659 1661 1669 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.615e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3345 1669 1196 1659 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.499e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.06 
m3346 1 1206 1669 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3347 1 1671 1670 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.484e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.47 
m3348 1672 1345 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m3349 1671 1327 1672 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.372e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.44 nrd=0.15 
m3350 1 1673 1661 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.226e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.32 
m3351 1664 1659 1674 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.447e-11 ad=1.386e-11 ps=1.722e-05 pd=1.719e-05 
+ nrs=0.1 nrd=0.1 
m3352 1675 1196 1664 1 penh l=1.1e-06 w=1.88e-05 
+ as=1.621e-11 ad=2.267e-11 ps=2.153e-05 pd=2.698e-05 
+ nrs=0.05 nrd=0.06 
m3353 1676 1206 1675 1 penh l=1.1e-06 w=2.12e-05 
+ as=1.814e-11 ad=1.827e-11 ps=2.344e-05 pd=2.427e-05 
+ nrs=0.04 nrd=0.04 
m3354 1674 1661 1676 1 penh l=1.1e-06 w=2.24e-05 
+ as=2.588e-11 ad=1.916e-11 ps=3.21e-05 pd=2.476e-05 
+ nrs=0.05 nrd=0.04 
m3355 1 1196 1674 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.664e-11 ps=2.718e-05 pd=2.063e-05 
+ nrs=0.15 nrd=0.08 
m3356 1674 1661 1 1 penh l=1.1e-06 w=1.52e-05 
+ as=1.756e-11 ad=3.384e-11 ps=2.178e-05 pd=2.869e-05 
+ nrs=0.08 nrd=0.15 
m3357 1 1206 1674 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.386e-11 ps=2.265e-05 pd=1.719e-05 
+ nrs=0.19 nrd=0.1 
m3358 1667 1664 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.04e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.08 nrd=0.12 
m3359 1673 1677 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.298e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.48 nrd=0.43 
m3360 0 1671 1670 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m3361 1671 1345 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=5.55e-12 ps=6.1e-06 pd=5.25e-06 
+ nrs=0.59 nrd=0.71 
m3362 0 1327 1671 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=4.62e-12 ps=5.25e-06 pd=6.1e-06 
+ nrs=0.71 nrd=0.59 
m3363 0 1673 1661 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.52e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.37 
m3364 0 1677 1673 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3365 0 1331 1677 0 nenh l=1.1e-06 w=3.2e-06 
+ as=6.34e-12 ad=6.09e-12 ps=6e-06 pd=7.29e-06 
+ nrs=0.62 nrd=0.6 
m3366 1677 1345 1 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.098e-11 ps=8.2e-06 pd=1.406e-05 
+ nrs=0.53 nrd=0.85 
m3367 0 1321 1677 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.86e-12 ps=6.75e-06 pd=8.2e-06 
+ nrs=0.55 nrd=0.53 
m3368 1677 1343 858 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.036e-11 ps=8.2e-06 pd=1.246e-05 
+ nrs=0.53 nrd=0.8 
m3369 852 1327 1677 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.86e-12 ps=1.202e-05 pd=8.2e-06 
+ nrs=0.77 nrd=0.53 
m3370 0 1679 1678 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.427e-11 ad=2.196e-11 ps=1.35e-05 pd=2.05e-05 
+ nrs=0.28 nrd=0.42 
m3371 1679 1680 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m3372 0 1682 1681 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.22e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.76 
m3373 1682 1683 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.22e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.76 nrd=0.5 
m3374 1 1679 1678 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m3375 1679 1680 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3376 1684 1685 0 0 nenh l=1.1e-06 w=4e-06 
+ as=6.6e-12 ad=7.93e-12 ps=7.3e-06 pd=7.5e-06 
+ nrs=0.41 nrd=0.5 
m3377 0 1685 1684 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=6.6e-12 ps=7.5e-06 pd=7.3e-06 
+ nrs=0.5 nrd=0.41 
m3378 1686 1687 1685 0 nenh l=1.1e-06 w=8.8e-06 
+ as=7.66e-12 ad=1.964e-11 ps=1.122e-05 pd=2.37e-05 
+ nrs=0.1 nrd=0.25 
m3379 1688 1689 1686 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.4e-12 ps=1.25e-05 pd=1.378e-05 
+ nrs=0.08 nrd=0.08 
m3380 0 1335 1688 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m3381 1690 1687 0 0 nenh l=1.1e-06 w=8.8e-06 
+ as=9.24e-12 ad=1.744e-11 ps=1.13e-05 pd=1.65e-05 
+ nrs=0.12 nrd=0.23 
m3382 0 1691 1690 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.744e-11 ad=9.24e-12 ps=1.65e-05 pd=1.13e-05 
+ nrs=0.23 nrd=0.12 
m3383 1692 1693 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=1.665e-11 ps=1.01e-05 pd=1.575e-05 
+ nrs=0.1 nrd=0.24 
m3384 1694 1695 1692 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.89e-11 ad=7.14e-12 ps=2.29e-05 pd=1.01e-05 
+ nrs=0.27 nrd=0.1 
m3385 1 1682 1681 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=2.358e-11 ps=1.737e-05 pd=2.29e-05 
+ nrs=0.24 nrd=0.28 
m3386 1682 1683 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.358e-11 ad=2.048e-11 ps=2.29e-05 pd=1.737e-05 
+ nrs=0.28 nrd=0.24 
m3387 1684 1685 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.128e-11 ad=2.494e-11 ps=1.37e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m3388 1 1685 1684 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.128e-11 ps=2.114e-05 pd=1.37e-05 
+ nrs=0.2 nrd=0.09 
m3389 1696 1689 1695 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.27e-12 ad=2.16e-11 ps=1.176e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.23 
m3390 1697 1335 1696 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.31e-12 ps=1.25e-05 pd=1.324e-05 
+ nrs=0.08 nrd=0.08 
m3391 0 1698 1697 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m3392 1699 1687 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m3393 1700 1701 1699 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.31e-12 ad=9.18e-12 ps=1.324e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m3394 1693 1324 1700 0 nenh l=1.1e-06 w=9.6e-06 
+ as=2.16e-11 ad=8.27e-12 ps=2.53e-05 pd=1.176e-05 
+ nrs=0.23 nrd=0.09 
m3395 1 1687 1685 1 penh l=1.1e-06 w=9.6e-06 
+ as=2.137e-11 ad=1.315e-11 ps=1.812e-05 pd=1.587e-05 
+ nrs=0.23 nrd=0.14 
m3396 1685 1689 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.26e-11 ad=2.048e-11 ps=1.521e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m3397 1 1335 1685 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.26e-11 ps=1.737e-05 pd=1.521e-05 
+ nrs=0.24 nrd=0.15 
m3398 1702 1687 1 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.194e-11 ad=2.939e-11 ps=1.49e-05 pd=2.492e-05 
+ nrs=0.07 nrd=0.17 
m3399 1690 1691 1702 1 penh l=1.1e-06 w=1.32e-05 
+ as=2.586e-11 ad=1.194e-11 ps=3.01e-05 pd=1.49e-05 
+ nrs=0.15 nrd=0.07 
m3400 1694 1693 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.466e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.07 nrd=0.15 
m3401 1 1695 1694 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.466e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.07 
m3402 1 1689 1695 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m3403 1695 1335 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m3404 1 1698 1695 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m3405 1693 1687 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m3406 1 1701 1693 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m3407 1693 1324 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m3408 1683 1703 1 1 penh l=1.1e-06 w=1e-05 
+ as=2.346e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.23 nrd=0.22 
m3409 1703 1704 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3410 1680 1694 1 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=8.54e-12 ps=7.22e-06 pd=1.094e-05 
+ nrs=0.69 nrd=1.09 
m3411 910 1684 1680 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m3412 1705 1691 1706 1 penh l=1.1e-06 w=1.04e-05 
+ as=8.84e-12 ad=2.596e-11 ps=1.21e-05 pd=2.69e-05 
+ nrs=0.08 nrd=0.24 
m3413 1 1698 1705 1 penh l=1.1e-06 w=1.04e-05 
+ as=2.316e-11 ad=8.84e-12 ps=1.963e-05 pd=1.21e-05 
+ nrs=0.21 nrd=0.08 
m3414 1707 1324 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m3415 1 1701 1707 1 penh l=1.1e-06 w=8e-06 
+ as=1.781e-11 ad=1.075e-11 ps=1.51e-05 pd=1.383e-05 
+ nrs=0.28 nrd=0.17 
m3416 1707 1698 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m3417 1708 1707 1 1 penh l=1.1e-06 w=1e-05 
+ as=1.058e-11 ad=2.227e-11 ps=1.25e-05 pd=1.888e-05 
+ nrs=0.11 nrd=0.22 
m3418 1 1707 1708 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=1.058e-11 ps=1.888e-05 pd=1.25e-05 
+ nrs=0.22 nrd=0.11 
m3419 1704 1708 595 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.74e-12 ps=7.22e-06 pd=9.64e-06 
+ nrs=0.69 nrd=0.99 
m3420 602 1684 1704 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=5.4e-12 ps=9.87e-06 pd=7.22e-06 
+ nrs=1.04 nrd=0.69 
m3421 1704 1690 910 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.88e-12 ps=7.22e-06 pd=1.048e-05 
+ nrs=0.69 nrd=1 
m3422 911 1706 1704 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m3423 0 1694 1704 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.4e-12 ps=5.25e-06 pd=7.22e-06 
+ nrs=0.71 nrd=0.69 
m3424 1709 1701 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=2.405e-11 ps=1.41e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m3425 1691 1324 1709 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.046e-11 ad=1.014e-11 ps=1.25e-05 pd=1.41e-05 
+ nrs=0.09 nrd=0.09 
m3426 1710 1335 1691 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=1.046e-11 ps=1.41e-05 pd=1.25e-05 
+ nrs=0.09 nrd=0.09 
m3427 1 1689 1710 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.014e-11 ps=2.039e-05 pd=1.41e-05 
+ nrs=0.21 nrd=0.09 
m3428 911 1708 1680 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m3429 1680 1690 911 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.91e-12 ps=7.22e-06 pd=1.05e-05 
+ nrs=0.69 nrd=1.01 
m3430 910 1706 1680 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m3431 0 1703 1683 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m3432 0 1704 1703 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m3433 1706 1691 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m3434 0 1698 1706 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m3435 1711 1324 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m3436 1712 1701 1711 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.4e-12 ad=9.18e-12 ps=1.378e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m3437 1707 1698 1712 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.964e-11 ad=7.66e-12 ps=2.37e-05 pd=1.122e-05 
+ nrs=0.25 nrd=0.1 
m3438 1708 1707 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m3439 0 1707 1708 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m3440 1713 1701 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=9.84e-12 ad=2.061e-11 ps=1.319e-05 pd=1.949e-05 
+ nrs=0.09 nrd=0.19 
m3441 1691 1335 1713 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.06e-11 ps=1.29e-05 pd=1.421e-05 
+ nrs=0.09 nrd=0.08 
m3442 1714 1324 1691 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.062e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.08 nrd=0.09 
m3443 0 1689 1714 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.024e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m3444 0 1716 1715 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3445 1717 1718 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3446 0 1315 1717 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3447 1719 1718 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3448 1716 1315 1719 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3449 1717 1318 1716 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3450 1720 1318 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3451 1721 1716 1720 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3452 1 1716 1715 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3453 1722 1315 1721 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3454 1723 1318 1722 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3455 0 1718 1723 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3456 1720 1315 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3457 0 1718 1720 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3458 1724 1718 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3459 1725 1315 1724 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3460 1716 1718 1725 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3461 1725 1315 1716 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3462 1726 1721 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3463 1 1318 1725 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3464 1721 1716 1727 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3465 1728 1315 1721 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3466 1729 1318 1728 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3467 1718 1730 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3468 1730 1731 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3469 1727 1718 1729 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3470 1 1315 1727 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3471 1727 1718 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3472 1 1318 1727 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3473 1726 1721 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3474 0 1730 1718 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3475 0 1731 1730 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3476 0 1694 1731 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3477 1731 1708 612 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3478 601 1684 1731 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3479 1731 1706 602 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.045e-11 ps=8.18e-06 pd=1.269e-05 
+ nrs=0.54 nrd=0.81 
m3480 595 1690 1731 0 nenh l=1.1e-06 w=3.6e-06 
+ as=9.95e-12 ad=6.95e-12 ps=1.239e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3481 0 1733 1732 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3482 1734 1735 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3483 0 1319 1734 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3484 1736 1735 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3485 1733 1319 1736 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3486 1734 1352 1733 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3487 1737 1352 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3488 1738 1733 1737 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3489 1 1733 1732 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3490 1739 1319 1738 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3491 1740 1352 1739 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3492 0 1735 1740 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3493 1737 1319 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3494 0 1735 1737 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3495 1741 1735 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3496 1742 1319 1741 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3497 1733 1735 1742 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3498 1742 1319 1733 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3499 1743 1738 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3500 1 1352 1742 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3501 1738 1733 1744 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3502 1745 1319 1738 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3503 1746 1352 1745 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3504 1735 1747 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3505 1747 1748 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3506 1744 1735 1746 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3507 1 1319 1744 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3508 1744 1735 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3509 1 1352 1744 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3510 1743 1738 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3511 0 1747 1735 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3512 0 1748 1747 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3513 0 1694 1748 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3514 1748 1708 627 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3515 617 1684 1748 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3516 1748 1706 601 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3517 612 1690 1748 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3518 0 1750 1749 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3519 1751 1752 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3520 0 1363 1751 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3521 1753 1752 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3522 1750 1363 1753 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3523 1751 1369 1750 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3524 1754 1369 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3525 1755 1750 1754 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3526 1 1750 1749 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3527 1756 1363 1755 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3528 1757 1369 1756 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3529 0 1752 1757 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3530 1754 1363 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3531 0 1752 1754 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3532 1758 1752 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3533 1759 1363 1758 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3534 1750 1752 1759 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3535 1759 1363 1750 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3536 1760 1755 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3537 1 1369 1759 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3538 1755 1750 1761 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3539 1762 1363 1755 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3540 1763 1369 1762 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3541 1752 1764 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3542 1764 1765 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3543 1761 1752 1763 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3544 1 1363 1761 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3545 1761 1752 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3546 1 1369 1761 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3547 1760 1755 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3548 0 1764 1752 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3549 0 1765 1764 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3550 0 1694 1765 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3551 1765 1708 642 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3552 632 1684 1765 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3553 1765 1706 617 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3554 627 1690 1765 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3555 0 1767 1766 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3556 1768 1769 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3557 0 1380 1768 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3558 1770 1769 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3559 1767 1380 1770 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3560 1768 1386 1767 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3561 1771 1386 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3562 1772 1767 1771 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3563 1 1767 1766 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3564 1773 1380 1772 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3565 1774 1386 1773 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3566 0 1769 1774 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3567 1771 1380 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3568 0 1769 1771 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3569 1775 1769 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3570 1776 1380 1775 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3571 1767 1769 1776 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3572 1776 1380 1767 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3573 1777 1772 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3574 1 1386 1776 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3575 1772 1767 1778 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3576 1779 1380 1772 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3577 1780 1386 1779 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3578 1769 1781 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3579 1781 1782 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3580 1778 1769 1780 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3581 1 1380 1778 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3582 1778 1769 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3583 1 1386 1778 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3584 1777 1772 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3585 0 1781 1769 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3586 0 1782 1781 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3587 0 1694 1782 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3588 1782 1708 657 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3589 647 1684 1782 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3590 1782 1706 632 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3591 642 1690 1782 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3592 0 1784 1783 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3593 1785 1786 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3594 0 1397 1785 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3595 1787 1786 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3596 1784 1397 1787 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3597 1785 1403 1784 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3598 1788 1403 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3599 1789 1784 1788 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3600 1 1784 1783 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3601 1790 1397 1789 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3602 1791 1403 1790 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3603 0 1786 1791 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3604 1788 1397 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3605 0 1786 1788 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3606 1792 1786 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3607 1793 1397 1792 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3608 1784 1786 1793 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3609 1793 1397 1784 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3610 1794 1789 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3611 1 1403 1793 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3612 1789 1784 1795 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3613 1796 1397 1789 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3614 1797 1403 1796 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3615 1786 1798 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3616 1798 1799 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3617 1795 1786 1797 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3618 1 1397 1795 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3619 1795 1786 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3620 1 1403 1795 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3621 1794 1789 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3622 0 1798 1786 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3623 0 1799 1798 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3624 0 1694 1799 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3625 1799 1708 672 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3626 662 1684 1799 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3627 1799 1706 647 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3628 657 1690 1799 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3629 0 1801 1800 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3630 1802 1803 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3631 0 1414 1802 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3632 1804 1803 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3633 1801 1414 1804 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3634 1802 1420 1801 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3635 1805 1420 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3636 1806 1801 1805 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3637 1 1801 1800 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3638 1807 1414 1806 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3639 1808 1420 1807 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3640 0 1803 1808 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3641 1805 1414 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3642 0 1803 1805 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3643 1809 1803 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3644 1810 1414 1809 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3645 1801 1803 1810 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3646 1810 1414 1801 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3647 1811 1806 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3648 1 1420 1810 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3649 1806 1801 1812 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3650 1813 1414 1806 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3651 1814 1420 1813 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3652 1803 1815 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3653 1815 1816 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3654 1812 1803 1814 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3655 1 1414 1812 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3656 1812 1803 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3657 1 1420 1812 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3658 1811 1806 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3659 0 1815 1803 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3660 0 1816 1815 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3661 0 1694 1816 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3662 1816 1708 687 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3663 677 1684 1816 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3664 1816 1706 662 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3665 672 1690 1816 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3666 0 1818 1817 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3667 1819 1820 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3668 0 1431 1819 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3669 1821 1820 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3670 1818 1431 1821 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3671 1819 1437 1818 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3672 1822 1437 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3673 1823 1818 1822 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3674 1 1818 1817 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3675 1824 1431 1823 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3676 1825 1437 1824 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3677 0 1820 1825 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3678 1822 1431 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3679 0 1820 1822 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3680 1826 1820 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3681 1827 1431 1826 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3682 1818 1820 1827 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3683 1827 1431 1818 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3684 1828 1823 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3685 1 1437 1827 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3686 1823 1818 1829 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3687 1830 1431 1823 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3688 1831 1437 1830 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3689 1820 1832 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3690 1832 1833 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3691 1829 1820 1831 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3692 1 1431 1829 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3693 1829 1820 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3694 1 1437 1829 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3695 1828 1823 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3696 0 1832 1820 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3697 0 1833 1832 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3698 0 1694 1833 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3699 1833 1708 702 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3700 692 1684 1833 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3701 1833 1706 677 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3702 687 1690 1833 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3703 0 1835 1834 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3704 1836 1837 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3705 0 1448 1836 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3706 1838 1837 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3707 1835 1448 1838 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3708 1836 1454 1835 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3709 1839 1454 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3710 1840 1835 1839 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3711 1 1835 1834 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3712 1841 1448 1840 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3713 1842 1454 1841 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3714 0 1837 1842 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3715 1839 1448 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3716 0 1837 1839 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3717 1843 1837 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3718 1844 1448 1843 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3719 1835 1837 1844 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3720 1844 1448 1835 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3721 1845 1840 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3722 1 1454 1844 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3723 1840 1835 1846 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3724 1847 1448 1840 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3725 1848 1454 1847 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3726 1837 1849 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3727 1849 1850 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3728 1846 1837 1848 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3729 1 1448 1846 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3730 1846 1837 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3731 1 1454 1846 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3732 1845 1840 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3733 0 1849 1837 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3734 0 1850 1849 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3735 0 1694 1850 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3736 1850 1708 717 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3737 707 1684 1850 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3738 1850 1706 692 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3739 702 1690 1850 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3740 0 1852 1851 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3741 1853 1854 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3742 0 1465 1853 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3743 1855 1854 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3744 1852 1465 1855 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3745 1853 1471 1852 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3746 1856 1471 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3747 1857 1852 1856 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3748 1 1852 1851 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3749 1858 1465 1857 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3750 1859 1471 1858 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3751 0 1854 1859 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3752 1856 1465 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3753 0 1854 1856 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3754 1860 1854 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3755 1861 1465 1860 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3756 1852 1854 1861 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3757 1861 1465 1852 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3758 1862 1857 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3759 1 1471 1861 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3760 1857 1852 1863 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3761 1864 1465 1857 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3762 1865 1471 1864 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3763 1854 1866 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3764 1866 1867 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3765 1863 1854 1865 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3766 1 1465 1863 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3767 1863 1854 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3768 1 1471 1863 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3769 1862 1857 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3770 0 1866 1854 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3771 0 1867 1866 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3772 0 1694 1867 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3773 1867 1708 732 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3774 722 1684 1867 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3775 1867 1706 707 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3776 717 1690 1867 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3777 0 1869 1868 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3778 1870 1871 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3779 0 1482 1870 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3780 1872 1871 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3781 1869 1482 1872 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3782 1870 1488 1869 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3783 1873 1488 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3784 1874 1869 1873 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3785 1 1869 1868 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3786 1875 1482 1874 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3787 1876 1488 1875 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3788 0 1871 1876 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3789 1873 1482 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3790 0 1871 1873 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3791 1877 1871 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3792 1878 1482 1877 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3793 1869 1871 1878 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3794 1878 1482 1869 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3795 1879 1874 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3796 1 1488 1878 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3797 1874 1869 1880 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3798 1881 1482 1874 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3799 1882 1488 1881 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3800 1871 1883 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3801 1883 1884 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3802 1880 1871 1882 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3803 1 1482 1880 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3804 1880 1871 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3805 1 1488 1880 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3806 1879 1874 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3807 0 1883 1871 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3808 0 1884 1883 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3809 0 1694 1884 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3810 1884 1708 747 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3811 737 1684 1884 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3812 1884 1706 722 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3813 732 1690 1884 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3814 0 1886 1885 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3815 1887 1888 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3816 0 1499 1887 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3817 1889 1888 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3818 1886 1499 1889 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3819 1887 1505 1886 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3820 1890 1505 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3821 1891 1886 1890 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3822 1 1886 1885 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3823 1892 1499 1891 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3824 1893 1505 1892 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3825 0 1888 1893 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3826 1890 1499 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3827 0 1888 1890 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3828 1894 1888 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3829 1895 1499 1894 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3830 1886 1888 1895 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3831 1895 1499 1886 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3832 1896 1891 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3833 1 1505 1895 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3834 1891 1886 1897 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3835 1898 1499 1891 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3836 1899 1505 1898 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3837 1888 1900 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3838 1900 1901 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3839 1897 1888 1899 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3840 1 1499 1897 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3841 1897 1888 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3842 1 1505 1897 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3843 1896 1891 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3844 0 1900 1888 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3845 0 1901 1900 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3846 0 1694 1901 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3847 1901 1708 762 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3848 752 1684 1901 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3849 1901 1706 737 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3850 747 1690 1901 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3851 0 1903 1902 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3852 1904 1905 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3853 0 1516 1904 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3854 1906 1905 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3855 1903 1516 1906 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3856 1904 1522 1903 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3857 1907 1522 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3858 1908 1903 1907 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3859 1 1903 1902 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3860 1909 1516 1908 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3861 1910 1522 1909 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3862 0 1905 1910 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3863 1907 1516 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3864 0 1905 1907 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3865 1911 1905 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3866 1912 1516 1911 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3867 1903 1905 1912 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3868 1912 1516 1903 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3869 1913 1908 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3870 1 1522 1912 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3871 1908 1903 1914 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3872 1915 1516 1908 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3873 1916 1522 1915 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3874 1905 1917 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3875 1917 1918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3876 1914 1905 1916 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3877 1 1516 1914 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3878 1914 1905 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3879 1 1522 1914 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3880 1913 1908 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3881 0 1917 1905 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3882 0 1918 1917 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3883 0 1694 1918 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3884 1918 1708 777 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3885 767 1684 1918 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3886 1918 1706 752 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3887 762 1690 1918 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3888 0 1920 1919 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3889 1921 1922 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3890 0 1533 1921 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3891 1923 1922 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3892 1920 1533 1923 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3893 1921 1539 1920 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3894 1924 1539 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3895 1925 1920 1924 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3896 1 1920 1919 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3897 1926 1533 1925 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3898 1927 1539 1926 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3899 0 1922 1927 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3900 1924 1533 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3901 0 1922 1924 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3902 1928 1922 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3903 1929 1533 1928 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3904 1920 1922 1929 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3905 1929 1533 1920 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3906 1930 1925 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3907 1 1539 1929 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3908 1925 1920 1931 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3909 1932 1533 1925 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3910 1933 1539 1932 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3911 1922 1934 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3912 1934 1935 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3913 1931 1922 1933 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3914 1 1533 1931 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3915 1931 1922 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3916 1 1539 1931 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3917 1930 1925 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3918 0 1934 1922 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3919 0 1935 1934 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3920 0 1694 1935 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3921 1935 1708 792 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3922 782 1684 1935 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3923 1935 1706 767 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3924 777 1690 1935 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3925 0 1937 1936 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3926 1938 1939 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3927 0 1550 1938 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3928 1940 1939 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3929 1937 1550 1940 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3930 1938 1556 1937 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3931 1941 1556 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3932 1942 1937 1941 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3933 1 1937 1936 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3934 1943 1550 1942 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3935 1944 1556 1943 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3936 0 1939 1944 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3937 1941 1550 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3938 0 1939 1941 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3939 1945 1939 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3940 1946 1550 1945 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3941 1937 1939 1946 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3942 1946 1550 1937 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3943 1947 1942 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3944 1 1556 1946 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3945 1942 1937 1948 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3946 1949 1550 1942 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3947 1950 1556 1949 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3948 1939 1951 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3949 1951 1952 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3950 1948 1939 1950 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3951 1 1550 1948 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3952 1948 1939 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3953 1 1556 1948 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3954 1947 1942 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3955 0 1951 1939 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3956 0 1952 1951 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3957 0 1694 1952 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3958 1952 1708 807 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3959 797 1684 1952 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3960 1952 1706 782 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3961 792 1690 1952 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3962 0 1954 1953 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m3963 1955 1956 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m3964 0 1567 1955 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m3965 1957 1956 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m3966 1954 1567 1957 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m3967 1955 1573 1954 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m3968 1958 1573 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m3969 1959 1954 1958 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m3970 1 1954 1953 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m3971 1960 1567 1959 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m3972 1961 1573 1960 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m3973 0 1956 1961 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m3974 1958 1567 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m3975 0 1956 1958 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m3976 1962 1956 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m3977 1963 1567 1962 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m3978 1954 1956 1963 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m3979 1963 1567 1954 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m3980 1964 1959 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m3981 1 1573 1963 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m3982 1959 1954 1965 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m3983 1966 1567 1959 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m3984 1967 1573 1966 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m3985 1956 1968 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m3986 1968 1969 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m3987 1965 1956 1967 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m3988 1 1567 1965 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m3989 1965 1956 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m3990 1 1573 1965 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m3991 1964 1959 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m3992 0 1968 1956 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m3993 0 1969 1968 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m3994 0 1694 1969 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m3995 1969 1708 822 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m3996 812 1684 1969 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m3997 1969 1706 797 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m3998 807 1690 1969 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m3999 0 1971 1970 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4000 1972 1973 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4001 0 1584 1972 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4002 1974 1973 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4003 1971 1584 1974 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4004 1972 1590 1971 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4005 1975 1590 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4006 1976 1971 1975 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4007 1 1971 1970 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4008 1977 1584 1976 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4009 1978 1590 1977 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4010 0 1973 1978 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4011 1975 1584 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4012 0 1973 1975 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4013 1979 1973 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4014 1980 1584 1979 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4015 1971 1973 1980 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4016 1980 1584 1971 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4017 1981 1976 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4018 1 1590 1980 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4019 1976 1971 1982 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4020 1983 1584 1976 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4021 1984 1590 1983 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4022 1973 1985 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4023 1985 1986 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4024 1982 1973 1984 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4025 1 1584 1982 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4026 1982 1973 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4027 1 1590 1982 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4028 1981 1976 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4029 0 1985 1973 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4030 0 1986 1985 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4031 0 1694 1986 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4032 1986 1708 837 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4033 827 1684 1986 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4034 1986 1706 812 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4035 822 1690 1986 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4036 0 1988 1987 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4037 1989 1990 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4038 0 1601 1989 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4039 1991 1990 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4040 1988 1601 1991 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4041 1989 1607 1988 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4042 1992 1607 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4043 1993 1988 1992 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4044 1 1988 1987 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4045 1994 1601 1993 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4046 1995 1607 1994 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4047 0 1990 1995 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4048 1992 1601 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4049 0 1990 1992 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4050 1996 1990 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4051 1997 1601 1996 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4052 1988 1990 1997 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4053 1997 1601 1988 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4054 1998 1993 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4055 1 1607 1997 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4056 1993 1988 1999 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4057 2000 1601 1993 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4058 2001 1607 2000 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4059 1990 2002 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4060 2002 2003 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4061 1999 1990 2001 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4062 1 1601 1999 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4063 1999 1990 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4064 1 1607 1999 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4065 1998 1993 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4066 0 2002 1990 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4067 0 2003 2002 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4068 0 1694 2003 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4069 2003 1708 868 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4070 842 1684 2003 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4071 2003 1706 827 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4072 837 1690 2003 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4073 0 2005 2004 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4074 2006 2007 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4075 0 1618 2006 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4076 2008 2007 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4077 2005 1618 2008 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4078 2006 1624 2005 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4079 2009 1624 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4080 2010 2005 2009 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4081 1 2005 2004 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4082 2011 1618 2010 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4083 2012 1624 2011 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4084 0 2007 2012 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4085 2009 1618 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4086 0 2007 2009 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4087 2013 2007 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4088 2014 1618 2013 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4089 2005 2007 2014 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4090 2014 1618 2005 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4091 2015 2010 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4092 1 1624 2014 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4093 2010 2005 2016 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4094 2017 1618 2010 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4095 2018 1624 2017 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4096 2007 2019 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4097 2019 2020 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4098 2016 2007 2018 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4099 1 1618 2016 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4100 2016 2007 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4101 1 1624 2016 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4102 2015 2010 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4103 0 2019 2007 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4104 0 2020 2019 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4105 0 1694 2020 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4106 2020 1708 852 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4107 858 1684 2020 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.036e-11 ad=6.95e-12 ps=1.246e-05 pd=8.18e-06 
+ nrs=0.8 nrd=0.54 
m4108 2020 1706 842 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4109 868 1690 2020 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4110 2021 2022 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=5.99e-12 ad=1.348e-11 ps=9.58e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m4111 236 2023 2021 0 nenh l=1.1e-06 w=6.4e-06 
+ as=7.52e-12 ad=5.63e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.14 
m4112 2024 2025 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m4113 2023 2026 2024 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m4114 2027 2028 2023 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m4115 0 2029 2027 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m4116 2025 2029 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m4117 0 2031 2030 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m4118 2032 2026 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m4119 2033 2030 2032 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m4120 2034 2031 2033 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m4121 0 2028 2034 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m4122 2026 2028 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m4123 2035 2033 236 0 nenh l=1.1e-06 w=6.4e-06 
+ as=5.63e-12 ad=7.52e-12 ps=9.02e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m4124 0 2036 2035 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.99e-12 ps=1.275e-05 pd=9.58e-06 
+ nrs=0.29 nrd=0.13 
m4125 2037 2022 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m4126 236 2033 2037 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m4127 2038 2023 236 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m4128 1 2036 2038 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m4129 2039 2025 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m4130 2023 2028 2039 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m4131 2040 2026 2023 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m4132 1 2029 2040 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m4133 2025 2029 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4134 2041 2029 2042 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.57e-11 ps=1.429e-05 pd=2.04e-05 
+ nrs=0.11 nrd=0.12 
m4135 2043 2044 2041 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m4136 2042 2045 2043 0 nenh l=1.1e-06 w=1e-05 
+ as=1.354e-11 ad=8.5e-12 ps=1.759e-05 pd=1.17e-05 
+ nrs=0.14 nrd=0.08 
m4137 0 2045 2042 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m4138 2042 2044 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m4139 0 2044 2046 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m4140 2046 2045 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m4141 2047 2045 2046 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.354e-11 ps=1.17e-05 pd=1.759e-05 
+ nrs=0.08 nrd=0.14 
m4142 2048 2044 2047 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m4143 0 2049 2045 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m4144 2050 2045 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m4145 2028 2044 2050 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m4146 2051 2015 2028 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m4147 0 2049 2051 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m4148 2044 2015 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m4149 2046 2031 2048 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=1.416e-11 ps=2.04e-05 pd=1.429e-05 
+ nrs=0.12 nrd=0.11 
m4150 1 2031 2030 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m4151 2052 2026 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m4152 2033 2031 2052 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m4153 2053 2030 2033 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m4154 1 2028 2053 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m4155 2026 2028 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m4156 2041 2029 2054 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m4157 2055 2044 2041 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m4158 1 2045 2055 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m4159 2054 2045 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m4160 1 2044 2054 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m4161 2056 2044 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m4162 1 2045 2056 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m4163 2057 2045 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m4164 2048 2044 2057 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m4165 2056 2031 2048 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m4166 1 2049 2045 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=3.262e-11 ps=2.039e-05 pd=2.77e-05 
+ nrs=0.21 nrd=0.28 
m4167 2058 2045 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.23e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m4168 2028 2015 2058 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.067e-11 ad=7.27e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.1 
m4169 2059 2044 2028 1 penh l=1.1e-06 w=7.6e-06 
+ as=6.5e-12 ad=9.65e-12 ps=9.55e-06 pd=9.97e-06 
+ nrs=0.11 nrd=0.17 
m4170 1 2049 2059 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.16e-12 ps=1.359e-05 pd=9.05e-06 
+ nrs=0.31 nrd=0.12 
m4171 2044 2015 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.67e-11 ad=2.405e-11 ps=2.77e-05 pd=2.039e-05 
+ nrs=0.23 nrd=0.21 
m4172 1 2060 207 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m4173 2061 2022 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m4174 2060 2062 2061 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m4175 2063 2064 2060 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m4176 1 2036 2063 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m4177 2065 2066 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m4178 2064 2067 2065 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m4179 2068 2069 2064 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m4180 1 2070 2068 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m4181 2066 2070 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4182 1 2072 2071 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m4183 2073 2069 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m4184 2062 2072 2073 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m4185 2074 2071 2062 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m4186 1 2067 2074 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m4187 2069 2067 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m4188 0 2060 207 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m4189 2075 2022 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=7.37e-12 ad=1.506e-11 ps=1.097e-05 pd=1.425e-05 
+ nrs=0.13 nrd=0.26 
m4190 2060 2064 2075 0 nenh l=1.1e-06 w=6.4e-06 
+ as=8.77e-12 ad=6.21e-12 ps=9.49e-06 pd=9.23e-06 
+ nrs=0.21 nrd=0.15 
m4191 2076 2062 2060 0 nenh l=1.1e-06 w=5.6e-06 
+ as=5.09e-12 ad=7.67e-12 ps=7.68e-06 pd=8.31e-06 
+ nrs=0.16 nrd=0.24 
m4192 0 2036 2076 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=6.17e-12 ps=1.275e-05 pd=9.32e-06 
+ nrs=0.29 nrd=0.13 
m4193 1 2078 2077 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=2.67e-11 ps=2.039e-05 pd=2.77e-05 
+ nrs=0.21 nrd=0.23 
m4194 2079 2080 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=9.84e-12 ad=1.959e-11 ps=1.17e-05 pd=1.661e-05 
+ nrs=0.13 nrd=0.25 
m4195 2067 2078 2079 1 penh l=1.1e-06 w=7.6e-06 
+ as=8.13e-12 ad=8.5e-12 ps=9.97e-06 pd=1.01e-05 
+ nrs=0.14 nrd=0.15 
m4196 2081 2077 2067 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.015e-11 ad=8.99e-12 ps=1.143e-05 pd=1.103e-05 
+ nrs=0.14 nrd=0.13 
m4197 1 2082 2081 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=1.063e-11 ps=1.661e-05 pd=1.197e-05 
+ nrs=0.25 nrd=0.14 
m4198 2080 2082 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m4199 2083 2070 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.55e-11 ad=2.672e-11 ps=1.478e-05 pd=2.265e-05 
+ nrs=0.11 nrd=0.19 
m4200 2029 2078 2083 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.151e-11 ad=1.498e-11 ps=1.394e-05 pd=1.428e-05 
+ nrs=0.09 nrd=0.11 
m4201 2083 2082 2029 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.705e-11 ad=1.309e-11 ps=1.625e-05 pd=1.586e-05 
+ nrs=0.1 nrd=0.08 
m4202 2084 2082 2083 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.498e-11 ps=1.33e-05 pd=1.428e-05 
+ nrs=0.07 nrd=0.11 
m4203 1 2078 2084 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m4204 2085 2078 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m4205 2086 2082 2085 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=9.86e-12 ps=1.428e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m4206 2031 2082 2086 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.309e-11 ad=1.705e-11 ps=1.586e-05 pd=1.625e-05 
+ nrs=0.08 nrd=0.1 
m4207 2086 2078 2031 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=1.151e-11 ps=1.428e-05 pd=1.394e-05 
+ nrs=0.11 nrd=0.09 
m4208 1 2072 2086 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.55e-11 ps=2.265e-05 pd=1.478e-05 
+ nrs=0.19 nrd=0.11 
m4209 2087 2066 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m4210 2064 2069 2087 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m4211 2088 2067 2064 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m4212 0 2070 2088 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m4213 2066 2070 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m4214 0 2072 2071 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m4215 2089 2069 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m4216 2062 2071 2089 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m4217 2090 2072 2062 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m4218 0 2067 2090 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m4219 2069 2067 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m4220 0 2078 2077 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m4221 2091 2080 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m4222 2067 2077 2091 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m4223 2092 2078 2067 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m4224 0 2082 2092 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m4225 2080 2082 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.468e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.47 nrd=0.35 
m4226 2029 2070 2093 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.175e-11 ad=1.755e-11 ps=1.429e-05 pd=1.841e-05 
+ nrs=0.09 nrd=0.13 
m4227 2094 2078 2029 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.013e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.1 
m4228 0 2082 2094 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=8.5e-12 ps=1.874e-05 pd=1.17e-05 
+ nrs=0.2 nrd=0.08 
m4229 2093 2082 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=2.299e-11 ps=1.841e-05 pd=2.174e-05 
+ nrs=0.13 nrd=0.17 
m4230 0 2078 2093 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=1.513e-11 ps=1.874e-05 pd=1.587e-05 
+ nrs=0.2 nrd=0.15 
m4231 2095 2078 0 0 nenh l=1.1e-06 w=1e-05 
+ as=1.513e-11 ad=1.982e-11 ps=1.587e-05 pd=1.874e-05 
+ nrs=0.15 nrd=0.2 
m4232 0 2082 2095 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.755e-11 ps=2.174e-05 pd=1.841e-05 
+ nrs=0.17 nrd=0.13 
m4233 2096 2082 0 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.982e-11 ps=1.17e-05 pd=1.874e-05 
+ nrs=0.08 nrd=0.2 
m4234 2031 2078 2096 0 nenh l=1.1e-06 w=1e-05 
+ as=1.013e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.1 nrd=0.08 
m4235 2095 2072 2031 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=1.175e-11 ps=1.841e-05 pd=1.429e-05 
+ nrs=0.13 nrd=0.09 
m4236 2097 2022 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.04e-12 ad=1.348e-11 ps=9.88e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m4237 178 2098 2097 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=5.33e-12 ps=8.5e-06 pd=8.72e-06 
+ nrs=0.19 nrd=0.15 
m4238 2099 2100 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m4239 2098 2101 2099 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m4240 2102 2103 2098 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m4241 0 2104 2102 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m4242 2100 2104 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m4243 0 2106 2105 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m4244 2107 2101 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m4245 2108 2105 2107 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m4246 2109 2106 2108 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m4247 0 2103 2109 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m4248 2101 2103 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m4249 2110 2108 178 0 nenh l=1.1e-06 w=6e-06 
+ as=5.29e-12 ad=6.86e-12 ps=8.61e-06 pd=8.5e-06 
+ nrs=0.15 nrd=0.19 
m4250 0 2036 2110 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=5.65e-12 ps=1.2e-05 pd=9.19e-06 
+ nrs=0.31 nrd=0.14 
m4251 2111 2022 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m4252 178 2108 2111 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m4253 2112 2098 178 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m4254 1 2036 2112 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m4255 2113 2100 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m4256 2098 2103 2113 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m4257 2114 2101 2098 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m4258 1 2104 2114 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m4259 2100 2104 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.308e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.42 nrd=0.4 
m4260 2070 2104 2115 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.57e-11 ps=1.429e-05 pd=2.04e-05 
+ nrs=0.11 nrd=0.12 
m4261 2116 2117 2070 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m4262 2115 2118 2116 0 nenh l=1.1e-06 w=1e-05 
+ as=1.354e-11 ad=8.5e-12 ps=1.759e-05 pd=1.17e-05 
+ nrs=0.14 nrd=0.08 
m4263 0 2118 2115 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m4264 2115 2117 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m4265 0 2117 2119 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m4266 2119 2118 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m4267 2120 2118 2119 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.354e-11 ps=1.17e-05 pd=1.759e-05 
+ nrs=0.08 nrd=0.14 
m4268 2072 2117 2120 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m4269 2119 2106 2072 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=1.416e-11 ps=2.04e-05 pd=1.429e-05 
+ nrs=0.12 nrd=0.11 
m4270 0 1658 2118 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.42e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.45 
m4271 2121 2118 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m4272 2103 2117 2121 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m4273 2122 1652 2103 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m4274 0 1658 2122 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m4275 2117 1652 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.372e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.44 nrd=0.35 
m4276 1 2106 2105 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m4277 2123 2101 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m4278 2108 2106 2123 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m4279 2124 2105 2108 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m4280 1 2103 2124 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m4281 2101 2103 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m4282 2070 2104 2125 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m4283 2126 2117 2070 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m4284 1 2118 2126 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m4285 2125 2118 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m4286 1 2117 2125 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m4287 2127 2117 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m4288 1 2118 2127 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m4289 2128 2118 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m4290 2072 2117 2128 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m4291 2127 2106 2072 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m4292 1 1658 2118 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=2.67e-11 ps=2.039e-05 pd=2.77e-05 
+ nrs=0.21 nrd=0.23 
m4293 2129 2118 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.45e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m4294 2103 1652 2129 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.033e-11 ad=7.53e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.11 
m4295 2130 2117 2103 1 penh l=1.1e-06 w=7.6e-06 
+ as=7.02e-12 ad=9.35e-12 ps=1.01e-05 pd=9.97e-06 
+ nrs=0.12 nrd=0.16 
m4296 1 1658 2130 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=8.12e-12 ps=1.661e-05 pd=1.17e-05 
+ nrs=0.25 nrd=0.1 
m4297 2117 1652 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.67e-11 ad=2.405e-11 ps=2.77e-05 pd=2.039e-05 
+ nrs=0.23 nrd=0.21 
m4298 1 2131 149 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m4299 2132 2022 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m4300 2131 2133 2132 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m4301 2134 2135 2131 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m4302 1 2036 2134 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m4303 2022 2036 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.484e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m4304 1 2036 2022 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.484e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m4305 2036 2136 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m4306 1 2136 2036 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m4307 2135 2133 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.596e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.51 nrd=0.4 
m4308 1 1667 2137 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m4309 2138 2139 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m4310 2133 1667 2138 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m4311 2140 2137 2133 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m4312 1 1670 2140 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m4313 2139 1670 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m4314 0 2131 149 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m4315 2141 2022 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=7.37e-12 ad=1.506e-11 ps=1.097e-05 pd=1.425e-05 
+ nrs=0.13 nrd=0.26 
m4316 2131 2135 2141 0 nenh l=1.1e-06 w=6.4e-06 
+ as=8.77e-12 ad=6.21e-12 ps=9.49e-06 pd=9.23e-06 
+ nrs=0.21 nrd=0.15 
m4317 2142 2133 2131 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=7.67e-12 ps=7.3e-06 pd=8.31e-06 
+ nrs=0.15 nrd=0.24 
m4318 0 2036 2142 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m4319 2022 2036 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.254e-11 ad=1.506e-11 ps=1.09e-05 pd=1.425e-05 
+ nrs=0.22 nrd=0.26 
m4320 0 2036 2022 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.506e-11 ad=1.254e-11 ps=1.425e-05 pd=1.09e-05 
+ nrs=0.26 nrd=0.22 
m4321 2036 2136 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m4322 0 2136 2036 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m4323 2135 2133 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m4324 2143 1667 2104 1 penh l=1.1e-06 w=1.44e-05 
+ as=1.224e-11 ad=4.04e-11 ps=1.61e-05 pd=3.49e-05 
+ nrs=0.06 nrd=0.19 
m4325 1 1670 2143 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.224e-11 ps=2.718e-05 pd=1.61e-05 
+ nrs=0.15 nrd=0.06 
m4326 2136 2144 1 1 penh l=1.1e-06 w=1.44e-05 
+ as=2.376e-11 ad=3.206e-11 ps=1.77e-05 pd=2.718e-05 
+ nrs=0.11 nrd=0.15 
m4327 1 2144 2136 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=2.376e-11 ps=2.718e-05 pd=1.77e-05 
+ nrs=0.15 nrd=0.11 
m4328 2144 1249 1 1 penh l=1.1e-06 w=1.28e-05 
+ as=1.616e-11 ad=2.85e-11 ps=1.53e-05 pd=2.416e-05 
+ nrs=0.1 nrd=0.17 
m4329 1 1257 2144 1 penh l=1.1e-06 w=1.28e-05 
+ as=2.85e-11 ad=1.616e-11 ps=2.416e-05 pd=1.53e-05 
+ nrs=0.17 nrd=0.1 
m4330 2106 1667 1 1 penh l=1.1e-06 w=1.28e-05 
+ as=1.264e-11 ad=2.85e-11 ps=1.53e-05 pd=2.416e-05 
+ nrs=0.08 nrd=0.17 
m4331 1 1670 2106 1 penh l=1.1e-06 w=1.28e-05 
+ as=2.85e-11 ad=1.264e-11 ps=2.416e-05 pd=1.53e-05 
+ nrs=0.17 nrd=0.08 
m4332 0 1667 2137 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.031e-11 ad=1.586e-11 ps=9.75e-06 pd=1.65e-05 
+ nrs=0.38 nrd=0.59 
m4333 2145 2139 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.32e-12 ad=1.348e-11 ps=9.63e-06 pd=1.275e-05 
+ nrs=0.14 nrd=0.29 
m4334 2133 2137 2145 0 nenh l=1.1e-06 w=5.2e-06 
+ as=8.58e-12 ad=4.84e-12 ps=8.5e-06 pd=7.37e-06 
+ nrs=0.32 nrd=0.18 
m4335 2146 1667 2133 0 nenh l=1.1e-06 w=5.2e-06 
+ as=4.56e-12 ad=8.58e-12 ps=7.37e-06 pd=8.5e-06 
+ nrs=0.17 nrd=0.32 
m4336 0 1670 2146 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.96e-12 ps=1.275e-05 pd=9.63e-06 
+ nrs=0.29 nrd=0.13 
m4337 2139 1670 0 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.031e-11 ps=1.65e-05 pd=9.75e-06 
+ nrs=0.59 nrd=0.38 
m4338 2104 1667 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=1.06e-11 ad=2.061e-11 ps=1.29e-05 pd=1.949e-05 
+ nrs=0.1 nrd=0.19 
m4339 0 1670 2104 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.061e-11 ad=1.06e-11 ps=1.949e-05 pd=1.29e-05 
+ nrs=0.19 nrd=0.1 
m4340 2136 2144 0 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.584e-11 ad=1.903e-11 ps=1.29e-05 pd=1.799e-05 
+ nrs=0.17 nrd=0.21 
m4341 0 2144 2136 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=1.584e-11 ps=1.799e-05 pd=1.29e-05 
+ nrs=0.21 nrd=0.17 
m4342 2147 1249 0 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.16e-12 ad=1.903e-11 ps=1.13e-05 pd=1.799e-05 
+ nrs=0.09 nrd=0.21 
m4343 2144 1257 2147 0 nenh l=1.1e-06 w=9.6e-06 
+ as=2.928e-11 ad=8.16e-12 ps=2.53e-05 pd=1.13e-05 
+ nrs=0.32 nrd=0.09 
m4344 2148 1667 2106 0 nenh l=1.1e-06 w=1.28e-05 
+ as=1.088e-11 ad=3.904e-11 ps=1.45e-05 pd=3.17e-05 
+ nrs=0.07 nrd=0.24 
m4345 0 1670 2148 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.088e-11 ps=2.399e-05 pd=1.45e-05 
+ nrs=0.15 nrd=0.07 
m4346 0 2149 2049 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=3.144e-11 ps=2.699e-05 pd=3.25e-05 
+ nrs=0.14 nrd=0.15 
m4347 2150 2151 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.083e-11 ad=3.013e-11 ps=2.27e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m4348 0 1635 2150 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.083e-11 ps=2.849e-05 pd=2.27e-05 
+ nrs=0.13 nrd=0.09 
m4349 2152 2151 0 0 nenh l=1.1e-06 w=1.68e-05 
+ as=1.454e-11 ad=3.33e-11 ps=1.992e-05 pd=3.149e-05 
+ nrs=0.05 nrd=0.12 
m4350 2149 1635 2152 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.246e-11 ps=1.795e-05 pd=1.708e-05 
+ nrs=0.07 nrd=0.06 
m4351 2150 1641 2149 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.919e-11 ad=1.383e-11 ps=2.091e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m4352 2153 1641 0 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.352e-11 ad=2.854e-11 ps=1.61e-05 pd=2.699e-05 
+ nrs=0.07 nrd=0.14 
m4353 2154 2149 2153 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.449e-11 ad=1.352e-11 ps=1.785e-05 pd=1.61e-05 
+ nrs=0.07 nrd=0.07 
m4354 2155 1635 2154 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.489e-11 ps=1.701e-05 pd=1.835e-05 
+ nrs=0.06 nrd=0.07 
m4355 2156 1641 2155 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4356 0 2151 2156 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4357 2153 1635 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.502e-11 ad=3.171e-11 ps=1.789e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4358 0 2151 2153 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.202e-11 ps=2.399e-05 pd=1.431e-05 
+ nrs=0.15 nrd=0.07 
m4359 1 2149 2049 1 penh l=1.1e-06 w=1.8e-05 
+ as=4.008e-11 ad=3.314e-11 ps=3.398e-05 pd=3.89e-05 
+ nrs=0.12 nrd=0.1 
m4360 2078 2154 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4361 2157 2151 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m4362 2158 1635 2157 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m4363 2149 2151 2158 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.615e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4364 2158 1635 2149 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.499e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.06 
m4365 1 1641 2158 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4366 1 2159 2082 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.484e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.47 
m4367 2160 1708 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m4368 2159 1690 2160 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.372e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.44 nrd=0.15 
m4369 1 2161 2151 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.226e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.32 
m4370 2154 2149 2162 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.447e-11 ad=1.386e-11 ps=1.722e-05 pd=1.719e-05 
+ nrs=0.1 nrd=0.1 
m4371 2163 1635 2154 1 penh l=1.1e-06 w=1.88e-05 
+ as=1.621e-11 ad=2.267e-11 ps=2.153e-05 pd=2.698e-05 
+ nrs=0.05 nrd=0.06 
m4372 2164 1641 2163 1 penh l=1.1e-06 w=2.12e-05 
+ as=1.814e-11 ad=1.827e-11 ps=2.344e-05 pd=2.427e-05 
+ nrs=0.04 nrd=0.04 
m4373 2162 2151 2164 1 penh l=1.1e-06 w=2.24e-05 
+ as=2.588e-11 ad=1.916e-11 ps=3.21e-05 pd=2.476e-05 
+ nrs=0.05 nrd=0.04 
m4374 1 1635 2162 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.664e-11 ps=2.718e-05 pd=2.063e-05 
+ nrs=0.15 nrd=0.08 
m4375 2162 2151 1 1 penh l=1.1e-06 w=1.52e-05 
+ as=1.756e-11 ad=3.384e-11 ps=2.178e-05 pd=2.869e-05 
+ nrs=0.08 nrd=0.15 
m4376 1 1641 2162 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.386e-11 ps=2.265e-05 pd=1.719e-05 
+ nrs=0.19 nrd=0.1 
m4377 2078 2154 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.04e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.08 nrd=0.12 
m4378 2161 2165 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.298e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.48 nrd=0.43 
m4379 0 2159 2082 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m4380 2159 1708 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=5.55e-12 ps=6.1e-06 pd=5.25e-06 
+ nrs=0.59 nrd=0.71 
m4381 0 1690 2159 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=4.62e-12 ps=5.25e-06 pd=6.1e-06 
+ nrs=0.71 nrd=0.59 
m4382 0 2161 2151 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.52e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.37 
m4383 0 2165 2161 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4384 0 1694 2165 0 nenh l=1.1e-06 w=3.2e-06 
+ as=6.34e-12 ad=6.09e-12 ps=6e-06 pd=7.29e-06 
+ nrs=0.62 nrd=0.6 
m4385 2165 1708 1 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.098e-11 ps=8.2e-06 pd=1.406e-05 
+ nrs=0.53 nrd=0.85 
m4386 0 1684 2165 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.86e-12 ps=6.75e-06 pd=8.2e-06 
+ nrs=0.55 nrd=0.53 
m4387 2165 1706 858 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.036e-11 ps=8.2e-06 pd=1.246e-05 
+ nrs=0.53 nrd=0.8 
m4388 852 1690 2165 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.86e-12 ps=1.202e-05 pd=8.2e-06 
+ nrs=0.77 nrd=0.53 
m4389 0 2167 2166 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.427e-11 ad=2.196e-11 ps=1.35e-05 pd=2.05e-05 
+ nrs=0.28 nrd=0.42 
m4390 2167 2168 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m4391 0 2170 2169 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.22e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.76 
m4392 2170 2171 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.22e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.76 nrd=0.5 
m4393 1 2167 2166 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m4394 2167 2168 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4395 2172 2173 0 0 nenh l=1.1e-06 w=4e-06 
+ as=6.6e-12 ad=7.93e-12 ps=7.3e-06 pd=7.5e-06 
+ nrs=0.41 nrd=0.5 
m4396 0 2173 2172 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=6.6e-12 ps=7.5e-06 pd=7.3e-06 
+ nrs=0.5 nrd=0.41 
m4397 2174 2175 2173 0 nenh l=1.1e-06 w=8.8e-06 
+ as=7.66e-12 ad=1.964e-11 ps=1.122e-05 pd=2.37e-05 
+ nrs=0.1 nrd=0.25 
m4398 2176 2177 2174 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.4e-12 ps=1.25e-05 pd=1.378e-05 
+ nrs=0.08 nrd=0.08 
m4399 0 1698 2176 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m4400 2178 2175 0 0 nenh l=1.1e-06 w=8.8e-06 
+ as=9.24e-12 ad=1.744e-11 ps=1.13e-05 pd=1.65e-05 
+ nrs=0.12 nrd=0.23 
m4401 0 2179 2178 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.744e-11 ad=9.24e-12 ps=1.65e-05 pd=1.13e-05 
+ nrs=0.23 nrd=0.12 
m4402 2180 2181 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=1.665e-11 ps=1.01e-05 pd=1.575e-05 
+ nrs=0.1 nrd=0.24 
m4403 2182 2183 2180 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.89e-11 ad=7.14e-12 ps=2.29e-05 pd=1.01e-05 
+ nrs=0.27 nrd=0.1 
m4404 1 2170 2169 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=2.358e-11 ps=1.737e-05 pd=2.29e-05 
+ nrs=0.24 nrd=0.28 
m4405 2170 2171 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.358e-11 ad=2.048e-11 ps=2.29e-05 pd=1.737e-05 
+ nrs=0.28 nrd=0.24 
m4406 2172 2173 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.128e-11 ad=2.494e-11 ps=1.37e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m4407 1 2173 2172 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.128e-11 ps=2.114e-05 pd=1.37e-05 
+ nrs=0.2 nrd=0.09 
m4408 2184 2177 2183 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.27e-12 ad=2.16e-11 ps=1.176e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.23 
m4409 2185 1698 2184 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.31e-12 ps=1.25e-05 pd=1.324e-05 
+ nrs=0.08 nrd=0.08 
m4410 0 2186 2185 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m4411 2187 2175 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m4412 2188 2189 2187 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.31e-12 ad=9.18e-12 ps=1.324e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m4413 2181 1687 2188 0 nenh l=1.1e-06 w=9.6e-06 
+ as=2.16e-11 ad=8.27e-12 ps=2.53e-05 pd=1.176e-05 
+ nrs=0.23 nrd=0.09 
m4414 1 2175 2173 1 penh l=1.1e-06 w=9.6e-06 
+ as=2.137e-11 ad=1.315e-11 ps=1.812e-05 pd=1.587e-05 
+ nrs=0.23 nrd=0.14 
m4415 2173 2177 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.26e-11 ad=2.048e-11 ps=1.521e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m4416 1 1698 2173 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.26e-11 ps=1.737e-05 pd=1.521e-05 
+ nrs=0.24 nrd=0.15 
m4417 2190 2175 1 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.194e-11 ad=2.939e-11 ps=1.49e-05 pd=2.492e-05 
+ nrs=0.07 nrd=0.17 
m4418 2178 2179 2190 1 penh l=1.1e-06 w=1.32e-05 
+ as=2.586e-11 ad=1.194e-11 ps=3.01e-05 pd=1.49e-05 
+ nrs=0.15 nrd=0.07 
m4419 2182 2181 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.466e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.07 nrd=0.15 
m4420 1 2183 2182 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.466e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.07 
m4421 1 2177 2183 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m4422 2183 1698 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m4423 1 2186 2183 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m4424 2181 2175 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m4425 1 2189 2181 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m4426 2181 1687 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m4427 2171 2191 1 1 penh l=1.1e-06 w=1e-05 
+ as=2.346e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.23 nrd=0.22 
m4428 2191 2192 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4429 2168 2182 1 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=8.54e-12 ps=7.22e-06 pd=1.094e-05 
+ nrs=0.69 nrd=1.09 
m4430 910 2172 2168 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m4431 2193 2179 2194 1 penh l=1.1e-06 w=1.04e-05 
+ as=8.84e-12 ad=2.596e-11 ps=1.21e-05 pd=2.69e-05 
+ nrs=0.08 nrd=0.24 
m4432 1 2186 2193 1 penh l=1.1e-06 w=1.04e-05 
+ as=2.316e-11 ad=8.84e-12 ps=1.963e-05 pd=1.21e-05 
+ nrs=0.21 nrd=0.08 
m4433 2195 1687 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m4434 1 2189 2195 1 penh l=1.1e-06 w=8e-06 
+ as=1.781e-11 ad=1.075e-11 ps=1.51e-05 pd=1.383e-05 
+ nrs=0.28 nrd=0.17 
m4435 2195 2186 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m4436 2196 2195 1 1 penh l=1.1e-06 w=1e-05 
+ as=1.058e-11 ad=2.227e-11 ps=1.25e-05 pd=1.888e-05 
+ nrs=0.11 nrd=0.22 
m4437 1 2195 2196 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=1.058e-11 ps=1.888e-05 pd=1.25e-05 
+ nrs=0.22 nrd=0.11 
m4438 2192 2196 595 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.74e-12 ps=7.22e-06 pd=9.64e-06 
+ nrs=0.69 nrd=0.99 
m4439 602 2172 2192 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=5.4e-12 ps=9.87e-06 pd=7.22e-06 
+ nrs=1.04 nrd=0.69 
m4440 2192 2178 910 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.88e-12 ps=7.22e-06 pd=1.048e-05 
+ nrs=0.69 nrd=1 
m4441 911 2194 2192 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m4442 0 2182 2192 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.4e-12 ps=5.25e-06 pd=7.22e-06 
+ nrs=0.71 nrd=0.69 
m4443 2197 2189 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=2.405e-11 ps=1.41e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m4444 2179 1687 2197 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.046e-11 ad=1.014e-11 ps=1.25e-05 pd=1.41e-05 
+ nrs=0.09 nrd=0.09 
m4445 2198 1698 2179 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=1.046e-11 ps=1.41e-05 pd=1.25e-05 
+ nrs=0.09 nrd=0.09 
m4446 1 2177 2198 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.014e-11 ps=2.039e-05 pd=1.41e-05 
+ nrs=0.21 nrd=0.09 
m4447 911 2196 2168 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m4448 2168 2178 911 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.91e-12 ps=7.22e-06 pd=1.05e-05 
+ nrs=0.69 nrd=1.01 
m4449 910 2194 2168 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m4450 0 2191 2171 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m4451 0 2192 2191 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m4452 2194 2179 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m4453 0 2186 2194 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m4454 2199 1687 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m4455 2200 2189 2199 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.4e-12 ad=9.18e-12 ps=1.378e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m4456 2195 2186 2200 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.964e-11 ad=7.66e-12 ps=2.37e-05 pd=1.122e-05 
+ nrs=0.25 nrd=0.1 
m4457 2196 2195 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m4458 0 2195 2196 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m4459 2201 2189 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=9.84e-12 ad=2.061e-11 ps=1.319e-05 pd=1.949e-05 
+ nrs=0.09 nrd=0.19 
m4460 2179 1698 2201 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.06e-11 ps=1.29e-05 pd=1.421e-05 
+ nrs=0.09 nrd=0.08 
m4461 2202 1687 2179 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.062e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.08 nrd=0.09 
m4462 0 2177 2202 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.024e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m4463 0 2204 2203 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4464 2205 2206 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4465 0 1678 2205 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4466 2207 2206 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4467 2204 1678 2207 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4468 2205 1681 2204 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4469 2208 1681 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4470 2209 2204 2208 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4471 1 2204 2203 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4472 2210 1678 2209 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4473 2211 1681 2210 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4474 0 2206 2211 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4475 2208 1678 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4476 0 2206 2208 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4477 2212 2206 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4478 2213 1678 2212 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4479 2204 2206 2213 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4480 2213 1678 2204 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4481 2214 2209 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4482 1 1681 2213 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4483 2209 2204 2215 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4484 2216 1678 2209 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4485 2217 1681 2216 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4486 2206 2218 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4487 2218 2219 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4488 2215 2206 2217 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4489 1 1678 2215 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4490 2215 2206 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4491 1 1681 2215 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4492 2214 2209 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4493 0 2218 2206 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4494 0 2219 2218 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4495 0 2182 2219 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4496 2219 2196 612 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4497 601 2172 2219 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4498 2219 2194 602 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.045e-11 ps=8.18e-06 pd=1.269e-05 
+ nrs=0.54 nrd=0.81 
m4499 595 2178 2219 0 nenh l=1.1e-06 w=3.6e-06 
+ as=9.95e-12 ad=6.95e-12 ps=1.239e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4500 0 2221 2220 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4501 2222 2223 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4502 0 1682 2222 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4503 2224 2223 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4504 2221 1682 2224 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4505 2222 1715 2221 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4506 2225 1715 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4507 2226 2221 2225 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4508 1 2221 2220 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4509 2227 1682 2226 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4510 2228 1715 2227 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4511 0 2223 2228 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4512 2225 1682 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4513 0 2223 2225 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4514 2229 2223 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4515 2230 1682 2229 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4516 2221 2223 2230 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4517 2230 1682 2221 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4518 2231 2226 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4519 1 1715 2230 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4520 2226 2221 2232 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4521 2233 1682 2226 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4522 2234 1715 2233 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4523 2223 2235 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4524 2235 2236 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4525 2232 2223 2234 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4526 1 1682 2232 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4527 2232 2223 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4528 1 1715 2232 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4529 2231 2226 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4530 0 2235 2223 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4531 0 2236 2235 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4532 0 2182 2236 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4533 2236 2196 627 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4534 617 2172 2236 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4535 2236 2194 601 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4536 612 2178 2236 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4537 0 2238 2237 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4538 2239 2240 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4539 0 1726 2239 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4540 2241 2240 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4541 2238 1726 2241 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4542 2239 1732 2238 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4543 2242 1732 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4544 2243 2238 2242 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4545 1 2238 2237 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4546 2244 1726 2243 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4547 2245 1732 2244 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4548 0 2240 2245 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4549 2242 1726 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4550 0 2240 2242 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4551 2246 2240 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4552 2247 1726 2246 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4553 2238 2240 2247 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4554 2247 1726 2238 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4555 2248 2243 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4556 1 1732 2247 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4557 2243 2238 2249 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4558 2250 1726 2243 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4559 2251 1732 2250 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4560 2240 2252 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4561 2252 2253 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4562 2249 2240 2251 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4563 1 1726 2249 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4564 2249 2240 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4565 1 1732 2249 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4566 2248 2243 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4567 0 2252 2240 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4568 0 2253 2252 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4569 0 2182 2253 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4570 2253 2196 642 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4571 632 2172 2253 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4572 2253 2194 617 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4573 627 2178 2253 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4574 0 2255 2254 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4575 2256 2257 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4576 0 1743 2256 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4577 2258 2257 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4578 2255 1743 2258 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4579 2256 1749 2255 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4580 2259 1749 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4581 2260 2255 2259 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4582 1 2255 2254 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4583 2261 1743 2260 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4584 2262 1749 2261 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4585 0 2257 2262 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4586 2259 1743 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4587 0 2257 2259 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4588 2263 2257 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4589 2264 1743 2263 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4590 2255 2257 2264 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4591 2264 1743 2255 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4592 2265 2260 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4593 1 1749 2264 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4594 2260 2255 2266 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4595 2267 1743 2260 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4596 2268 1749 2267 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4597 2257 2269 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4598 2269 2270 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4599 2266 2257 2268 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4600 1 1743 2266 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4601 2266 2257 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4602 1 1749 2266 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4603 2265 2260 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4604 0 2269 2257 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4605 0 2270 2269 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4606 0 2182 2270 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4607 2270 2196 657 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4608 647 2172 2270 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4609 2270 2194 632 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4610 642 2178 2270 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4611 0 2272 2271 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4612 2273 2274 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4613 0 1760 2273 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4614 2275 2274 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4615 2272 1760 2275 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4616 2273 1766 2272 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4617 2276 1766 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4618 2277 2272 2276 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4619 1 2272 2271 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4620 2278 1760 2277 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4621 2279 1766 2278 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4622 0 2274 2279 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4623 2276 1760 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4624 0 2274 2276 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4625 2280 2274 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4626 2281 1760 2280 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4627 2272 2274 2281 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4628 2281 1760 2272 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4629 2282 2277 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4630 1 1766 2281 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4631 2277 2272 2283 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4632 2284 1760 2277 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4633 2285 1766 2284 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4634 2274 2286 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4635 2286 2287 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4636 2283 2274 2285 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4637 1 1760 2283 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4638 2283 2274 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4639 1 1766 2283 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4640 2282 2277 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4641 0 2286 2274 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4642 0 2287 2286 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4643 0 2182 2287 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4644 2287 2196 672 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4645 662 2172 2287 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4646 2287 2194 647 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4647 657 2178 2287 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4648 0 2289 2288 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4649 2290 2291 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4650 0 1777 2290 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4651 2292 2291 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4652 2289 1777 2292 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4653 2290 1783 2289 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4654 2293 1783 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4655 2294 2289 2293 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4656 1 2289 2288 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4657 2295 1777 2294 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4658 2296 1783 2295 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4659 0 2291 2296 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4660 2293 1777 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4661 0 2291 2293 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4662 2297 2291 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4663 2298 1777 2297 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4664 2289 2291 2298 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4665 2298 1777 2289 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4666 2299 2294 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4667 1 1783 2298 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4668 2294 2289 2300 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4669 2301 1777 2294 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4670 2302 1783 2301 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4671 2291 2303 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4672 2303 2304 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4673 2300 2291 2302 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4674 1 1777 2300 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4675 2300 2291 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4676 1 1783 2300 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4677 2299 2294 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4678 0 2303 2291 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4679 0 2304 2303 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4680 0 2182 2304 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4681 2304 2196 687 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4682 677 2172 2304 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4683 2304 2194 662 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4684 672 2178 2304 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4685 0 2306 2305 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4686 2307 2308 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4687 0 1794 2307 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4688 2309 2308 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4689 2306 1794 2309 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4690 2307 1800 2306 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4691 2310 1800 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4692 2311 2306 2310 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4693 1 2306 2305 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4694 2312 1794 2311 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4695 2313 1800 2312 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4696 0 2308 2313 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4697 2310 1794 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4698 0 2308 2310 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4699 2314 2308 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4700 2315 1794 2314 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4701 2306 2308 2315 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4702 2315 1794 2306 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4703 2316 2311 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4704 1 1800 2315 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4705 2311 2306 2317 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4706 2318 1794 2311 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4707 2319 1800 2318 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4708 2308 2320 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4709 2320 2321 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4710 2317 2308 2319 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4711 1 1794 2317 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4712 2317 2308 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4713 1 1800 2317 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4714 2316 2311 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4715 0 2320 2308 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4716 0 2321 2320 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4717 0 2182 2321 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4718 2321 2196 702 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4719 692 2172 2321 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4720 2321 2194 677 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4721 687 2178 2321 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4722 0 2323 2322 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4723 2324 2325 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4724 0 1811 2324 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4725 2326 2325 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4726 2323 1811 2326 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4727 2324 1817 2323 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4728 2327 1817 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4729 2328 2323 2327 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4730 1 2323 2322 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4731 2329 1811 2328 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4732 2330 1817 2329 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4733 0 2325 2330 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4734 2327 1811 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4735 0 2325 2327 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4736 2331 2325 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4737 2332 1811 2331 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4738 2323 2325 2332 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4739 2332 1811 2323 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4740 2333 2328 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4741 1 1817 2332 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4742 2328 2323 2334 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4743 2335 1811 2328 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4744 2336 1817 2335 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4745 2325 2337 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4746 2337 2338 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4747 2334 2325 2336 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4748 1 1811 2334 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4749 2334 2325 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4750 1 1817 2334 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4751 2333 2328 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4752 0 2337 2325 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4753 0 2338 2337 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4754 0 2182 2338 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4755 2338 2196 717 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4756 707 2172 2338 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4757 2338 2194 692 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4758 702 2178 2338 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4759 0 2340 2339 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4760 2341 2342 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4761 0 1828 2341 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4762 2343 2342 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4763 2340 1828 2343 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4764 2341 1834 2340 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4765 2344 1834 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4766 2345 2340 2344 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4767 1 2340 2339 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4768 2346 1828 2345 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4769 2347 1834 2346 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4770 0 2342 2347 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4771 2344 1828 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4772 0 2342 2344 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4773 2348 2342 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4774 2349 1828 2348 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4775 2340 2342 2349 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4776 2349 1828 2340 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4777 2350 2345 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4778 1 1834 2349 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4779 2345 2340 2351 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4780 2352 1828 2345 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4781 2353 1834 2352 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4782 2342 2354 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4783 2354 2355 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4784 2351 2342 2353 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4785 1 1828 2351 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4786 2351 2342 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4787 1 1834 2351 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4788 2350 2345 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4789 0 2354 2342 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4790 0 2355 2354 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4791 0 2182 2355 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4792 2355 2196 732 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4793 722 2172 2355 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4794 2355 2194 707 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4795 717 2178 2355 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4796 0 2357 2356 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4797 2358 2359 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4798 0 1845 2358 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4799 2360 2359 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4800 2357 1845 2360 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4801 2358 1851 2357 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4802 2361 1851 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4803 2362 2357 2361 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4804 1 2357 2356 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4805 2363 1845 2362 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4806 2364 1851 2363 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4807 0 2359 2364 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4808 2361 1845 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4809 0 2359 2361 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4810 2365 2359 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4811 2366 1845 2365 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4812 2357 2359 2366 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4813 2366 1845 2357 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4814 2367 2362 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4815 1 1851 2366 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4816 2362 2357 2368 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4817 2369 1845 2362 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4818 2370 1851 2369 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4819 2359 2371 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4820 2371 2372 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4821 2368 2359 2370 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4822 1 1845 2368 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4823 2368 2359 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4824 1 1851 2368 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4825 2367 2362 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4826 0 2371 2359 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4827 0 2372 2371 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4828 0 2182 2372 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4829 2372 2196 747 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4830 737 2172 2372 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4831 2372 2194 722 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4832 732 2178 2372 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4833 0 2374 2373 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4834 2375 2376 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4835 0 1862 2375 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4836 2377 2376 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4837 2374 1862 2377 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4838 2375 1868 2374 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4839 2378 1868 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4840 2379 2374 2378 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4841 1 2374 2373 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4842 2380 1862 2379 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4843 2381 1868 2380 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4844 0 2376 2381 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4845 2378 1862 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4846 0 2376 2378 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4847 2382 2376 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4848 2383 1862 2382 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4849 2374 2376 2383 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4850 2383 1862 2374 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4851 2384 2379 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4852 1 1868 2383 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4853 2379 2374 2385 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4854 2386 1862 2379 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4855 2387 1868 2386 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4856 2376 2388 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4857 2388 2389 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4858 2385 2376 2387 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4859 1 1862 2385 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4860 2385 2376 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4861 1 1868 2385 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4862 2384 2379 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4863 0 2388 2376 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4864 0 2389 2388 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4865 0 2182 2389 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4866 2389 2196 762 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4867 752 2172 2389 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4868 2389 2194 737 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4869 747 2178 2389 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4870 0 2391 2390 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4871 2392 2393 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4872 0 1879 2392 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4873 2394 2393 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4874 2391 1879 2394 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4875 2392 1885 2391 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4876 2395 1885 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4877 2396 2391 2395 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4878 1 2391 2390 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4879 2397 1879 2396 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4880 2398 1885 2397 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4881 0 2393 2398 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4882 2395 1879 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4883 0 2393 2395 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4884 2399 2393 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4885 2400 1879 2399 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4886 2391 2393 2400 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4887 2400 1879 2391 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4888 2401 2396 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4889 1 1885 2400 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4890 2396 2391 2402 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4891 2403 1879 2396 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4892 2404 1885 2403 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4893 2393 2405 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4894 2405 2406 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4895 2402 2393 2404 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4896 1 1879 2402 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4897 2402 2393 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4898 1 1885 2402 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4899 2401 2396 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4900 0 2405 2393 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4901 0 2406 2405 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4902 0 2182 2406 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4903 2406 2196 777 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4904 767 2172 2406 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4905 2406 2194 752 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4906 762 2178 2406 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4907 0 2408 2407 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4908 2409 2410 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4909 0 1896 2409 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4910 2411 2410 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4911 2408 1896 2411 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4912 2409 1902 2408 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4913 2412 1902 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4914 2413 2408 2412 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4915 1 2408 2407 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4916 2414 1896 2413 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4917 2415 1902 2414 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4918 0 2410 2415 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4919 2412 1896 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4920 0 2410 2412 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4921 2416 2410 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4922 2417 1896 2416 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4923 2408 2410 2417 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4924 2417 1896 2408 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4925 2418 2413 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4926 1 1902 2417 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4927 2413 2408 2419 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4928 2420 1896 2413 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4929 2421 1902 2420 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4930 2410 2422 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4931 2422 2423 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4932 2419 2410 2421 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4933 1 1896 2419 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4934 2419 2410 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4935 1 1902 2419 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4936 2418 2413 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4937 0 2422 2410 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4938 0 2423 2422 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4939 0 2182 2423 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4940 2423 2196 792 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4941 782 2172 2423 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4942 2423 2194 767 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4943 777 2178 2423 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4944 0 2425 2424 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4945 2426 2427 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4946 0 1913 2426 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4947 2428 2427 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4948 2425 1913 2428 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4949 2426 1919 2425 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4950 2429 1919 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4951 2430 2425 2429 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4952 1 2425 2424 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4953 2431 1913 2430 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4954 2432 1919 2431 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4955 0 2427 2432 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4956 2429 1913 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4957 0 2427 2429 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4958 2433 2427 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4959 2434 1913 2433 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4960 2425 2427 2434 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4961 2434 1913 2425 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4962 2435 2430 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m4963 1 1919 2434 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m4964 2430 2425 2436 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m4965 2437 1913 2430 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m4966 2438 1919 2437 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m4967 2427 2439 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m4968 2439 2440 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m4969 2436 2427 2438 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m4970 1 1913 2436 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m4971 2436 2427 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m4972 1 1919 2436 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m4973 2435 2430 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m4974 0 2439 2427 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m4975 0 2440 2439 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m4976 0 2182 2440 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m4977 2440 2196 807 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m4978 797 2172 2440 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m4979 2440 2194 782 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m4980 792 2178 2440 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m4981 0 2442 2441 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m4982 2443 2444 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m4983 0 1930 2443 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m4984 2445 2444 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m4985 2442 1930 2445 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m4986 2443 1936 2442 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m4987 2446 1936 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m4988 2447 2442 2446 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m4989 1 2442 2441 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m4990 2448 1930 2447 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m4991 2449 1936 2448 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m4992 0 2444 2449 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m4993 2446 1930 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m4994 0 2444 2446 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m4995 2450 2444 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m4996 2451 1930 2450 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m4997 2442 2444 2451 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m4998 2451 1930 2442 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m4999 2452 2447 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5000 1 1936 2451 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5001 2447 2442 2453 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5002 2454 1930 2447 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5003 2455 1936 2454 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5004 2444 2456 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5005 2456 2457 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5006 2453 2444 2455 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5007 1 1930 2453 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5008 2453 2444 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5009 1 1936 2453 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5010 2452 2447 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5011 0 2456 2444 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5012 0 2457 2456 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5013 0 2182 2457 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5014 2457 2196 822 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5015 812 2172 2457 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5016 2457 2194 797 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5017 807 2178 2457 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5018 0 2459 2458 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5019 2460 2461 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5020 0 1947 2460 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5021 2462 2461 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5022 2459 1947 2462 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5023 2460 1953 2459 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5024 2463 1953 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5025 2464 2459 2463 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5026 1 2459 2458 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5027 2465 1947 2464 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5028 2466 1953 2465 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5029 0 2461 2466 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5030 2463 1947 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5031 0 2461 2463 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5032 2467 2461 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5033 2468 1947 2467 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5034 2459 2461 2468 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5035 2468 1947 2459 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5036 2469 2464 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5037 1 1953 2468 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5038 2464 2459 2470 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5039 2471 1947 2464 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5040 2472 1953 2471 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5041 2461 2473 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5042 2473 2474 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5043 2470 2461 2472 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5044 1 1947 2470 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5045 2470 2461 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5046 1 1953 2470 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5047 2469 2464 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5048 0 2473 2461 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5049 0 2474 2473 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5050 0 2182 2474 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5051 2474 2196 837 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5052 827 2172 2474 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5053 2474 2194 812 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5054 822 2178 2474 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5055 0 2476 2475 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5056 2477 2478 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5057 0 1964 2477 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5058 2479 2478 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5059 2476 1964 2479 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5060 2477 1970 2476 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5061 2480 1970 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5062 2481 2476 2480 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5063 1 2476 2475 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5064 2482 1964 2481 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5065 2483 1970 2482 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5066 0 2478 2483 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5067 2480 1964 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5068 0 2478 2480 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5069 2484 2478 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5070 2485 1964 2484 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5071 2476 2478 2485 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5072 2485 1964 2476 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5073 2486 2481 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5074 1 1970 2485 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5075 2481 2476 2487 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5076 2488 1964 2481 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5077 2489 1970 2488 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5078 2478 2490 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5079 2490 2491 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5080 2487 2478 2489 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5081 1 1964 2487 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5082 2487 2478 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5083 1 1970 2487 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5084 2486 2481 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5085 0 2490 2478 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5086 0 2491 2490 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5087 0 2182 2491 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5088 2491 2196 868 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5089 842 2172 2491 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5090 2491 2194 827 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5091 837 2178 2491 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5092 0 2493 2492 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5093 2494 2495 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5094 0 1981 2494 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5095 2496 2495 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5096 2493 1981 2496 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5097 2494 1987 2493 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5098 2497 1987 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5099 2498 2493 2497 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5100 1 2493 2492 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5101 2499 1981 2498 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5102 2500 1987 2499 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5103 0 2495 2500 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5104 2497 1981 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5105 0 2495 2497 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5106 2501 2495 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5107 2502 1981 2501 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5108 2493 2495 2502 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5109 2502 1981 2493 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5110 2503 2498 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5111 1 1987 2502 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5112 2498 2493 2504 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5113 2505 1981 2498 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5114 2506 1987 2505 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5115 2495 2507 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5116 2507 2508 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5117 2504 2495 2506 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5118 1 1981 2504 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5119 2504 2495 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5120 1 1987 2504 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5121 2503 2498 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5122 0 2507 2495 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5123 0 2508 2507 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5124 0 2182 2508 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5125 2508 2196 852 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5126 858 2172 2508 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.036e-11 ad=6.95e-12 ps=1.246e-05 pd=8.18e-06 
+ nrs=0.8 nrd=0.54 
m5127 2508 2194 842 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5128 868 2178 2508 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5129 0 2510 2509 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=3.144e-11 ps=2.699e-05 pd=3.25e-05 
+ nrs=0.14 nrd=0.15 
m5130 2511 2512 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.083e-11 ad=3.013e-11 ps=2.27e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m5131 0 1998 2511 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.083e-11 ps=2.849e-05 pd=2.27e-05 
+ nrs=0.13 nrd=0.09 
m5132 2513 2512 0 0 nenh l=1.1e-06 w=1.68e-05 
+ as=1.454e-11 ad=3.33e-11 ps=1.992e-05 pd=3.149e-05 
+ nrs=0.05 nrd=0.12 
m5133 2510 1998 2513 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.246e-11 ps=1.795e-05 pd=1.708e-05 
+ nrs=0.07 nrd=0.06 
m5134 2511 2004 2510 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.919e-11 ad=1.383e-11 ps=2.091e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m5135 2514 2004 0 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.352e-11 ad=2.854e-11 ps=1.61e-05 pd=2.699e-05 
+ nrs=0.07 nrd=0.14 
m5136 2515 2510 2514 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.449e-11 ad=1.352e-11 ps=1.785e-05 pd=1.61e-05 
+ nrs=0.07 nrd=0.07 
m5137 2516 1998 2515 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.489e-11 ps=1.701e-05 pd=1.835e-05 
+ nrs=0.06 nrd=0.07 
m5138 2517 2004 2516 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5139 0 2512 2517 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5140 2514 1998 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.502e-11 ad=3.171e-11 ps=1.789e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5141 0 2512 2514 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.202e-11 ps=2.399e-05 pd=1.431e-05 
+ nrs=0.15 nrd=0.07 
m5142 1 2510 2509 1 penh l=1.1e-06 w=1.8e-05 
+ as=4.008e-11 ad=3.314e-11 ps=3.398e-05 pd=3.89e-05 
+ nrs=0.12 nrd=0.1 
m5143 2518 2515 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5144 2519 2512 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m5145 2520 1998 2519 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m5146 2510 2512 2520 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.615e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5147 2520 1998 2510 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.499e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.06 
m5148 1 2004 2520 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5149 1 2522 2521 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.484e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.47 
m5150 2523 2196 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m5151 2522 2178 2523 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.372e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.44 nrd=0.15 
m5152 1 2524 2512 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.226e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.32 
m5153 2515 2510 2525 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.447e-11 ad=1.386e-11 ps=1.722e-05 pd=1.719e-05 
+ nrs=0.1 nrd=0.1 
m5154 2526 1998 2515 1 penh l=1.1e-06 w=1.88e-05 
+ as=1.621e-11 ad=2.267e-11 ps=2.153e-05 pd=2.698e-05 
+ nrs=0.05 nrd=0.06 
m5155 2527 2004 2526 1 penh l=1.1e-06 w=2.12e-05 
+ as=1.814e-11 ad=1.827e-11 ps=2.344e-05 pd=2.427e-05 
+ nrs=0.04 nrd=0.04 
m5156 2525 2512 2527 1 penh l=1.1e-06 w=2.24e-05 
+ as=2.588e-11 ad=1.916e-11 ps=3.21e-05 pd=2.476e-05 
+ nrs=0.05 nrd=0.04 
m5157 1 1998 2525 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.664e-11 ps=2.718e-05 pd=2.063e-05 
+ nrs=0.15 nrd=0.08 
m5158 2525 2512 1 1 penh l=1.1e-06 w=1.52e-05 
+ as=1.756e-11 ad=3.384e-11 ps=2.178e-05 pd=2.869e-05 
+ nrs=0.08 nrd=0.15 
m5159 1 2004 2525 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.386e-11 ps=2.265e-05 pd=1.719e-05 
+ nrs=0.19 nrd=0.1 
m5160 2518 2515 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.04e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.08 nrd=0.12 
m5161 2524 2528 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.298e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.48 nrd=0.43 
m5162 0 2522 2521 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m5163 2522 2196 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=5.55e-12 ps=6.1e-06 pd=5.25e-06 
+ nrs=0.59 nrd=0.71 
m5164 0 2178 2522 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=4.62e-12 ps=5.25e-06 pd=6.1e-06 
+ nrs=0.71 nrd=0.59 
m5165 0 2524 2512 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.52e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.37 
m5166 0 2528 2524 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5167 0 2182 2528 0 nenh l=1.1e-06 w=3.2e-06 
+ as=6.34e-12 ad=6.09e-12 ps=6e-06 pd=7.29e-06 
+ nrs=0.62 nrd=0.6 
m5168 2528 2196 1 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.098e-11 ps=8.2e-06 pd=1.406e-05 
+ nrs=0.53 nrd=0.85 
m5169 0 2172 2528 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.86e-12 ps=6.75e-06 pd=8.2e-06 
+ nrs=0.55 nrd=0.53 
m5170 2528 2194 858 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.036e-11 ps=8.2e-06 pd=1.246e-05 
+ nrs=0.53 nrd=0.8 
m5171 852 2178 2528 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.86e-12 ps=1.202e-05 pd=8.2e-06 
+ nrs=0.77 nrd=0.53 
m5172 0 2530 2529 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.427e-11 ad=2.196e-11 ps=1.35e-05 pd=2.05e-05 
+ nrs=0.28 nrd=0.42 
m5173 2530 2531 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m5174 0 2533 2532 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.22e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.76 
m5175 2533 2534 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.22e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.76 nrd=0.5 
m5176 1 2530 2529 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m5177 2530 2531 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5178 2535 2536 0 0 nenh l=1.1e-06 w=4e-06 
+ as=6.6e-12 ad=7.93e-12 ps=7.3e-06 pd=7.5e-06 
+ nrs=0.41 nrd=0.5 
m5179 0 2536 2535 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=6.6e-12 ps=7.5e-06 pd=7.3e-06 
+ nrs=0.5 nrd=0.41 
m5180 2537 2538 2536 0 nenh l=1.1e-06 w=8.8e-06 
+ as=7.66e-12 ad=1.964e-11 ps=1.122e-05 pd=2.37e-05 
+ nrs=0.1 nrd=0.25 
m5181 2539 2540 2537 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.4e-12 ps=1.25e-05 pd=1.378e-05 
+ nrs=0.08 nrd=0.08 
m5182 0 2186 2539 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m5183 2541 2538 0 0 nenh l=1.1e-06 w=8.8e-06 
+ as=9.24e-12 ad=1.744e-11 ps=1.13e-05 pd=1.65e-05 
+ nrs=0.12 nrd=0.23 
m5184 0 2542 2541 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.744e-11 ad=9.24e-12 ps=1.65e-05 pd=1.13e-05 
+ nrs=0.23 nrd=0.12 
m5185 2543 2544 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=1.665e-11 ps=1.01e-05 pd=1.575e-05 
+ nrs=0.1 nrd=0.24 
m5186 2545 2546 2543 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.89e-11 ad=7.14e-12 ps=2.29e-05 pd=1.01e-05 
+ nrs=0.27 nrd=0.1 
m5187 1 2533 2532 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=2.358e-11 ps=1.737e-05 pd=2.29e-05 
+ nrs=0.24 nrd=0.28 
m5188 2533 2534 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.358e-11 ad=2.048e-11 ps=2.29e-05 pd=1.737e-05 
+ nrs=0.28 nrd=0.24 
m5189 2535 2536 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.128e-11 ad=2.494e-11 ps=1.37e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m5190 1 2536 2535 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.128e-11 ps=2.114e-05 pd=1.37e-05 
+ nrs=0.2 nrd=0.09 
m5191 2547 2540 2546 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.27e-12 ad=2.16e-11 ps=1.176e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.23 
m5192 2548 2186 2547 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.31e-12 ps=1.25e-05 pd=1.324e-05 
+ nrs=0.08 nrd=0.08 
m5193 0 2549 2548 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m5194 2550 2538 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m5195 2551 2552 2550 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.31e-12 ad=9.18e-12 ps=1.324e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m5196 2544 2175 2551 0 nenh l=1.1e-06 w=9.6e-06 
+ as=2.16e-11 ad=8.27e-12 ps=2.53e-05 pd=1.176e-05 
+ nrs=0.23 nrd=0.09 
m5197 1 2538 2536 1 penh l=1.1e-06 w=9.6e-06 
+ as=2.137e-11 ad=1.315e-11 ps=1.812e-05 pd=1.587e-05 
+ nrs=0.23 nrd=0.14 
m5198 2536 2540 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.26e-11 ad=2.048e-11 ps=1.521e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m5199 1 2186 2536 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.26e-11 ps=1.737e-05 pd=1.521e-05 
+ nrs=0.24 nrd=0.15 
m5200 2553 2538 1 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.194e-11 ad=2.939e-11 ps=1.49e-05 pd=2.492e-05 
+ nrs=0.07 nrd=0.17 
m5201 2541 2542 2553 1 penh l=1.1e-06 w=1.32e-05 
+ as=2.586e-11 ad=1.194e-11 ps=3.01e-05 pd=1.49e-05 
+ nrs=0.15 nrd=0.07 
m5202 2545 2544 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.466e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.07 nrd=0.15 
m5203 1 2546 2545 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.466e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.07 
m5204 1 2540 2546 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m5205 2546 2186 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m5206 1 2549 2546 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m5207 2544 2538 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m5208 1 2552 2544 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m5209 2544 2175 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m5210 2534 2554 1 1 penh l=1.1e-06 w=1e-05 
+ as=2.346e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.23 nrd=0.22 
m5211 2554 2555 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5212 2531 2545 1 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=8.54e-12 ps=7.22e-06 pd=1.094e-05 
+ nrs=0.69 nrd=1.09 
m5213 910 2535 2531 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m5214 2556 2542 2557 1 penh l=1.1e-06 w=1.04e-05 
+ as=8.84e-12 ad=2.596e-11 ps=1.21e-05 pd=2.69e-05 
+ nrs=0.08 nrd=0.24 
m5215 1 2549 2556 1 penh l=1.1e-06 w=1.04e-05 
+ as=2.316e-11 ad=8.84e-12 ps=1.963e-05 pd=1.21e-05 
+ nrs=0.21 nrd=0.08 
m5216 2558 2175 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m5217 1 2552 2558 1 penh l=1.1e-06 w=8e-06 
+ as=1.781e-11 ad=1.075e-11 ps=1.51e-05 pd=1.383e-05 
+ nrs=0.28 nrd=0.17 
m5218 2558 2549 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m5219 2559 2558 1 1 penh l=1.1e-06 w=1e-05 
+ as=1.058e-11 ad=2.227e-11 ps=1.25e-05 pd=1.888e-05 
+ nrs=0.11 nrd=0.22 
m5220 1 2558 2559 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=1.058e-11 ps=1.888e-05 pd=1.25e-05 
+ nrs=0.22 nrd=0.11 
m5221 2555 2559 595 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.74e-12 ps=7.22e-06 pd=9.64e-06 
+ nrs=0.69 nrd=0.99 
m5222 602 2535 2555 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=5.4e-12 ps=9.87e-06 pd=7.22e-06 
+ nrs=1.04 nrd=0.69 
m5223 2555 2541 910 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.88e-12 ps=7.22e-06 pd=1.048e-05 
+ nrs=0.69 nrd=1 
m5224 911 2557 2555 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m5225 0 2545 2555 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.4e-12 ps=5.25e-06 pd=7.22e-06 
+ nrs=0.71 nrd=0.69 
m5226 2560 2552 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=2.405e-11 ps=1.41e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m5227 2542 2175 2560 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.046e-11 ad=1.014e-11 ps=1.25e-05 pd=1.41e-05 
+ nrs=0.09 nrd=0.09 
m5228 2561 2186 2542 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=1.046e-11 ps=1.41e-05 pd=1.25e-05 
+ nrs=0.09 nrd=0.09 
m5229 1 2540 2561 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.014e-11 ps=2.039e-05 pd=1.41e-05 
+ nrs=0.21 nrd=0.09 
m5230 911 2559 2531 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m5231 2531 2541 911 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.91e-12 ps=7.22e-06 pd=1.05e-05 
+ nrs=0.69 nrd=1.01 
m5232 910 2557 2531 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m5233 0 2554 2534 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m5234 0 2555 2554 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m5235 2557 2542 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m5236 0 2549 2557 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m5237 2562 2175 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m5238 2563 2552 2562 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.4e-12 ad=9.18e-12 ps=1.378e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m5239 2558 2549 2563 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.964e-11 ad=7.66e-12 ps=2.37e-05 pd=1.122e-05 
+ nrs=0.25 nrd=0.1 
m5240 2559 2558 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m5241 0 2558 2559 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m5242 2564 2552 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=9.84e-12 ad=2.061e-11 ps=1.319e-05 pd=1.949e-05 
+ nrs=0.09 nrd=0.19 
m5243 2542 2186 2564 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.06e-11 ps=1.29e-05 pd=1.421e-05 
+ nrs=0.09 nrd=0.08 
m5244 2565 2175 2542 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.062e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.08 nrd=0.09 
m5245 0 2540 2565 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.024e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m5246 0 2567 2566 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5247 2568 2569 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5248 0 2166 2568 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5249 2570 2569 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5250 2567 2166 2570 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5251 2568 2169 2567 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5252 2571 2169 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5253 2572 2567 2571 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5254 1 2567 2566 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5255 2573 2166 2572 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5256 2574 2169 2573 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5257 0 2569 2574 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5258 2571 2166 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5259 0 2569 2571 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5260 2575 2569 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5261 2576 2166 2575 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5262 2567 2569 2576 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5263 2576 2166 2567 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5264 2577 2572 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5265 1 2169 2576 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5266 2572 2567 2578 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5267 2579 2166 2572 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5268 2580 2169 2579 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5269 2569 2581 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5270 2581 2582 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5271 2578 2569 2580 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5272 1 2166 2578 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5273 2578 2569 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5274 1 2169 2578 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5275 2577 2572 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5276 0 2581 2569 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5277 0 2582 2581 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5278 0 2545 2582 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5279 2582 2559 612 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5280 601 2535 2582 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5281 2582 2557 602 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.045e-11 ps=8.18e-06 pd=1.269e-05 
+ nrs=0.54 nrd=0.81 
m5282 595 2541 2582 0 nenh l=1.1e-06 w=3.6e-06 
+ as=9.95e-12 ad=6.95e-12 ps=1.239e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5283 0 2584 2583 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5284 2585 2586 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5285 0 2170 2585 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5286 2587 2586 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5287 2584 2170 2587 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5288 2585 2203 2584 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5289 2588 2203 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5290 2589 2584 2588 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5291 1 2584 2583 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5292 2590 2170 2589 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5293 2591 2203 2590 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5294 0 2586 2591 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5295 2588 2170 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5296 0 2586 2588 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5297 2592 2586 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5298 2593 2170 2592 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5299 2584 2586 2593 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5300 2593 2170 2584 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5301 2594 2589 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5302 1 2203 2593 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5303 2589 2584 2595 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5304 2596 2170 2589 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5305 2597 2203 2596 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5306 2586 2598 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5307 2598 2599 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5308 2595 2586 2597 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5309 1 2170 2595 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5310 2595 2586 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5311 1 2203 2595 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5312 2594 2589 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5313 0 2598 2586 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5314 0 2599 2598 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5315 0 2545 2599 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5316 2599 2559 627 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5317 617 2535 2599 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5318 2599 2557 601 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5319 612 2541 2599 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5320 0 2601 2600 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5321 2602 2603 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5322 0 2214 2602 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5323 2604 2603 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5324 2601 2214 2604 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5325 2602 2220 2601 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5326 2605 2220 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5327 2606 2601 2605 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5328 1 2601 2600 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5329 2607 2214 2606 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5330 2608 2220 2607 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5331 0 2603 2608 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5332 2605 2214 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5333 0 2603 2605 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5334 2609 2603 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5335 2610 2214 2609 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5336 2601 2603 2610 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5337 2610 2214 2601 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5338 2611 2606 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5339 1 2220 2610 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5340 2606 2601 2612 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5341 2613 2214 2606 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5342 2614 2220 2613 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5343 2603 2615 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5344 2615 2616 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5345 2612 2603 2614 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5346 1 2214 2612 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5347 2612 2603 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5348 1 2220 2612 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5349 2611 2606 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5350 0 2615 2603 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5351 0 2616 2615 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5352 0 2545 2616 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5353 2616 2559 642 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5354 632 2535 2616 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5355 2616 2557 617 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5356 627 2541 2616 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5357 0 2618 2617 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5358 2619 2620 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5359 0 2231 2619 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5360 2621 2620 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5361 2618 2231 2621 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5362 2619 2237 2618 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5363 2622 2237 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5364 2623 2618 2622 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5365 1 2618 2617 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5366 2624 2231 2623 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5367 2625 2237 2624 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5368 0 2620 2625 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5369 2622 2231 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5370 0 2620 2622 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5371 2626 2620 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5372 2627 2231 2626 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5373 2618 2620 2627 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5374 2627 2231 2618 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5375 2628 2623 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5376 1 2237 2627 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5377 2623 2618 2629 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5378 2630 2231 2623 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5379 2631 2237 2630 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5380 2620 2632 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5381 2632 2633 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5382 2629 2620 2631 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5383 1 2231 2629 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5384 2629 2620 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5385 1 2237 2629 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5386 2628 2623 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5387 0 2632 2620 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5388 0 2633 2632 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5389 0 2545 2633 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5390 2633 2559 657 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5391 647 2535 2633 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5392 2633 2557 632 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5393 642 2541 2633 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5394 0 2635 2634 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5395 2636 2637 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5396 0 2248 2636 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5397 2638 2637 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5398 2635 2248 2638 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5399 2636 2254 2635 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5400 2639 2254 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5401 2640 2635 2639 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5402 1 2635 2634 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5403 2641 2248 2640 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5404 2642 2254 2641 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5405 0 2637 2642 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5406 2639 2248 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5407 0 2637 2639 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5408 2643 2637 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5409 2644 2248 2643 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5410 2635 2637 2644 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5411 2644 2248 2635 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5412 2645 2640 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5413 1 2254 2644 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5414 2640 2635 2646 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5415 2647 2248 2640 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5416 2648 2254 2647 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5417 2637 2649 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5418 2649 2650 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5419 2646 2637 2648 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5420 1 2248 2646 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5421 2646 2637 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5422 1 2254 2646 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5423 2645 2640 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5424 0 2649 2637 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5425 0 2650 2649 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5426 0 2545 2650 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5427 2650 2559 672 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5428 662 2535 2650 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5429 2650 2557 647 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5430 657 2541 2650 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5431 0 2652 2651 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5432 2653 2654 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5433 0 2265 2653 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5434 2655 2654 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5435 2652 2265 2655 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5436 2653 2271 2652 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5437 2656 2271 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5438 2657 2652 2656 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5439 1 2652 2651 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5440 2658 2265 2657 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5441 2659 2271 2658 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5442 0 2654 2659 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5443 2656 2265 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5444 0 2654 2656 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5445 2660 2654 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5446 2661 2265 2660 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5447 2652 2654 2661 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5448 2661 2265 2652 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5449 2662 2657 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5450 1 2271 2661 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5451 2657 2652 2663 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5452 2664 2265 2657 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5453 2665 2271 2664 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5454 2654 2666 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5455 2666 2667 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5456 2663 2654 2665 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5457 1 2265 2663 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5458 2663 2654 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5459 1 2271 2663 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5460 2662 2657 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5461 0 2666 2654 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5462 0 2667 2666 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5463 0 2545 2667 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5464 2667 2559 687 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5465 677 2535 2667 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5466 2667 2557 662 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5467 672 2541 2667 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5468 0 2669 2668 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5469 2670 2671 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5470 0 2282 2670 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5471 2672 2671 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5472 2669 2282 2672 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5473 2670 2288 2669 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5474 2673 2288 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5475 2674 2669 2673 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5476 1 2669 2668 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5477 2675 2282 2674 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5478 2676 2288 2675 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5479 0 2671 2676 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5480 2673 2282 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5481 0 2671 2673 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5482 2677 2671 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5483 2678 2282 2677 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5484 2669 2671 2678 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5485 2678 2282 2669 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5486 2679 2674 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5487 1 2288 2678 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5488 2674 2669 2680 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5489 2681 2282 2674 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5490 2682 2288 2681 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5491 2671 2683 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5492 2683 2684 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5493 2680 2671 2682 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5494 1 2282 2680 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5495 2680 2671 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5496 1 2288 2680 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5497 2679 2674 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5498 0 2683 2671 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5499 0 2684 2683 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5500 0 2545 2684 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5501 2684 2559 702 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5502 692 2535 2684 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5503 2684 2557 677 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5504 687 2541 2684 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5505 0 2686 2685 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5506 2687 2688 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5507 0 2299 2687 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5508 2689 2688 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5509 2686 2299 2689 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5510 2687 2305 2686 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5511 2690 2305 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5512 2691 2686 2690 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5513 1 2686 2685 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5514 2692 2299 2691 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5515 2693 2305 2692 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5516 0 2688 2693 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5517 2690 2299 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5518 0 2688 2690 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5519 2694 2688 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5520 2695 2299 2694 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5521 2686 2688 2695 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5522 2695 2299 2686 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5523 2696 2691 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5524 1 2305 2695 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5525 2691 2686 2697 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5526 2698 2299 2691 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5527 2699 2305 2698 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5528 2688 2700 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5529 2700 2701 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5530 2697 2688 2699 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5531 1 2299 2697 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5532 2697 2688 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5533 1 2305 2697 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5534 2696 2691 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5535 0 2700 2688 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5536 0 2701 2700 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5537 0 2545 2701 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5538 2701 2559 717 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5539 707 2535 2701 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5540 2701 2557 692 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5541 702 2541 2701 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5542 0 2703 2702 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5543 2704 2705 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5544 0 2316 2704 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5545 2706 2705 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5546 2703 2316 2706 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5547 2704 2322 2703 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5548 2707 2322 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5549 2708 2703 2707 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5550 1 2703 2702 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5551 2709 2316 2708 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5552 2710 2322 2709 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5553 0 2705 2710 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5554 2707 2316 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5555 0 2705 2707 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5556 2711 2705 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5557 2712 2316 2711 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5558 2703 2705 2712 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5559 2712 2316 2703 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5560 2713 2708 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5561 1 2322 2712 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5562 2708 2703 2714 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5563 2715 2316 2708 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5564 2716 2322 2715 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5565 2705 2717 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5566 2717 2718 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5567 2714 2705 2716 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5568 1 2316 2714 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5569 2714 2705 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5570 1 2322 2714 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5571 2713 2708 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5572 0 2717 2705 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5573 0 2718 2717 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5574 0 2545 2718 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5575 2718 2559 732 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5576 722 2535 2718 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5577 2718 2557 707 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5578 717 2541 2718 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5579 0 2720 2719 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5580 2721 2722 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5581 0 2333 2721 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5582 2723 2722 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5583 2720 2333 2723 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5584 2721 2339 2720 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5585 2724 2339 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5586 2725 2720 2724 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5587 1 2720 2719 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5588 2726 2333 2725 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5589 2727 2339 2726 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5590 0 2722 2727 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5591 2724 2333 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5592 0 2722 2724 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5593 2728 2722 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5594 2729 2333 2728 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5595 2720 2722 2729 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5596 2729 2333 2720 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5597 2730 2725 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5598 1 2339 2729 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5599 2725 2720 2731 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5600 2732 2333 2725 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5601 2733 2339 2732 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5602 2722 2734 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5603 2734 2735 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5604 2731 2722 2733 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5605 1 2333 2731 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5606 2731 2722 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5607 1 2339 2731 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5608 2730 2725 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5609 0 2734 2722 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5610 0 2735 2734 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5611 0 2545 2735 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5612 2735 2559 747 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5613 737 2535 2735 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5614 2735 2557 722 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5615 732 2541 2735 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5616 0 2737 2736 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5617 2738 2739 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5618 0 2350 2738 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5619 2740 2739 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5620 2737 2350 2740 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5621 2738 2356 2737 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5622 2741 2356 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5623 2742 2737 2741 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5624 1 2737 2736 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5625 2743 2350 2742 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5626 2744 2356 2743 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5627 0 2739 2744 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5628 2741 2350 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5629 0 2739 2741 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5630 2745 2739 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5631 2746 2350 2745 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5632 2737 2739 2746 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5633 2746 2350 2737 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5634 2747 2742 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5635 1 2356 2746 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5636 2742 2737 2748 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5637 2749 2350 2742 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5638 2750 2356 2749 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5639 2739 2751 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5640 2751 2752 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5641 2748 2739 2750 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5642 1 2350 2748 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5643 2748 2739 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5644 1 2356 2748 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5645 2747 2742 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5646 0 2751 2739 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5647 0 2752 2751 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5648 0 2545 2752 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5649 2752 2559 762 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5650 752 2535 2752 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5651 2752 2557 737 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5652 747 2541 2752 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5653 0 2754 2753 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5654 2755 2756 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5655 0 2367 2755 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5656 2757 2756 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5657 2754 2367 2757 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5658 2755 2373 2754 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5659 2758 2373 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5660 2759 2754 2758 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5661 1 2754 2753 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5662 2760 2367 2759 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5663 2761 2373 2760 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5664 0 2756 2761 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5665 2758 2367 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5666 0 2756 2758 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5667 2762 2756 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5668 2763 2367 2762 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5669 2754 2756 2763 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5670 2763 2367 2754 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5671 2764 2759 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5672 1 2373 2763 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5673 2759 2754 2765 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5674 2766 2367 2759 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5675 2767 2373 2766 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5676 2756 2768 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5677 2768 2769 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5678 2765 2756 2767 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5679 1 2367 2765 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5680 2765 2756 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5681 1 2373 2765 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5682 2764 2759 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5683 0 2768 2756 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5684 0 2769 2768 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5685 0 2545 2769 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5686 2769 2559 777 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5687 767 2535 2769 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5688 2769 2557 752 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5689 762 2541 2769 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5690 0 2771 2770 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5691 2772 2773 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5692 0 2384 2772 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5693 2774 2773 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5694 2771 2384 2774 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5695 2772 2390 2771 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5696 2775 2390 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5697 2776 2771 2775 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5698 1 2771 2770 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5699 2777 2384 2776 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5700 2778 2390 2777 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5701 0 2773 2778 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5702 2775 2384 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5703 0 2773 2775 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5704 2779 2773 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5705 2780 2384 2779 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5706 2771 2773 2780 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5707 2780 2384 2771 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5708 2781 2776 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5709 1 2390 2780 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5710 2776 2771 2782 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5711 2783 2384 2776 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5712 2784 2390 2783 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5713 2773 2785 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5714 2785 2786 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5715 2782 2773 2784 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5716 1 2384 2782 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5717 2782 2773 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5718 1 2390 2782 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5719 2781 2776 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5720 0 2785 2773 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5721 0 2786 2785 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5722 0 2545 2786 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5723 2786 2559 792 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5724 782 2535 2786 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5725 2786 2557 767 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5726 777 2541 2786 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5727 0 2788 2787 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5728 2789 2790 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5729 0 2401 2789 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5730 2791 2790 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5731 2788 2401 2791 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5732 2789 2407 2788 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5733 2792 2407 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5734 2793 2788 2792 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5735 1 2788 2787 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5736 2794 2401 2793 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5737 2795 2407 2794 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5738 0 2790 2795 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5739 2792 2401 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5740 0 2790 2792 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5741 2796 2790 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5742 2797 2401 2796 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5743 2788 2790 2797 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5744 2797 2401 2788 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5745 2798 2793 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5746 1 2407 2797 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5747 2793 2788 2799 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5748 2800 2401 2793 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5749 2801 2407 2800 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5750 2790 2802 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5751 2802 2803 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5752 2799 2790 2801 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5753 1 2401 2799 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5754 2799 2790 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5755 1 2407 2799 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5756 2798 2793 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5757 0 2802 2790 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5758 0 2803 2802 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5759 0 2545 2803 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5760 2803 2559 807 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5761 797 2535 2803 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5762 2803 2557 782 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5763 792 2541 2803 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5764 0 2805 2804 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5765 2806 2807 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5766 0 2418 2806 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5767 2808 2807 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5768 2805 2418 2808 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5769 2806 2424 2805 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5770 2809 2424 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5771 2810 2805 2809 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5772 1 2805 2804 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5773 2811 2418 2810 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5774 2812 2424 2811 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5775 0 2807 2812 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5776 2809 2418 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5777 0 2807 2809 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5778 2813 2807 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5779 2814 2418 2813 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5780 2805 2807 2814 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5781 2814 2418 2805 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5782 2815 2810 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5783 1 2424 2814 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5784 2810 2805 2816 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5785 2817 2418 2810 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5786 2818 2424 2817 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5787 2807 2819 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5788 2819 2820 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5789 2816 2807 2818 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5790 1 2418 2816 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5791 2816 2807 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5792 1 2424 2816 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5793 2815 2810 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5794 0 2819 2807 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5795 0 2820 2819 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5796 0 2545 2820 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5797 2820 2559 822 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5798 812 2535 2820 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5799 2820 2557 797 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5800 807 2541 2820 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5801 0 2822 2821 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5802 2823 2824 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5803 0 2435 2823 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5804 2825 2824 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5805 2822 2435 2825 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5806 2823 2441 2822 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5807 2826 2441 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5808 2827 2822 2826 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5809 1 2822 2821 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5810 2828 2435 2827 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5811 2829 2441 2828 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5812 0 2824 2829 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5813 2826 2435 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5814 0 2824 2826 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5815 2830 2824 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5816 2831 2435 2830 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5817 2822 2824 2831 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5818 2831 2435 2822 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5819 2832 2827 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5820 1 2441 2831 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5821 2827 2822 2833 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5822 2834 2435 2827 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5823 2835 2441 2834 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5824 2824 2836 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5825 2836 2837 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5826 2833 2824 2835 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5827 1 2435 2833 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5828 2833 2824 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5829 1 2441 2833 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5830 2832 2827 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5831 0 2836 2824 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5832 0 2837 2836 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5833 0 2545 2837 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5834 2837 2559 837 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5835 827 2535 2837 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5836 2837 2557 812 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5837 822 2541 2837 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5838 0 2839 2838 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5839 2840 2841 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5840 0 2452 2840 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5841 2842 2841 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5842 2839 2452 2842 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5843 2840 2458 2839 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5844 2843 2458 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5845 2844 2839 2843 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5846 1 2839 2838 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5847 2845 2452 2844 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5848 2846 2458 2845 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5849 0 2841 2846 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5850 2843 2452 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5851 0 2841 2843 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5852 2847 2841 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5853 2848 2452 2847 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5854 2839 2841 2848 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5855 2848 2452 2839 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5856 2849 2844 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5857 1 2458 2848 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5858 2844 2839 2850 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5859 2851 2452 2844 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5860 2852 2458 2851 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5861 2841 2853 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5862 2853 2854 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5863 2850 2841 2852 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5864 1 2452 2850 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5865 2850 2841 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5866 1 2458 2850 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5867 2849 2844 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5868 0 2853 2841 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5869 0 2854 2853 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5870 0 2545 2854 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5871 2854 2559 868 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5872 842 2535 2854 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m5873 2854 2557 827 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5874 837 2541 2854 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5875 0 2856 2855 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m5876 2857 2858 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m5877 0 2469 2857 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m5878 2859 2858 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m5879 2856 2469 2859 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m5880 2857 2475 2856 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m5881 2860 2475 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m5882 2861 2856 2860 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m5883 1 2856 2855 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m5884 2862 2469 2861 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m5885 2863 2475 2862 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m5886 0 2858 2863 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m5887 2860 2469 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m5888 0 2858 2860 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m5889 2864 2858 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m5890 2865 2469 2864 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m5891 2856 2858 2865 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m5892 2865 2469 2856 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m5893 2866 2861 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m5894 1 2475 2865 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m5895 2861 2856 2867 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m5896 2868 2469 2861 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m5897 2869 2475 2868 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m5898 2858 2870 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m5899 2870 2871 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5900 2867 2858 2869 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m5901 1 2469 2867 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m5902 2867 2858 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m5903 1 2475 2867 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m5904 2866 2861 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m5905 0 2870 2858 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m5906 0 2871 2870 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m5907 0 2545 2871 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m5908 2871 2559 852 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m5909 858 2535 2871 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.036e-11 ad=6.95e-12 ps=1.246e-05 pd=8.18e-06 
+ nrs=0.8 nrd=0.54 
m5910 2871 2557 842 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m5911 868 2541 2871 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m5912 2872 2873 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=5.99e-12 ad=1.348e-11 ps=9.58e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m5913 352 2874 2872 0 nenh l=1.1e-06 w=6.4e-06 
+ as=7.52e-12 ad=5.63e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.14 
m5914 2875 2876 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m5915 2874 2877 2875 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m5916 2878 2879 2874 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m5917 0 2880 2878 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m5918 2876 2880 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m5919 0 2882 2881 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m5920 2883 2877 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m5921 2884 2881 2883 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m5922 2885 2882 2884 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m5923 0 2879 2885 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m5924 2877 2879 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m5925 2886 2884 352 0 nenh l=1.1e-06 w=6.4e-06 
+ as=5.63e-12 ad=7.52e-12 ps=9.02e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m5926 0 2887 2886 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.99e-12 ps=1.275e-05 pd=9.58e-06 
+ nrs=0.29 nrd=0.13 
m5927 2888 2873 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m5928 352 2884 2888 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m5929 2889 2874 352 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m5930 1 2887 2889 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m5931 2890 2876 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m5932 2874 2879 2890 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m5933 2891 2877 2874 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m5934 1 2880 2891 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m5935 2876 2880 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5936 2892 2880 2893 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.57e-11 ps=1.429e-05 pd=2.04e-05 
+ nrs=0.11 nrd=0.12 
m5937 2894 2895 2892 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m5938 2893 2896 2894 0 nenh l=1.1e-06 w=1e-05 
+ as=1.354e-11 ad=8.5e-12 ps=1.759e-05 pd=1.17e-05 
+ nrs=0.14 nrd=0.08 
m5939 0 2896 2893 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m5940 2893 2895 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m5941 0 2895 2897 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m5942 2897 2896 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m5943 2898 2896 2897 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.354e-11 ps=1.17e-05 pd=1.759e-05 
+ nrs=0.08 nrd=0.14 
m5944 2899 2895 2898 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m5945 0 2900 2896 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m5946 2901 2896 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m5947 2879 2895 2901 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m5948 2902 2866 2879 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m5949 0 2900 2902 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m5950 2895 2866 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m5951 2897 2882 2899 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=1.416e-11 ps=2.04e-05 pd=1.429e-05 
+ nrs=0.12 nrd=0.11 
m5952 1 2882 2881 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m5953 2903 2877 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m5954 2884 2882 2903 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m5955 2904 2881 2884 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m5956 1 2879 2904 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m5957 2877 2879 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m5958 2892 2880 2905 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m5959 2906 2895 2892 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m5960 1 2896 2906 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m5961 2905 2896 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m5962 1 2895 2905 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m5963 2907 2895 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m5964 1 2896 2907 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m5965 2908 2896 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m5966 2899 2895 2908 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m5967 2907 2882 2899 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m5968 1 2900 2896 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=3.262e-11 ps=2.039e-05 pd=2.77e-05 
+ nrs=0.21 nrd=0.28 
m5969 2909 2896 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.23e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m5970 2879 2866 2909 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.067e-11 ad=7.27e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.1 
m5971 2910 2895 2879 1 penh l=1.1e-06 w=7.6e-06 
+ as=6.5e-12 ad=9.65e-12 ps=9.55e-06 pd=9.97e-06 
+ nrs=0.11 nrd=0.17 
m5972 1 2900 2910 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.16e-12 ps=1.359e-05 pd=9.05e-06 
+ nrs=0.31 nrd=0.12 
m5973 2895 2866 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.67e-11 ad=2.405e-11 ps=2.77e-05 pd=2.039e-05 
+ nrs=0.23 nrd=0.21 
m5974 1 2911 323 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m5975 2912 2873 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m5976 2911 2913 2912 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m5977 2914 2915 2911 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m5978 1 2887 2914 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m5979 2916 2917 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m5980 2915 2918 2916 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m5981 2919 2920 2915 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m5982 1 2921 2919 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m5983 2917 2921 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m5984 1 2923 2922 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m5985 2924 2920 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m5986 2913 2923 2924 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m5987 2925 2922 2913 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m5988 1 2918 2925 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m5989 2920 2918 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m5990 0 2911 323 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m5991 2926 2873 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=7.37e-12 ad=1.506e-11 ps=1.097e-05 pd=1.425e-05 
+ nrs=0.13 nrd=0.26 
m5992 2911 2915 2926 0 nenh l=1.1e-06 w=6.4e-06 
+ as=8.77e-12 ad=6.21e-12 ps=9.49e-06 pd=9.23e-06 
+ nrs=0.21 nrd=0.15 
m5993 2927 2913 2911 0 nenh l=1.1e-06 w=5.6e-06 
+ as=5.09e-12 ad=7.67e-12 ps=7.68e-06 pd=8.31e-06 
+ nrs=0.16 nrd=0.24 
m5994 0 2887 2927 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=6.17e-12 ps=1.275e-05 pd=9.32e-06 
+ nrs=0.29 nrd=0.13 
m5995 1 2929 2928 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=2.67e-11 ps=2.039e-05 pd=2.77e-05 
+ nrs=0.21 nrd=0.23 
m5996 2930 2931 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=9.84e-12 ad=1.959e-11 ps=1.17e-05 pd=1.661e-05 
+ nrs=0.13 nrd=0.25 
m5997 2918 2929 2930 1 penh l=1.1e-06 w=7.6e-06 
+ as=8.13e-12 ad=8.5e-12 ps=9.97e-06 pd=1.01e-05 
+ nrs=0.14 nrd=0.15 
m5998 2932 2928 2918 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.015e-11 ad=8.99e-12 ps=1.143e-05 pd=1.103e-05 
+ nrs=0.14 nrd=0.13 
m5999 1 2933 2932 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=1.063e-11 ps=1.661e-05 pd=1.197e-05 
+ nrs=0.25 nrd=0.14 
m6000 2931 2933 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m6001 2934 2921 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.55e-11 ad=2.672e-11 ps=1.478e-05 pd=2.265e-05 
+ nrs=0.11 nrd=0.19 
m6002 2880 2929 2934 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.151e-11 ad=1.498e-11 ps=1.394e-05 pd=1.428e-05 
+ nrs=0.09 nrd=0.11 
m6003 2934 2933 2880 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.705e-11 ad=1.309e-11 ps=1.625e-05 pd=1.586e-05 
+ nrs=0.1 nrd=0.08 
m6004 2935 2933 2934 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.498e-11 ps=1.33e-05 pd=1.428e-05 
+ nrs=0.07 nrd=0.11 
m6005 1 2929 2935 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m6006 2936 2929 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m6007 2937 2933 2936 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=9.86e-12 ps=1.428e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m6008 2882 2933 2937 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.309e-11 ad=1.705e-11 ps=1.586e-05 pd=1.625e-05 
+ nrs=0.08 nrd=0.1 
m6009 2937 2929 2882 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=1.151e-11 ps=1.428e-05 pd=1.394e-05 
+ nrs=0.11 nrd=0.09 
m6010 1 2923 2937 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.55e-11 ps=2.265e-05 pd=1.478e-05 
+ nrs=0.19 nrd=0.11 
m6011 2938 2917 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m6012 2915 2920 2938 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m6013 2939 2918 2915 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m6014 0 2921 2939 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m6015 2917 2921 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m6016 0 2923 2922 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m6017 2940 2920 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m6018 2913 2922 2940 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m6019 2941 2923 2913 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m6020 0 2918 2941 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m6021 2920 2918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m6022 0 2929 2928 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m6023 2942 2931 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m6024 2918 2928 2942 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m6025 2943 2929 2918 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m6026 0 2933 2943 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m6027 2931 2933 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.468e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.47 nrd=0.35 
m6028 2880 2921 2944 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.175e-11 ad=1.755e-11 ps=1.429e-05 pd=1.841e-05 
+ nrs=0.09 nrd=0.13 
m6029 2945 2929 2880 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.013e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.1 
m6030 0 2933 2945 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=8.5e-12 ps=1.874e-05 pd=1.17e-05 
+ nrs=0.2 nrd=0.08 
m6031 2944 2933 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=2.299e-11 ps=1.841e-05 pd=2.174e-05 
+ nrs=0.13 nrd=0.17 
m6032 0 2929 2944 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=1.513e-11 ps=1.874e-05 pd=1.587e-05 
+ nrs=0.2 nrd=0.15 
m6033 2946 2929 0 0 nenh l=1.1e-06 w=1e-05 
+ as=1.513e-11 ad=1.982e-11 ps=1.587e-05 pd=1.874e-05 
+ nrs=0.15 nrd=0.2 
m6034 0 2933 2946 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.755e-11 ps=2.174e-05 pd=1.841e-05 
+ nrs=0.17 nrd=0.13 
m6035 2947 2933 0 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.982e-11 ps=1.17e-05 pd=1.874e-05 
+ nrs=0.08 nrd=0.2 
m6036 2882 2929 2947 0 nenh l=1.1e-06 w=1e-05 
+ as=1.013e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.1 nrd=0.08 
m6037 2946 2923 2882 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=1.175e-11 ps=1.841e-05 pd=1.429e-05 
+ nrs=0.13 nrd=0.09 
m6038 2948 2873 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.04e-12 ad=1.348e-11 ps=9.88e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m6039 294 2949 2948 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=5.33e-12 ps=8.5e-06 pd=8.72e-06 
+ nrs=0.19 nrd=0.15 
m6040 2950 2951 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m6041 2949 2952 2950 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m6042 2953 2954 2949 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m6043 0 2955 2953 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m6044 2951 2955 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m6045 0 2957 2956 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m6046 2958 2952 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m6047 2959 2956 2958 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m6048 2960 2957 2959 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m6049 0 2954 2960 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m6050 2952 2954 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m6051 2961 2959 294 0 nenh l=1.1e-06 w=6e-06 
+ as=5.29e-12 ad=6.86e-12 ps=8.61e-06 pd=8.5e-06 
+ nrs=0.15 nrd=0.19 
m6052 0 2887 2961 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=5.65e-12 ps=1.2e-05 pd=9.19e-06 
+ nrs=0.31 nrd=0.14 
m6053 2962 2873 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m6054 294 2959 2962 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m6055 2963 2949 294 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m6056 1 2887 2963 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m6057 2964 2951 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m6058 2949 2954 2964 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m6059 2965 2952 2949 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m6060 1 2955 2965 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m6061 2951 2955 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.308e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.42 nrd=0.4 
m6062 2921 2955 2966 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.57e-11 ps=1.429e-05 pd=2.04e-05 
+ nrs=0.11 nrd=0.12 
m6063 2967 2968 2921 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m6064 2966 2969 2967 0 nenh l=1.1e-06 w=1e-05 
+ as=1.354e-11 ad=8.5e-12 ps=1.759e-05 pd=1.17e-05 
+ nrs=0.14 nrd=0.08 
m6065 0 2969 2966 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m6066 2966 2968 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m6067 0 2968 2970 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m6068 2970 2969 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m6069 2971 2969 2970 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.354e-11 ps=1.17e-05 pd=1.759e-05 
+ nrs=0.08 nrd=0.14 
m6070 2923 2968 2971 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m6071 2970 2957 2923 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=1.416e-11 ps=2.04e-05 pd=1.429e-05 
+ nrs=0.12 nrd=0.11 
m6072 0 2509 2969 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.42e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.45 
m6073 2972 2969 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m6074 2954 2968 2972 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m6075 2973 2503 2954 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m6076 0 2509 2973 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m6077 2968 2503 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.372e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.44 nrd=0.35 
m6078 1 2957 2956 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m6079 2974 2952 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m6080 2959 2957 2974 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m6081 2975 2956 2959 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m6082 1 2954 2975 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m6083 2952 2954 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m6084 2921 2955 2976 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m6085 2977 2968 2921 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m6086 1 2969 2977 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m6087 2976 2969 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m6088 1 2968 2976 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m6089 2978 2968 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m6090 1 2969 2978 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m6091 2979 2969 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m6092 2923 2968 2979 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m6093 2978 2957 2923 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m6094 1 2509 2969 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=2.67e-11 ps=2.039e-05 pd=2.77e-05 
+ nrs=0.21 nrd=0.23 
m6095 2980 2969 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.45e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m6096 2954 2503 2980 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.033e-11 ad=7.53e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.11 
m6097 2981 2968 2954 1 penh l=1.1e-06 w=7.6e-06 
+ as=7.02e-12 ad=9.35e-12 ps=1.01e-05 pd=9.97e-06 
+ nrs=0.12 nrd=0.16 
m6098 1 2509 2981 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=8.12e-12 ps=1.661e-05 pd=1.17e-05 
+ nrs=0.25 nrd=0.1 
m6099 2968 2503 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.67e-11 ad=2.405e-11 ps=2.77e-05 pd=2.039e-05 
+ nrs=0.23 nrd=0.21 
m6100 1 2982 265 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m6101 2983 2873 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m6102 2982 2984 2983 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m6103 2985 2986 2982 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m6104 1 2887 2985 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m6105 2873 2887 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.484e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m6106 1 2887 2873 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.484e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m6107 2887 2987 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m6108 1 2987 2887 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m6109 2986 2984 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.596e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.51 nrd=0.4 
m6110 1 2518 2988 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m6111 2989 2990 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m6112 2984 2518 2989 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m6113 2991 2988 2984 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m6114 1 2521 2991 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m6115 2990 2521 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m6116 0 2982 265 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m6117 2992 2873 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=7.37e-12 ad=1.506e-11 ps=1.097e-05 pd=1.425e-05 
+ nrs=0.13 nrd=0.26 
m6118 2982 2986 2992 0 nenh l=1.1e-06 w=6.4e-06 
+ as=8.77e-12 ad=6.21e-12 ps=9.49e-06 pd=9.23e-06 
+ nrs=0.21 nrd=0.15 
m6119 2993 2984 2982 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=7.67e-12 ps=7.3e-06 pd=8.31e-06 
+ nrs=0.15 nrd=0.24 
m6120 0 2887 2993 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m6121 2873 2887 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.254e-11 ad=1.506e-11 ps=1.09e-05 pd=1.425e-05 
+ nrs=0.22 nrd=0.26 
m6122 0 2887 2873 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.506e-11 ad=1.254e-11 ps=1.425e-05 pd=1.09e-05 
+ nrs=0.26 nrd=0.22 
m6123 2887 2987 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m6124 0 2987 2887 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m6125 2986 2984 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m6126 2994 2518 2955 1 penh l=1.1e-06 w=1.44e-05 
+ as=1.224e-11 ad=4.04e-11 ps=1.61e-05 pd=3.49e-05 
+ nrs=0.06 nrd=0.19 
m6127 1 2521 2994 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.224e-11 ps=2.718e-05 pd=1.61e-05 
+ nrs=0.15 nrd=0.06 
m6128 2987 2995 1 1 penh l=1.1e-06 w=1.44e-05 
+ as=2.376e-11 ad=3.206e-11 ps=1.77e-05 pd=2.718e-05 
+ nrs=0.11 nrd=0.15 
m6129 1 2995 2987 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=2.376e-11 ps=2.718e-05 pd=1.77e-05 
+ nrs=0.15 nrd=0.11 
m6130 2995 2041 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.98e-11 ad=2.672e-11 ps=1.53e-05 pd=2.265e-05 
+ nrs=0.14 nrd=0.19 
m6131 2996 2136 2995 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.02e-11 ad=1.98e-11 ps=1.37e-05 pd=1.53e-05 
+ nrs=0.07 nrd=0.14 
m6132 1 2048 2996 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.02e-11 ps=2.265e-05 pd=1.37e-05 
+ nrs=0.19 nrd=0.07 
m6133 2957 2518 1 1 penh l=1.1e-06 w=1.28e-05 
+ as=1.264e-11 ad=2.85e-11 ps=1.53e-05 pd=2.416e-05 
+ nrs=0.08 nrd=0.17 
m6134 1 2521 2957 1 penh l=1.1e-06 w=1.28e-05 
+ as=2.85e-11 ad=1.264e-11 ps=2.416e-05 pd=1.53e-05 
+ nrs=0.17 nrd=0.08 
m6135 0 2518 2988 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.031e-11 ad=1.586e-11 ps=9.75e-06 pd=1.65e-05 
+ nrs=0.38 nrd=0.59 
m6136 2997 2990 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.32e-12 ad=1.348e-11 ps=9.63e-06 pd=1.275e-05 
+ nrs=0.14 nrd=0.29 
m6137 2984 2988 2997 0 nenh l=1.1e-06 w=5.2e-06 
+ as=8.58e-12 ad=4.84e-12 ps=8.5e-06 pd=7.37e-06 
+ nrs=0.32 nrd=0.18 
m6138 2998 2518 2984 0 nenh l=1.1e-06 w=5.2e-06 
+ as=4.56e-12 ad=8.58e-12 ps=7.37e-06 pd=8.5e-06 
+ nrs=0.17 nrd=0.32 
m6139 0 2521 2998 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.96e-12 ps=1.275e-05 pd=9.63e-06 
+ nrs=0.29 nrd=0.13 
m6140 2990 2521 0 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.031e-11 ps=1.65e-05 pd=9.75e-06 
+ nrs=0.59 nrd=0.38 
m6141 2955 2518 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=1.06e-11 ad=2.061e-11 ps=1.29e-05 pd=1.949e-05 
+ nrs=0.1 nrd=0.19 
m6142 0 2521 2955 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.061e-11 ad=1.06e-11 ps=1.949e-05 pd=1.29e-05 
+ nrs=0.19 nrd=0.1 
m6143 2987 2995 0 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.584e-11 ad=1.903e-11 ps=1.29e-05 pd=1.799e-05 
+ nrs=0.17 nrd=0.21 
m6144 0 2995 2987 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=1.584e-11 ps=1.799e-05 pd=1.29e-05 
+ nrs=0.21 nrd=0.17 
m6145 2999 2041 0 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.955e-11 ad=1.903e-11 ps=1.68e-05 pd=1.799e-05 
+ nrs=0.21 nrd=0.21 
m6146 2995 2136 2999 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.604e-11 ad=1.955e-11 ps=1.303e-05 pd=1.68e-05 
+ nrs=0.17 nrd=0.21 
m6147 2999 2048 2995 0 nenh l=1.1e-06 w=1e-05 
+ as=2.036e-11 ad=1.67e-11 ps=1.75e-05 pd=1.357e-05 
+ nrs=0.2 nrd=0.17 
m6148 3000 2518 2957 0 nenh l=1.1e-06 w=1.28e-05 
+ as=1.088e-11 ad=3.904e-11 ps=1.45e-05 pd=3.17e-05 
+ nrs=0.07 nrd=0.24 
m6149 0 2521 3000 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.088e-11 ps=2.399e-05 pd=1.45e-05 
+ nrs=0.15 nrd=0.07 
m6150 0 3001 2900 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=3.144e-11 ps=2.699e-05 pd=3.25e-05 
+ nrs=0.14 nrd=0.15 
m6151 3002 3003 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.083e-11 ad=3.013e-11 ps=2.27e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m6152 0 2486 3002 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.083e-11 ps=2.849e-05 pd=2.27e-05 
+ nrs=0.13 nrd=0.09 
m6153 3004 3003 0 0 nenh l=1.1e-06 w=1.68e-05 
+ as=1.454e-11 ad=3.33e-11 ps=1.992e-05 pd=3.149e-05 
+ nrs=0.05 nrd=0.12 
m6154 3001 2486 3004 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.246e-11 ps=1.795e-05 pd=1.708e-05 
+ nrs=0.07 nrd=0.06 
m6155 3002 2492 3001 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.919e-11 ad=1.383e-11 ps=2.091e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m6156 3005 2492 0 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.352e-11 ad=2.854e-11 ps=1.61e-05 pd=2.699e-05 
+ nrs=0.07 nrd=0.14 
m6157 3006 3001 3005 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.449e-11 ad=1.352e-11 ps=1.785e-05 pd=1.61e-05 
+ nrs=0.07 nrd=0.07 
m6158 3007 2486 3006 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.489e-11 ps=1.701e-05 pd=1.835e-05 
+ nrs=0.06 nrd=0.07 
m6159 3008 2492 3007 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6160 0 3003 3008 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6161 3005 2486 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.502e-11 ad=3.171e-11 ps=1.789e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6162 0 3003 3005 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.202e-11 ps=2.399e-05 pd=1.431e-05 
+ nrs=0.15 nrd=0.07 
m6163 1 3001 2900 1 penh l=1.1e-06 w=1.8e-05 
+ as=4.008e-11 ad=3.314e-11 ps=3.398e-05 pd=3.89e-05 
+ nrs=0.12 nrd=0.1 
m6164 2929 3006 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6165 3009 3003 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m6166 3010 2486 3009 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m6167 3001 3003 3010 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.615e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6168 3010 2486 3001 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.499e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.06 
m6169 1 2492 3010 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6170 1 3011 2933 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.484e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.47 
m6171 3012 2559 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m6172 3011 2541 3012 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.372e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.44 nrd=0.15 
m6173 1 3013 3003 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.226e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.32 
m6174 3006 3001 3014 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.447e-11 ad=1.386e-11 ps=1.722e-05 pd=1.719e-05 
+ nrs=0.1 nrd=0.1 
m6175 3015 2486 3006 1 penh l=1.1e-06 w=1.88e-05 
+ as=1.621e-11 ad=2.267e-11 ps=2.153e-05 pd=2.698e-05 
+ nrs=0.05 nrd=0.06 
m6176 3016 2492 3015 1 penh l=1.1e-06 w=2.12e-05 
+ as=1.814e-11 ad=1.827e-11 ps=2.344e-05 pd=2.427e-05 
+ nrs=0.04 nrd=0.04 
m6177 3014 3003 3016 1 penh l=1.1e-06 w=2.24e-05 
+ as=2.588e-11 ad=1.916e-11 ps=3.21e-05 pd=2.476e-05 
+ nrs=0.05 nrd=0.04 
m6178 1 2486 3014 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.664e-11 ps=2.718e-05 pd=2.063e-05 
+ nrs=0.15 nrd=0.08 
m6179 3014 3003 1 1 penh l=1.1e-06 w=1.52e-05 
+ as=1.756e-11 ad=3.384e-11 ps=2.178e-05 pd=2.869e-05 
+ nrs=0.08 nrd=0.15 
m6180 1 2492 3014 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.386e-11 ps=2.265e-05 pd=1.719e-05 
+ nrs=0.19 nrd=0.1 
m6181 2929 3006 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.04e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.08 nrd=0.12 
m6182 3013 3017 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.298e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.48 nrd=0.43 
m6183 0 3011 2933 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m6184 3011 2559 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=5.55e-12 ps=6.1e-06 pd=5.25e-06 
+ nrs=0.59 nrd=0.71 
m6185 0 2541 3011 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=4.62e-12 ps=5.25e-06 pd=6.1e-06 
+ nrs=0.71 nrd=0.59 
m6186 0 3013 3003 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.52e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.37 
m6187 0 3017 3013 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6188 0 2545 3017 0 nenh l=1.1e-06 w=3.2e-06 
+ as=6.34e-12 ad=6.09e-12 ps=6e-06 pd=7.29e-06 
+ nrs=0.62 nrd=0.6 
m6189 3017 2559 1 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.098e-11 ps=8.2e-06 pd=1.406e-05 
+ nrs=0.53 nrd=0.85 
m6190 0 2535 3017 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.86e-12 ps=6.75e-06 pd=8.2e-06 
+ nrs=0.55 nrd=0.53 
m6191 3017 2557 858 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.036e-11 ps=8.2e-06 pd=1.246e-05 
+ nrs=0.53 nrd=0.8 
m6192 852 2541 3017 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.86e-12 ps=1.202e-05 pd=8.2e-06 
+ nrs=0.77 nrd=0.53 
m6193 0 3019 3018 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.427e-11 ad=2.196e-11 ps=1.35e-05 pd=2.05e-05 
+ nrs=0.28 nrd=0.42 
m6194 3019 3020 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m6195 0 3022 3021 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.22e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.76 
m6196 3022 3023 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.22e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.76 nrd=0.5 
m6197 1 3019 3018 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m6198 3019 3020 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6199 3024 3025 0 0 nenh l=1.1e-06 w=4e-06 
+ as=6.6e-12 ad=7.93e-12 ps=7.3e-06 pd=7.5e-06 
+ nrs=0.41 nrd=0.5 
m6200 0 3025 3024 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=6.6e-12 ps=7.5e-06 pd=7.3e-06 
+ nrs=0.5 nrd=0.41 
m6201 3026 3027 3025 0 nenh l=1.1e-06 w=8.8e-06 
+ as=7.66e-12 ad=1.964e-11 ps=1.122e-05 pd=2.37e-05 
+ nrs=0.1 nrd=0.25 
m6202 3028 3029 3026 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.4e-12 ps=1.25e-05 pd=1.378e-05 
+ nrs=0.08 nrd=0.08 
m6203 0 2549 3028 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m6204 3030 3027 0 0 nenh l=1.1e-06 w=8.8e-06 
+ as=9.24e-12 ad=1.744e-11 ps=1.13e-05 pd=1.65e-05 
+ nrs=0.12 nrd=0.23 
m6205 0 3031 3030 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.744e-11 ad=9.24e-12 ps=1.65e-05 pd=1.13e-05 
+ nrs=0.23 nrd=0.12 
m6206 3032 3033 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=1.665e-11 ps=1.01e-05 pd=1.575e-05 
+ nrs=0.1 nrd=0.24 
m6207 3034 3035 3032 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.89e-11 ad=7.14e-12 ps=2.29e-05 pd=1.01e-05 
+ nrs=0.27 nrd=0.1 
m6208 1 3022 3021 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=2.358e-11 ps=1.737e-05 pd=2.29e-05 
+ nrs=0.24 nrd=0.28 
m6209 3022 3023 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.358e-11 ad=2.048e-11 ps=2.29e-05 pd=1.737e-05 
+ nrs=0.28 nrd=0.24 
m6210 3024 3025 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.128e-11 ad=2.494e-11 ps=1.37e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m6211 1 3025 3024 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.128e-11 ps=2.114e-05 pd=1.37e-05 
+ nrs=0.2 nrd=0.09 
m6212 3036 3029 3035 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.27e-12 ad=2.16e-11 ps=1.176e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.23 
m6213 3037 2549 3036 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.31e-12 ps=1.25e-05 pd=1.324e-05 
+ nrs=0.08 nrd=0.08 
m6214 0 3038 3037 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m6215 3039 3027 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m6216 3040 3041 3039 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.31e-12 ad=9.18e-12 ps=1.324e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m6217 3033 2538 3040 0 nenh l=1.1e-06 w=9.6e-06 
+ as=2.16e-11 ad=8.27e-12 ps=2.53e-05 pd=1.176e-05 
+ nrs=0.23 nrd=0.09 
m6218 1 3027 3025 1 penh l=1.1e-06 w=9.6e-06 
+ as=2.137e-11 ad=1.315e-11 ps=1.812e-05 pd=1.587e-05 
+ nrs=0.23 nrd=0.14 
m6219 3025 3029 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.26e-11 ad=2.048e-11 ps=1.521e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m6220 1 2549 3025 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.26e-11 ps=1.737e-05 pd=1.521e-05 
+ nrs=0.24 nrd=0.15 
m6221 3042 3027 1 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.194e-11 ad=2.939e-11 ps=1.49e-05 pd=2.492e-05 
+ nrs=0.07 nrd=0.17 
m6222 3030 3031 3042 1 penh l=1.1e-06 w=1.32e-05 
+ as=2.586e-11 ad=1.194e-11 ps=3.01e-05 pd=1.49e-05 
+ nrs=0.15 nrd=0.07 
m6223 3034 3033 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.466e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.07 nrd=0.15 
m6224 1 3035 3034 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.466e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.07 
m6225 1 3029 3035 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m6226 3035 2549 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m6227 1 3038 3035 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m6228 3033 3027 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m6229 1 3041 3033 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m6230 3033 2538 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m6231 3023 3043 1 1 penh l=1.1e-06 w=1e-05 
+ as=2.346e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.23 nrd=0.22 
m6232 3043 3044 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6233 3020 3034 1 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=8.54e-12 ps=7.22e-06 pd=1.094e-05 
+ nrs=0.69 nrd=1.09 
m6234 910 3024 3020 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m6235 3045 3031 3046 1 penh l=1.1e-06 w=1.04e-05 
+ as=8.84e-12 ad=2.596e-11 ps=1.21e-05 pd=2.69e-05 
+ nrs=0.08 nrd=0.24 
m6236 1 3038 3045 1 penh l=1.1e-06 w=1.04e-05 
+ as=2.316e-11 ad=8.84e-12 ps=1.963e-05 pd=1.21e-05 
+ nrs=0.21 nrd=0.08 
m6237 3047 2538 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m6238 1 3041 3047 1 penh l=1.1e-06 w=8e-06 
+ as=1.781e-11 ad=1.075e-11 ps=1.51e-05 pd=1.383e-05 
+ nrs=0.28 nrd=0.17 
m6239 3047 3038 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m6240 3048 3047 1 1 penh l=1.1e-06 w=1e-05 
+ as=1.058e-11 ad=2.227e-11 ps=1.25e-05 pd=1.888e-05 
+ nrs=0.11 nrd=0.22 
m6241 1 3047 3048 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=1.058e-11 ps=1.888e-05 pd=1.25e-05 
+ nrs=0.22 nrd=0.11 
m6242 3044 3048 595 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.74e-12 ps=7.22e-06 pd=9.64e-06 
+ nrs=0.69 nrd=0.99 
m6243 602 3024 3044 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=5.4e-12 ps=9.87e-06 pd=7.22e-06 
+ nrs=1.04 nrd=0.69 
m6244 3044 3030 910 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.88e-12 ps=7.22e-06 pd=1.048e-05 
+ nrs=0.69 nrd=1 
m6245 911 3046 3044 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m6246 0 3034 3044 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.4e-12 ps=5.25e-06 pd=7.22e-06 
+ nrs=0.71 nrd=0.69 
m6247 3049 3041 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=2.405e-11 ps=1.41e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m6248 3031 2538 3049 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.046e-11 ad=1.014e-11 ps=1.25e-05 pd=1.41e-05 
+ nrs=0.09 nrd=0.09 
m6249 3050 2549 3031 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=1.046e-11 ps=1.41e-05 pd=1.25e-05 
+ nrs=0.09 nrd=0.09 
m6250 1 3029 3050 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.014e-11 ps=2.039e-05 pd=1.41e-05 
+ nrs=0.21 nrd=0.09 
m6251 911 3048 3020 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m6252 3020 3030 911 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.91e-12 ps=7.22e-06 pd=1.05e-05 
+ nrs=0.69 nrd=1.01 
m6253 910 3046 3020 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m6254 0 3043 3023 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m6255 0 3044 3043 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m6256 3046 3031 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m6257 0 3038 3046 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m6258 3051 2538 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m6259 3052 3041 3051 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.4e-12 ad=9.18e-12 ps=1.378e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m6260 3047 3038 3052 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.964e-11 ad=7.66e-12 ps=2.37e-05 pd=1.122e-05 
+ nrs=0.25 nrd=0.1 
m6261 3048 3047 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m6262 0 3047 3048 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m6263 3053 3041 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=9.84e-12 ad=2.061e-11 ps=1.319e-05 pd=1.949e-05 
+ nrs=0.09 nrd=0.19 
m6264 3031 2549 3053 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.06e-11 ps=1.29e-05 pd=1.421e-05 
+ nrs=0.09 nrd=0.08 
m6265 3054 2538 3031 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.062e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.08 nrd=0.09 
m6266 0 3029 3054 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.024e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m6267 0 3056 3055 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6268 3057 3058 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6269 0 2529 3057 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6270 3059 3058 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6271 3056 2529 3059 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6272 3057 2532 3056 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6273 3060 2532 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6274 3061 3056 3060 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6275 1 3056 3055 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6276 3062 2529 3061 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6277 3063 2532 3062 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6278 0 3058 3063 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6279 3060 2529 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6280 0 3058 3060 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6281 3064 3058 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6282 3065 2529 3064 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6283 3056 3058 3065 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6284 3065 2529 3056 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6285 3066 3061 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6286 1 2532 3065 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6287 3061 3056 3067 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6288 3068 2529 3061 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6289 3069 2532 3068 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6290 3058 3070 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6291 3070 3071 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6292 3067 3058 3069 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6293 1 2529 3067 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6294 3067 3058 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6295 1 2532 3067 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6296 3066 3061 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6297 0 3070 3058 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6298 0 3071 3070 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6299 0 3034 3071 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6300 3071 3048 612 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6301 601 3024 3071 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6302 3071 3046 602 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.045e-11 ps=8.18e-06 pd=1.269e-05 
+ nrs=0.54 nrd=0.81 
m6303 595 3030 3071 0 nenh l=1.1e-06 w=3.6e-06 
+ as=9.95e-12 ad=6.95e-12 ps=1.239e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6304 0 3073 3072 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6305 3074 3075 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6306 0 2533 3074 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6307 3076 3075 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6308 3073 2533 3076 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6309 3074 2566 3073 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6310 3077 2566 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6311 3078 3073 3077 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6312 1 3073 3072 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6313 3079 2533 3078 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6314 3080 2566 3079 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6315 0 3075 3080 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6316 3077 2533 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6317 0 3075 3077 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6318 3081 3075 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6319 3082 2533 3081 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6320 3073 3075 3082 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6321 3082 2533 3073 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6322 3083 3078 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6323 1 2566 3082 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6324 3078 3073 3084 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6325 3085 2533 3078 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6326 3086 2566 3085 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6327 3075 3087 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6328 3087 3088 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6329 3084 3075 3086 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6330 1 2533 3084 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6331 3084 3075 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6332 1 2566 3084 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6333 3083 3078 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6334 0 3087 3075 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6335 0 3088 3087 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6336 0 3034 3088 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6337 3088 3048 627 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6338 617 3024 3088 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6339 3088 3046 601 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6340 612 3030 3088 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6341 0 3090 3089 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6342 3091 3092 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6343 0 2577 3091 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6344 3093 3092 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6345 3090 2577 3093 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6346 3091 2583 3090 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6347 3094 2583 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6348 3095 3090 3094 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6349 1 3090 3089 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6350 3096 2577 3095 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6351 3097 2583 3096 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6352 0 3092 3097 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6353 3094 2577 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6354 0 3092 3094 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6355 3098 3092 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6356 3099 2577 3098 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6357 3090 3092 3099 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6358 3099 2577 3090 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6359 3100 3095 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6360 1 2583 3099 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6361 3095 3090 3101 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6362 3102 2577 3095 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6363 3103 2583 3102 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6364 3092 3104 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6365 3104 3105 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6366 3101 3092 3103 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6367 1 2577 3101 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6368 3101 3092 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6369 1 2583 3101 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6370 3100 3095 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6371 0 3104 3092 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6372 0 3105 3104 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6373 0 3034 3105 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6374 3105 3048 642 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6375 632 3024 3105 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6376 3105 3046 617 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6377 627 3030 3105 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6378 0 3107 3106 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6379 3108 3109 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6380 0 2594 3108 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6381 3110 3109 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6382 3107 2594 3110 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6383 3108 2600 3107 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6384 3111 2600 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6385 3112 3107 3111 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6386 1 3107 3106 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6387 3113 2594 3112 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6388 3114 2600 3113 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6389 0 3109 3114 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6390 3111 2594 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6391 0 3109 3111 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6392 3115 3109 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6393 3116 2594 3115 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6394 3107 3109 3116 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6395 3116 2594 3107 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6396 3117 3112 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6397 1 2600 3116 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6398 3112 3107 3118 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6399 3119 2594 3112 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6400 3120 2600 3119 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6401 3109 3121 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6402 3121 3122 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6403 3118 3109 3120 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6404 1 2594 3118 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6405 3118 3109 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6406 1 2600 3118 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6407 3117 3112 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6408 0 3121 3109 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6409 0 3122 3121 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6410 0 3034 3122 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6411 3122 3048 657 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6412 647 3024 3122 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6413 3122 3046 632 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6414 642 3030 3122 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6415 0 3124 3123 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6416 3125 3126 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6417 0 2611 3125 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6418 3127 3126 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6419 3124 2611 3127 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6420 3125 2617 3124 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6421 3128 2617 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6422 3129 3124 3128 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6423 1 3124 3123 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6424 3130 2611 3129 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6425 3131 2617 3130 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6426 0 3126 3131 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6427 3128 2611 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6428 0 3126 3128 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6429 3132 3126 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6430 3133 2611 3132 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6431 3124 3126 3133 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6432 3133 2611 3124 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6433 3134 3129 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6434 1 2617 3133 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6435 3129 3124 3135 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6436 3136 2611 3129 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6437 3137 2617 3136 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6438 3126 3138 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6439 3138 3139 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6440 3135 3126 3137 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6441 1 2611 3135 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6442 3135 3126 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6443 1 2617 3135 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6444 3134 3129 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6445 0 3138 3126 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6446 0 3139 3138 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6447 0 3034 3139 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6448 3139 3048 672 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6449 662 3024 3139 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6450 3139 3046 647 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6451 657 3030 3139 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6452 0 3141 3140 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6453 3142 3143 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6454 0 2628 3142 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6455 3144 3143 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6456 3141 2628 3144 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6457 3142 2634 3141 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6458 3145 2634 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6459 3146 3141 3145 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6460 1 3141 3140 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6461 3147 2628 3146 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6462 3148 2634 3147 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6463 0 3143 3148 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6464 3145 2628 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6465 0 3143 3145 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6466 3149 3143 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6467 3150 2628 3149 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6468 3141 3143 3150 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6469 3150 2628 3141 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6470 3151 3146 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6471 1 2634 3150 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6472 3146 3141 3152 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6473 3153 2628 3146 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6474 3154 2634 3153 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6475 3143 3155 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6476 3155 3156 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6477 3152 3143 3154 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6478 1 2628 3152 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6479 3152 3143 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6480 1 2634 3152 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6481 3151 3146 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6482 0 3155 3143 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6483 0 3156 3155 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6484 0 3034 3156 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6485 3156 3048 687 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6486 677 3024 3156 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6487 3156 3046 662 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6488 672 3030 3156 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6489 0 3158 3157 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6490 3159 3160 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6491 0 2645 3159 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6492 3161 3160 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6493 3158 2645 3161 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6494 3159 2651 3158 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6495 3162 2651 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6496 3163 3158 3162 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6497 1 3158 3157 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6498 3164 2645 3163 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6499 3165 2651 3164 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6500 0 3160 3165 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6501 3162 2645 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6502 0 3160 3162 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6503 3166 3160 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6504 3167 2645 3166 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6505 3158 3160 3167 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6506 3167 2645 3158 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6507 3168 3163 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6508 1 2651 3167 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6509 3163 3158 3169 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6510 3170 2645 3163 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6511 3171 2651 3170 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6512 3160 3172 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6513 3172 3173 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6514 3169 3160 3171 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6515 1 2645 3169 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6516 3169 3160 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6517 1 2651 3169 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6518 3168 3163 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6519 0 3172 3160 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6520 0 3173 3172 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6521 0 3034 3173 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6522 3173 3048 702 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6523 692 3024 3173 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6524 3173 3046 677 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6525 687 3030 3173 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6526 0 3175 3174 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6527 3176 3177 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6528 0 2662 3176 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6529 3178 3177 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6530 3175 2662 3178 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6531 3176 2668 3175 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6532 3179 2668 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6533 3180 3175 3179 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6534 1 3175 3174 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6535 3181 2662 3180 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6536 3182 2668 3181 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6537 0 3177 3182 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6538 3179 2662 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6539 0 3177 3179 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6540 3183 3177 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6541 3184 2662 3183 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6542 3175 3177 3184 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6543 3184 2662 3175 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6544 3185 3180 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6545 1 2668 3184 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6546 3180 3175 3186 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6547 3187 2662 3180 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6548 3188 2668 3187 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6549 3177 3189 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6550 3189 3190 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6551 3186 3177 3188 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6552 1 2662 3186 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6553 3186 3177 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6554 1 2668 3186 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6555 3185 3180 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6556 0 3189 3177 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6557 0 3190 3189 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6558 0 3034 3190 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6559 3190 3048 717 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6560 707 3024 3190 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6561 3190 3046 692 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6562 702 3030 3190 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6563 0 3192 3191 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6564 3193 3194 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6565 0 2679 3193 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6566 3195 3194 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6567 3192 2679 3195 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6568 3193 2685 3192 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6569 3196 2685 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6570 3197 3192 3196 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6571 1 3192 3191 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6572 3198 2679 3197 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6573 3199 2685 3198 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6574 0 3194 3199 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6575 3196 2679 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6576 0 3194 3196 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6577 3200 3194 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6578 3201 2679 3200 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6579 3192 3194 3201 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6580 3201 2679 3192 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6581 3202 3197 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6582 1 2685 3201 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6583 3197 3192 3203 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6584 3204 2679 3197 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6585 3205 2685 3204 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6586 3194 3206 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6587 3206 3207 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6588 3203 3194 3205 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6589 1 2679 3203 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6590 3203 3194 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6591 1 2685 3203 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6592 3202 3197 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6593 0 3206 3194 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6594 0 3207 3206 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6595 0 3034 3207 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6596 3207 3048 732 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6597 722 3024 3207 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6598 3207 3046 707 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6599 717 3030 3207 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6600 0 3209 3208 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6601 3210 3211 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6602 0 2696 3210 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6603 3212 3211 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6604 3209 2696 3212 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6605 3210 2702 3209 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6606 3213 2702 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6607 3214 3209 3213 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6608 1 3209 3208 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6609 3215 2696 3214 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6610 3216 2702 3215 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6611 0 3211 3216 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6612 3213 2696 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6613 0 3211 3213 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6614 3217 3211 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6615 3218 2696 3217 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6616 3209 3211 3218 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6617 3218 2696 3209 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6618 3219 3214 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6619 1 2702 3218 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6620 3214 3209 3220 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6621 3221 2696 3214 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6622 3222 2702 3221 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6623 3211 3223 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6624 3223 3224 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6625 3220 3211 3222 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6626 1 2696 3220 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6627 3220 3211 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6628 1 2702 3220 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6629 3219 3214 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6630 0 3223 3211 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6631 0 3224 3223 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6632 0 3034 3224 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6633 3224 3048 747 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6634 737 3024 3224 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6635 3224 3046 722 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6636 732 3030 3224 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6637 0 3226 3225 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6638 3227 3228 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6639 0 2713 3227 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6640 3229 3228 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6641 3226 2713 3229 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6642 3227 2719 3226 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6643 3230 2719 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6644 3231 3226 3230 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6645 1 3226 3225 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6646 3232 2713 3231 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6647 3233 2719 3232 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6648 0 3228 3233 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6649 3230 2713 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6650 0 3228 3230 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6651 3234 3228 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6652 3235 2713 3234 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6653 3226 3228 3235 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6654 3235 2713 3226 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6655 3236 3231 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6656 1 2719 3235 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6657 3231 3226 3237 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6658 3238 2713 3231 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6659 3239 2719 3238 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6660 3228 3240 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6661 3240 3241 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6662 3237 3228 3239 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6663 1 2713 3237 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6664 3237 3228 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6665 1 2719 3237 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6666 3236 3231 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6667 0 3240 3228 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6668 0 3241 3240 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6669 0 3034 3241 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6670 3241 3048 762 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6671 752 3024 3241 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6672 3241 3046 737 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6673 747 3030 3241 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6674 0 3243 3242 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6675 3244 3245 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6676 0 2730 3244 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6677 3246 3245 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6678 3243 2730 3246 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6679 3244 2736 3243 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6680 3247 2736 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6681 3248 3243 3247 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6682 1 3243 3242 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6683 3249 2730 3248 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6684 3250 2736 3249 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6685 0 3245 3250 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6686 3247 2730 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6687 0 3245 3247 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6688 3251 3245 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6689 3252 2730 3251 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6690 3243 3245 3252 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6691 3252 2730 3243 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6692 3253 3248 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6693 1 2736 3252 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6694 3248 3243 3254 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6695 3255 2730 3248 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6696 3256 2736 3255 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6697 3245 3257 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6698 3257 3258 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6699 3254 3245 3256 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6700 1 2730 3254 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6701 3254 3245 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6702 1 2736 3254 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6703 3253 3248 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6704 0 3257 3245 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6705 0 3258 3257 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6706 0 3034 3258 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6707 3258 3048 777 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6708 767 3024 3258 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6709 3258 3046 752 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6710 762 3030 3258 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6711 0 3260 3259 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6712 3261 3262 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6713 0 2747 3261 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6714 3263 3262 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6715 3260 2747 3263 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6716 3261 2753 3260 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6717 3264 2753 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6718 3265 3260 3264 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6719 1 3260 3259 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6720 3266 2747 3265 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6721 3267 2753 3266 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6722 0 3262 3267 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6723 3264 2747 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6724 0 3262 3264 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6725 3268 3262 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6726 3269 2747 3268 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6727 3260 3262 3269 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6728 3269 2747 3260 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6729 3270 3265 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6730 1 2753 3269 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6731 3265 3260 3271 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6732 3272 2747 3265 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6733 3273 2753 3272 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6734 3262 3274 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6735 3274 3275 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6736 3271 3262 3273 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6737 1 2747 3271 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6738 3271 3262 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6739 1 2753 3271 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6740 3270 3265 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6741 0 3274 3262 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6742 0 3275 3274 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6743 0 3034 3275 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6744 3275 3048 792 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6745 782 3024 3275 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6746 3275 3046 767 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6747 777 3030 3275 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6748 0 3277 3276 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6749 3278 3279 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6750 0 2764 3278 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6751 3280 3279 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6752 3277 2764 3280 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6753 3278 2770 3277 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6754 3281 2770 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6755 3282 3277 3281 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6756 1 3277 3276 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6757 3283 2764 3282 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6758 3284 2770 3283 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6759 0 3279 3284 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6760 3281 2764 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6761 0 3279 3281 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6762 3285 3279 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6763 3286 2764 3285 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6764 3277 3279 3286 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6765 3286 2764 3277 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6766 3287 3282 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6767 1 2770 3286 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6768 3282 3277 3288 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6769 3289 2764 3282 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6770 3290 2770 3289 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6771 3279 3291 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6772 3291 3292 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6773 3288 3279 3290 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6774 1 2764 3288 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6775 3288 3279 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6776 1 2770 3288 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6777 3287 3282 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6778 0 3291 3279 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6779 0 3292 3291 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6780 0 3034 3292 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6781 3292 3048 807 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6782 797 3024 3292 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6783 3292 3046 782 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6784 792 3030 3292 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6785 0 3294 3293 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6786 3295 3296 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6787 0 2781 3295 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6788 3297 3296 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6789 3294 2781 3297 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6790 3295 2787 3294 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6791 3298 2787 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6792 3299 3294 3298 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6793 1 3294 3293 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6794 3300 2781 3299 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6795 3301 2787 3300 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6796 0 3296 3301 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6797 3298 2781 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6798 0 3296 3298 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6799 3302 3296 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6800 3303 2781 3302 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6801 3294 3296 3303 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6802 3303 2781 3294 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6803 3304 3299 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6804 1 2787 3303 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6805 3299 3294 3305 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6806 3306 2781 3299 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6807 3307 2787 3306 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6808 3296 3308 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6809 3308 3309 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6810 3305 3296 3307 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6811 1 2781 3305 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6812 3305 3296 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6813 1 2787 3305 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6814 3304 3299 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6815 0 3308 3296 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6816 0 3309 3308 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6817 0 3034 3309 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6818 3309 3048 822 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6819 812 3024 3309 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6820 3309 3046 797 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6821 807 3030 3309 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6822 0 3311 3310 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6823 3312 3313 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6824 0 2798 3312 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6825 3314 3313 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6826 3311 2798 3314 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6827 3312 2804 3311 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6828 3315 2804 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6829 3316 3311 3315 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6830 1 3311 3310 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6831 3317 2798 3316 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6832 3318 2804 3317 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6833 0 3313 3318 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6834 3315 2798 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6835 0 3313 3315 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6836 3319 3313 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6837 3320 2798 3319 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6838 3311 3313 3320 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6839 3320 2798 3311 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6840 3321 3316 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6841 1 2804 3320 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6842 3316 3311 3322 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6843 3323 2798 3316 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6844 3324 2804 3323 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6845 3313 3325 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6846 3325 3326 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6847 3322 3313 3324 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6848 1 2798 3322 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6849 3322 3313 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6850 1 2804 3322 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6851 3321 3316 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6852 0 3325 3313 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6853 0 3326 3325 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6854 0 3034 3326 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6855 3326 3048 837 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6856 827 3024 3326 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6857 3326 3046 812 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6858 822 3030 3326 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6859 0 3328 3327 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6860 3329 3330 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6861 0 2815 3329 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6862 3331 3330 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6863 3328 2815 3331 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6864 3329 2821 3328 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6865 3332 2821 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6866 3333 3328 3332 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6867 1 3328 3327 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6868 3334 2815 3333 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6869 3335 2821 3334 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6870 0 3330 3335 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6871 3332 2815 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6872 0 3330 3332 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6873 3336 3330 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6874 3337 2815 3336 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6875 3328 3330 3337 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6876 3337 2815 3328 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6877 3338 3333 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6878 1 2821 3337 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6879 3333 3328 3339 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6880 3340 2815 3333 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6881 3341 2821 3340 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6882 3330 3342 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6883 3342 3343 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6884 3339 3330 3341 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6885 1 2815 3339 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6886 3339 3330 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6887 1 2821 3339 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6888 3338 3333 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6889 0 3342 3330 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6890 0 3343 3342 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6891 0 3034 3343 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6892 3343 3048 868 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6893 842 3024 3343 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m6894 3343 3046 827 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6895 837 3030 3343 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6896 0 3345 3344 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m6897 3346 3347 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m6898 0 2832 3346 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m6899 3348 3347 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m6900 3345 2832 3348 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m6901 3346 2838 3345 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m6902 3349 2838 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m6903 3350 3345 3349 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m6904 1 3345 3344 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m6905 3351 2832 3350 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m6906 3352 2838 3351 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6907 0 3347 3352 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6908 3349 2832 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6909 0 3347 3349 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m6910 3353 3347 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m6911 3354 2832 3353 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m6912 3345 3347 3354 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6913 3354 2832 3345 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m6914 3355 3350 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6915 1 2838 3354 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6916 3350 3345 3356 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m6917 3357 2832 3350 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m6918 3358 2838 3357 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m6919 3347 3359 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m6920 3359 3360 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6921 3356 3347 3358 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m6922 1 2832 3356 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m6923 3356 3347 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m6924 1 2838 3356 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m6925 3355 3350 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m6926 0 3359 3347 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m6927 0 3360 3359 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6928 0 3034 3360 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m6929 3360 3048 852 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m6930 858 3024 3360 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.036e-11 ad=6.95e-12 ps=1.246e-05 pd=8.18e-06 
+ nrs=0.8 nrd=0.54 
m6931 3360 3046 842 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m6932 868 3030 3360 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m6933 0 3362 3361 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=3.144e-11 ps=2.699e-05 pd=3.25e-05 
+ nrs=0.14 nrd=0.15 
m6934 3363 3364 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.083e-11 ad=3.013e-11 ps=2.27e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m6935 0 2849 3363 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.083e-11 ps=2.849e-05 pd=2.27e-05 
+ nrs=0.13 nrd=0.09 
m6936 3365 3364 0 0 nenh l=1.1e-06 w=1.68e-05 
+ as=1.454e-11 ad=3.33e-11 ps=1.992e-05 pd=3.149e-05 
+ nrs=0.05 nrd=0.12 
m6937 3362 2849 3365 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.246e-11 ps=1.795e-05 pd=1.708e-05 
+ nrs=0.07 nrd=0.06 
m6938 3363 2855 3362 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.919e-11 ad=1.383e-11 ps=2.091e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m6939 3366 2855 0 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.352e-11 ad=2.854e-11 ps=1.61e-05 pd=2.699e-05 
+ nrs=0.07 nrd=0.14 
m6940 3367 3362 3366 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.449e-11 ad=1.352e-11 ps=1.785e-05 pd=1.61e-05 
+ nrs=0.07 nrd=0.07 
m6941 3368 2849 3367 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.489e-11 ps=1.701e-05 pd=1.835e-05 
+ nrs=0.06 nrd=0.07 
m6942 3369 2855 3368 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m6943 0 3364 3369 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m6944 3366 2849 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.502e-11 ad=3.171e-11 ps=1.789e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m6945 0 3364 3366 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.202e-11 ps=2.399e-05 pd=1.431e-05 
+ nrs=0.15 nrd=0.07 
m6946 1 3362 3361 1 penh l=1.1e-06 w=1.8e-05 
+ as=4.008e-11 ad=3.314e-11 ps=3.398e-05 pd=3.89e-05 
+ nrs=0.12 nrd=0.1 
m6947 3370 3367 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m6948 3371 3364 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m6949 3372 2849 3371 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m6950 3362 3364 3372 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.615e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m6951 3372 2849 3362 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.499e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.06 
m6952 1 2855 3372 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m6953 1 3374 3373 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.484e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.47 
m6954 3375 3048 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m6955 3374 3030 3375 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.372e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.44 nrd=0.15 
m6956 1 3376 3364 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.226e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.32 
m6957 3367 3362 3377 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.447e-11 ad=1.386e-11 ps=1.722e-05 pd=1.719e-05 
+ nrs=0.1 nrd=0.1 
m6958 3378 2849 3367 1 penh l=1.1e-06 w=1.88e-05 
+ as=1.621e-11 ad=2.267e-11 ps=2.153e-05 pd=2.698e-05 
+ nrs=0.05 nrd=0.06 
m6959 3379 2855 3378 1 penh l=1.1e-06 w=2.12e-05 
+ as=1.814e-11 ad=1.827e-11 ps=2.344e-05 pd=2.427e-05 
+ nrs=0.04 nrd=0.04 
m6960 3377 3364 3379 1 penh l=1.1e-06 w=2.24e-05 
+ as=2.588e-11 ad=1.916e-11 ps=3.21e-05 pd=2.476e-05 
+ nrs=0.05 nrd=0.04 
m6961 1 2849 3377 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.664e-11 ps=2.718e-05 pd=2.063e-05 
+ nrs=0.15 nrd=0.08 
m6962 3377 3364 1 1 penh l=1.1e-06 w=1.52e-05 
+ as=1.756e-11 ad=3.384e-11 ps=2.178e-05 pd=2.869e-05 
+ nrs=0.08 nrd=0.15 
m6963 1 2855 3377 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.386e-11 ps=2.265e-05 pd=1.719e-05 
+ nrs=0.19 nrd=0.1 
m6964 3370 3367 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.04e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.08 nrd=0.12 
m6965 3376 3380 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.298e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.48 nrd=0.43 
m6966 0 3374 3373 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m6967 3374 3048 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=5.55e-12 ps=6.1e-06 pd=5.25e-06 
+ nrs=0.59 nrd=0.71 
m6968 0 3030 3374 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=4.62e-12 ps=5.25e-06 pd=6.1e-06 
+ nrs=0.71 nrd=0.59 
m6969 0 3376 3364 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.52e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.37 
m6970 0 3380 3376 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m6971 0 3034 3380 0 nenh l=1.1e-06 w=3.2e-06 
+ as=6.34e-12 ad=6.09e-12 ps=6e-06 pd=7.29e-06 
+ nrs=0.62 nrd=0.6 
m6972 3380 3048 1 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.098e-11 ps=8.2e-06 pd=1.406e-05 
+ nrs=0.53 nrd=0.85 
m6973 0 3024 3380 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.86e-12 ps=6.75e-06 pd=8.2e-06 
+ nrs=0.55 nrd=0.53 
m6974 3380 3046 858 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.036e-11 ps=8.2e-06 pd=1.246e-05 
+ nrs=0.53 nrd=0.8 
m6975 852 3030 3380 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.86e-12 ps=1.202e-05 pd=8.2e-06 
+ nrs=0.77 nrd=0.53 
m6976 0 3382 3381 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.427e-11 ad=2.196e-11 ps=1.35e-05 pd=2.05e-05 
+ nrs=0.28 nrd=0.42 
m6977 3382 3383 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m6978 0 3385 3384 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.22e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.76 
m6979 3385 3386 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.22e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.76 nrd=0.5 
m6980 1 3382 3381 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m6981 3382 3383 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m6982 3387 3388 0 0 nenh l=1.1e-06 w=4e-06 
+ as=6.6e-12 ad=7.93e-12 ps=7.3e-06 pd=7.5e-06 
+ nrs=0.41 nrd=0.5 
m6983 0 3388 3387 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=6.6e-12 ps=7.5e-06 pd=7.3e-06 
+ nrs=0.5 nrd=0.41 
m6984 3389 3390 3388 0 nenh l=1.1e-06 w=8.8e-06 
+ as=7.66e-12 ad=1.964e-11 ps=1.122e-05 pd=2.37e-05 
+ nrs=0.1 nrd=0.25 
m6985 3391 3392 3389 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.4e-12 ps=1.25e-05 pd=1.378e-05 
+ nrs=0.08 nrd=0.08 
m6986 0 3038 3391 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m6987 3393 3390 0 0 nenh l=1.1e-06 w=8.8e-06 
+ as=9.24e-12 ad=1.744e-11 ps=1.13e-05 pd=1.65e-05 
+ nrs=0.12 nrd=0.23 
m6988 0 3394 3393 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.744e-11 ad=9.24e-12 ps=1.65e-05 pd=1.13e-05 
+ nrs=0.23 nrd=0.12 
m6989 3395 3396 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=1.665e-11 ps=1.01e-05 pd=1.575e-05 
+ nrs=0.1 nrd=0.24 
m6990 3397 3398 3395 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.89e-11 ad=7.14e-12 ps=2.29e-05 pd=1.01e-05 
+ nrs=0.27 nrd=0.1 
m6991 1 3385 3384 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=2.358e-11 ps=1.737e-05 pd=2.29e-05 
+ nrs=0.24 nrd=0.28 
m6992 3385 3386 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.358e-11 ad=2.048e-11 ps=2.29e-05 pd=1.737e-05 
+ nrs=0.28 nrd=0.24 
m6993 3387 3388 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.128e-11 ad=2.494e-11 ps=1.37e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m6994 1 3388 3387 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.128e-11 ps=2.114e-05 pd=1.37e-05 
+ nrs=0.2 nrd=0.09 
m6995 3399 3392 3398 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.27e-12 ad=2.16e-11 ps=1.176e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.23 
m6996 3400 3038 3399 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.31e-12 ps=1.25e-05 pd=1.324e-05 
+ nrs=0.08 nrd=0.08 
m6997 0 3401 3400 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m6998 3402 3390 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m6999 3403 3404 3402 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.31e-12 ad=9.18e-12 ps=1.324e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m7000 3396 3027 3403 0 nenh l=1.1e-06 w=9.6e-06 
+ as=2.16e-11 ad=8.27e-12 ps=2.53e-05 pd=1.176e-05 
+ nrs=0.23 nrd=0.09 
m7001 1 3390 3388 1 penh l=1.1e-06 w=9.6e-06 
+ as=2.137e-11 ad=1.315e-11 ps=1.812e-05 pd=1.587e-05 
+ nrs=0.23 nrd=0.14 
m7002 3388 3392 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.26e-11 ad=2.048e-11 ps=1.521e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m7003 1 3038 3388 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.26e-11 ps=1.737e-05 pd=1.521e-05 
+ nrs=0.24 nrd=0.15 
m7004 3405 3390 1 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.194e-11 ad=2.939e-11 ps=1.49e-05 pd=2.492e-05 
+ nrs=0.07 nrd=0.17 
m7005 3393 3394 3405 1 penh l=1.1e-06 w=1.32e-05 
+ as=2.586e-11 ad=1.194e-11 ps=3.01e-05 pd=1.49e-05 
+ nrs=0.15 nrd=0.07 
m7006 3397 3396 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.466e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.07 nrd=0.15 
m7007 1 3398 3397 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.466e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.07 
m7008 1 3392 3398 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m7009 3398 3038 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m7010 1 3401 3398 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m7011 3396 3390 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m7012 1 3404 3396 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m7013 3396 3027 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m7014 3386 3406 1 1 penh l=1.1e-06 w=1e-05 
+ as=2.346e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.23 nrd=0.22 
m7015 3406 3407 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7016 3383 3397 1 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=8.54e-12 ps=7.22e-06 pd=1.094e-05 
+ nrs=0.69 nrd=1.09 
m7017 910 3387 3383 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m7018 3408 3394 3409 1 penh l=1.1e-06 w=1.04e-05 
+ as=8.84e-12 ad=2.596e-11 ps=1.21e-05 pd=2.69e-05 
+ nrs=0.08 nrd=0.24 
m7019 1 3401 3408 1 penh l=1.1e-06 w=1.04e-05 
+ as=2.316e-11 ad=8.84e-12 ps=1.963e-05 pd=1.21e-05 
+ nrs=0.21 nrd=0.08 
m7020 3410 3027 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m7021 1 3404 3410 1 penh l=1.1e-06 w=8e-06 
+ as=1.781e-11 ad=1.075e-11 ps=1.51e-05 pd=1.383e-05 
+ nrs=0.28 nrd=0.17 
m7022 3410 3401 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m7023 3411 3410 1 1 penh l=1.1e-06 w=1e-05 
+ as=1.058e-11 ad=2.227e-11 ps=1.25e-05 pd=1.888e-05 
+ nrs=0.11 nrd=0.22 
m7024 1 3410 3411 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=1.058e-11 ps=1.888e-05 pd=1.25e-05 
+ nrs=0.22 nrd=0.11 
m7025 3407 3411 595 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.74e-12 ps=7.22e-06 pd=9.64e-06 
+ nrs=0.69 nrd=0.99 
m7026 602 3387 3407 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=5.4e-12 ps=9.87e-06 pd=7.22e-06 
+ nrs=1.04 nrd=0.69 
m7027 3407 3393 910 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.88e-12 ps=7.22e-06 pd=1.048e-05 
+ nrs=0.69 nrd=1 
m7028 911 3409 3407 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m7029 0 3397 3407 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.4e-12 ps=5.25e-06 pd=7.22e-06 
+ nrs=0.71 nrd=0.69 
m7030 3412 3404 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=2.405e-11 ps=1.41e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m7031 3394 3027 3412 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.046e-11 ad=1.014e-11 ps=1.25e-05 pd=1.41e-05 
+ nrs=0.09 nrd=0.09 
m7032 3413 3038 3394 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=1.046e-11 ps=1.41e-05 pd=1.25e-05 
+ nrs=0.09 nrd=0.09 
m7033 1 3392 3413 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.014e-11 ps=2.039e-05 pd=1.41e-05 
+ nrs=0.21 nrd=0.09 
m7034 911 3411 3383 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m7035 3383 3393 911 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.91e-12 ps=7.22e-06 pd=1.05e-05 
+ nrs=0.69 nrd=1.01 
m7036 910 3409 3383 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m7037 0 3406 3386 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m7038 0 3407 3406 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m7039 3409 3394 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m7040 0 3401 3409 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m7041 3414 3027 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m7042 3415 3404 3414 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.4e-12 ad=9.18e-12 ps=1.378e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m7043 3410 3401 3415 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.964e-11 ad=7.66e-12 ps=2.37e-05 pd=1.122e-05 
+ nrs=0.25 nrd=0.1 
m7044 3411 3410 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m7045 0 3410 3411 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m7046 3416 3404 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=9.84e-12 ad=2.061e-11 ps=1.319e-05 pd=1.949e-05 
+ nrs=0.09 nrd=0.19 
m7047 3394 3038 3416 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.06e-11 ps=1.29e-05 pd=1.421e-05 
+ nrs=0.09 nrd=0.08 
m7048 3417 3027 3394 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.062e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.08 nrd=0.09 
m7049 0 3392 3417 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.024e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m7050 0 3419 3418 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7051 3420 3421 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7052 0 3018 3420 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7053 3422 3421 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7054 3419 3018 3422 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7055 3420 3021 3419 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7056 3423 3021 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7057 3424 3419 3423 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7058 1 3419 3418 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7059 3425 3018 3424 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7060 3426 3021 3425 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7061 0 3421 3426 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7062 3423 3018 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7063 0 3421 3423 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7064 3427 3421 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7065 3428 3018 3427 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7066 3419 3421 3428 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7067 3428 3018 3419 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7068 3429 3424 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7069 1 3021 3428 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7070 3424 3419 3430 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7071 3431 3018 3424 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7072 3432 3021 3431 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7073 3421 3433 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7074 3433 3434 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7075 3430 3421 3432 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7076 1 3018 3430 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7077 3430 3421 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7078 1 3021 3430 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7079 3429 3424 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7080 0 3433 3421 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7081 0 3434 3433 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7082 0 3397 3434 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7083 3434 3411 612 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7084 601 3387 3434 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7085 3434 3409 602 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.045e-11 ps=8.18e-06 pd=1.269e-05 
+ nrs=0.54 nrd=0.81 
m7086 595 3393 3434 0 nenh l=1.1e-06 w=3.6e-06 
+ as=9.95e-12 ad=6.95e-12 ps=1.239e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7087 0 3436 3435 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7088 3437 3438 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7089 0 3022 3437 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7090 3439 3438 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7091 3436 3022 3439 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7092 3437 3055 3436 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7093 3440 3055 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7094 3441 3436 3440 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7095 1 3436 3435 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7096 3442 3022 3441 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7097 3443 3055 3442 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7098 0 3438 3443 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7099 3440 3022 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7100 0 3438 3440 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7101 3444 3438 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7102 3445 3022 3444 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7103 3436 3438 3445 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7104 3445 3022 3436 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7105 3446 3441 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7106 1 3055 3445 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7107 3441 3436 3447 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7108 3448 3022 3441 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7109 3449 3055 3448 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7110 3438 3450 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7111 3450 3451 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7112 3447 3438 3449 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7113 1 3022 3447 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7114 3447 3438 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7115 1 3055 3447 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7116 3446 3441 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7117 0 3450 3438 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7118 0 3451 3450 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7119 0 3397 3451 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7120 3451 3411 627 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7121 617 3387 3451 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7122 3451 3409 601 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7123 612 3393 3451 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7124 0 3453 3452 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7125 3454 3455 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7126 0 3066 3454 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7127 3456 3455 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7128 3453 3066 3456 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7129 3454 3072 3453 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7130 3457 3072 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7131 3458 3453 3457 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7132 1 3453 3452 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7133 3459 3066 3458 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7134 3460 3072 3459 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7135 0 3455 3460 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7136 3457 3066 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7137 0 3455 3457 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7138 3461 3455 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7139 3462 3066 3461 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7140 3453 3455 3462 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7141 3462 3066 3453 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7142 3463 3458 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7143 1 3072 3462 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7144 3458 3453 3464 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7145 3465 3066 3458 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7146 3466 3072 3465 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7147 3455 3467 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7148 3467 3468 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7149 3464 3455 3466 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7150 1 3066 3464 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7151 3464 3455 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7152 1 3072 3464 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7153 3463 3458 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7154 0 3467 3455 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7155 0 3468 3467 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7156 0 3397 3468 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7157 3468 3411 642 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7158 632 3387 3468 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7159 3468 3409 617 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7160 627 3393 3468 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7161 0 3470 3469 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7162 3471 3472 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7163 0 3083 3471 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7164 3473 3472 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7165 3470 3083 3473 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7166 3471 3089 3470 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7167 3474 3089 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7168 3475 3470 3474 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7169 1 3470 3469 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7170 3476 3083 3475 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7171 3477 3089 3476 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7172 0 3472 3477 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7173 3474 3083 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7174 0 3472 3474 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7175 3478 3472 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7176 3479 3083 3478 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7177 3470 3472 3479 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7178 3479 3083 3470 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7179 3480 3475 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7180 1 3089 3479 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7181 3475 3470 3481 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7182 3482 3083 3475 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7183 3483 3089 3482 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7184 3472 3484 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7185 3484 3485 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7186 3481 3472 3483 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7187 1 3083 3481 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7188 3481 3472 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7189 1 3089 3481 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7190 3480 3475 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7191 0 3484 3472 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7192 0 3485 3484 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7193 0 3397 3485 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7194 3485 3411 657 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7195 647 3387 3485 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7196 3485 3409 632 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7197 642 3393 3485 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7198 0 3487 3486 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7199 3488 3489 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7200 0 3100 3488 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7201 3490 3489 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7202 3487 3100 3490 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7203 3488 3106 3487 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7204 3491 3106 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7205 3492 3487 3491 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7206 1 3487 3486 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7207 3493 3100 3492 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7208 3494 3106 3493 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7209 0 3489 3494 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7210 3491 3100 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7211 0 3489 3491 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7212 3495 3489 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7213 3496 3100 3495 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7214 3487 3489 3496 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7215 3496 3100 3487 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7216 3497 3492 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7217 1 3106 3496 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7218 3492 3487 3498 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7219 3499 3100 3492 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7220 3500 3106 3499 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7221 3489 3501 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7222 3501 3502 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7223 3498 3489 3500 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7224 1 3100 3498 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7225 3498 3489 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7226 1 3106 3498 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7227 3497 3492 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7228 0 3501 3489 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7229 0 3502 3501 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7230 0 3397 3502 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7231 3502 3411 672 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7232 662 3387 3502 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7233 3502 3409 647 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7234 657 3393 3502 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7235 0 3504 3503 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7236 3505 3506 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7237 0 3117 3505 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7238 3507 3506 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7239 3504 3117 3507 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7240 3505 3123 3504 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7241 3508 3123 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7242 3509 3504 3508 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7243 1 3504 3503 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7244 3510 3117 3509 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7245 3511 3123 3510 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7246 0 3506 3511 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7247 3508 3117 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7248 0 3506 3508 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7249 3512 3506 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7250 3513 3117 3512 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7251 3504 3506 3513 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7252 3513 3117 3504 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7253 3514 3509 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7254 1 3123 3513 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7255 3509 3504 3515 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7256 3516 3117 3509 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7257 3517 3123 3516 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7258 3506 3518 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7259 3518 3519 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7260 3515 3506 3517 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7261 1 3117 3515 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7262 3515 3506 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7263 1 3123 3515 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7264 3514 3509 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7265 0 3518 3506 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7266 0 3519 3518 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7267 0 3397 3519 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7268 3519 3411 687 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7269 677 3387 3519 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7270 3519 3409 662 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7271 672 3393 3519 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7272 0 3521 3520 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7273 3522 3523 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7274 0 3134 3522 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7275 3524 3523 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7276 3521 3134 3524 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7277 3522 3140 3521 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7278 3525 3140 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7279 3526 3521 3525 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7280 1 3521 3520 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7281 3527 3134 3526 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7282 3528 3140 3527 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7283 0 3523 3528 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7284 3525 3134 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7285 0 3523 3525 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7286 3529 3523 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7287 3530 3134 3529 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7288 3521 3523 3530 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7289 3530 3134 3521 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7290 3531 3526 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7291 1 3140 3530 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7292 3526 3521 3532 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7293 3533 3134 3526 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7294 3534 3140 3533 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7295 3523 3535 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7296 3535 3536 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7297 3532 3523 3534 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7298 1 3134 3532 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7299 3532 3523 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7300 1 3140 3532 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7301 3531 3526 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7302 0 3535 3523 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7303 0 3536 3535 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7304 0 3397 3536 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7305 3536 3411 702 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7306 692 3387 3536 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7307 3536 3409 677 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7308 687 3393 3536 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7309 0 3538 3537 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7310 3539 3540 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7311 0 3151 3539 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7312 3541 3540 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7313 3538 3151 3541 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7314 3539 3157 3538 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7315 3542 3157 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7316 3543 3538 3542 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7317 1 3538 3537 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7318 3544 3151 3543 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7319 3545 3157 3544 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7320 0 3540 3545 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7321 3542 3151 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7322 0 3540 3542 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7323 3546 3540 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7324 3547 3151 3546 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7325 3538 3540 3547 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7326 3547 3151 3538 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7327 3548 3543 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7328 1 3157 3547 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7329 3543 3538 3549 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7330 3550 3151 3543 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7331 3551 3157 3550 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7332 3540 3552 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7333 3552 3553 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7334 3549 3540 3551 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7335 1 3151 3549 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7336 3549 3540 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7337 1 3157 3549 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7338 3548 3543 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7339 0 3552 3540 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7340 0 3553 3552 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7341 0 3397 3553 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7342 3553 3411 717 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7343 707 3387 3553 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7344 3553 3409 692 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7345 702 3393 3553 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7346 0 3555 3554 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7347 3556 3557 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7348 0 3168 3556 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7349 3558 3557 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7350 3555 3168 3558 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7351 3556 3174 3555 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7352 3559 3174 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7353 3560 3555 3559 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7354 1 3555 3554 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7355 3561 3168 3560 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7356 3562 3174 3561 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7357 0 3557 3562 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7358 3559 3168 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7359 0 3557 3559 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7360 3563 3557 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7361 3564 3168 3563 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7362 3555 3557 3564 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7363 3564 3168 3555 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7364 3565 3560 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7365 1 3174 3564 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7366 3560 3555 3566 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7367 3567 3168 3560 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7368 3568 3174 3567 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7369 3557 3569 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7370 3569 3570 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7371 3566 3557 3568 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7372 1 3168 3566 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7373 3566 3557 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7374 1 3174 3566 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7375 3565 3560 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7376 0 3569 3557 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7377 0 3570 3569 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7378 0 3397 3570 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7379 3570 3411 732 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7380 722 3387 3570 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7381 3570 3409 707 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7382 717 3393 3570 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7383 0 3572 3571 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7384 3573 3574 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7385 0 3185 3573 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7386 3575 3574 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7387 3572 3185 3575 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7388 3573 3191 3572 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7389 3576 3191 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7390 3577 3572 3576 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7391 1 3572 3571 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7392 3578 3185 3577 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7393 3579 3191 3578 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7394 0 3574 3579 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7395 3576 3185 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7396 0 3574 3576 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7397 3580 3574 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7398 3581 3185 3580 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7399 3572 3574 3581 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7400 3581 3185 3572 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7401 3582 3577 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7402 1 3191 3581 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7403 3577 3572 3583 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7404 3584 3185 3577 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7405 3585 3191 3584 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7406 3574 3586 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7407 3586 3587 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7408 3583 3574 3585 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7409 1 3185 3583 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7410 3583 3574 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7411 1 3191 3583 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7412 3582 3577 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7413 0 3586 3574 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7414 0 3587 3586 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7415 0 3397 3587 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7416 3587 3411 747 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7417 737 3387 3587 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7418 3587 3409 722 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7419 732 3393 3587 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7420 0 3589 3588 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7421 3590 3591 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7422 0 3202 3590 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7423 3592 3591 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7424 3589 3202 3592 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7425 3590 3208 3589 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7426 3593 3208 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7427 3594 3589 3593 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7428 1 3589 3588 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7429 3595 3202 3594 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7430 3596 3208 3595 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7431 0 3591 3596 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7432 3593 3202 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7433 0 3591 3593 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7434 3597 3591 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7435 3598 3202 3597 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7436 3589 3591 3598 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7437 3598 3202 3589 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7438 3599 3594 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7439 1 3208 3598 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7440 3594 3589 3600 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7441 3601 3202 3594 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7442 3602 3208 3601 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7443 3591 3603 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7444 3603 3604 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7445 3600 3591 3602 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7446 1 3202 3600 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7447 3600 3591 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7448 1 3208 3600 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7449 3599 3594 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7450 0 3603 3591 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7451 0 3604 3603 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7452 0 3397 3604 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7453 3604 3411 762 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7454 752 3387 3604 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7455 3604 3409 737 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7456 747 3393 3604 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7457 0 3606 3605 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7458 3607 3608 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7459 0 3219 3607 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7460 3609 3608 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7461 3606 3219 3609 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7462 3607 3225 3606 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7463 3610 3225 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7464 3611 3606 3610 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7465 1 3606 3605 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7466 3612 3219 3611 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7467 3613 3225 3612 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7468 0 3608 3613 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7469 3610 3219 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7470 0 3608 3610 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7471 3614 3608 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7472 3615 3219 3614 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7473 3606 3608 3615 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7474 3615 3219 3606 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7475 3616 3611 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7476 1 3225 3615 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7477 3611 3606 3617 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7478 3618 3219 3611 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7479 3619 3225 3618 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7480 3608 3620 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7481 3620 3621 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7482 3617 3608 3619 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7483 1 3219 3617 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7484 3617 3608 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7485 1 3225 3617 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7486 3616 3611 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7487 0 3620 3608 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7488 0 3621 3620 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7489 0 3397 3621 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7490 3621 3411 777 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7491 767 3387 3621 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7492 3621 3409 752 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7493 762 3393 3621 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7494 0 3623 3622 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7495 3624 3625 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7496 0 3236 3624 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7497 3626 3625 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7498 3623 3236 3626 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7499 3624 3242 3623 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7500 3627 3242 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7501 3628 3623 3627 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7502 1 3623 3622 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7503 3629 3236 3628 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7504 3630 3242 3629 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7505 0 3625 3630 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7506 3627 3236 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7507 0 3625 3627 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7508 3631 3625 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7509 3632 3236 3631 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7510 3623 3625 3632 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7511 3632 3236 3623 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7512 3633 3628 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7513 1 3242 3632 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7514 3628 3623 3634 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7515 3635 3236 3628 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7516 3636 3242 3635 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7517 3625 3637 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7518 3637 3638 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7519 3634 3625 3636 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7520 1 3236 3634 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7521 3634 3625 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7522 1 3242 3634 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7523 3633 3628 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7524 0 3637 3625 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7525 0 3638 3637 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7526 0 3397 3638 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7527 3638 3411 792 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7528 782 3387 3638 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7529 3638 3409 767 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7530 777 3393 3638 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7531 0 3640 3639 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7532 3641 3642 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7533 0 3253 3641 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7534 3643 3642 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7535 3640 3253 3643 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7536 3641 3259 3640 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7537 3644 3259 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7538 3645 3640 3644 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7539 1 3640 3639 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7540 3646 3253 3645 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7541 3647 3259 3646 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7542 0 3642 3647 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7543 3644 3253 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7544 0 3642 3644 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7545 3648 3642 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7546 3649 3253 3648 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7547 3640 3642 3649 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7548 3649 3253 3640 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7549 3650 3645 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7550 1 3259 3649 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7551 3645 3640 3651 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7552 3652 3253 3645 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7553 3653 3259 3652 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7554 3642 3654 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7555 3654 3655 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7556 3651 3642 3653 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7557 1 3253 3651 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7558 3651 3642 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7559 1 3259 3651 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7560 3650 3645 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7561 0 3654 3642 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7562 0 3655 3654 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7563 0 3397 3655 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7564 3655 3411 807 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7565 797 3387 3655 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7566 3655 3409 782 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7567 792 3393 3655 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7568 0 3657 3656 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7569 3658 3659 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7570 0 3270 3658 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7571 3660 3659 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7572 3657 3270 3660 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7573 3658 3276 3657 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7574 3661 3276 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7575 3662 3657 3661 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7576 1 3657 3656 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7577 3663 3270 3662 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7578 3664 3276 3663 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7579 0 3659 3664 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7580 3661 3270 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7581 0 3659 3661 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7582 3665 3659 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7583 3666 3270 3665 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7584 3657 3659 3666 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7585 3666 3270 3657 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7586 3667 3662 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7587 1 3276 3666 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7588 3662 3657 3668 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7589 3669 3270 3662 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7590 3670 3276 3669 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7591 3659 3671 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7592 3671 3672 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7593 3668 3659 3670 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7594 1 3270 3668 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7595 3668 3659 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7596 1 3276 3668 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7597 3667 3662 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7598 0 3671 3659 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7599 0 3672 3671 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7600 0 3397 3672 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7601 3672 3411 822 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7602 812 3387 3672 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7603 3672 3409 797 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7604 807 3393 3672 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7605 0 3674 3673 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7606 3675 3676 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7607 0 3287 3675 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7608 3677 3676 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7609 3674 3287 3677 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7610 3675 3293 3674 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7611 3678 3293 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7612 3679 3674 3678 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7613 1 3674 3673 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7614 3680 3287 3679 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7615 3681 3293 3680 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7616 0 3676 3681 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7617 3678 3287 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7618 0 3676 3678 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7619 3682 3676 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7620 3683 3287 3682 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7621 3674 3676 3683 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7622 3683 3287 3674 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7623 3684 3679 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7624 1 3293 3683 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7625 3679 3674 3685 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7626 3686 3287 3679 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7627 3687 3293 3686 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7628 3676 3688 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7629 3688 3689 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7630 3685 3676 3687 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7631 1 3287 3685 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7632 3685 3676 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7633 1 3293 3685 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7634 3684 3679 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7635 0 3688 3676 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7636 0 3689 3688 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7637 0 3397 3689 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7638 3689 3411 837 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7639 827 3387 3689 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7640 3689 3409 812 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7641 822 3393 3689 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7642 0 3691 3690 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7643 3692 3693 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7644 0 3304 3692 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7645 3694 3693 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7646 3691 3304 3694 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7647 3692 3310 3691 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7648 3695 3310 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7649 3696 3691 3695 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7650 1 3691 3690 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7651 3697 3304 3696 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7652 3698 3310 3697 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7653 0 3693 3698 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7654 3695 3304 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7655 0 3693 3695 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7656 3699 3693 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7657 3700 3304 3699 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7658 3691 3693 3700 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7659 3700 3304 3691 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7660 3701 3696 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7661 1 3310 3700 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7662 3696 3691 3702 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7663 3703 3304 3696 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7664 3704 3310 3703 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7665 3693 3705 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7666 3705 3706 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7667 3702 3693 3704 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7668 1 3304 3702 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7669 3702 3693 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7670 1 3310 3702 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7671 3701 3696 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7672 0 3705 3693 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7673 0 3706 3705 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7674 0 3397 3706 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7675 3706 3411 868 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7676 842 3387 3706 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m7677 3706 3409 827 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7678 837 3393 3706 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7679 0 3708 3707 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m7680 3709 3710 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m7681 0 3321 3709 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m7682 3711 3710 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m7683 3708 3321 3711 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m7684 3709 3327 3708 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m7685 3712 3327 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m7686 3713 3708 3712 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m7687 1 3708 3707 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m7688 3714 3321 3713 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m7689 3715 3327 3714 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7690 0 3710 3715 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7691 3712 3321 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7692 0 3710 3712 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m7693 3716 3710 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m7694 3717 3321 3716 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m7695 3708 3710 3717 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7696 3717 3321 3708 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m7697 3718 3713 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7698 1 3327 3717 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7699 3713 3708 3719 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m7700 3720 3321 3713 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m7701 3721 3327 3720 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m7702 3710 3722 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m7703 3722 3723 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7704 3719 3710 3721 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m7705 1 3321 3719 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m7706 3719 3710 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m7707 1 3327 3719 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m7708 3718 3713 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m7709 0 3722 3710 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m7710 0 3723 3722 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7711 0 3397 3723 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m7712 3723 3411 852 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m7713 858 3387 3723 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.036e-11 ad=6.95e-12 ps=1.246e-05 pd=8.18e-06 
+ nrs=0.8 nrd=0.54 
m7714 3723 3409 842 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m7715 868 3393 3723 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m7716 3724 3725 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=5.99e-12 ad=1.348e-11 ps=9.58e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m7717 468 3726 3724 0 nenh l=1.1e-06 w=6.4e-06 
+ as=7.52e-12 ad=5.63e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.14 
m7718 3727 3728 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m7719 3726 3729 3727 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m7720 3730 3731 3726 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m7721 0 3732 3730 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m7722 3728 3732 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m7723 0 3734 3733 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m7724 3735 3729 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m7725 3736 3733 3735 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m7726 3737 3734 3736 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m7727 0 3731 3737 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m7728 3729 3731 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m7729 3738 3736 468 0 nenh l=1.1e-06 w=6.4e-06 
+ as=5.63e-12 ad=7.52e-12 ps=9.02e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m7730 0 3739 3738 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.99e-12 ps=1.275e-05 pd=9.58e-06 
+ nrs=0.29 nrd=0.13 
m7731 3740 3725 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m7732 468 3736 3740 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m7733 3741 3726 468 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m7734 1 3739 3741 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m7735 3742 3728 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m7736 3726 3731 3742 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m7737 3743 3729 3726 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m7738 1 3732 3743 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m7739 3728 3732 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7740 3744 3732 3745 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.57e-11 ps=1.429e-05 pd=2.04e-05 
+ nrs=0.11 nrd=0.12 
m7741 3746 3747 3744 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m7742 3745 3748 3746 0 nenh l=1.1e-06 w=1e-05 
+ as=1.354e-11 ad=8.5e-12 ps=1.759e-05 pd=1.17e-05 
+ nrs=0.14 nrd=0.08 
m7743 0 3748 3745 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m7744 3745 3747 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m7745 0 3747 3749 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m7746 3749 3748 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m7747 3750 3748 3749 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.354e-11 ps=1.17e-05 pd=1.759e-05 
+ nrs=0.08 nrd=0.14 
m7748 3751 3747 3750 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m7749 0 3752 3748 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m7750 3753 3748 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m7751 3731 3747 3753 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m7752 3754 3718 3731 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m7753 0 3752 3754 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m7754 3747 3718 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m7755 3749 3734 3751 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=1.416e-11 ps=2.04e-05 pd=1.429e-05 
+ nrs=0.12 nrd=0.11 
m7756 1 3734 3733 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m7757 3755 3729 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m7758 3736 3734 3755 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m7759 3756 3733 3736 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m7760 1 3731 3756 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m7761 3729 3731 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m7762 3744 3732 3757 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m7763 3758 3747 3744 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m7764 1 3748 3758 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m7765 3757 3748 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m7766 1 3747 3757 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m7767 3759 3747 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m7768 1 3748 3759 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m7769 3760 3748 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m7770 3751 3747 3760 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m7771 3759 3734 3751 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m7772 1 3752 3748 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=3.262e-11 ps=2.039e-05 pd=2.77e-05 
+ nrs=0.21 nrd=0.28 
m7773 3761 3748 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.23e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m7774 3731 3718 3761 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.067e-11 ad=7.27e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.1 
m7775 3762 3747 3731 1 penh l=1.1e-06 w=7.6e-06 
+ as=6.5e-12 ad=9.65e-12 ps=9.55e-06 pd=9.97e-06 
+ nrs=0.11 nrd=0.17 
m7776 1 3752 3762 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.16e-12 ps=1.359e-05 pd=9.05e-06 
+ nrs=0.31 nrd=0.12 
m7777 3747 3718 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.67e-11 ad=2.405e-11 ps=2.77e-05 pd=2.039e-05 
+ nrs=0.23 nrd=0.21 
m7778 1 3763 439 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m7779 3764 3725 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m7780 3763 3765 3764 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m7781 3766 3767 3763 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m7782 1 3739 3766 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m7783 3768 3769 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m7784 3767 3770 3768 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m7785 3771 3772 3767 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m7786 1 3773 3771 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m7787 3769 3773 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m7788 1 3775 3774 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m7789 3776 3772 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m7790 3765 3775 3776 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m7791 3777 3774 3765 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m7792 1 3770 3777 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m7793 3772 3770 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m7794 0 3763 439 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m7795 3778 3725 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=7.37e-12 ad=1.506e-11 ps=1.097e-05 pd=1.425e-05 
+ nrs=0.13 nrd=0.26 
m7796 3763 3767 3778 0 nenh l=1.1e-06 w=6.4e-06 
+ as=8.77e-12 ad=6.21e-12 ps=9.49e-06 pd=9.23e-06 
+ nrs=0.21 nrd=0.15 
m7797 3779 3765 3763 0 nenh l=1.1e-06 w=5.6e-06 
+ as=5.09e-12 ad=7.67e-12 ps=7.68e-06 pd=8.31e-06 
+ nrs=0.16 nrd=0.24 
m7798 0 3739 3779 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=6.17e-12 ps=1.275e-05 pd=9.32e-06 
+ nrs=0.29 nrd=0.13 
m7799 1 3781 3780 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=2.67e-11 ps=2.039e-05 pd=2.77e-05 
+ nrs=0.21 nrd=0.23 
m7800 3782 3783 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=9.84e-12 ad=1.959e-11 ps=1.17e-05 pd=1.661e-05 
+ nrs=0.13 nrd=0.25 
m7801 3770 3781 3782 1 penh l=1.1e-06 w=7.6e-06 
+ as=8.13e-12 ad=8.5e-12 ps=9.97e-06 pd=1.01e-05 
+ nrs=0.14 nrd=0.15 
m7802 3784 3780 3770 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.015e-11 ad=8.99e-12 ps=1.143e-05 pd=1.103e-05 
+ nrs=0.14 nrd=0.13 
m7803 1 3785 3784 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=1.063e-11 ps=1.661e-05 pd=1.197e-05 
+ nrs=0.25 nrd=0.14 
m7804 3783 3785 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.744e-11 ad=2.494e-11 ps=2.85e-05 pd=2.114e-05 
+ nrs=0.22 nrd=0.2 
m7805 3786 3773 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.55e-11 ad=2.672e-11 ps=1.478e-05 pd=2.265e-05 
+ nrs=0.11 nrd=0.19 
m7806 3732 3781 3786 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.151e-11 ad=1.498e-11 ps=1.394e-05 pd=1.428e-05 
+ nrs=0.09 nrd=0.11 
m7807 3786 3785 3732 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.705e-11 ad=1.309e-11 ps=1.625e-05 pd=1.586e-05 
+ nrs=0.1 nrd=0.08 
m7808 3787 3785 3786 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.498e-11 ps=1.33e-05 pd=1.428e-05 
+ nrs=0.07 nrd=0.11 
m7809 1 3781 3787 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m7810 3788 3781 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m7811 3789 3785 3788 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=9.86e-12 ps=1.428e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m7812 3734 3785 3789 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.309e-11 ad=1.705e-11 ps=1.586e-05 pd=1.625e-05 
+ nrs=0.08 nrd=0.1 
m7813 3789 3781 3734 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=1.151e-11 ps=1.428e-05 pd=1.394e-05 
+ nrs=0.11 nrd=0.09 
m7814 1 3775 3789 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.55e-11 ps=2.265e-05 pd=1.478e-05 
+ nrs=0.19 nrd=0.11 
m7815 3790 3769 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m7816 3767 3772 3790 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m7817 3791 3770 3767 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m7818 0 3773 3791 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m7819 3769 3773 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m7820 0 3775 3774 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m7821 3792 3772 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m7822 3765 3774 3792 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m7823 3793 3775 3765 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m7824 0 3770 3793 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m7825 3772 3770 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m7826 0 3781 3780 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m7827 3794 3783 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m7828 3770 3780 3794 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m7829 3795 3781 3770 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m7830 0 3785 3795 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m7831 3783 3785 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.468e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.47 nrd=0.35 
m7832 3732 3773 3796 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.175e-11 ad=1.755e-11 ps=1.429e-05 pd=1.841e-05 
+ nrs=0.09 nrd=0.13 
m7833 3797 3781 3732 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.013e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.1 
m7834 0 3785 3797 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=8.5e-12 ps=1.874e-05 pd=1.17e-05 
+ nrs=0.2 nrd=0.08 
m7835 3796 3785 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=2.299e-11 ps=1.841e-05 pd=2.174e-05 
+ nrs=0.13 nrd=0.17 
m7836 0 3781 3796 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=1.513e-11 ps=1.874e-05 pd=1.587e-05 
+ nrs=0.2 nrd=0.15 
m7837 3798 3781 0 0 nenh l=1.1e-06 w=1e-05 
+ as=1.513e-11 ad=1.982e-11 ps=1.587e-05 pd=1.874e-05 
+ nrs=0.15 nrd=0.2 
m7838 0 3785 3798 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.755e-11 ps=2.174e-05 pd=1.841e-05 
+ nrs=0.17 nrd=0.13 
m7839 3799 3785 0 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.982e-11 ps=1.17e-05 pd=1.874e-05 
+ nrs=0.08 nrd=0.2 
m7840 3734 3781 3799 0 nenh l=1.1e-06 w=1e-05 
+ as=1.013e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.1 nrd=0.08 
m7841 3798 3775 3734 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=1.175e-11 ps=1.841e-05 pd=1.429e-05 
+ nrs=0.13 nrd=0.09 
m7842 3800 3725 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.04e-12 ad=1.348e-11 ps=9.88e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m7843 410 3801 3800 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=5.33e-12 ps=8.5e-06 pd=8.72e-06 
+ nrs=0.19 nrd=0.15 
m7844 3802 3803 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m7845 3801 3804 3802 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m7846 3805 3806 3801 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m7847 0 3807 3805 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m7848 3803 3807 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m7849 0 3809 3808 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m7850 3810 3804 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m7851 3811 3808 3810 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m7852 3812 3809 3811 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m7853 0 3806 3812 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m7854 3804 3806 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m7855 3813 3811 410 0 nenh l=1.1e-06 w=6e-06 
+ as=5.29e-12 ad=6.86e-12 ps=8.61e-06 pd=8.5e-06 
+ nrs=0.15 nrd=0.19 
m7856 0 3739 3813 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=5.65e-12 ps=1.2e-05 pd=9.19e-06 
+ nrs=0.31 nrd=0.14 
m7857 3814 3725 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m7858 410 3811 3814 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m7859 3815 3801 410 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m7860 1 3739 3815 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m7861 3816 3803 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m7862 3801 3806 3816 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m7863 3817 3804 3801 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m7864 1 3807 3817 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m7865 3803 3807 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.308e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.42 nrd=0.4 
m7866 3773 3807 3818 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.57e-11 ps=1.429e-05 pd=2.04e-05 
+ nrs=0.11 nrd=0.12 
m7867 3819 3820 3773 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m7868 3818 3821 3819 0 nenh l=1.1e-06 w=1e-05 
+ as=1.354e-11 ad=8.5e-12 ps=1.759e-05 pd=1.17e-05 
+ nrs=0.14 nrd=0.08 
m7869 0 3821 3818 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m7870 3818 3820 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m7871 0 3820 3822 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m7872 3822 3821 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m7873 3823 3821 3822 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.354e-11 ps=1.17e-05 pd=1.759e-05 
+ nrs=0.08 nrd=0.14 
m7874 3775 3820 3823 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m7875 3822 3809 3775 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=1.416e-11 ps=2.04e-05 pd=1.429e-05 
+ nrs=0.12 nrd=0.11 
m7876 0 3361 3821 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.42e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.45 
m7877 3824 3821 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m7878 3806 3820 3824 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m7879 3825 3355 3806 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m7880 0 3361 3825 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m7881 3820 3355 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.372e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.44 nrd=0.35 
m7882 1 3809 3808 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m7883 3826 3804 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m7884 3811 3809 3826 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m7885 3827 3808 3811 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m7886 1 3806 3827 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m7887 3804 3806 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m7888 3773 3807 3828 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m7889 3829 3820 3773 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m7890 1 3821 3829 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m7891 3828 3821 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m7892 1 3820 3828 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m7893 3830 3820 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m7894 1 3821 3830 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m7895 3831 3821 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m7896 3775 3820 3831 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m7897 3830 3809 3775 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m7898 1 3361 3821 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=2.67e-11 ps=2.039e-05 pd=2.77e-05 
+ nrs=0.21 nrd=0.23 
m7899 3832 3821 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.45e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m7900 3806 3355 3832 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.033e-11 ad=7.53e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.11 
m7901 3833 3820 3806 1 penh l=1.1e-06 w=7.6e-06 
+ as=7.02e-12 ad=9.35e-12 ps=1.01e-05 pd=9.97e-06 
+ nrs=0.12 nrd=0.16 
m7902 1 3361 3833 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=8.12e-12 ps=1.661e-05 pd=1.17e-05 
+ nrs=0.25 nrd=0.1 
m7903 3820 3355 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.67e-11 ad=2.405e-11 ps=2.77e-05 pd=2.039e-05 
+ nrs=0.23 nrd=0.21 
m7904 1 3834 381 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m7905 3835 3725 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m7906 3834 3836 3835 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m7907 3837 3838 3834 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m7908 1 3739 3837 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m7909 3725 3739 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.484e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m7910 1 3739 3725 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.484e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m7911 3739 3839 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m7912 1 3839 3739 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m7913 3838 3836 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.596e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.51 nrd=0.4 
m7914 1 3370 3840 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m7915 3841 3842 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m7916 3836 3370 3841 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m7917 3843 3840 3836 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m7918 1 3373 3843 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m7919 3842 3373 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m7920 0 3834 381 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m7921 3844 3725 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=7.37e-12 ad=1.506e-11 ps=1.097e-05 pd=1.425e-05 
+ nrs=0.13 nrd=0.26 
m7922 3834 3838 3844 0 nenh l=1.1e-06 w=6.4e-06 
+ as=8.77e-12 ad=6.21e-12 ps=9.49e-06 pd=9.23e-06 
+ nrs=0.21 nrd=0.15 
m7923 3845 3836 3834 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=7.67e-12 ps=7.3e-06 pd=8.31e-06 
+ nrs=0.15 nrd=0.24 
m7924 0 3739 3845 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m7925 3725 3739 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.254e-11 ad=1.506e-11 ps=1.09e-05 pd=1.425e-05 
+ nrs=0.22 nrd=0.26 
m7926 0 3739 3725 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.506e-11 ad=1.254e-11 ps=1.425e-05 pd=1.09e-05 
+ nrs=0.26 nrd=0.22 
m7927 3739 3839 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m7928 0 3839 3739 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m7929 3838 3836 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m7930 3846 3370 3807 1 penh l=1.1e-06 w=1.44e-05 
+ as=1.224e-11 ad=4.04e-11 ps=1.61e-05 pd=3.49e-05 
+ nrs=0.06 nrd=0.19 
m7931 1 3373 3846 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.224e-11 ps=2.718e-05 pd=1.61e-05 
+ nrs=0.15 nrd=0.06 
m7932 3839 3847 1 1 penh l=1.1e-06 w=1.44e-05 
+ as=2.376e-11 ad=3.206e-11 ps=1.77e-05 pd=2.718e-05 
+ nrs=0.11 nrd=0.15 
m7933 1 3847 3839 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=2.376e-11 ps=2.718e-05 pd=1.77e-05 
+ nrs=0.15 nrd=0.11 
m7934 3847 2892 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.98e-11 ad=2.672e-11 ps=1.53e-05 pd=2.265e-05 
+ nrs=0.14 nrd=0.19 
m7935 3848 2987 3847 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.02e-11 ad=1.98e-11 ps=1.37e-05 pd=1.53e-05 
+ nrs=0.07 nrd=0.14 
m7936 1 2899 3848 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.02e-11 ps=2.265e-05 pd=1.37e-05 
+ nrs=0.19 nrd=0.07 
m7937 3809 3370 1 1 penh l=1.1e-06 w=1.28e-05 
+ as=1.264e-11 ad=2.85e-11 ps=1.53e-05 pd=2.416e-05 
+ nrs=0.08 nrd=0.17 
m7938 1 3373 3809 1 penh l=1.1e-06 w=1.28e-05 
+ as=2.85e-11 ad=1.264e-11 ps=2.416e-05 pd=1.53e-05 
+ nrs=0.17 nrd=0.08 
m7939 0 3370 3840 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.031e-11 ad=1.586e-11 ps=9.75e-06 pd=1.65e-05 
+ nrs=0.38 nrd=0.59 
m7940 3849 3842 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.32e-12 ad=1.348e-11 ps=9.63e-06 pd=1.275e-05 
+ nrs=0.14 nrd=0.29 
m7941 3836 3840 3849 0 nenh l=1.1e-06 w=5.2e-06 
+ as=8.58e-12 ad=4.84e-12 ps=8.5e-06 pd=7.37e-06 
+ nrs=0.32 nrd=0.18 
m7942 3850 3370 3836 0 nenh l=1.1e-06 w=5.2e-06 
+ as=4.56e-12 ad=8.58e-12 ps=7.37e-06 pd=8.5e-06 
+ nrs=0.17 nrd=0.32 
m7943 0 3373 3850 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.96e-12 ps=1.275e-05 pd=9.63e-06 
+ nrs=0.29 nrd=0.13 
m7944 3842 3373 0 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.031e-11 ps=1.65e-05 pd=9.75e-06 
+ nrs=0.59 nrd=0.38 
m7945 3807 3370 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=1.06e-11 ad=2.061e-11 ps=1.29e-05 pd=1.949e-05 
+ nrs=0.1 nrd=0.19 
m7946 0 3373 3807 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.061e-11 ad=1.06e-11 ps=1.949e-05 pd=1.29e-05 
+ nrs=0.19 nrd=0.1 
m7947 3839 3847 0 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.584e-11 ad=1.903e-11 ps=1.29e-05 pd=1.799e-05 
+ nrs=0.17 nrd=0.21 
m7948 0 3847 3839 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=1.584e-11 ps=1.799e-05 pd=1.29e-05 
+ nrs=0.21 nrd=0.17 
m7949 3851 2892 0 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.955e-11 ad=1.903e-11 ps=1.68e-05 pd=1.799e-05 
+ nrs=0.21 nrd=0.21 
m7950 3847 2987 3851 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.604e-11 ad=1.955e-11 ps=1.303e-05 pd=1.68e-05 
+ nrs=0.17 nrd=0.21 
m7951 3851 2899 3847 0 nenh l=1.1e-06 w=1e-05 
+ as=2.036e-11 ad=1.67e-11 ps=1.75e-05 pd=1.357e-05 
+ nrs=0.2 nrd=0.17 
m7952 3852 3370 3809 0 nenh l=1.1e-06 w=1.28e-05 
+ as=1.088e-11 ad=3.904e-11 ps=1.45e-05 pd=3.17e-05 
+ nrs=0.07 nrd=0.24 
m7953 0 3373 3852 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.088e-11 ps=2.399e-05 pd=1.45e-05 
+ nrs=0.15 nrd=0.07 
m7954 0 3853 3752 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=3.144e-11 ps=2.699e-05 pd=3.25e-05 
+ nrs=0.14 nrd=0.15 
m7955 3854 3855 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.083e-11 ad=3.013e-11 ps=2.27e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m7956 0 3338 3854 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.083e-11 ps=2.849e-05 pd=2.27e-05 
+ nrs=0.13 nrd=0.09 
m7957 3856 3855 0 0 nenh l=1.1e-06 w=1.68e-05 
+ as=1.454e-11 ad=3.33e-11 ps=1.992e-05 pd=3.149e-05 
+ nrs=0.05 nrd=0.12 
m7958 3853 3338 3856 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.246e-11 ps=1.795e-05 pd=1.708e-05 
+ nrs=0.07 nrd=0.06 
m7959 3854 3344 3853 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.919e-11 ad=1.383e-11 ps=2.091e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m7960 3857 3344 0 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.352e-11 ad=2.854e-11 ps=1.61e-05 pd=2.699e-05 
+ nrs=0.07 nrd=0.14 
m7961 3858 3853 3857 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.449e-11 ad=1.352e-11 ps=1.785e-05 pd=1.61e-05 
+ nrs=0.07 nrd=0.07 
m7962 3859 3338 3858 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.489e-11 ps=1.701e-05 pd=1.835e-05 
+ nrs=0.06 nrd=0.07 
m7963 3860 3344 3859 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m7964 0 3855 3860 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m7965 3857 3338 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.502e-11 ad=3.171e-11 ps=1.789e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m7966 0 3855 3857 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.202e-11 ps=2.399e-05 pd=1.431e-05 
+ nrs=0.15 nrd=0.07 
m7967 1 3853 3752 1 penh l=1.1e-06 w=1.8e-05 
+ as=4.008e-11 ad=3.314e-11 ps=3.398e-05 pd=3.89e-05 
+ nrs=0.12 nrd=0.1 
m7968 3781 3858 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m7969 3861 3855 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m7970 3862 3338 3861 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m7971 3853 3855 3862 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.615e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m7972 3862 3338 3853 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.499e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.06 
m7973 1 3344 3862 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m7974 1 3863 3785 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.484e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.47 
m7975 3864 3411 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m7976 3863 3393 3864 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.372e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.44 nrd=0.15 
m7977 1 3865 3855 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.226e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.32 
m7978 3858 3853 3866 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.447e-11 ad=1.386e-11 ps=1.722e-05 pd=1.719e-05 
+ nrs=0.1 nrd=0.1 
m7979 3867 3338 3858 1 penh l=1.1e-06 w=1.88e-05 
+ as=1.621e-11 ad=2.267e-11 ps=2.153e-05 pd=2.698e-05 
+ nrs=0.05 nrd=0.06 
m7980 3868 3344 3867 1 penh l=1.1e-06 w=2.12e-05 
+ as=1.814e-11 ad=1.827e-11 ps=2.344e-05 pd=2.427e-05 
+ nrs=0.04 nrd=0.04 
m7981 3866 3855 3868 1 penh l=1.1e-06 w=2.24e-05 
+ as=2.588e-11 ad=1.916e-11 ps=3.21e-05 pd=2.476e-05 
+ nrs=0.05 nrd=0.04 
m7982 1 3338 3866 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.664e-11 ps=2.718e-05 pd=2.063e-05 
+ nrs=0.15 nrd=0.08 
m7983 3866 3855 1 1 penh l=1.1e-06 w=1.52e-05 
+ as=1.756e-11 ad=3.384e-11 ps=2.178e-05 pd=2.869e-05 
+ nrs=0.08 nrd=0.15 
m7984 1 3344 3866 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.386e-11 ps=2.265e-05 pd=1.719e-05 
+ nrs=0.19 nrd=0.1 
m7985 3781 3858 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.04e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.08 nrd=0.12 
m7986 3865 3869 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.298e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.48 nrd=0.43 
m7987 0 3863 3785 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m7988 3863 3411 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=5.55e-12 ps=6.1e-06 pd=5.25e-06 
+ nrs=0.59 nrd=0.71 
m7989 0 3393 3863 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=4.62e-12 ps=5.25e-06 pd=6.1e-06 
+ nrs=0.71 nrd=0.59 
m7990 0 3865 3855 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.52e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.37 
m7991 0 3869 3865 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m7992 0 3397 3869 0 nenh l=1.1e-06 w=3.2e-06 
+ as=6.34e-12 ad=6.09e-12 ps=6e-06 pd=7.29e-06 
+ nrs=0.62 nrd=0.6 
m7993 3869 3411 1 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.098e-11 ps=8.2e-06 pd=1.406e-05 
+ nrs=0.53 nrd=0.85 
m7994 0 3387 3869 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.86e-12 ps=6.75e-06 pd=8.2e-06 
+ nrs=0.55 nrd=0.53 
m7995 3869 3409 858 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.036e-11 ps=8.2e-06 pd=1.246e-05 
+ nrs=0.53 nrd=0.8 
m7996 852 3393 3869 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.86e-12 ps=1.202e-05 pd=8.2e-06 
+ nrs=0.77 nrd=0.53 
m7997 0 3871 3870 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.427e-11 ad=2.196e-11 ps=1.35e-05 pd=2.05e-05 
+ nrs=0.28 nrd=0.42 
m7998 3871 3872 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m7999 0 3874 3873 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.22e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.76 
m8000 3874 3875 0 0 nenh l=1.1e-06 w=4e-06 
+ as=1.22e-11 ad=7.93e-12 ps=1.41e-05 pd=7.5e-06 
+ nrs=0.76 nrd=0.5 
m8001 1 3871 3870 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m8002 3871 3872 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8003 3876 3877 0 0 nenh l=1.1e-06 w=4e-06 
+ as=6.6e-12 ad=7.93e-12 ps=7.3e-06 pd=7.5e-06 
+ nrs=0.41 nrd=0.5 
m8004 0 3877 3876 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=6.6e-12 ps=7.5e-06 pd=7.3e-06 
+ nrs=0.5 nrd=0.41 
m8005 3878 3879 3877 0 nenh l=1.1e-06 w=8.8e-06 
+ as=7.66e-12 ad=1.964e-11 ps=1.122e-05 pd=2.37e-05 
+ nrs=0.1 nrd=0.25 
m8006 3880 3881 3878 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.4e-12 ps=1.25e-05 pd=1.378e-05 
+ nrs=0.08 nrd=0.08 
m8007 0 3401 3880 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m8008 3882 3879 0 0 nenh l=1.1e-06 w=8.8e-06 
+ as=9.24e-12 ad=1.744e-11 ps=1.13e-05 pd=1.65e-05 
+ nrs=0.12 nrd=0.23 
m8009 0 3883 3882 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.744e-11 ad=9.24e-12 ps=1.65e-05 pd=1.13e-05 
+ nrs=0.23 nrd=0.12 
m8010 3884 3885 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=1.665e-11 ps=1.01e-05 pd=1.575e-05 
+ nrs=0.1 nrd=0.24 
m8011 3886 3887 3884 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.89e-11 ad=7.14e-12 ps=2.29e-05 pd=1.01e-05 
+ nrs=0.27 nrd=0.1 
m8012 1 3874 3873 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=2.358e-11 ps=1.737e-05 pd=2.29e-05 
+ nrs=0.24 nrd=0.28 
m8013 3874 3875 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.358e-11 ad=2.048e-11 ps=2.29e-05 pd=1.737e-05 
+ nrs=0.28 nrd=0.24 
m8014 3876 3877 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.128e-11 ad=2.494e-11 ps=1.37e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8015 1 3877 3876 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.128e-11 ps=2.114e-05 pd=1.37e-05 
+ nrs=0.2 nrd=0.09 
m8016 3888 3881 3887 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.27e-12 ad=2.16e-11 ps=1.176e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.23 
m8017 3889 3401 3888 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.31e-12 ps=1.25e-05 pd=1.324e-05 
+ nrs=0.08 nrd=0.08 
m8018 0 3890 3889 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m8019 3891 3879 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m8020 3892 3893 3891 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.31e-12 ad=9.18e-12 ps=1.324e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m8021 3885 3390 3892 0 nenh l=1.1e-06 w=9.6e-06 
+ as=2.16e-11 ad=8.27e-12 ps=2.53e-05 pd=1.176e-05 
+ nrs=0.23 nrd=0.09 
m8022 1 3879 3877 1 penh l=1.1e-06 w=9.6e-06 
+ as=2.137e-11 ad=1.315e-11 ps=1.812e-05 pd=1.587e-05 
+ nrs=0.23 nrd=0.14 
m8023 3877 3881 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.26e-11 ad=2.048e-11 ps=1.521e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m8024 1 3401 3877 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.26e-11 ps=1.737e-05 pd=1.521e-05 
+ nrs=0.24 nrd=0.15 
m8025 3894 3879 1 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.194e-11 ad=2.939e-11 ps=1.49e-05 pd=2.492e-05 
+ nrs=0.07 nrd=0.17 
m8026 3882 3883 3894 1 penh l=1.1e-06 w=1.32e-05 
+ as=2.586e-11 ad=1.194e-11 ps=3.01e-05 pd=1.49e-05 
+ nrs=0.15 nrd=0.07 
m8027 3886 3885 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.466e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.07 nrd=0.15 
m8028 1 3887 3886 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.466e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.07 
m8029 1 3881 3887 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m8030 3887 3401 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m8031 1 3890 3887 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m8032 3885 3879 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m8033 1 3893 3885 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m8034 3885 3390 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m8035 3875 3895 1 1 penh l=1.1e-06 w=1e-05 
+ as=2.346e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.23 nrd=0.22 
m8036 3895 3896 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8037 3872 3886 1 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=8.54e-12 ps=7.22e-06 pd=1.094e-05 
+ nrs=0.69 nrd=1.09 
m8038 910 3876 3872 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m8039 3897 3883 3898 1 penh l=1.1e-06 w=1.04e-05 
+ as=8.84e-12 ad=2.596e-11 ps=1.21e-05 pd=2.69e-05 
+ nrs=0.08 nrd=0.24 
m8040 1 3890 3897 1 penh l=1.1e-06 w=1.04e-05 
+ as=2.316e-11 ad=8.84e-12 ps=1.963e-05 pd=1.21e-05 
+ nrs=0.21 nrd=0.08 
m8041 3899 3390 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m8042 1 3893 3899 1 penh l=1.1e-06 w=8e-06 
+ as=1.781e-11 ad=1.075e-11 ps=1.51e-05 pd=1.383e-05 
+ nrs=0.28 nrd=0.17 
m8043 3899 3890 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m8044 3900 3899 1 1 penh l=1.1e-06 w=1e-05 
+ as=1.058e-11 ad=2.227e-11 ps=1.25e-05 pd=1.888e-05 
+ nrs=0.11 nrd=0.22 
m8045 1 3899 3900 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=1.058e-11 ps=1.888e-05 pd=1.25e-05 
+ nrs=0.22 nrd=0.11 
m8046 3896 3900 595 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.74e-12 ps=7.22e-06 pd=9.64e-06 
+ nrs=0.69 nrd=0.99 
m8047 602 3876 3896 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=5.4e-12 ps=9.87e-06 pd=7.22e-06 
+ nrs=1.04 nrd=0.69 
m8048 3896 3882 910 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.88e-12 ps=7.22e-06 pd=1.048e-05 
+ nrs=0.69 nrd=1 
m8049 911 3898 3896 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m8050 0 3886 3896 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.4e-12 ps=5.25e-06 pd=7.22e-06 
+ nrs=0.71 nrd=0.69 
m8051 3901 3893 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=2.405e-11 ps=1.41e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m8052 3883 3390 3901 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.046e-11 ad=1.014e-11 ps=1.25e-05 pd=1.41e-05 
+ nrs=0.09 nrd=0.09 
m8053 3902 3401 3883 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=1.046e-11 ps=1.41e-05 pd=1.25e-05 
+ nrs=0.09 nrd=0.09 
m8054 1 3881 3902 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.014e-11 ps=2.039e-05 pd=1.41e-05 
+ nrs=0.21 nrd=0.09 
m8055 911 3900 3872 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m8056 3872 3882 911 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.91e-12 ps=7.22e-06 pd=1.05e-05 
+ nrs=0.69 nrd=1.01 
m8057 910 3898 3872 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m8058 0 3895 3875 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m8059 0 3896 3895 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m8060 3898 3883 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m8061 0 3890 3898 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m8062 3903 3390 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m8063 3904 3893 3903 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.4e-12 ad=9.18e-12 ps=1.378e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m8064 3899 3890 3904 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.964e-11 ad=7.66e-12 ps=2.37e-05 pd=1.122e-05 
+ nrs=0.25 nrd=0.1 
m8065 3900 3899 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m8066 0 3899 3900 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m8067 3905 3893 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=9.84e-12 ad=2.061e-11 ps=1.319e-05 pd=1.949e-05 
+ nrs=0.09 nrd=0.19 
m8068 3883 3401 3905 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.06e-11 ps=1.29e-05 pd=1.421e-05 
+ nrs=0.09 nrd=0.08 
m8069 3906 3390 3883 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.062e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.08 nrd=0.09 
m8070 0 3881 3906 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.024e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m8071 898 886 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8072 0 886 898 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8073 886 3907 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8074 0 3907 886 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8075 0 3908 3907 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8076 3909 3907 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8077 3910 19 3908 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8078 0 3911 3910 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8079 3911 37 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=5.55e-12 ps=6.74e-06 pd=5.25e-06 
+ nrs=0.78 nrd=0.71 
m8080 3912 3910 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8081 3911 19 3912 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8082 898 886 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8083 1 886 898 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8084 886 3907 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8085 1 3907 886 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8086 1 3908 3907 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8087 3913 3914 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8088 3915 3909 3913 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8089 3916 3917 3915 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8090 0 3918 3916 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8091 3914 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8092 3911 25 3919 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8093 3915 26 3911 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8094 3908 19 3909 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.31e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8095 0 3920 3917 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8096 3909 3907 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.227e-11 ad=2.761e-11 ps=2.43e-05 pd=2.341e-05 
+ nrs=0.14 nrd=0.18 
m8097 1 3911 3910 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.114e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.3 
m8098 3921 3910 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8099 3922 25 3921 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8100 3911 26 3922 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8101 3923 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8102 3915 3909 3923 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8103 3924 3917 3915 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8104 1 3914 3924 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8105 3914 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8106 1 3920 3917 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8107 888 901 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8108 1 901 888 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8109 901 3919 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8110 1 3919 901 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8111 1 3925 3919 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8112 3926 3919 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.227e-11 ad=2.761e-11 ps=2.43e-05 pd=2.341e-05 
+ nrs=0.14 nrd=0.18 
m8113 1 3928 3927 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.114e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.3 
m8114 3925 19 3926 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.31e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8115 888 901 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8116 0 901 888 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8117 901 3919 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8118 0 3919 901 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8119 3929 3927 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8120 3930 25 3929 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8121 3928 26 3930 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8122 0 3925 3919 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8123 3931 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8124 3932 3926 3931 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8125 3933 3934 3932 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8126 1 3935 3933 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8127 3935 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8128 3927 19 3925 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8129 3926 3919 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8130 0 3928 3927 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8131 3936 3927 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8132 3928 19 3936 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8133 3928 25 3937 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8134 3932 26 3928 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8135 1 3938 3934 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8136 0 37 3928 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m8137 3939 3935 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8138 3932 3926 3939 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8139 3940 3934 3932 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8140 0 3918 3940 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8141 3935 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8142 0 3938 3934 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8143 889 902 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8144 0 902 889 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8145 902 3937 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8146 0 3937 902 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8147 0 3941 3937 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8148 3942 3937 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8149 3943 19 3941 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8150 0 3944 3943 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8151 3944 37 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=5.55e-12 ps=6.74e-06 pd=5.25e-06 
+ nrs=0.78 nrd=0.71 
m8152 3945 3943 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8153 3944 19 3945 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8154 889 902 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8155 1 902 889 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8156 902 3937 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8157 1 3937 902 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8158 1 3941 3937 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8159 3946 3947 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8160 3948 3942 3946 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8161 3949 3950 3948 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8162 0 3918 3949 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8163 3947 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8164 3944 25 3951 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8165 3948 26 3944 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8166 3941 19 3942 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.31e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8167 0 3952 3950 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8168 3942 3937 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.227e-11 ad=2.761e-11 ps=2.43e-05 pd=2.341e-05 
+ nrs=0.14 nrd=0.18 
m8169 1 3944 3943 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=1.89e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.27 
m8170 3953 3943 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8171 3954 25 3953 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8172 3944 26 3954 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8173 3955 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8174 3948 3942 3955 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8175 3956 3950 3948 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8176 1 3947 3956 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8177 3947 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8178 1 3952 3950 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8179 929 943 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8180 1 943 929 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8181 943 3951 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8182 1 3951 943 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8183 1 3957 3951 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8184 3958 3951 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.227e-11 ad=2.761e-11 ps=2.43e-05 pd=2.341e-05 
+ nrs=0.14 nrd=0.18 
m8185 1 3960 3959 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=1.89e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.27 
m8186 3957 19 3958 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.31e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8187 929 943 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8188 0 943 929 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8189 943 3951 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8190 0 3951 943 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8191 3961 3959 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8192 3962 25 3961 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8193 3960 26 3962 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8194 0 3957 3951 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8195 3963 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8196 3964 3958 3963 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8197 3965 3966 3964 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8198 1 3967 3965 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8199 3967 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8200 3959 19 3957 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8201 3958 3951 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8202 0 3960 3959 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8203 3968 3959 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8204 3960 19 3968 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8205 3960 25 36 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=1.098e-11 ps=8.66e-06 pd=1.33e-05 
+ nrs=0.6 nrd=0.85 
m8206 3964 26 3960 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8207 1 3969 3966 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8208 0 37 3960 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m8209 3970 3967 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8210 3964 3958 3970 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8211 3971 3966 3964 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8212 0 3918 3971 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8213 3967 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8214 0 3969 3966 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8215 1335 1324 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8216 0 1324 1335 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8217 1324 3972 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8218 0 3972 1324 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8219 0 3973 3972 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8220 3974 3972 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8221 3975 19 3973 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8222 0 3976 3975 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8223 3976 37 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=5.55e-12 ps=6.74e-06 pd=5.25e-06 
+ nrs=0.78 nrd=0.71 
m8224 3977 3975 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8225 3976 19 3977 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8226 1335 1324 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8227 1 1324 1335 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8228 1324 3972 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8229 1 3972 1324 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8230 1 3973 3972 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8231 3978 3979 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8232 3980 3974 3978 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8233 3981 3982 3980 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8234 0 3918 3981 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8235 3979 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8236 3976 25 3983 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8237 3980 26 3976 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8238 3973 19 3974 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8239 0 3984 3982 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8240 3974 3972 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8241 1 3976 3975 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.562e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m8242 3985 3975 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8243 3986 25 3985 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8244 3976 26 3986 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8245 3987 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8246 3980 3974 3987 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8247 3988 3982 3980 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8248 1 3979 3988 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8249 3979 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8250 1 3984 3982 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8251 1326 1338 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8252 1 1338 1326 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8253 1338 3983 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8254 1 3983 1338 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8255 1 3989 3983 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8256 3990 3983 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8257 1 3992 3991 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.114e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.3 
m8258 3989 19 3990 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8259 1326 1338 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8260 0 1338 1326 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8261 1338 3983 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8262 0 3983 1338 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8263 3993 3991 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8264 3994 25 3993 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8265 3992 26 3994 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8266 0 3989 3983 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8267 3995 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8268 3996 3990 3995 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8269 3997 3998 3996 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8270 1 3999 3997 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8271 3999 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8272 3991 19 3989 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8273 3990 3983 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8274 0 3992 3991 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8275 4000 3991 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8276 3992 19 4000 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8277 3992 25 3907 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8278 3996 26 3992 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8279 1 4001 3998 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8280 0 37 3992 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m8281 4002 3999 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8282 3996 3990 4002 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8283 4003 3998 3996 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8284 0 3918 4003 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8285 3999 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8286 0 4001 3998 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8287 1698 1687 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8288 0 1687 1698 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8289 1687 4004 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8290 0 4004 1687 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8291 0 4005 4004 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8292 4006 4004 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8293 4007 19 4005 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8294 0 4008 4007 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8295 4008 37 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=5.55e-12 ps=6.74e-06 pd=5.25e-06 
+ nrs=0.78 nrd=0.71 
m8296 4009 4007 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8297 4008 19 4009 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8298 1698 1687 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8299 1 1687 1698 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8300 1687 4004 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8301 1 4004 1687 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8302 1 4005 4004 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8303 4010 4011 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8304 4012 4006 4010 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8305 4013 4014 4012 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8306 0 3918 4013 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8307 4011 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8308 4008 25 4015 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8309 4012 26 4008 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8310 4005 19 4006 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8311 0 4016 4014 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8312 4006 4004 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8313 1 4008 4007 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.562e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m8314 4017 4007 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8315 4018 25 4017 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8316 4008 26 4018 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8317 4019 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8318 4012 4006 4019 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8319 4020 4014 4012 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8320 1 4011 4020 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8321 4011 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8322 1 4016 4014 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8323 1689 1701 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8324 1 1701 1689 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8325 1701 4015 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8326 1 4015 1701 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8327 1 4021 4015 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8328 4022 4015 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8329 1 4024 4023 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.114e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.3 
m8330 4021 19 4022 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8331 1689 1701 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8332 0 1701 1689 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8333 1701 4015 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8334 0 4015 1701 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8335 4025 4023 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8336 4026 25 4025 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8337 4024 26 4026 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8338 0 4021 4015 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8339 4027 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8340 4028 4022 4027 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8341 4029 4030 4028 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8342 1 4031 4029 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8343 4031 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8344 4023 19 4021 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8345 4022 4015 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8346 0 4024 4023 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8347 4032 4023 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8348 4024 19 4032 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8349 4024 25 3972 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8350 4028 26 4024 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8351 1 4033 4030 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8352 0 37 4024 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m8353 4034 4031 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8354 4028 4022 4034 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8355 4035 4030 4028 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8356 0 3918 4035 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8357 4031 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8358 0 4033 4030 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8359 2186 2175 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8360 0 2175 2186 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8361 2175 4036 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8362 0 4036 2175 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8363 0 4037 4036 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8364 4038 4036 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8365 4039 19 4037 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8366 0 4040 4039 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8367 4040 37 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=5.55e-12 ps=6.74e-06 pd=5.25e-06 
+ nrs=0.78 nrd=0.71 
m8368 4041 4039 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8369 4040 19 4041 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8370 2186 2175 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8371 1 2175 2186 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8372 2175 4036 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8373 1 4036 2175 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8374 1 4037 4036 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8375 4042 4043 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8376 4044 4038 4042 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8377 4045 4046 4044 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8378 0 3918 4045 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8379 4043 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8380 4040 25 4047 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8381 4044 26 4040 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8382 4037 19 4038 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8383 0 4048 4046 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8384 4038 4036 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8385 1 4040 4039 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.562e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m8386 4049 4039 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8387 4050 25 4049 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8388 4040 26 4050 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8389 4051 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8390 4044 4038 4051 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8391 4052 4046 4044 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8392 1 4043 4052 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8393 4043 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8394 1 4048 4046 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8395 2177 2189 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8396 1 2189 2177 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8397 2189 4047 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8398 1 4047 2189 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8399 1 4053 4047 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8400 4054 4047 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8401 1 4056 4055 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.114e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.3 
m8402 4053 19 4054 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8403 2177 2189 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8404 0 2189 2177 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8405 2189 4047 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8406 0 4047 2189 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8407 4057 4055 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8408 4058 25 4057 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8409 4056 26 4058 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8410 0 4053 4047 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8411 4059 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8412 4060 4054 4059 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8413 4061 4062 4060 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8414 1 4063 4061 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8415 4063 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8416 4055 19 4053 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8417 4054 4047 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8418 0 4056 4055 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8419 4064 4055 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8420 4056 19 4064 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8421 4056 25 4004 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8422 4060 26 4056 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8423 1 4065 4062 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8424 0 37 4056 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m8425 4066 4063 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8426 4060 4054 4066 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8427 4067 4062 4060 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8428 0 3918 4067 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8429 4063 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8430 0 4065 4062 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8431 2549 2538 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8432 0 2538 2549 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8433 2538 4068 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8434 0 4068 2538 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8435 0 4069 4068 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8436 4070 4068 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8437 4071 19 4069 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8438 0 4072 4071 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8439 4072 37 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=5.55e-12 ps=6.74e-06 pd=5.25e-06 
+ nrs=0.78 nrd=0.71 
m8440 4073 4071 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8441 4072 19 4073 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8442 2549 2538 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8443 1 2538 2549 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8444 2538 4068 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8445 1 4068 2538 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8446 1 4069 4068 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8447 4074 4075 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8448 4076 4070 4074 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8449 4077 4078 4076 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8450 0 3918 4077 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8451 4075 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8452 4072 25 4079 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8453 4076 26 4072 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8454 4069 19 4070 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8455 0 4080 4078 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8456 4070 4068 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8457 1 4072 4071 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.562e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m8458 4081 4071 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8459 4082 25 4081 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8460 4072 26 4082 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8461 4083 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8462 4076 4070 4083 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8463 4084 4078 4076 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8464 1 4075 4084 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8465 4075 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8466 1 4080 4078 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8467 2540 2552 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8468 1 2552 2540 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8469 2552 4079 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8470 1 4079 2552 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8471 1 4085 4079 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8472 4086 4079 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8473 1 4088 4087 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.114e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.3 
m8474 4085 19 4086 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8475 2540 2552 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8476 0 2552 2540 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8477 2552 4079 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8478 0 4079 2552 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8479 4089 4087 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8480 4090 25 4089 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8481 4088 26 4090 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8482 0 4085 4079 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8483 4091 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8484 4092 4086 4091 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8485 4093 4094 4092 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8486 1 4095 4093 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8487 4095 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8488 4087 19 4085 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8489 4086 4079 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8490 0 4088 4087 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8491 4096 4087 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8492 4088 19 4096 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8493 4088 25 4036 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8494 4092 26 4088 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8495 1 4097 4094 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8496 0 37 4088 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m8497 4098 4095 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8498 4092 4086 4098 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8499 4099 4094 4092 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8500 0 3918 4099 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8501 4095 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8502 0 4097 4094 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8503 3038 3027 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8504 0 3027 3038 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8505 3027 4100 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8506 0 4100 3027 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8507 0 4101 4100 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8508 4102 4100 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8509 4103 19 4101 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8510 0 4104 4103 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8511 4104 37 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=5.55e-12 ps=6.74e-06 pd=5.25e-06 
+ nrs=0.78 nrd=0.71 
m8512 4105 4103 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8513 4104 19 4105 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8514 3038 3027 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8515 1 3027 3038 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8516 3027 4100 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8517 1 4100 3027 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8518 1 4101 4100 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8519 4106 4107 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8520 4108 4102 4106 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8521 4109 4110 4108 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8522 0 3918 4109 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8523 4107 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8524 4104 25 4111 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8525 4108 26 4104 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8526 4101 19 4102 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8527 0 4112 4110 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8528 4102 4100 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8529 1 4104 4103 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.562e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m8530 4113 4103 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8531 4114 25 4113 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8532 4104 26 4114 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8533 4115 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8534 4108 4102 4115 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8535 4116 4110 4108 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8536 1 4107 4116 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8537 4107 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8538 1 4112 4110 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8539 3029 3041 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8540 1 3041 3029 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8541 3041 4111 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8542 1 4111 3041 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8543 1 4117 4111 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8544 4118 4111 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8545 1 4120 4119 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.114e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.3 
m8546 4117 19 4118 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8547 3029 3041 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8548 0 3041 3029 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8549 3041 4111 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8550 0 4111 3041 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8551 4121 4119 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8552 4122 25 4121 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8553 4120 26 4122 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8554 0 4117 4111 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8555 4123 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8556 4124 4118 4123 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8557 4125 4126 4124 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8558 1 4127 4125 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8559 4127 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8560 4119 19 4117 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8561 4118 4111 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8562 0 4120 4119 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8563 4128 4119 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8564 4120 19 4128 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8565 4120 25 4068 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8566 4124 26 4120 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8567 1 4129 4126 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8568 0 37 4120 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m8569 4130 4127 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8570 4124 4118 4130 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8571 4131 4126 4124 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8572 0 3918 4131 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8573 4127 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8574 0 4129 4126 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8575 3401 3390 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8576 0 3390 3401 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8577 3390 4132 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8578 0 4132 3390 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8579 0 4133 4132 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8580 4134 4132 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8581 4135 19 4133 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8582 0 4136 4135 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8583 4136 37 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=5.55e-12 ps=6.74e-06 pd=5.25e-06 
+ nrs=0.78 nrd=0.71 
m8584 4137 4135 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8585 4136 19 4137 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8586 3401 3390 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8587 1 3390 3401 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8588 3390 4132 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8589 1 4132 3390 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8590 1 4133 4132 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8591 4138 4139 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8592 4140 4134 4138 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8593 4141 4142 4140 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8594 0 3918 4141 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8595 4139 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8596 4136 25 4143 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8597 4140 26 4136 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8598 4133 19 4134 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8599 0 4144 4142 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8600 4134 4132 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8601 1 4136 4135 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.562e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m8602 4145 4135 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8603 4146 25 4145 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8604 4136 26 4146 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8605 4147 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8606 4140 4134 4147 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8607 4148 4142 4140 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8608 1 4139 4148 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8609 4139 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8610 1 4144 4142 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8611 3392 3404 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8612 1 3404 3392 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8613 3404 4143 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8614 1 4143 3404 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8615 1 4149 4143 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8616 4150 4143 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8617 1 4152 4151 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.114e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.3 
m8618 4149 19 4150 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8619 3392 3404 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8620 0 3404 3392 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8621 3404 4143 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8622 0 4143 3404 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8623 4153 4151 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8624 4154 25 4153 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8625 4152 26 4154 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8626 0 4149 4143 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8627 4155 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8628 4156 4150 4155 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8629 4157 4158 4156 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8630 1 4159 4157 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8631 4159 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8632 4151 19 4149 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8633 4150 4143 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8634 0 4152 4151 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8635 4160 4151 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8636 4152 19 4160 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8637 4152 25 4100 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8638 4156 26 4152 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8639 1 4161 4158 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8640 0 37 4152 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m8641 4162 4159 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8642 4156 4150 4162 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8643 4163 4158 4156 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8644 0 3918 4163 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8645 4159 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8646 0 4161 4158 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8647 3890 3879 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8648 0 3879 3890 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8649 3879 4164 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8650 0 4164 3879 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8651 0 4165 4164 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8652 4166 4164 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8653 4167 19 4165 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8654 0 4168 4167 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8655 4168 37 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=5.55e-12 ps=6.74e-06 pd=5.25e-06 
+ nrs=0.78 nrd=0.71 
m8656 4169 4167 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8657 4168 19 4169 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8658 3890 3879 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8659 1 3879 3890 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8660 3879 4164 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8661 1 4164 3879 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8662 1 4165 4164 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8663 4170 4171 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8664 4172 4166 4170 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8665 4173 4174 4172 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8666 0 3918 4173 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8667 4171 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8668 4168 25 4175 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8669 4172 26 4168 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8670 4165 19 4166 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8671 0 4176 4174 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8672 4166 4164 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8673 1 4168 4167 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.562e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m8674 4177 4167 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8675 4178 25 4177 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8676 4168 26 4178 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8677 4179 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8678 4172 4166 4179 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8679 4180 4174 4172 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8680 1 4171 4180 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8681 4171 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8682 1 4176 4174 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8683 3881 3893 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8684 1 3893 3881 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8685 3893 4175 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8686 1 4175 3893 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8687 1 4181 4175 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8688 4182 4175 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8689 1 4184 4183 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.114e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.3 
m8690 4181 19 4182 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8691 3881 3893 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8692 0 3893 3881 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8693 3893 4175 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8694 0 4175 3893 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8695 4185 4183 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8696 4186 25 4185 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8697 4184 26 4186 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8698 0 4181 4175 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8699 4187 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8700 4188 4182 4187 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8701 4189 4190 4188 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8702 1 4191 4189 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8703 4191 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8704 4183 19 4181 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8705 4182 4175 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8706 0 4184 4183 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8707 4192 4183 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8708 4184 19 4192 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8709 4184 25 4132 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8710 4188 26 4184 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8711 1 4193 4190 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8712 0 37 4184 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m8713 4194 4191 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8714 4188 4182 4194 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8715 4195 4190 4188 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8716 0 3918 4195 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8717 4191 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8718 0 4193 4190 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8719 4196 4197 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8720 0 4197 4196 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8721 4197 857 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8722 0 857 4197 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8723 0 4198 857 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.893e-11 ps=2.099e-05 pd=3.189e-05 
+ nrs=0.18 nrd=0.23 
m8724 4199 857 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8725 4200 19 4198 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8726 0 4201 4200 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8727 4201 37 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=5.55e-12 ps=6.74e-06 pd=5.25e-06 
+ nrs=0.78 nrd=0.71 
m8728 4202 4200 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8729 4201 19 4202 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8730 4196 4197 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8731 1 4197 4196 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8732 4197 857 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8733 1 857 4197 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8734 1 4198 857 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8735 4203 4204 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8736 4205 4199 4203 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8737 4206 4207 4205 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8738 0 3918 4206 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8739 4204 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8740 4201 25 4208 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8741 4205 26 4201 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8742 4198 19 4199 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8743 0 4209 4207 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8744 4199 857 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8745 1 4201 4200 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.562e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.36 
m8746 4210 4200 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8747 4211 25 4210 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8748 4201 26 4211 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8749 4212 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8750 4205 4199 4212 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8751 4213 4207 4205 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8752 1 4204 4213 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8753 4204 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8754 1 4209 4207 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8755 4214 4215 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8756 1 4215 4214 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8757 4215 4208 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.658e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.08 nrd=0.15 
m8758 1 4208 4215 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.658e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.08 
m8759 1 4216 4208 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=2.978e-11 ps=2.794e-05 pd=3.25e-05 
+ nrs=0.15 nrd=0.14 
m8760 4217 4208 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.167e-11 ad=2.672e-11 ps=2.35e-05 pd=2.265e-05 
+ nrs=0.15 nrd=0.19 
m8761 1 4219 4218 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.114e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.3 
m8762 4216 19 4217 1 penh l=1.1e-06 w=2.4e-06 
+ as=9.4e-12 ad=4.33e-12 ps=1.25e-05 pd=4.7e-06 
+ nrs=1.63 nrd=0.75 
m8763 4214 4215 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8764 0 4215 4214 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8765 4215 4208 0 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.182e-11 ad=1.823e-11 ps=1.17e-05 pd=1.724e-05 
+ nrs=0.14 nrd=0.22 
m8766 0 4208 4215 0 nenh l=1.1e-06 w=9.2e-06 
+ as=1.823e-11 ad=1.182e-11 ps=1.724e-05 pd=1.17e-05 
+ nrs=0.22 nrd=0.14 
m8767 4220 4218 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m8768 4221 25 4220 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=4.76e-12 ps=7.3e-06 pd=7.3e-06 
+ nrs=0.15 nrd=0.15 
m8769 4219 26 4221 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.54 nrd=0.15 
m8770 0 4216 4208 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=2.907e-11 ps=2.099e-05 pd=3.163e-05 
+ nrs=0.18 nrd=0.23 
m8771 4222 3918 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.083e-11 ad=2.494e-11 ps=1.323e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m8772 4223 4217 4222 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=1.161e-11 ps=1.45e-05 pd=1.417e-05 
+ nrs=0.1 nrd=0.08 
m8773 4224 4225 4223 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.161e-11 ad=1.42e-11 ps=1.417e-05 pd=1.45e-05 
+ nrs=0.08 nrd=0.1 
m8774 1 4226 4224 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.083e-11 ps=2.114e-05 pd=1.323e-05 
+ nrs=0.2 nrd=0.09 
m8775 4226 3918 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8776 4218 19 4216 0 nenh l=1.1e-06 w=3.6e-06 
+ as=8.39e-12 ad=1.098e-11 ps=7.26e-06 pd=1.33e-05 
+ nrs=0.65 nrd=0.85 
m8777 4217 4208 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.276e-11 ad=2.061e-11 ps=2.37e-05 pd=1.949e-05 
+ nrs=0.21 nrd=0.19 
m8778 0 4219 4218 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.957e-11 ps=1.575e-05 pd=1.694e-05 
+ nrs=0.24 nrd=0.28 
m8779 4227 4218 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m8780 4219 19 4227 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.09e-12 ad=2.38e-12 ps=6.74e-06 pd=4.5e-06 
+ nrs=0.78 nrd=0.3 
m8781 4219 25 4164 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.83e-12 ad=9.35e-12 ps=8.66e-06 pd=1.017e-05 
+ nrs=0.6 nrd=0.72 
m8782 4223 26 4219 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.52e-12 ad=7.83e-12 ps=7.76e-06 pd=8.66e-06 
+ nrs=0.58 nrd=0.6 
m8783 1 4228 4225 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=3.08e-11 ps=2.114e-05 pd=2.85e-05 
+ nrs=0.2 nrd=0.25 
m8784 0 37 4219 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=6.09e-12 ps=5.25e-06 pd=6.74e-06 
+ nrs=0.71 nrd=0.78 
m8785 4229 4226 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m8786 4223 4217 4229 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.169e-11 ad=4.76e-12 ps=1.207e-05 pd=7.3e-06 
+ nrs=0.37 nrd=0.15 
m8787 4230 4225 4223 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.169e-11 ps=7.3e-06 pd=1.207e-05 
+ nrs=0.15 nrd=0.37 
m8788 0 3918 4230 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m8789 4226 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m8790 0 4228 4225 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m8791 0 4232 4231 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m8792 4233 4234 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m8793 0 3381 4233 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m8794 4235 4234 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m8795 4232 3381 4235 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m8796 4233 3384 4232 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m8797 4236 3384 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m8798 4237 4232 4236 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m8799 1 4232 4231 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m8800 4238 3381 4237 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m8801 4239 3384 4238 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m8802 0 4234 4239 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m8803 4236 3381 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m8804 0 4234 4236 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m8805 4240 4234 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m8806 4241 3381 4240 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m8807 4232 4234 4241 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m8808 4241 3381 4232 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m8809 4242 4237 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m8810 1 3384 4241 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m8811 4237 4232 4243 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m8812 4244 3381 4237 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m8813 4245 3384 4244 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m8814 4234 4246 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m8815 4246 4247 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8816 4243 4234 4245 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m8817 1 3381 4243 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m8818 4243 4234 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m8819 1 3384 4243 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m8820 4242 4237 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m8821 0 4246 4234 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m8822 0 4247 4246 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m8823 0 3886 4247 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m8824 4247 3900 612 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m8825 601 3876 4247 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m8826 4247 3898 602 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.045e-11 ps=8.18e-06 pd=1.269e-05 
+ nrs=0.54 nrd=0.81 
m8827 595 3882 4247 0 nenh l=1.1e-06 w=3.6e-06 
+ as=9.95e-12 ad=6.95e-12 ps=1.239e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m8828 0 4249 4248 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m8829 4250 4251 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m8830 0 3385 4250 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m8831 4252 4251 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m8832 4249 3385 4252 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m8833 4250 3418 4249 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m8834 4253 3418 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m8835 4254 4249 4253 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m8836 1 4249 4248 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m8837 4255 3385 4254 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m8838 4256 3418 4255 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m8839 0 4251 4256 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m8840 4253 3385 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m8841 0 4251 4253 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m8842 4257 4251 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m8843 4258 3385 4257 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m8844 4249 4251 4258 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m8845 4258 3385 4249 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m8846 4259 4254 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m8847 1 3418 4258 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m8848 4254 4249 4260 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m8849 4261 3385 4254 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m8850 4262 3418 4261 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m8851 4251 4263 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m8852 4263 4264 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8853 4260 4251 4262 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m8854 1 3385 4260 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m8855 4260 4251 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m8856 1 3418 4260 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m8857 4259 4254 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m8858 0 4263 4251 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m8859 0 4264 4263 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m8860 0 3886 4264 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m8861 4264 3900 627 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m8862 617 3876 4264 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m8863 4264 3898 601 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m8864 612 3882 4264 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m8865 0 4266 4265 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m8866 4267 4268 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m8867 0 3429 4267 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m8868 4269 4268 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m8869 4266 3429 4269 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m8870 4267 3435 4266 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m8871 4270 3435 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m8872 4271 4266 4270 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m8873 1 4266 4265 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m8874 4272 3429 4271 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m8875 4273 3435 4272 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m8876 0 4268 4273 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m8877 4270 3429 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m8878 0 4268 4270 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m8879 4274 4268 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m8880 4275 3429 4274 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m8881 4266 4268 4275 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m8882 4275 3429 4266 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m8883 4276 4271 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m8884 1 3435 4275 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m8885 4271 4266 4277 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m8886 4278 3429 4271 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m8887 4279 3435 4278 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m8888 4268 4280 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m8889 4280 4281 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8890 4277 4268 4279 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m8891 1 3429 4277 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m8892 4277 4268 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m8893 1 3435 4277 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m8894 4276 4271 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m8895 0 4280 4268 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m8896 0 4281 4280 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m8897 0 3886 4281 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m8898 4281 3900 642 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m8899 632 3876 4281 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m8900 4281 3898 617 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m8901 627 3882 4281 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m8902 0 4283 4282 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m8903 4284 4285 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m8904 0 3446 4284 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m8905 4286 4285 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m8906 4283 3446 4286 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m8907 4284 3452 4283 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m8908 4287 3452 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m8909 4288 4283 4287 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m8910 1 4283 4282 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m8911 4289 3446 4288 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m8912 4290 3452 4289 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m8913 0 4285 4290 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m8914 4287 3446 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m8915 0 4285 4287 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m8916 4291 4285 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m8917 4292 3446 4291 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m8918 4283 4285 4292 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m8919 4292 3446 4283 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m8920 4293 4288 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m8921 1 3452 4292 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m8922 4288 4283 4294 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m8923 4295 3446 4288 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m8924 4296 3452 4295 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m8925 4285 4297 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m8926 4297 4298 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8927 4294 4285 4296 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m8928 1 3446 4294 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m8929 4294 4285 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m8930 1 3452 4294 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m8931 4293 4288 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m8932 0 4297 4285 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m8933 0 4298 4297 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m8934 0 3886 4298 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m8935 4298 3900 657 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m8936 647 3876 4298 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m8937 4298 3898 632 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m8938 642 3882 4298 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m8939 0 4300 4299 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m8940 4301 4302 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m8941 0 3463 4301 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m8942 4303 4302 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m8943 4300 3463 4303 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m8944 4301 3469 4300 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m8945 4304 3469 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m8946 4305 4300 4304 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m8947 1 4300 4299 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m8948 4306 3463 4305 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m8949 4307 3469 4306 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m8950 0 4302 4307 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m8951 4304 3463 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m8952 0 4302 4304 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m8953 4308 4302 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m8954 4309 3463 4308 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m8955 4300 4302 4309 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m8956 4309 3463 4300 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m8957 4310 4305 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m8958 1 3469 4309 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m8959 4305 4300 4311 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m8960 4312 3463 4305 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m8961 4313 3469 4312 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m8962 4302 4314 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m8963 4314 4315 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m8964 4311 4302 4313 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m8965 1 3463 4311 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m8966 4311 4302 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m8967 1 3469 4311 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m8968 4310 4305 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m8969 0 4314 4302 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m8970 0 4315 4314 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m8971 0 3886 4315 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m8972 4315 3900 672 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m8973 662 3876 4315 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m8974 4315 3898 647 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m8975 657 3882 4315 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m8976 0 4317 4316 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m8977 4318 4319 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m8978 0 3480 4318 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m8979 4320 4319 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m8980 4317 3480 4320 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m8981 4318 3486 4317 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m8982 4321 3486 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m8983 4322 4317 4321 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m8984 1 4317 4316 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m8985 4323 3480 4322 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m8986 4324 3486 4323 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m8987 0 4319 4324 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m8988 4321 3480 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m8989 0 4319 4321 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m8990 4325 4319 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m8991 4326 3480 4325 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m8992 4317 4319 4326 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m8993 4326 3480 4317 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m8994 4327 4322 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m8995 1 3486 4326 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m8996 4322 4317 4328 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m8997 4329 3480 4322 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m8998 4330 3486 4329 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m8999 4319 4331 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9000 4331 4332 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9001 4328 4319 4330 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9002 1 3480 4328 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9003 4328 4319 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9004 1 3486 4328 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9005 4327 4322 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m9006 0 4331 4319 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9007 0 4332 4331 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9008 0 3886 4332 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9009 4332 3900 687 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9010 677 3876 4332 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9011 4332 3898 662 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9012 672 3882 4332 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9013 0 4334 4333 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m9014 4335 4336 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m9015 0 3497 4335 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m9016 4337 4336 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m9017 4334 3497 4337 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m9018 4335 3503 4334 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m9019 4338 3503 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9020 4339 4334 4338 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9021 1 4334 4333 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m9022 4340 3497 4339 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m9023 4341 3503 4340 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m9024 0 4336 4341 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m9025 4338 3497 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9026 0 4336 4338 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9027 4342 4336 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m9028 4343 3497 4342 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m9029 4334 4336 4343 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9030 4343 3497 4334 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9031 4344 4339 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m9032 1 3503 4343 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9033 4339 4334 4345 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9034 4346 3497 4339 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9035 4347 3503 4346 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9036 4336 4348 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9037 4348 4349 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9038 4345 4336 4347 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9039 1 3497 4345 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9040 4345 4336 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9041 1 3503 4345 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9042 4344 4339 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m9043 0 4348 4336 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9044 0 4349 4348 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9045 0 3886 4349 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9046 4349 3900 702 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9047 692 3876 4349 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9048 4349 3898 677 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9049 687 3882 4349 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9050 0 4351 4350 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m9051 4352 4353 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m9052 0 3514 4352 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m9053 4354 4353 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m9054 4351 3514 4354 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m9055 4352 3520 4351 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m9056 4355 3520 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9057 4356 4351 4355 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9058 1 4351 4350 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m9059 4357 3514 4356 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m9060 4358 3520 4357 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m9061 0 4353 4358 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m9062 4355 3514 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9063 0 4353 4355 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9064 4359 4353 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m9065 4360 3514 4359 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m9066 4351 4353 4360 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9067 4360 3514 4351 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9068 4361 4356 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m9069 1 3520 4360 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9070 4356 4351 4362 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9071 4363 3514 4356 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9072 4364 3520 4363 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9073 4353 4365 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9074 4365 4366 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9075 4362 4353 4364 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9076 1 3514 4362 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9077 4362 4353 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9078 1 3520 4362 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9079 4361 4356 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m9080 0 4365 4353 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9081 0 4366 4365 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9082 0 3886 4366 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9083 4366 3900 717 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9084 707 3876 4366 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9085 4366 3898 692 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9086 702 3882 4366 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9087 0 4368 4367 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m9088 4369 4370 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m9089 0 3531 4369 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m9090 4371 4370 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m9091 4368 3531 4371 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m9092 4369 3537 4368 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m9093 4372 3537 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9094 4373 4368 4372 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9095 1 4368 4367 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m9096 4374 3531 4373 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m9097 4375 3537 4374 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m9098 0 4370 4375 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m9099 4372 3531 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9100 0 4370 4372 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9101 4376 4370 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m9102 4377 3531 4376 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m9103 4368 4370 4377 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9104 4377 3531 4368 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9105 4378 4373 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m9106 1 3537 4377 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9107 4373 4368 4379 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9108 4380 3531 4373 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9109 4381 3537 4380 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9110 4370 4382 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9111 4382 4383 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9112 4379 4370 4381 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9113 1 3531 4379 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9114 4379 4370 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9115 1 3537 4379 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9116 4378 4373 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m9117 0 4382 4370 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9118 0 4383 4382 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9119 0 3886 4383 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9120 4383 3900 732 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9121 722 3876 4383 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9122 4383 3898 707 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9123 717 3882 4383 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9124 0 4385 4384 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m9125 4386 4387 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m9126 0 3548 4386 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m9127 4388 4387 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m9128 4385 3548 4388 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m9129 4386 3554 4385 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m9130 4389 3554 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9131 4390 4385 4389 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9132 1 4385 4384 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m9133 4391 3548 4390 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m9134 4392 3554 4391 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m9135 0 4387 4392 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m9136 4389 3548 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9137 0 4387 4389 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9138 4393 4387 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m9139 4394 3548 4393 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m9140 4385 4387 4394 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9141 4394 3548 4385 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9142 4395 4390 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m9143 1 3554 4394 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9144 4390 4385 4396 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9145 4397 3548 4390 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9146 4398 3554 4397 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9147 4387 4399 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9148 4399 4400 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9149 4396 4387 4398 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9150 1 3548 4396 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9151 4396 4387 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9152 1 3554 4396 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9153 4395 4390 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m9154 0 4399 4387 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9155 0 4400 4399 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9156 0 3886 4400 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9157 4400 3900 747 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9158 737 3876 4400 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9159 4400 3898 722 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9160 732 3882 4400 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9161 0 4402 4401 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m9162 4403 4404 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m9163 0 3565 4403 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m9164 4405 4404 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m9165 4402 3565 4405 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m9166 4403 3571 4402 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m9167 4406 3571 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9168 4407 4402 4406 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9169 1 4402 4401 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m9170 4408 3565 4407 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m9171 4409 3571 4408 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m9172 0 4404 4409 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m9173 4406 3565 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9174 0 4404 4406 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9175 4410 4404 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m9176 4411 3565 4410 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m9177 4402 4404 4411 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9178 4411 3565 4402 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9179 4412 4407 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m9180 1 3571 4411 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9181 4407 4402 4413 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9182 4414 3565 4407 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9183 4415 3571 4414 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9184 4404 4416 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9185 4416 4417 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9186 4413 4404 4415 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9187 1 3565 4413 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9188 4413 4404 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9189 1 3571 4413 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9190 4412 4407 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m9191 0 4416 4404 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9192 0 4417 4416 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9193 0 3886 4417 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9194 4417 3900 762 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9195 752 3876 4417 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9196 4417 3898 737 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9197 747 3882 4417 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9198 0 4419 4418 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m9199 4420 4421 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m9200 0 3582 4420 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m9201 4422 4421 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m9202 4419 3582 4422 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m9203 4420 3588 4419 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m9204 4423 3588 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9205 4424 4419 4423 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9206 1 4419 4418 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m9207 4425 3582 4424 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m9208 4426 3588 4425 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m9209 0 4421 4426 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m9210 4423 3582 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9211 0 4421 4423 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9212 4427 4421 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m9213 4428 3582 4427 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m9214 4419 4421 4428 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9215 4428 3582 4419 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9216 4429 4424 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m9217 1 3588 4428 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9218 4424 4419 4430 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9219 4431 3582 4424 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9220 4432 3588 4431 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9221 4421 4433 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9222 4433 4434 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9223 4430 4421 4432 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9224 1 3582 4430 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9225 4430 4421 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9226 1 3588 4430 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9227 4429 4424 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m9228 0 4433 4421 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9229 0 4434 4433 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9230 0 3886 4434 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9231 4434 3900 777 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9232 767 3876 4434 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9233 4434 3898 752 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9234 762 3882 4434 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9235 0 4436 4435 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m9236 4437 4438 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m9237 0 3599 4437 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m9238 4439 4438 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m9239 4436 3599 4439 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m9240 4437 3605 4436 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m9241 4440 3605 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9242 4441 4436 4440 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9243 1 4436 4435 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m9244 4442 3599 4441 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m9245 4443 3605 4442 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m9246 0 4438 4443 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m9247 4440 3599 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9248 0 4438 4440 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9249 4444 4438 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m9250 4445 3599 4444 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m9251 4436 4438 4445 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9252 4445 3599 4436 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9253 4446 4441 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m9254 1 3605 4445 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9255 4441 4436 4447 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9256 4448 3599 4441 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9257 4449 3605 4448 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9258 4438 4450 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9259 4450 4451 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9260 4447 4438 4449 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9261 1 3599 4447 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9262 4447 4438 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9263 1 3605 4447 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9264 4446 4441 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m9265 0 4450 4438 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9266 0 4451 4450 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9267 0 3886 4451 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9268 4451 3900 792 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9269 782 3876 4451 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9270 4451 3898 767 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9271 777 3882 4451 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9272 0 4453 4452 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m9273 4454 4455 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m9274 0 3616 4454 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m9275 4456 4455 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m9276 4453 3616 4456 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m9277 4454 3622 4453 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m9278 4457 3622 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9279 4458 4453 4457 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9280 1 4453 4452 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m9281 4459 3616 4458 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m9282 4460 3622 4459 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m9283 0 4455 4460 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m9284 4457 3616 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9285 0 4455 4457 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9286 4461 4455 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m9287 4462 3616 4461 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m9288 4453 4455 4462 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9289 4462 3616 4453 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9290 4463 4458 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m9291 1 3622 4462 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9292 4458 4453 4464 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9293 4465 3616 4458 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9294 4466 3622 4465 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9295 4455 4467 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9296 4467 4468 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9297 4464 4455 4466 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9298 1 3616 4464 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9299 4464 4455 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9300 1 3622 4464 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9301 4463 4458 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m9302 0 4467 4455 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9303 0 4468 4467 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9304 0 3886 4468 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9305 4468 3900 807 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9306 797 3876 4468 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9307 4468 3898 782 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9308 792 3882 4468 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9309 0 4470 4469 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m9310 4471 4472 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m9311 0 3633 4471 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m9312 4473 4472 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m9313 4470 3633 4473 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m9314 4471 3639 4470 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m9315 4474 3639 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9316 4475 4470 4474 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9317 1 4470 4469 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m9318 4476 3633 4475 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m9319 4477 3639 4476 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m9320 0 4472 4477 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m9321 4474 3633 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9322 0 4472 4474 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9323 4478 4472 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m9324 4479 3633 4478 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m9325 4470 4472 4479 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9326 4479 3633 4470 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9327 4480 4475 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m9328 1 3639 4479 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9329 4475 4470 4481 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9330 4482 3633 4475 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9331 4483 3639 4482 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9332 4472 4484 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9333 4484 4485 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9334 4481 4472 4483 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9335 1 3633 4481 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9336 4481 4472 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9337 1 3639 4481 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9338 4480 4475 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m9339 0 4484 4472 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9340 0 4485 4484 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9341 0 3886 4485 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9342 4485 3900 822 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9343 812 3876 4485 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9344 4485 3898 797 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9345 807 3882 4485 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9346 0 4487 4486 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m9347 4488 4489 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m9348 0 3650 4488 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m9349 4490 4489 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m9350 4487 3650 4490 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m9351 4488 3656 4487 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m9352 4491 3656 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9353 4492 4487 4491 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9354 1 4487 4486 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m9355 4493 3650 4492 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m9356 4494 3656 4493 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m9357 0 4489 4494 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m9358 4491 3650 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9359 0 4489 4491 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9360 4495 4489 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m9361 4496 3650 4495 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m9362 4487 4489 4496 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9363 4496 3650 4487 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9364 4497 4492 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m9365 1 3656 4496 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9366 4492 4487 4498 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9367 4499 3650 4492 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9368 4500 3656 4499 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9369 4489 4501 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9370 4501 4502 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9371 4498 4489 4500 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9372 1 3650 4498 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9373 4498 4489 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9374 1 3656 4498 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9375 4497 4492 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m9376 0 4501 4489 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9377 0 4502 4501 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9378 0 3886 4502 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9379 4502 3900 837 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9380 827 3876 4502 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9381 4502 3898 812 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9382 822 3882 4502 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9383 0 4504 4503 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m9384 4505 4506 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m9385 0 3667 4505 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m9386 4507 4506 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m9387 4504 3667 4507 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m9388 4505 3673 4504 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m9389 4508 3673 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9390 4509 4504 4508 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9391 1 4504 4503 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m9392 4510 3667 4509 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m9393 4511 3673 4510 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m9394 0 4506 4511 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m9395 4508 3667 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9396 0 4506 4508 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9397 4512 4506 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m9398 4513 3667 4512 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m9399 4504 4506 4513 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9400 4513 3667 4504 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9401 4514 4509 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m9402 1 3673 4513 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9403 4509 4504 4515 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9404 4516 3667 4509 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9405 4517 3673 4516 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9406 4506 4518 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9407 4518 4519 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9408 4515 4506 4517 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9409 1 3667 4515 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9410 4515 4506 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9411 1 3673 4515 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9412 4514 4509 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m9413 0 4518 4506 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9414 0 4519 4518 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9415 0 3886 4519 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9416 4519 3900 868 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9417 842 3876 4519 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9418 4519 3898 827 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9419 837 3882 4519 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9420 0 4521 4520 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m9421 4522 4523 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.249e-11 ad=2.933e-11 ps=2.223e-05 pd=2.774e-05 
+ nrs=0.1 nrd=0.13 
m9422 0 3684 4522 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=2.249e-11 ps=2.774e-05 pd=2.223e-05 
+ nrs=0.13 nrd=0.1 
m9423 4524 4523 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.377e-11 ad=3.171e-11 ps=1.863e-05 pd=2.999e-05 
+ nrs=0.05 nrd=0.12 
m9424 4521 3684 4524 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.239e-11 ps=1.795e-05 pd=1.677e-05 
+ nrs=0.07 nrd=0.06 
m9425 4522 3690 4521 0 nenh l=1.1e-06 w=1.4e-05 
+ as=2.128e-11 ad=1.383e-11 ps=2.103e-05 pd=1.745e-05 
+ nrs=0.11 nrd=0.07 
m9426 4525 3690 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9427 4526 4521 4525 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.53e-11 ad=1.404e-11 ps=1.85e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9428 1 4521 4520 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.288e-11 ps=3.323e-05 pd=3.73e-05 
+ nrs=0.13 nrd=0.11 
m9429 4527 3684 4526 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.53e-11 ps=1.701e-05 pd=1.85e-05 
+ nrs=0.06 nrd=0.07 
m9430 4528 3690 4527 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m9431 0 4523 4528 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m9432 4525 3684 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9433 0 4523 4525 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9434 4529 4523 1 1 penh l=1.1e-06 w=1.76e-05 
+ as=1.504e-11 ad=3.919e-11 ps=1.975e-05 pd=3.323e-05 
+ nrs=0.05 nrd=0.13 
m9435 4530 3684 4529 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.436e-11 ps=1.967e-05 pd=1.885e-05 
+ nrs=0.06 nrd=0.05 
m9436 4521 4523 4530 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9437 4530 3684 4521 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9438 4531 4526 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m9439 1 3690 4530 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9440 4526 4521 4532 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9441 4533 3684 4526 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9442 4534 3690 4533 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9443 4523 4535 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9444 4535 4536 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9445 4532 4523 4534 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9446 1 3684 4532 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9447 4532 4523 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9448 1 3690 4532 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9449 4531 4526 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.488e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.09 nrd=0.12 
m9450 0 4535 4523 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.824e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9451 0 4536 4535 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9452 0 3886 4536 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9453 4536 3900 852 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9454 858 3876 4536 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.036e-11 ad=6.95e-12 ps=1.246e-05 pd=8.18e-06 
+ nrs=0.8 nrd=0.54 
m9455 4536 3898 842 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9456 868 3882 4536 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9457 0 4538 4537 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=3.144e-11 ps=2.699e-05 pd=3.25e-05 
+ nrs=0.14 nrd=0.15 
m9458 4539 4540 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.083e-11 ad=3.013e-11 ps=2.27e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m9459 0 3701 4539 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.083e-11 ps=2.849e-05 pd=2.27e-05 
+ nrs=0.13 nrd=0.09 
m9460 4541 4540 0 0 nenh l=1.1e-06 w=1.68e-05 
+ as=1.454e-11 ad=3.33e-11 ps=1.992e-05 pd=3.149e-05 
+ nrs=0.05 nrd=0.12 
m9461 4538 3701 4541 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.246e-11 ps=1.795e-05 pd=1.708e-05 
+ nrs=0.07 nrd=0.06 
m9462 4539 3707 4538 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.919e-11 ad=1.383e-11 ps=2.091e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m9463 4542 3707 0 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.352e-11 ad=2.854e-11 ps=1.61e-05 pd=2.699e-05 
+ nrs=0.07 nrd=0.14 
m9464 4543 4538 4542 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.449e-11 ad=1.352e-11 ps=1.785e-05 pd=1.61e-05 
+ nrs=0.07 nrd=0.07 
m9465 4544 3701 4543 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.489e-11 ps=1.701e-05 pd=1.835e-05 
+ nrs=0.06 nrd=0.07 
m9466 4545 3707 4544 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m9467 0 4540 4545 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m9468 4542 3701 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.502e-11 ad=3.171e-11 ps=1.789e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9469 0 4540 4542 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.202e-11 ps=2.399e-05 pd=1.431e-05 
+ nrs=0.15 nrd=0.07 
m9470 1 4538 4537 1 penh l=1.1e-06 w=1.8e-05 
+ as=4.008e-11 ad=3.314e-11 ps=3.398e-05 pd=3.89e-05 
+ nrs=0.12 nrd=0.1 
m9471 4546 4543 0 0 nenh l=1.1e-06 w=2.12e-05 
+ as=3.138e-11 ad=4.202e-11 ps=4.21e-05 pd=3.974e-05 
+ nrs=0.07 nrd=0.09 
m9472 4547 4540 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m9473 4548 3701 4547 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m9474 4538 4540 4548 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.615e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9475 4548 3701 4538 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.499e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.06 
m9476 1 3707 4548 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9477 1 4550 4549 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.484e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.47 
m9478 4551 3900 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m9479 4550 3882 4551 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.372e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.44 nrd=0.15 
m9480 1 4552 4540 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=2.226e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.32 
m9481 4543 4538 4553 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.447e-11 ad=1.386e-11 ps=1.722e-05 pd=1.719e-05 
+ nrs=0.1 nrd=0.1 
m9482 4554 3701 4543 1 penh l=1.1e-06 w=1.88e-05 
+ as=1.621e-11 ad=2.267e-11 ps=2.153e-05 pd=2.698e-05 
+ nrs=0.05 nrd=0.06 
m9483 4555 3707 4554 1 penh l=1.1e-06 w=2.12e-05 
+ as=1.814e-11 ad=1.827e-11 ps=2.344e-05 pd=2.427e-05 
+ nrs=0.04 nrd=0.04 
m9484 4553 4540 4555 1 penh l=1.1e-06 w=2.24e-05 
+ as=2.588e-11 ad=1.916e-11 ps=3.21e-05 pd=2.476e-05 
+ nrs=0.05 nrd=0.04 
m9485 1 3701 4553 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.664e-11 ps=2.718e-05 pd=2.063e-05 
+ nrs=0.15 nrd=0.08 
m9486 4553 4540 1 1 penh l=1.1e-06 w=1.52e-05 
+ as=1.756e-11 ad=3.384e-11 ps=2.178e-05 pd=2.869e-05 
+ nrs=0.08 nrd=0.15 
m9487 1 3707 4553 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.386e-11 ps=2.265e-05 pd=1.719e-05 
+ nrs=0.19 nrd=0.1 
m9488 4546 4543 1 1 penh l=1.1e-06 w=1.92e-05 
+ as=3.04e-11 ad=4.275e-11 ps=4.13e-05 pd=3.625e-05 
+ nrs=0.08 nrd=0.12 
m9489 4552 4556 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.298e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.48 nrd=0.43 
m9490 0 4550 4549 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m9491 4550 3900 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=5.55e-12 ps=6.1e-06 pd=5.25e-06 
+ nrs=0.59 nrd=0.71 
m9492 0 3882 4550 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=4.62e-12 ps=5.25e-06 pd=6.1e-06 
+ nrs=0.71 nrd=0.59 
m9493 0 4552 4540 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.52e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.37 
m9494 0 4556 4552 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9495 0 3886 4556 0 nenh l=1.1e-06 w=3.2e-06 
+ as=6.34e-12 ad=6.09e-12 ps=6e-06 pd=7.29e-06 
+ nrs=0.62 nrd=0.6 
m9496 4556 3900 1 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.098e-11 ps=8.2e-06 pd=1.406e-05 
+ nrs=0.53 nrd=0.85 
m9497 0 3876 4556 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.86e-12 ps=6.75e-06 pd=8.2e-06 
+ nrs=0.55 nrd=0.53 
m9498 4556 3898 858 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.036e-11 ps=8.2e-06 pd=1.246e-05 
+ nrs=0.53 nrd=0.8 
m9499 852 3882 4556 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.86e-12 ps=1.202e-05 pd=8.2e-06 
+ nrs=0.77 nrd=0.53 
m9500 0 4558 4557 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.427e-11 ad=2.196e-11 ps=1.35e-05 pd=2.05e-05 
+ nrs=0.28 nrd=0.42 
m9501 4558 4559 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m9502 4560 4197 4561 0 nenh l=1.1e-06 w=8.8e-06 
+ as=7.66e-12 ad=1.964e-11 ps=1.122e-05 pd=2.37e-05 
+ nrs=0.1 nrd=0.25 
m9503 4562 4214 4560 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.4e-12 ps=1.25e-05 pd=1.378e-05 
+ nrs=0.08 nrd=0.08 
m9504 0 3890 4562 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m9505 4563 4197 0 0 nenh l=1.1e-06 w=8.8e-06 
+ as=9.24e-12 ad=1.744e-11 ps=1.13e-05 pd=1.65e-05 
+ nrs=0.12 nrd=0.23 
m9506 0 4564 4563 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.744e-11 ad=9.24e-12 ps=1.65e-05 pd=1.13e-05 
+ nrs=0.23 nrd=0.12 
m9507 4565 4566 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=1.665e-11 ps=1.01e-05 pd=1.575e-05 
+ nrs=0.1 nrd=0.24 
m9508 4567 4568 4565 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.89e-11 ad=7.14e-12 ps=2.29e-05 pd=1.01e-05 
+ nrs=0.27 nrd=0.1 
m9509 0 4570 4569 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=1.22e-11 ps=7.5e-06 pd=1.41e-05 
+ nrs=0.5 nrd=0.76 
m9510 4571 4561 0 0 nenh l=1.1e-06 w=4e-06 
+ as=6.6e-12 ad=7.93e-12 ps=7.3e-06 pd=7.5e-06 
+ nrs=0.41 nrd=0.5 
m9511 0 4561 4571 0 nenh l=1.1e-06 w=4e-06 
+ as=7.93e-12 ad=6.6e-12 ps=7.5e-06 pd=7.3e-06 
+ nrs=0.5 nrd=0.41 
m9512 1 4558 4557 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m9513 4558 4559 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9514 1 4570 4569 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=2.358e-11 ps=1.737e-05 pd=2.29e-05 
+ nrs=0.24 nrd=0.28 
m9515 4571 4561 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.128e-11 ad=2.494e-11 ps=1.37e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m9516 1 4561 4571 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.128e-11 ps=2.114e-05 pd=1.37e-05 
+ nrs=0.2 nrd=0.09 
m9517 4572 4214 4568 0 nenh l=1.1e-06 w=9.6e-06 
+ as=8.27e-12 ad=2.16e-11 ps=1.176e-05 pd=2.53e-05 
+ nrs=0.09 nrd=0.23 
m9518 4573 3890 4572 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=9.31e-12 ps=1.25e-05 pd=1.324e-05 
+ nrs=0.08 nrd=0.08 
m9519 0 4196 4573 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=9.18e-12 ps=2.024e-05 pd=1.25e-05 
+ nrs=0.18 nrd=0.08 
m9520 4574 4197 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m9521 4575 4215 4574 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.31e-12 ad=9.18e-12 ps=1.324e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m9522 4566 3879 4575 0 nenh l=1.1e-06 w=9.6e-06 
+ as=2.16e-11 ad=8.27e-12 ps=2.53e-05 pd=1.176e-05 
+ nrs=0.23 nrd=0.09 
m9523 1 4197 4561 1 penh l=1.1e-06 w=9.6e-06 
+ as=2.137e-11 ad=1.315e-11 ps=1.812e-05 pd=1.587e-05 
+ nrs=0.23 nrd=0.14 
m9524 4561 4214 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.26e-11 ad=2.048e-11 ps=1.521e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m9525 1 3890 4561 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.26e-11 ps=1.737e-05 pd=1.521e-05 
+ nrs=0.24 nrd=0.15 
m9526 4576 4197 1 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.194e-11 ad=2.939e-11 ps=1.49e-05 pd=2.492e-05 
+ nrs=0.07 nrd=0.17 
m9527 4563 4564 4576 1 penh l=1.1e-06 w=1.32e-05 
+ as=2.586e-11 ad=1.194e-11 ps=3.01e-05 pd=1.49e-05 
+ nrs=0.15 nrd=0.07 
m9528 4567 4566 1 1 penh l=1.1e-06 w=1.48e-05 
+ as=1.466e-11 ad=3.295e-11 ps=1.73e-05 pd=2.794e-05 
+ nrs=0.07 nrd=0.15 
m9529 1 4568 4567 1 penh l=1.1e-06 w=1.48e-05 
+ as=3.295e-11 ad=1.466e-11 ps=2.794e-05 pd=1.73e-05 
+ nrs=0.15 nrd=0.07 
m9530 1 4214 4568 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m9531 4568 3890 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m9532 1 4196 4568 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m9533 4566 4197 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m9534 1 4215 4566 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.275e-11 ps=1.737e-05 pd=1.543e-05 
+ nrs=0.24 nrd=0.15 
m9535 4566 3879 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.275e-11 ad=2.048e-11 ps=1.543e-05 pd=1.737e-05 
+ nrs=0.15 nrd=0.24 
m9536 4570 4577 1 1 penh l=1.1e-06 w=1e-05 
+ as=2.346e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.23 nrd=0.22 
m9537 4577 4578 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.26e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.4 nrd=0.4 
m9538 4559 4567 1 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=8.54e-12 ps=7.22e-06 pd=1.094e-05 
+ nrs=0.69 nrd=1.09 
m9539 910 4571 4559 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m9540 4579 4564 4580 1 penh l=1.1e-06 w=1.04e-05 
+ as=8.84e-12 ad=2.276e-11 ps=1.21e-05 pd=2.69e-05 
+ nrs=0.08 nrd=0.21 
m9541 1 4196 4579 1 penh l=1.1e-06 w=1.04e-05 
+ as=2.316e-11 ad=8.84e-12 ps=1.963e-05 pd=1.21e-05 
+ nrs=0.21 nrd=0.08 
m9542 4581 3879 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m9543 1 4215 4581 1 penh l=1.1e-06 w=8e-06 
+ as=1.781e-11 ad=1.075e-11 ps=1.51e-05 pd=1.383e-05 
+ nrs=0.28 nrd=0.17 
m9544 4581 4196 1 1 penh l=1.1e-06 w=8e-06 
+ as=1.075e-11 ad=1.781e-11 ps=1.383e-05 pd=1.51e-05 
+ nrs=0.17 nrd=0.28 
m9545 4582 4581 1 1 penh l=1.1e-06 w=1e-05 
+ as=1.058e-11 ad=2.227e-11 ps=1.25e-05 pd=1.888e-05 
+ nrs=0.11 nrd=0.22 
m9546 1 4581 4582 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=1.058e-11 ps=1.888e-05 pd=1.25e-05 
+ nrs=0.22 nrd=0.11 
m9547 911 4582 4559 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m9548 4559 4563 911 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.91e-12 ps=7.22e-06 pd=1.05e-05 
+ nrs=0.69 nrd=1.01 
m9549 910 4580 4559 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.88e-12 ad=5.4e-12 ps=1.048e-05 pd=7.22e-06 
+ nrs=1 nrd=0.69 
m9550 4578 4582 595 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.74e-12 ps=7.22e-06 pd=9.64e-06 
+ nrs=0.69 nrd=0.99 
m9551 602 4571 4578 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=5.4e-12 ps=9.87e-06 pd=7.22e-06 
+ nrs=1.04 nrd=0.69 
m9552 4578 4563 910 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.4e-12 ad=7.88e-12 ps=7.22e-06 pd=1.048e-05 
+ nrs=0.69 nrd=1 
m9553 911 4580 4578 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.91e-12 ad=5.4e-12 ps=1.05e-05 pd=7.22e-06 
+ nrs=1.01 nrd=0.69 
m9554 0 4567 4578 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=5.4e-12 ps=5.25e-06 pd=7.22e-06 
+ nrs=0.71 nrd=0.69 
m9555 4583 4215 1 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=2.405e-11 ps=1.41e-05 pd=2.039e-05 
+ nrs=0.09 nrd=0.21 
m9556 4564 3879 4583 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.046e-11 ad=1.014e-11 ps=1.25e-05 pd=1.41e-05 
+ nrs=0.09 nrd=0.09 
m9557 4584 3890 4564 1 penh l=1.1e-06 w=1.08e-05 
+ as=1.014e-11 ad=1.046e-11 ps=1.41e-05 pd=1.25e-05 
+ nrs=0.09 nrd=0.09 
m9558 1 4214 4584 1 penh l=1.1e-06 w=1.08e-05 
+ as=2.405e-11 ad=1.014e-11 ps=2.039e-05 pd=1.41e-05 
+ nrs=0.21 nrd=0.09 
m9559 0 4577 4570 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.888e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.46 
m9560 0 4578 4577 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.372e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.44 
m9561 4580 4564 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m9562 0 4196 4580 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m9563 4585 3879 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.18e-12 ad=2.141e-11 ps=1.25e-05 pd=2.024e-05 
+ nrs=0.08 nrd=0.18 
m9564 4586 4215 4585 0 nenh l=1.1e-06 w=1.08e-05 
+ as=9.4e-12 ad=9.18e-12 ps=1.378e-05 pd=1.25e-05 
+ nrs=0.08 nrd=0.08 
m9565 4581 4196 4586 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.964e-11 ad=7.66e-12 ps=2.37e-05 pd=1.122e-05 
+ nrs=0.25 nrd=0.1 
m9566 4582 4581 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=7.54e-12 ad=1.348e-11 ps=9.3e-06 pd=1.275e-05 
+ nrs=0.16 nrd=0.29 
m9567 0 4581 4582 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=7.54e-12 ps=1.275e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.16 
m9568 4587 4215 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=9.84e-12 ad=2.061e-11 ps=1.319e-05 pd=1.949e-05 
+ nrs=0.09 nrd=0.19 
m9569 4564 3890 4587 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.08e-11 ad=1.06e-11 ps=1.29e-05 pd=1.421e-05 
+ nrs=0.09 nrd=0.08 
m9570 4588 3879 4564 0 nenh l=1.1e-06 w=1.12e-05 
+ as=1.062e-11 ad=1.08e-11 ps=1.436e-05 pd=1.29e-05 
+ nrs=0.08 nrd=0.09 
m9571 0 4214 4588 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.024e-11 ps=2.024e-05 pd=1.384e-05 
+ nrs=0.18 nrd=0.09 
m9572 0 4590 4589 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m9573 4591 4592 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m9574 0 3870 4591 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m9575 4593 4592 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m9576 4590 3870 4593 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m9577 4591 3873 4590 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m9578 4594 3873 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9579 4595 4590 4594 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9580 4596 3870 4595 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m9581 4597 3873 4596 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m9582 0 4592 4597 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m9583 4594 3870 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9584 0 4592 4594 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9585 1 4590 4589 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m9586 4598 4592 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m9587 4599 3870 4598 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m9588 4590 4592 4599 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9589 4599 3870 4590 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9590 4600 4595 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m9591 1 3873 4599 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9592 4595 4590 4601 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9593 4602 3870 4595 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9594 4603 3873 4602 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9595 4601 4592 4603 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9596 1 3870 4601 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9597 4601 4592 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9598 1 3873 4601 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9599 4592 4604 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9600 4604 4605 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9601 4600 4595 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m9602 0 4604 4592 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9603 0 4605 4604 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9604 0 4567 4605 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9605 4605 4582 612 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9606 601 4571 4605 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9607 4605 4580 602 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.045e-11 ps=8.18e-06 pd=1.269e-05 
+ nrs=0.54 nrd=0.81 
m9608 595 4563 4605 0 nenh l=1.1e-06 w=3.6e-06 
+ as=9.95e-12 ad=6.95e-12 ps=1.239e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9609 0 4607 4606 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m9610 4608 4609 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m9611 0 3874 4608 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m9612 4610 4609 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m9613 4607 3874 4610 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m9614 4608 4231 4607 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m9615 4611 4231 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9616 4612 4607 4611 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9617 4613 3874 4612 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m9618 4614 4231 4613 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m9619 0 4609 4614 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m9620 4611 3874 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9621 0 4609 4611 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9622 1 4607 4606 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m9623 4615 4609 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m9624 4616 3874 4615 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m9625 4607 4609 4616 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9626 4616 3874 4607 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9627 4617 4612 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m9628 1 4231 4616 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9629 4612 4607 4618 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9630 4619 3874 4612 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9631 4620 4231 4619 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9632 4618 4609 4620 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9633 1 3874 4618 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9634 4618 4609 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9635 1 4231 4618 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9636 4609 4621 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9637 4621 4622 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9638 4617 4612 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m9639 0 4621 4609 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9640 0 4622 4621 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9641 0 4567 4622 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9642 4622 4582 627 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9643 617 4571 4622 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9644 4622 4580 601 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9645 612 4563 4622 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9646 0 4624 4623 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m9647 4625 4626 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m9648 0 4242 4625 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m9649 4627 4626 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m9650 4624 4242 4627 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m9651 4625 4248 4624 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m9652 4628 4248 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9653 4629 4624 4628 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9654 4630 4242 4629 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m9655 4631 4248 4630 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m9656 0 4626 4631 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m9657 4628 4242 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9658 0 4626 4628 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9659 1 4624 4623 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m9660 4632 4626 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m9661 4633 4242 4632 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m9662 4624 4626 4633 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9663 4633 4242 4624 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9664 4634 4629 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m9665 1 4248 4633 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9666 4629 4624 4635 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9667 4636 4242 4629 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9668 4637 4248 4636 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9669 4635 4626 4637 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9670 1 4242 4635 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9671 4635 4626 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9672 1 4248 4635 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9673 4626 4638 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9674 4638 4639 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9675 4634 4629 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m9676 0 4638 4626 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9677 0 4639 4638 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9678 0 4567 4639 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9679 4639 4582 642 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9680 632 4571 4639 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9681 4639 4580 617 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9682 627 4563 4639 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9683 0 4641 4640 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m9684 4642 4643 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m9685 0 4259 4642 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m9686 4644 4643 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m9687 4641 4259 4644 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m9688 4642 4265 4641 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m9689 4645 4265 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9690 4646 4641 4645 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9691 4647 4259 4646 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m9692 4648 4265 4647 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m9693 0 4643 4648 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m9694 4645 4259 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9695 0 4643 4645 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9696 1 4641 4640 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m9697 4649 4643 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m9698 4650 4259 4649 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m9699 4641 4643 4650 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9700 4650 4259 4641 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9701 4651 4646 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m9702 1 4265 4650 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9703 4646 4641 4652 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9704 4653 4259 4646 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9705 4654 4265 4653 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9706 4652 4643 4654 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9707 1 4259 4652 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9708 4652 4643 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9709 1 4265 4652 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9710 4643 4655 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9711 4655 4656 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9712 4651 4646 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m9713 0 4655 4643 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9714 0 4656 4655 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9715 0 4567 4656 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9716 4656 4582 657 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9717 647 4571 4656 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9718 4656 4580 632 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9719 642 4563 4656 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9720 0 4658 4657 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m9721 4659 4660 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m9722 0 4276 4659 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m9723 4661 4660 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m9724 4658 4276 4661 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m9725 4659 4282 4658 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m9726 4662 4282 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9727 4663 4658 4662 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9728 4664 4276 4663 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m9729 4665 4282 4664 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m9730 0 4660 4665 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m9731 4662 4276 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9732 0 4660 4662 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9733 1 4658 4657 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m9734 4666 4660 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m9735 4667 4276 4666 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m9736 4658 4660 4667 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9737 4667 4276 4658 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9738 4668 4663 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m9739 1 4282 4667 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9740 4663 4658 4669 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9741 4670 4276 4663 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9742 4671 4282 4670 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9743 4669 4660 4671 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9744 1 4276 4669 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9745 4669 4660 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9746 1 4282 4669 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9747 4660 4672 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9748 4672 4673 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9749 4668 4663 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m9750 0 4672 4660 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9751 0 4673 4672 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9752 0 4567 4673 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9753 4673 4582 672 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9754 662 4571 4673 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9755 4673 4580 647 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9756 657 4563 4673 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9757 0 4675 4674 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m9758 4676 4677 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m9759 0 4293 4676 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m9760 4678 4677 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m9761 4675 4293 4678 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m9762 4676 4299 4675 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m9763 4679 4299 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9764 4680 4675 4679 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9765 4681 4293 4680 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m9766 4682 4299 4681 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m9767 0 4677 4682 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m9768 4679 4293 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9769 0 4677 4679 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9770 1 4675 4674 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m9771 4683 4677 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m9772 4684 4293 4683 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m9773 4675 4677 4684 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9774 4684 4293 4675 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9775 4685 4680 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m9776 1 4299 4684 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9777 4680 4675 4686 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9778 4687 4293 4680 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9779 4688 4299 4687 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9780 4686 4677 4688 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9781 1 4293 4686 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9782 4686 4677 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9783 1 4299 4686 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9784 4677 4689 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9785 4689 4690 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9786 4685 4680 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m9787 0 4689 4677 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9788 0 4690 4689 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9789 0 4567 4690 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9790 4690 4582 687 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9791 677 4571 4690 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9792 4690 4580 662 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9793 672 4563 4690 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9794 0 4692 4691 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m9795 4693 4694 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m9796 0 4310 4693 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m9797 4695 4694 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m9798 4692 4310 4695 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m9799 4693 4316 4692 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m9800 4696 4316 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9801 4697 4692 4696 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9802 4698 4310 4697 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m9803 4699 4316 4698 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m9804 0 4694 4699 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m9805 4696 4310 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9806 0 4694 4696 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9807 1 4692 4691 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m9808 4700 4694 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m9809 4701 4310 4700 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m9810 4692 4694 4701 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9811 4701 4310 4692 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9812 4702 4697 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m9813 1 4316 4701 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9814 4697 4692 4703 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9815 4704 4310 4697 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9816 4705 4316 4704 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9817 4703 4694 4705 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9818 1 4310 4703 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9819 4703 4694 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9820 1 4316 4703 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9821 4694 4706 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9822 4706 4707 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9823 4702 4697 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m9824 0 4706 4694 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9825 0 4707 4706 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9826 0 4567 4707 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9827 4707 4582 702 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9828 692 4571 4707 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9829 4707 4580 677 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9830 687 4563 4707 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9831 0 4709 4708 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m9832 4710 4711 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m9833 0 4327 4710 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m9834 4712 4711 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m9835 4709 4327 4712 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m9836 4710 4333 4709 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m9837 4713 4333 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9838 4714 4709 4713 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9839 4715 4327 4714 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m9840 4716 4333 4715 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m9841 0 4711 4716 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m9842 4713 4327 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9843 0 4711 4713 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9844 1 4709 4708 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m9845 4717 4711 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m9846 4718 4327 4717 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m9847 4709 4711 4718 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9848 4718 4327 4709 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9849 4719 4714 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m9850 1 4333 4718 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9851 4714 4709 4720 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9852 4721 4327 4714 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9853 4722 4333 4721 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9854 4720 4711 4722 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9855 1 4327 4720 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9856 4720 4711 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9857 1 4333 4720 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9858 4711 4723 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9859 4723 4724 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9860 4719 4714 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m9861 0 4723 4711 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9862 0 4724 4723 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9863 0 4567 4724 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9864 4724 4582 717 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9865 707 4571 4724 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9866 4724 4580 692 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9867 702 4563 4724 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9868 0 4726 4725 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m9869 4727 4728 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m9870 0 4344 4727 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m9871 4729 4728 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m9872 4726 4344 4729 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m9873 4727 4350 4726 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m9874 4730 4350 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9875 4731 4726 4730 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9876 4732 4344 4731 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m9877 4733 4350 4732 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m9878 0 4728 4733 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m9879 4730 4344 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9880 0 4728 4730 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9881 1 4726 4725 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m9882 4734 4728 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m9883 4735 4344 4734 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m9884 4726 4728 4735 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9885 4735 4344 4726 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9886 4736 4731 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m9887 1 4350 4735 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9888 4731 4726 4737 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9889 4738 4344 4731 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9890 4739 4350 4738 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9891 4737 4728 4739 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9892 1 4344 4737 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9893 4737 4728 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9894 1 4350 4737 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9895 4728 4740 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9896 4740 4741 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9897 4736 4731 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m9898 0 4740 4728 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9899 0 4741 4740 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9900 0 4567 4741 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9901 4741 4582 732 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9902 722 4571 4741 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9903 4741 4580 707 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9904 717 4563 4741 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9905 0 4743 4742 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m9906 4744 4745 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m9907 0 4361 4744 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m9908 4746 4745 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m9909 4743 4361 4746 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m9910 4744 4367 4743 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m9911 4747 4367 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9912 4748 4743 4747 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9913 4749 4361 4748 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m9914 4750 4367 4749 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m9915 0 4745 4750 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m9916 4747 4361 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9917 0 4745 4747 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9918 1 4743 4742 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m9919 4751 4745 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m9920 4752 4361 4751 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m9921 4743 4745 4752 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9922 4752 4361 4743 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9923 4753 4748 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m9924 1 4367 4752 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9925 4748 4743 4754 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9926 4755 4361 4748 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9927 4756 4367 4755 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9928 4754 4745 4756 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9929 1 4361 4754 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9930 4754 4745 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9931 1 4367 4754 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9932 4745 4757 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9933 4757 4758 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9934 4753 4748 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m9935 0 4757 4745 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9936 0 4758 4757 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9937 0 4567 4758 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9938 4758 4582 747 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9939 737 4571 4758 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9940 4758 4580 722 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9941 732 4563 4758 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9942 0 4760 4759 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m9943 4761 4762 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m9944 0 4378 4761 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m9945 4763 4762 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m9946 4760 4378 4763 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m9947 4761 4384 4760 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m9948 4764 4384 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9949 4765 4760 4764 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9950 4766 4378 4765 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m9951 4767 4384 4766 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m9952 0 4762 4767 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m9953 4764 4378 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9954 0 4762 4764 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9955 1 4760 4759 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m9956 4768 4762 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m9957 4769 4378 4768 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m9958 4760 4762 4769 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9959 4769 4378 4760 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9960 4770 4765 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m9961 1 4384 4769 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9962 4765 4760 4771 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m9963 4772 4378 4765 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m9964 4773 4384 4772 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m9965 4771 4762 4773 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m9966 1 4378 4771 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m9967 4771 4762 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m9968 1 4384 4771 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m9969 4762 4774 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m9970 4774 4775 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m9971 4770 4765 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m9972 0 4774 4762 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m9973 0 4775 4774 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m9974 0 4567 4775 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m9975 4775 4582 762 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m9976 752 4571 4775 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m9977 4775 4580 737 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m9978 747 4563 4775 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m9979 0 4777 4776 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m9980 4778 4779 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m9981 0 4395 4778 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m9982 4780 4779 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m9983 4777 4395 4780 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m9984 4778 4401 4777 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m9985 4781 4401 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m9986 4782 4777 4781 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m9987 4783 4395 4782 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m9988 4784 4401 4783 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m9989 0 4779 4784 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m9990 4781 4395 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m9991 0 4779 4781 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m9992 1 4777 4776 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m9993 4785 4779 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m9994 4786 4395 4785 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m9995 4777 4779 4786 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m9996 4786 4395 4777 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m9997 4787 4782 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m9998 1 4401 4786 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m9999 4782 4777 4788 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m10000 4789 4395 4782 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m10001 4790 4401 4789 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m10002 4788 4779 4790 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m10003 1 4395 4788 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m10004 4788 4779 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m10005 1 4401 4788 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m10006 4779 4791 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m10007 4791 4792 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10008 4787 4782 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m10009 0 4791 4779 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m10010 0 4792 4791 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m10011 0 4567 4792 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m10012 4792 4582 777 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m10013 767 4571 4792 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m10014 4792 4580 752 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m10015 762 4563 4792 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m10016 0 4794 4793 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m10017 4795 4796 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m10018 0 4412 4795 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m10019 4797 4796 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m10020 4794 4412 4797 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m10021 4795 4418 4794 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m10022 4798 4418 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m10023 4799 4794 4798 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m10024 4800 4412 4799 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m10025 4801 4418 4800 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m10026 0 4796 4801 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m10027 4798 4412 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m10028 0 4796 4798 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m10029 1 4794 4793 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m10030 4802 4796 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m10031 4803 4412 4802 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m10032 4794 4796 4803 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m10033 4803 4412 4794 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m10034 4804 4799 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m10035 1 4418 4803 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m10036 4799 4794 4805 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m10037 4806 4412 4799 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m10038 4807 4418 4806 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m10039 4805 4796 4807 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m10040 1 4412 4805 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m10041 4805 4796 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m10042 1 4418 4805 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m10043 4796 4808 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m10044 4808 4809 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10045 4804 4799 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m10046 0 4808 4796 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m10047 0 4809 4808 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m10048 0 4567 4809 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m10049 4809 4582 792 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m10050 782 4571 4809 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m10051 4809 4580 767 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m10052 777 4563 4809 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m10053 0 4811 4810 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m10054 4812 4813 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m10055 0 4429 4812 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m10056 4814 4813 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m10057 4811 4429 4814 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m10058 4812 4435 4811 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m10059 4815 4435 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m10060 4816 4811 4815 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m10061 4817 4429 4816 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m10062 4818 4435 4817 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m10063 0 4813 4818 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m10064 4815 4429 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m10065 0 4813 4815 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m10066 1 4811 4810 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m10067 4819 4813 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m10068 4820 4429 4819 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m10069 4811 4813 4820 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m10070 4820 4429 4811 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m10071 4821 4816 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m10072 1 4435 4820 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m10073 4816 4811 4822 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m10074 4823 4429 4816 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m10075 4824 4435 4823 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m10076 4822 4813 4824 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m10077 1 4429 4822 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m10078 4822 4813 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m10079 1 4435 4822 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m10080 4813 4825 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m10081 4825 4826 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10082 4821 4816 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m10083 0 4825 4813 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m10084 0 4826 4825 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m10085 0 4567 4826 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m10086 4826 4582 807 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m10087 797 4571 4826 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m10088 4826 4580 782 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m10089 792 4563 4826 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m10090 0 4828 4827 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m10091 4829 4830 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m10092 0 4446 4829 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m10093 4831 4830 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m10094 4828 4446 4831 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m10095 4829 4452 4828 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m10096 4832 4452 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m10097 4833 4828 4832 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m10098 4834 4446 4833 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m10099 4835 4452 4834 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m10100 0 4830 4835 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m10101 4832 4446 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m10102 0 4830 4832 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m10103 1 4828 4827 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m10104 4836 4830 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m10105 4837 4446 4836 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m10106 4828 4830 4837 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m10107 4837 4446 4828 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m10108 4838 4833 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m10109 1 4452 4837 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m10110 4833 4828 4839 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m10111 4840 4446 4833 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m10112 4841 4452 4840 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m10113 4839 4830 4841 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m10114 1 4446 4839 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m10115 4839 4830 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m10116 1 4452 4839 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m10117 4830 4842 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m10118 4842 4843 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10119 4838 4833 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m10120 0 4842 4830 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m10121 0 4843 4842 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m10122 0 4567 4843 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m10123 4843 4582 822 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m10124 812 4571 4843 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m10125 4843 4580 797 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m10126 807 4563 4843 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m10127 0 4845 4844 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m10128 4846 4847 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m10129 0 4463 4846 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m10130 4848 4847 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m10131 4845 4463 4848 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m10132 4846 4469 4845 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m10133 4849 4469 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m10134 4850 4845 4849 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m10135 4851 4463 4850 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m10136 4852 4469 4851 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m10137 0 4847 4852 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m10138 4849 4463 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m10139 0 4847 4849 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m10140 1 4845 4844 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m10141 4853 4847 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m10142 4854 4463 4853 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m10143 4845 4847 4854 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m10144 4854 4463 4845 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m10145 4855 4850 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m10146 1 4469 4854 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m10147 4850 4845 4856 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m10148 4857 4463 4850 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m10149 4858 4469 4857 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m10150 4856 4847 4858 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m10151 1 4463 4856 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m10152 4856 4847 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m10153 1 4469 4856 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m10154 4847 4859 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m10155 4859 4860 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10156 4855 4850 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m10157 0 4859 4847 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m10158 0 4860 4859 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m10159 0 4567 4860 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m10160 4860 4582 837 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m10161 827 4571 4860 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m10162 4860 4580 812 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m10163 822 4563 4860 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m10164 0 4862 4861 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=2.92e-11 ps=2.699e-05 pd=3.17e-05 
+ nrs=0.14 nrd=0.14 
m10165 4863 4864 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.04e-11 ad=3.013e-11 ps=2.215e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m10166 0 4480 4863 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.04e-11 ps=2.849e-05 pd=2.215e-05 
+ nrs=0.13 nrd=0.09 
m10167 4865 4864 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m10168 4862 4480 4865 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m10169 4863 4486 4862 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.879e-11 ad=1.383e-11 ps=2.04e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m10170 4866 4486 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m10171 4867 4862 4866 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m10172 4868 4480 4867 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m10173 4869 4486 4868 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m10174 0 4864 4869 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m10175 4866 4480 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m10176 0 4864 4866 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m10177 1 4862 4861 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m10178 4870 4864 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m10179 4871 4480 4870 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m10180 4862 4864 4871 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m10181 4871 4480 4862 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m10182 4872 4867 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m10183 1 4486 4871 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m10184 4867 4862 4873 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m10185 4874 4480 4867 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m10186 4875 4486 4874 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m10187 4873 4864 4875 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m10188 1 4480 4873 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m10189 4873 4864 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m10190 1 4486 4873 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m10191 4864 4876 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m10192 4876 4877 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10193 4872 4867 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m10194 0 4876 4864 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m10195 0 4877 4876 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.686e-11 ps=1.125e-05 pd=1.89e-05 
+ nrs=0.33 nrd=0.47 
m10196 0 4567 4877 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m10197 4877 4582 868 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m10198 842 4571 4877 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.048e-11 ad=6.95e-12 ps=1.23e-05 pd=8.18e-06 
+ nrs=0.81 nrd=0.54 
m10199 4877 4580 827 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m10200 837 4563 4877 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m10201 0 4879 4878 0 nenh l=1.1e-06 w=1.48e-05 
+ as=2.933e-11 ad=3.042e-11 ps=2.774e-05 pd=3.25e-05 
+ nrs=0.13 nrd=0.14 
m10202 4880 4881 0 0 nenh l=1.1e-06 w=1.56e-05 
+ as=2.08e-11 ad=3.092e-11 ps=2.261e-05 pd=2.924e-05 
+ nrs=0.09 nrd=0.13 
m10203 0 4497 4880 0 nenh l=1.1e-06 w=1.56e-05 
+ as=3.092e-11 ad=2.08e-11 ps=2.924e-05 pd=2.261e-05 
+ nrs=0.13 nrd=0.09 
m10204 4882 4881 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m10205 4879 4497 4882 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m10206 4880 4503 4879 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.866e-11 ad=1.383e-11 ps=2.029e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m10207 4883 4503 0 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.404e-11 ad=2.933e-11 ps=1.652e-05 pd=2.774e-05 
+ nrs=0.06 nrd=0.13 
m10208 4884 4879 4883 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.497e-11 ad=1.404e-11 ps=1.835e-05 pd=1.652e-05 
+ nrs=0.07 nrd=0.06 
m10209 4885 4497 4884 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.236e-11 ad=1.457e-11 ps=1.661e-05 pd=1.785e-05 
+ nrs=0.06 nrd=0.07 
m10210 4886 4503 4885 0 nenh l=1.1e-06 w=1.56e-05 
+ as=1.338e-11 ad=1.338e-11 ps=1.781e-05 pd=1.799e-05 
+ nrs=0.05 nrd=0.05 
m10211 0 4881 4886 0 nenh l=1.1e-06 w=1.68e-05 
+ as=3.33e-11 ad=1.44e-11 ps=3.149e-05 pd=1.919e-05 
+ nrs=0.12 nrd=0.05 
m10212 4883 4497 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.518e-11 ad=3.171e-11 ps=1.786e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m10213 0 4881 4883 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.214e-11 ps=2.399e-05 pd=1.429e-05 
+ nrs=0.15 nrd=0.07 
m10214 1 4879 4878 1 penh l=1.1e-06 w=1.76e-05 
+ as=3.919e-11 ad=3.16e-11 ps=3.323e-05 pd=3.89e-05 
+ nrs=0.13 nrd=0.1 
m10215 4887 4881 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m10216 4888 4497 4887 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m10217 4879 4881 4888 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.814e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m10218 4888 4497 4879 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.684e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.07 
m10219 4889 4884 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m10220 1 4503 4888 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m10221 4884 4879 4890 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.395e-11 ad=1.488e-11 ps=1.731e-05 pd=1.779e-05 
+ nrs=0.1 nrd=0.1 
m10222 4891 4497 4884 1 penh l=1.1e-06 w=1.92e-05 
+ as=1.655e-11 ad=2.233e-11 ps=2.193e-05 pd=2.769e-05 
+ nrs=0.04 nrd=0.06 
m10223 4892 4503 4891 1 penh l=1.1e-06 w=2.16e-05 
+ as=1.848e-11 ad=1.861e-11 ps=2.384e-05 pd=2.467e-05 
+ nrs=0.04 nrd=0.04 
m10224 4890 4881 4892 1 penh l=1.1e-06 w=2.28e-05 
+ as=2.828e-11 ad=1.95e-11 ps=3.38e-05 pd=2.516e-05 
+ nrs=0.05 nrd=0.04 
m10225 1 4497 4890 1 penh l=1.1e-06 w=1.36e-05 
+ as=3.028e-11 ad=1.687e-11 ps=2.567e-05 pd=2.016e-05 
+ nrs=0.16 nrd=0.09 
m10226 4890 4881 1 1 penh l=1.1e-06 w=1.36e-05 
+ as=1.687e-11 ad=3.028e-11 ps=2.016e-05 pd=2.567e-05 
+ nrs=0.09 nrd=0.16 
m10227 1 4503 4890 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.488e-11 ps=2.265e-05 pd=1.779e-05 
+ nrs=0.19 nrd=0.1 
m10228 4881 4893 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=2.172e-11 ad=1.959e-11 ps=2.37e-05 pd=1.661e-05 
+ nrs=0.28 nrd=0.25 
m10229 4893 4894 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10230 4889 4884 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m10231 0 4893 4881 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.856e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.45 
m10232 0 4894 4893 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.446e-11 ps=1.125e-05 pd=1.81e-05 
+ nrs=0.33 nrd=0.4 
m10233 0 4567 4894 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.95e-12 ps=6.75e-06 pd=8.18e-06 
+ nrs=0.55 nrd=0.54 
m10234 4894 4582 852 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.003e-11 ps=8.18e-06 pd=1.202e-05 
+ nrs=0.54 nrd=0.77 
m10235 858 4571 4894 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.036e-11 ad=6.95e-12 ps=1.246e-05 pd=8.18e-06 
+ nrs=0.8 nrd=0.54 
m10236 4894 4580 842 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.95e-12 ad=1.048e-11 ps=8.18e-06 pd=1.23e-05 
+ nrs=0.54 nrd=0.81 
m10237 868 4563 4894 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.95e-12 ps=1.202e-05 pd=8.18e-06 
+ nrs=0.77 nrd=0.54 
m10238 4895 4896 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=5.99e-12 ad=1.348e-11 ps=9.58e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m10239 64 4897 4895 0 nenh l=1.1e-06 w=6.4e-06 
+ as=7.52e-12 ad=5.63e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.14 
m10240 4898 4899 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10241 4897 4900 4898 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10242 4901 4902 4897 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10243 0 4903 4901 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10244 4899 4903 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10245 0 4905 4904 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m10246 4906 4900 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10247 4907 4904 4906 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10248 4908 4905 4907 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10249 0 4902 4908 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10250 4900 4902 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10251 4909 4907 64 0 nenh l=1.1e-06 w=6.4e-06 
+ as=5.63e-12 ad=7.52e-12 ps=9.02e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10252 0 4910 4909 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.99e-12 ps=1.275e-05 pd=9.58e-06 
+ nrs=0.29 nrd=0.13 
m10253 4911 4896 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m10254 64 4907 4911 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m10255 4912 4897 64 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10256 1 4910 4912 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m10257 4913 4899 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10258 4897 4902 4913 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m10259 4914 4900 4897 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m10260 1 4903 4914 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m10261 4899 4903 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10262 4915 4903 4916 0 nenh l=1.1e-06 w=8.8e-06 
+ as=9.42e-12 ad=1.37e-11 ps=1.155e-05 pd=1.663e-05 
+ nrs=0.12 nrd=0.18 
m10263 4917 4918 4915 0 nenh l=1.1e-06 w=7.2e-06 
+ as=6.12e-12 ad=7.7e-12 ps=8.9e-06 pd=9.45e-06 
+ nrs=0.12 nrd=0.15 
m10264 4916 4919 4917 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.121e-11 ad=6.12e-12 ps=1.361e-05 pd=8.9e-06 
+ nrs=0.22 nrd=0.12 
m10265 0 4919 4916 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.744e-11 ad=1.37e-11 ps=1.65e-05 pd=1.663e-05 
+ nrs=0.23 nrd=0.18 
m10266 4916 4918 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.246e-11 ad=1.586e-11 ps=1.512e-05 pd=1.5e-05 
+ nrs=0.19 nrd=0.25 
m10267 0 4918 4920 0 nenh l=1.1e-06 w=8e-06 
+ as=1.586e-11 ad=1.246e-11 ps=1.5e-05 pd=1.512e-05 
+ nrs=0.25 nrd=0.19 
m10268 4920 4919 0 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.37e-11 ad=1.744e-11 ps=1.663e-05 pd=1.65e-05 
+ nrs=0.18 nrd=0.23 
m10269 4921 4919 4920 0 nenh l=1.1e-06 w=7.2e-06 
+ as=6.12e-12 ad=1.121e-11 ps=8.9e-06 pd=1.361e-05 
+ nrs=0.12 nrd=0.22 
m10270 4922 4918 4921 0 nenh l=1.1e-06 w=7.2e-06 
+ as=7.7e-12 ad=6.12e-12 ps=9.45e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.12 
m10271 0 4923 4919 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m10272 4924 4919 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10273 4902 4918 4924 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10274 4925 4889 4902 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10275 0 4923 4925 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10276 4918 4889 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10277 4920 4905 4922 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.37e-11 ad=9.42e-12 ps=1.663e-05 pd=1.155e-05 
+ nrs=0.18 nrd=0.12 
m10278 1 4905 4904 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m10279 4926 4900 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m10280 4907 4905 4926 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m10281 4927 4904 4907 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m10282 1 4902 4927 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m10283 4900 4902 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m10284 4915 4903 4928 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.039e-11 ad=1.116e-11 ps=1.197e-05 pd=1.42e-05 
+ nrs=0.13 nrd=0.14 
m10285 4929 4918 4915 1 penh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=9.91e-12 ps=1.01e-05 pd=1.143e-05 
+ nrs=0.1 nrd=0.14 
m10286 1 4919 4929 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=7.14e-12 ps=1.586e-05 pd=1.01e-05 
+ nrs=0.27 nrd=0.1 
m10287 4928 4919 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.166e-11 ad=2.048e-11 ps=1.485e-05 pd=1.737e-05 
+ nrs=0.14 nrd=0.24 
m10288 1 4918 4928 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.166e-11 ps=1.737e-05 pd=1.485e-05 
+ nrs=0.24 nrd=0.14 
m10289 4930 4918 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.166e-11 ad=2.048e-11 ps=1.485e-05 pd=1.737e-05 
+ nrs=0.14 nrd=0.24 
m10290 1 4919 4930 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.166e-11 ps=1.737e-05 pd=1.485e-05 
+ nrs=0.24 nrd=0.14 
m10291 4931 4919 1 1 penh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=1.87e-11 ps=1.01e-05 pd=1.586e-05 
+ nrs=0.1 nrd=0.27 
m10292 4922 4918 4931 1 penh l=1.1e-06 w=8.4e-06 
+ as=9.91e-12 ad=7.14e-12 ps=1.143e-05 pd=1.01e-05 
+ nrs=0.14 nrd=0.1 
m10293 4930 4905 4922 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.116e-11 ad=1.039e-11 ps=1.42e-05 pd=1.197e-05 
+ nrs=0.14 nrd=0.13 
m10294 1 4923 4919 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m10295 4932 4919 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=4.53e-12 ad=1.158e-11 ps=7.26e-06 pd=9.82e-06 
+ nrs=0.17 nrd=0.43 
m10296 4902 4889 4932 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.32e-12 ad=5.57e-12 ps=9.07e-06 pd=8.94e-06 
+ nrs=0.18 nrd=0.14 
m10297 4933 4918 4902 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.8e-12 ad=6.4e-12 ps=7.57e-06 pd=7.93e-06 
+ nrs=0.15 nrd=0.2 
m10298 1 4923 4933 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=4.46e-12 ps=9.82e-06 pd=7.03e-06 
+ nrs=0.43 nrd=0.16 
m10299 4918 4889 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10300 1 4934 33 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m10301 4935 4896 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m10302 4934 4936 4935 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m10303 4937 4938 4934 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10304 1 4910 4937 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m10305 4939 4940 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10306 4938 4941 4939 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m10307 4942 4943 4938 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m10308 1 4944 4942 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m10309 4940 4944 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10310 1 4946 4945 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m10311 4947 4943 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m10312 4936 4946 4947 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m10313 4948 4945 4936 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m10314 1 4941 4948 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m10315 4943 4941 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m10316 1 4950 4949 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m10317 4951 4952 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m10318 4941 4950 4951 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m10319 4953 4949 4941 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m10320 1 4954 4953 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m10321 4952 4954 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m10322 0 4934 33 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m10323 4955 4896 0 0 nenh l=1.1e-06 w=7.2e-06 
+ as=6.43e-12 ad=1.427e-11 ps=1.058e-05 pd=1.35e-05 
+ nrs=0.12 nrd=0.28 
m10324 4934 4938 4955 0 nenh l=1.1e-06 w=6e-06 
+ as=8.27e-12 ad=5.35e-12 ps=9.11e-06 pd=8.82e-06 
+ nrs=0.23 nrd=0.15 
m10325 4956 4936 4934 0 nenh l=1.1e-06 w=5.2e-06 
+ as=4.53e-12 ad=7.17e-12 ps=7.26e-06 pd=7.89e-06 
+ nrs=0.17 nrd=0.27 
m10326 0 4910 4956 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=5.57e-12 ps=1.2e-05 pd=8.94e-06 
+ nrs=0.31 nrd=0.14 
m10327 4957 4944 1 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.023e-11 ad=1.959e-11 ps=1.157e-05 pd=1.661e-05 
+ nrs=0.13 nrd=0.25 
m10328 4903 4950 4957 1 penh l=1.1e-06 w=8.4e-06 
+ as=8.75e-12 ad=9.76e-12 ps=1.068e-05 pd=1.104e-05 
+ nrs=0.12 nrd=0.14 
m10329 4957 4954 4903 1 penh l=1.1e-06 w=1e-05 
+ as=1.162e-11 ad=1.041e-11 ps=1.315e-05 pd=1.272e-05 
+ nrs=0.12 nrd=0.1 
m10330 4958 4954 4957 1 penh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=9.76e-12 ps=1.01e-05 pd=1.104e-05 
+ nrs=0.1 nrd=0.14 
m10331 1 4950 4958 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=7.14e-12 ps=1.586e-05 pd=1.01e-05 
+ nrs=0.27 nrd=0.1 
m10332 4959 4950 1 1 penh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=1.87e-11 ps=1.01e-05 pd=1.586e-05 
+ nrs=0.1 nrd=0.27 
m10333 4960 4954 4959 1 penh l=1.1e-06 w=8.4e-06 
+ as=9.76e-12 ad=7.14e-12 ps=1.104e-05 pd=1.01e-05 
+ nrs=0.14 nrd=0.1 
m10334 4905 4954 4960 1 penh l=1.1e-06 w=1e-05 
+ as=1.041e-11 ad=1.162e-11 ps=1.272e-05 pd=1.315e-05 
+ nrs=0.1 nrd=0.12 
m10335 4960 4950 4905 1 penh l=1.1e-06 w=8.4e-06 
+ as=9.76e-12 ad=8.75e-12 ps=1.104e-05 pd=1.068e-05 
+ nrs=0.14 nrd=0.12 
m10336 1 4946 4960 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=1.023e-11 ps=1.661e-05 pd=1.157e-05 
+ nrs=0.25 nrd=0.13 
m10337 4961 4940 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10338 4938 4943 4961 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10339 4962 4941 4938 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10340 0 4944 4962 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10341 4940 4944 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10342 0 4946 4945 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m10343 4963 4943 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10344 4936 4945 4963 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10345 4964 4946 4936 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10346 0 4941 4964 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10347 4943 4941 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10348 0 4950 4949 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m10349 4965 4952 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10350 4941 4949 4965 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10351 4966 4950 4941 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10352 0 4954 4966 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10353 4952 4954 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10354 4903 4944 4967 0 nenh l=1.1e-06 w=8.8e-06 
+ as=9.42e-12 ad=1.151e-11 ps=1.155e-05 pd=1.473e-05 
+ nrs=0.12 nrd=0.15 
m10355 4968 4950 4903 0 nenh l=1.1e-06 w=7.2e-06 
+ as=6.12e-12 ad=7.7e-12 ps=8.9e-06 pd=9.45e-06 
+ nrs=0.12 nrd=0.15 
m10356 0 4954 4968 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.427e-11 ad=6.12e-12 ps=1.35e-05 pd=8.9e-06 
+ nrs=0.28 nrd=0.12 
m10357 4967 4954 0 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.151e-11 ad=1.744e-11 ps=1.473e-05 pd=1.65e-05 
+ nrs=0.15 nrd=0.23 
m10358 0 4950 4967 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.427e-11 ad=9.42e-12 ps=1.35e-05 pd=1.205e-05 
+ nrs=0.28 nrd=0.18 
m10359 4969 4950 0 0 nenh l=1.1e-06 w=7.2e-06 
+ as=9.42e-12 ad=1.427e-11 ps=1.205e-05 pd=1.35e-05 
+ nrs=0.18 nrd=0.28 
m10360 0 4954 4969 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.744e-11 ad=1.151e-11 ps=1.65e-05 pd=1.473e-05 
+ nrs=0.23 nrd=0.15 
m10361 4970 4954 0 0 nenh l=1.1e-06 w=7.2e-06 
+ as=6.12e-12 ad=1.427e-11 ps=8.9e-06 pd=1.35e-05 
+ nrs=0.12 nrd=0.28 
m10362 4905 4950 4970 0 nenh l=1.1e-06 w=7.2e-06 
+ as=7.7e-12 ad=6.12e-12 ps=9.45e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.12 
m10363 4969 4946 4905 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.151e-11 ad=9.42e-12 ps=1.473e-05 pd=1.155e-05 
+ nrs=0.15 nrd=0.12 
m10364 4971 4896 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.04e-12 ad=1.348e-11 ps=9.88e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m10365 526 4972 4971 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=5.33e-12 ps=8.5e-06 pd=8.72e-06 
+ nrs=0.19 nrd=0.15 
m10366 4973 4974 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10367 4972 4975 4973 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10368 4976 4977 4972 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10369 0 4978 4976 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10370 4974 4978 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10371 0 4980 4979 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m10372 4981 4975 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10373 4982 4979 4981 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10374 4983 4980 4982 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10375 0 4977 4983 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10376 4975 4977 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10377 4984 4982 526 0 nenh l=1.1e-06 w=6e-06 
+ as=5.29e-12 ad=6.86e-12 ps=8.61e-06 pd=8.5e-06 
+ nrs=0.15 nrd=0.19 
m10378 0 4910 4984 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=5.65e-12 ps=1.2e-05 pd=9.19e-06 
+ nrs=0.31 nrd=0.14 
m10379 4985 4896 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m10380 526 4982 4985 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m10381 4986 4972 526 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10382 1 4910 4986 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m10383 4987 4974 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10384 4972 4977 4987 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m10385 4988 4975 4972 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m10386 1 4978 4988 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m10387 4974 4978 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.308e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.42 nrd=0.4 
m10388 4944 4978 4989 0 nenh l=1.1e-06 w=8.8e-06 
+ as=9.42e-12 ad=1.37e-11 ps=1.155e-05 pd=1.663e-05 
+ nrs=0.12 nrd=0.18 
m10389 4990 4991 4944 0 nenh l=1.1e-06 w=7.2e-06 
+ as=6.12e-12 ad=7.7e-12 ps=8.9e-06 pd=9.45e-06 
+ nrs=0.12 nrd=0.15 
m10390 4989 4992 4990 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.121e-11 ad=6.12e-12 ps=1.361e-05 pd=8.9e-06 
+ nrs=0.22 nrd=0.12 
m10391 0 4992 4989 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.744e-11 ad=1.37e-11 ps=1.65e-05 pd=1.663e-05 
+ nrs=0.23 nrd=0.18 
m10392 4989 4991 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.246e-11 ad=1.586e-11 ps=1.512e-05 pd=1.5e-05 
+ nrs=0.19 nrd=0.25 
m10393 0 4991 4993 0 nenh l=1.1e-06 w=8e-06 
+ as=1.586e-11 ad=1.246e-11 ps=1.5e-05 pd=1.512e-05 
+ nrs=0.25 nrd=0.19 
m10394 4993 4992 0 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.37e-11 ad=1.744e-11 ps=1.663e-05 pd=1.65e-05 
+ nrs=0.18 nrd=0.23 
m10395 4994 4992 4993 0 nenh l=1.1e-06 w=7.2e-06 
+ as=6.12e-12 ad=1.121e-11 ps=8.9e-06 pd=1.361e-05 
+ nrs=0.12 nrd=0.22 
m10396 4946 4991 4994 0 nenh l=1.1e-06 w=7.2e-06 
+ as=7.7e-12 ad=6.12e-12 ps=9.45e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.12 
m10397 0 4537 4992 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m10398 4995 4992 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10399 4977 4991 4995 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10400 4996 4531 4977 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10401 0 4537 4996 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10402 4991 4531 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10403 4993 4980 4946 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.37e-11 ad=9.42e-12 ps=1.663e-05 pd=1.155e-05 
+ nrs=0.18 nrd=0.12 
m10404 1 4980 4979 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m10405 4997 4975 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m10406 4982 4980 4997 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m10407 4998 4979 4982 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m10408 1 4977 4998 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m10409 4975 4977 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m10410 4944 4978 4999 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.039e-11 ad=1.116e-11 ps=1.197e-05 pd=1.42e-05 
+ nrs=0.13 nrd=0.14 
m10411 5000 4991 4944 1 penh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=9.91e-12 ps=1.01e-05 pd=1.143e-05 
+ nrs=0.1 nrd=0.14 
m10412 1 4992 5000 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=7.14e-12 ps=1.586e-05 pd=1.01e-05 
+ nrs=0.27 nrd=0.1 
m10413 4999 4992 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.166e-11 ad=2.048e-11 ps=1.485e-05 pd=1.737e-05 
+ nrs=0.14 nrd=0.24 
m10414 1 4991 4999 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.166e-11 ps=1.737e-05 pd=1.485e-05 
+ nrs=0.24 nrd=0.14 
m10415 5001 4991 1 1 penh l=1.1e-06 w=9.2e-06 
+ as=1.166e-11 ad=2.048e-11 ps=1.485e-05 pd=1.737e-05 
+ nrs=0.14 nrd=0.24 
m10416 1 4992 5001 1 penh l=1.1e-06 w=9.2e-06 
+ as=2.048e-11 ad=1.166e-11 ps=1.737e-05 pd=1.485e-05 
+ nrs=0.24 nrd=0.14 
m10417 5002 4992 1 1 penh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=1.87e-11 ps=1.01e-05 pd=1.586e-05 
+ nrs=0.1 nrd=0.27 
m10418 4946 4991 5002 1 penh l=1.1e-06 w=8.4e-06 
+ as=9.91e-12 ad=7.14e-12 ps=1.143e-05 pd=1.01e-05 
+ nrs=0.14 nrd=0.1 
m10419 5001 4980 4946 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.116e-11 ad=1.039e-11 ps=1.42e-05 pd=1.197e-05 
+ nrs=0.14 nrd=0.13 
m10420 1 4537 4992 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m10421 5003 4992 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=4.53e-12 ad=1.158e-11 ps=7.26e-06 pd=9.82e-06 
+ nrs=0.17 nrd=0.43 
m10422 4977 4531 5003 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.32e-12 ad=5.57e-12 ps=9.07e-06 pd=8.94e-06 
+ nrs=0.18 nrd=0.14 
m10423 5004 4991 4977 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.94e-12 ad=6.4e-12 ps=8.04e-06 pd=7.93e-06 
+ nrs=0.16 nrd=0.2 
m10424 1 4537 5004 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6e-12 ps=1.284e-05 pd=9.76e-06 
+ nrs=0.33 nrd=0.13 
m10425 4991 4531 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.298e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.48 nrd=0.43 
m10426 1 5005 497 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m10427 5006 4896 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m10428 5005 5007 5006 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m10429 5008 5009 5005 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10430 1 4910 5008 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m10431 4896 4910 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=7.88e-12 ad=1.603e-11 ps=9.7e-06 pd=1.359e-05 
+ nrs=0.15 nrd=0.31 
m10432 1 4910 4896 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=7.88e-12 ps=1.359e-05 pd=9.7e-06 
+ nrs=0.31 nrd=0.15 
m10433 1 5010 4910 1 penh l=1.1e-06 w=1.28e-05 
+ as=2.85e-11 ad=3.568e-11 ps=2.416e-05 pd=3.17e-05 
+ nrs=0.17 nrd=0.22 
m10434 1 5007 5009 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m10435 1 4546 5011 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m10436 5012 5013 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10437 5007 4546 5012 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m10438 5014 5011 5007 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m10439 1 4549 5014 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m10440 5013 4549 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10441 0 5005 497 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m10442 5015 4896 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=7.37e-12 ad=1.506e-11 ps=1.097e-05 pd=1.425e-05 
+ nrs=0.13 nrd=0.26 
m10443 5005 5009 5015 0 nenh l=1.1e-06 w=6.4e-06 
+ as=8.77e-12 ad=6.21e-12 ps=9.49e-06 pd=9.23e-06 
+ nrs=0.21 nrd=0.15 
m10444 5016 5007 5005 0 nenh l=1.1e-06 w=5.6e-06 
+ as=5.09e-12 ad=7.67e-12 ps=7.68e-06 pd=8.31e-06 
+ nrs=0.16 nrd=0.24 
m10445 0 4910 5016 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=6.17e-12 ps=1.275e-05 pd=9.32e-06 
+ nrs=0.29 nrd=0.13 
m10446 4896 4910 0 0 nenh l=1.1e-06 w=3.2e-06 
+ as=5.28e-12 ad=6.34e-12 ps=6.5e-06 pd=6e-06 
+ nrs=0.52 nrd=0.62 
m10447 0 4910 4896 0 nenh l=1.1e-06 w=3.2e-06 
+ as=6.34e-12 ad=5.28e-12 ps=6e-06 pd=6.5e-06 
+ nrs=0.62 nrd=0.52 
m10448 0 5010 4910 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.952e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.48 
m10449 0 5007 5009 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m10450 5017 4549 1 1 penh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=1.87e-11 ps=1.01e-05 pd=1.586e-05 
+ nrs=0.1 nrd=0.27 
m10451 4978 4546 5017 1 penh l=1.1e-06 w=8.4e-06 
+ as=2.466e-11 ad=7.14e-12 ps=2.29e-05 pd=1.01e-05 
+ nrs=0.35 nrd=0.1 
m10452 1 5018 5010 1 penh l=1.1e-06 w=9.6e-06 
+ as=2.137e-11 ad=2.928e-11 ps=1.812e-05 pd=2.53e-05 
+ nrs=0.23 nrd=0.32 
m10453 5018 3744 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=9.41e-12 ad=1.247e-11 ps=9.25e-06 pd=1.057e-05 
+ nrs=0.3 nrd=0.4 
m10454 5019 3839 5018 1 penh l=1.1e-06 w=7.6e-06 
+ as=6.46e-12 ad=1.277e-11 ps=9.3e-06 pd=1.255e-05 
+ nrs=0.11 nrd=0.22 
m10455 1 3751 5019 1 penh l=1.1e-06 w=7.6e-06 
+ as=1.692e-11 ad=6.46e-12 ps=1.435e-05 pd=9.3e-06 
+ nrs=0.29 nrd=0.11 
m10456 4980 4546 1 1 penh l=1.1e-06 w=8e-06 
+ as=8.56e-12 ad=1.781e-11 ps=1.05e-05 pd=1.51e-05 
+ nrs=0.13 nrd=0.28 
m10457 1 4549 4980 1 penh l=1.1e-06 w=8e-06 
+ as=1.781e-11 ad=8.56e-12 ps=1.51e-05 pd=1.05e-05 
+ nrs=0.28 nrd=0.13 
m10458 0 4546 5011 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m10459 5020 5013 0 0 nenh l=1.1e-06 w=7.2e-06 
+ as=7.02e-12 ad=1.427e-11 ps=1.001e-05 pd=1.35e-05 
+ nrs=0.14 nrd=0.28 
m10460 5007 5011 5020 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=5.46e-12 ps=8.9e-06 pd=7.79e-06 
+ nrs=0.29 nrd=0.17 
m10461 5021 4546 5007 0 nenh l=1.1e-06 w=5.6e-06 
+ as=5.18e-12 ad=9.24e-12 ps=7.79e-06 pd=8.9e-06 
+ nrs=0.17 nrd=0.29 
m10462 0 4549 5021 0 nenh l=1.1e-06 w=7.2e-06 
+ as=1.427e-11 ad=6.66e-12 ps=1.35e-05 pd=1.001e-05 
+ nrs=0.28 nrd=0.13 
m10463 5013 4549 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m10464 4978 4549 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=8.22e-12 ad=1.506e-11 ps=1.01e-05 pd=1.425e-05 
+ nrs=0.14 nrd=0.26 
m10465 0 4546 4978 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.506e-11 ad=8.22e-12 ps=1.425e-05 pd=1.01e-05 
+ nrs=0.26 nrd=0.14 
m10466 0 5018 5010 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.506e-11 ad=1.358e-11 ps=1.425e-05 pd=1.81e-05 
+ nrs=0.26 nrd=0.24 
m10467 5022 3744 0 0 nenh l=1.1e-06 w=6e-06 
+ as=1.204e-11 ad=1.189e-11 ps=1.197e-05 pd=1.125e-05 
+ nrs=0.33 nrd=0.33 
m10468 5018 3839 5022 0 nenh l=1.1e-06 w=6e-06 
+ as=9.94e-12 ad=1.204e-11 ps=9.39e-06 pd=1.197e-05 
+ nrs=0.28 nrd=0.33 
m10469 5022 3751 5018 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.284e-11 ad=1.06e-11 ps=1.277e-05 pd=1.001e-05 
+ nrs=0.31 nrd=0.26 
m10470 5023 4546 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=7.14e-12 ad=1.665e-11 ps=1.01e-05 pd=1.575e-05 
+ nrs=0.1 nrd=0.24 
m10471 4980 4549 5023 0 nenh l=1.1e-06 w=8.4e-06 
+ as=2.562e-11 ad=7.14e-12 ps=2.29e-05 pd=1.01e-05 
+ nrs=0.36 nrd=0.1 
m10472 5024 5025 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=5.99e-12 ad=1.348e-11 ps=9.58e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m10473 180 5026 5024 0 nenh l=1.1e-06 w=6.4e-06 
+ as=7.52e-12 ad=5.63e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.14 
m10474 5027 5028 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10475 5026 5029 5027 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10476 5030 5031 5026 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10477 0 5032 5030 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10478 5028 5032 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10479 0 5034 5033 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m10480 5035 5029 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10481 5036 5033 5035 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10482 5037 5034 5036 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10483 0 5031 5037 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10484 5029 5031 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10485 5038 5036 180 0 nenh l=1.1e-06 w=6.4e-06 
+ as=5.63e-12 ad=7.52e-12 ps=9.02e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10486 0 5039 5038 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.99e-12 ps=1.275e-05 pd=9.58e-06 
+ nrs=0.29 nrd=0.13 
m10487 5040 5025 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m10488 180 5036 5040 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m10489 5041 5026 180 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10490 1 5039 5041 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m10491 5042 5028 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10492 5026 5031 5042 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m10493 5043 5029 5026 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m10494 1 5032 5043 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m10495 5028 5032 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10496 5044 5032 5045 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.745e-11 ps=1.429e-05 pd=2.077e-05 
+ nrs=0.11 nrd=0.13 
m10497 5046 5047 5044 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m10498 5045 5048 5046 0 nenh l=1.1e-06 w=1e-05 
+ as=1.505e-11 ad=8.5e-12 ps=1.791e-05 pd=1.17e-05 
+ nrs=0.15 nrd=0.08 
m10499 0 5048 5045 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.745e-11 ps=2.174e-05 pd=2.077e-05 
+ nrs=0.17 nrd=0.13 
m10500 5045 5047 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=1.625e-11 ad=2.141e-11 ps=1.934e-05 pd=2.024e-05 
+ nrs=0.14 nrd=0.18 
m10501 0 5047 5049 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.625e-11 ps=2.024e-05 pd=1.934e-05 
+ nrs=0.18 nrd=0.14 
m10502 5049 5048 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.745e-11 ad=2.299e-11 ps=2.077e-05 pd=2.174e-05 
+ nrs=0.13 nrd=0.17 
m10503 5050 5048 5049 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.505e-11 ps=1.17e-05 pd=1.791e-05 
+ nrs=0.08 nrd=0.15 
m10504 5051 5047 5050 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m10505 5049 5034 5051 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.745e-11 ad=1.416e-11 ps=2.077e-05 pd=1.429e-05 
+ nrs=0.13 nrd=0.11 
m10506 0 4827 5048 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m10507 5052 5048 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m10508 5031 5047 5052 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m10509 5053 4821 5031 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m10510 0 4827 5053 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m10511 5047 4821 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m10512 1 5034 5033 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m10513 5054 5029 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m10514 5036 5034 5054 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m10515 5055 5033 5036 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m10516 1 5031 5055 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m10517 5029 5031 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m10518 5044 5032 5056 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m10519 5057 5047 5044 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m10520 1 5048 5057 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m10521 5056 5048 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m10522 1 5047 5056 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m10523 5058 5047 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m10524 1 5048 5058 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m10525 5059 5048 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m10526 5051 5047 5059 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m10527 5058 5034 5051 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m10528 1 4827 5048 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m10529 5060 5048 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.45e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m10530 5031 4821 5060 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.033e-11 ad=7.53e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.11 
m10531 5061 5047 5031 1 penh l=1.1e-06 w=7.6e-06 
+ as=7.02e-12 ad=9.35e-12 ps=1.01e-05 pd=9.97e-06 
+ nrs=0.12 nrd=0.16 
m10532 1 4827 5061 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=8.12e-12 ps=1.661e-05 pd=1.17e-05 
+ nrs=0.25 nrd=0.1 
m10533 5047 4821 1 1 penh l=1.1e-06 w=1e-05 
+ as=3.05e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.31 nrd=0.22 
m10534 1 5062 151 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m10535 5063 5025 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m10536 5062 5064 5063 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m10537 5065 5066 5062 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10538 1 5039 5065 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m10539 5067 5068 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10540 5066 5069 5067 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m10541 5070 5071 5066 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m10542 1 5072 5070 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m10543 5068 5072 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10544 1 5074 5073 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m10545 5075 5071 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m10546 5064 5074 5075 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m10547 5076 5073 5064 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m10548 1 5069 5076 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m10549 5071 5069 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m10550 0 5062 151 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m10551 5077 5025 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=7.37e-12 ad=1.506e-11 ps=1.097e-05 pd=1.425e-05 
+ nrs=0.13 nrd=0.26 
m10552 5062 5066 5077 0 nenh l=1.1e-06 w=6.4e-06 
+ as=8.77e-12 ad=6.21e-12 ps=9.49e-06 pd=9.23e-06 
+ nrs=0.21 nrd=0.15 
m10553 5078 5064 5062 0 nenh l=1.1e-06 w=5.6e-06 
+ as=5.09e-12 ad=7.67e-12 ps=7.68e-06 pd=8.31e-06 
+ nrs=0.16 nrd=0.24 
m10554 0 5039 5078 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=6.17e-12 ps=1.275e-05 pd=9.32e-06 
+ nrs=0.29 nrd=0.13 
m10555 1 4838 5079 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=2.196e-11 ps=1.359e-05 pd=2.05e-05 
+ nrs=0.31 nrd=0.42 
m10556 5080 5081 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.55e-12 ad=1.603e-11 ps=9.05e-06 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10557 5069 4838 5080 1 penh l=1.1e-06 w=7.6e-06 
+ as=8.13e-12 ad=6.91e-12 ps=9.97e-06 pd=9.55e-06 
+ nrs=0.14 nrd=0.12 
m10558 5082 5079 5069 1 penh l=1.1e-06 w=8.4e-06 
+ as=8.56e-12 ad=8.99e-12 ps=1.088e-05 pd=1.103e-05 
+ nrs=0.12 nrd=0.13 
m10559 1 4844 5082 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=7.34e-12 ps=1.359e-05 pd=9.32e-06 
+ nrs=0.31 nrd=0.14 
m10560 5081 4844 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=2.196e-11 ad=1.603e-11 ps=2.05e-05 pd=1.359e-05 
+ nrs=0.42 nrd=0.31 
m10561 5083 5072 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.55e-11 ad=2.672e-11 ps=1.478e-05 pd=2.265e-05 
+ nrs=0.11 nrd=0.19 
m10562 5032 4838 5083 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.151e-11 ad=1.498e-11 ps=1.394e-05 pd=1.428e-05 
+ nrs=0.09 nrd=0.11 
m10563 5083 4844 5032 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.705e-11 ad=1.309e-11 ps=1.625e-05 pd=1.586e-05 
+ nrs=0.1 nrd=0.08 
m10564 5084 4844 5083 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.498e-11 ps=1.33e-05 pd=1.428e-05 
+ nrs=0.07 nrd=0.11 
m10565 1 4838 5084 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m10566 5085 4838 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m10567 5086 4844 5085 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=9.86e-12 ps=1.428e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m10568 5034 4844 5086 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.309e-11 ad=1.705e-11 ps=1.586e-05 pd=1.625e-05 
+ nrs=0.08 nrd=0.1 
m10569 5086 4838 5034 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=1.151e-11 ps=1.428e-05 pd=1.394e-05 
+ nrs=0.11 nrd=0.09 
m10570 1 5074 5086 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.55e-11 ps=2.265e-05 pd=1.478e-05 
+ nrs=0.19 nrd=0.11 
m10571 5087 5068 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10572 5066 5071 5087 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10573 5088 5069 5066 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10574 0 5072 5088 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10575 5068 5072 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10576 0 5074 5073 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m10577 5089 5071 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10578 5064 5073 5089 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10579 5090 5074 5064 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10580 0 5069 5090 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10581 5071 5069 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10582 0 4838 5079 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m10583 5091 5081 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m10584 5069 5079 5091 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m10585 5092 4838 5069 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m10586 0 4844 5092 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m10587 5081 4844 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m10588 5032 5072 5093 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.175e-11 ad=1.755e-11 ps=1.429e-05 pd=1.841e-05 
+ nrs=0.09 nrd=0.13 
m10589 5094 4838 5032 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.013e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.1 
m10590 0 4844 5094 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=8.5e-12 ps=1.874e-05 pd=1.17e-05 
+ nrs=0.2 nrd=0.08 
m10591 5093 4844 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=2.299e-11 ps=1.841e-05 pd=2.174e-05 
+ nrs=0.13 nrd=0.17 
m10592 0 4838 5093 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=1.513e-11 ps=1.874e-05 pd=1.587e-05 
+ nrs=0.2 nrd=0.15 
m10593 5095 4838 0 0 nenh l=1.1e-06 w=1e-05 
+ as=1.513e-11 ad=1.982e-11 ps=1.587e-05 pd=1.874e-05 
+ nrs=0.15 nrd=0.2 
m10594 0 4844 5095 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.755e-11 ps=2.174e-05 pd=1.841e-05 
+ nrs=0.17 nrd=0.13 
m10595 5096 4844 0 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.982e-11 ps=1.17e-05 pd=1.874e-05 
+ nrs=0.08 nrd=0.2 
m10596 5034 4838 5096 0 nenh l=1.1e-06 w=1e-05 
+ as=1.013e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.1 nrd=0.08 
m10597 5095 5074 5034 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=1.175e-11 ps=1.841e-05 pd=1.429e-05 
+ nrs=0.13 nrd=0.09 
m10598 5097 5025 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.04e-12 ad=1.348e-11 ps=9.88e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m10599 122 5098 5097 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=5.33e-12 ps=8.5e-06 pd=8.72e-06 
+ nrs=0.19 nrd=0.15 
m10600 5099 5100 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10601 5098 5101 5099 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10602 5102 5103 5098 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10603 0 5104 5102 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10604 5100 5104 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10605 0 5106 5105 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m10606 5107 5101 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10607 5108 5105 5107 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10608 5109 5106 5108 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10609 0 5103 5109 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10610 5101 5103 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10611 5110 5108 122 0 nenh l=1.1e-06 w=6e-06 
+ as=5.29e-12 ad=6.86e-12 ps=8.61e-06 pd=8.5e-06 
+ nrs=0.15 nrd=0.19 
m10612 0 5039 5110 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=5.65e-12 ps=1.2e-05 pd=9.19e-06 
+ nrs=0.31 nrd=0.14 
m10613 5072 5104 5111 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.57e-11 ps=1.429e-05 pd=2.04e-05 
+ nrs=0.11 nrd=0.12 
m10614 5112 5113 5072 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m10615 5111 5114 5112 0 nenh l=1.1e-06 w=1e-05 
+ as=1.354e-11 ad=8.5e-12 ps=1.759e-05 pd=1.17e-05 
+ nrs=0.14 nrd=0.08 
m10616 0 5114 5111 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m10617 5111 5113 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m10618 0 5113 5115 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m10619 5115 5114 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m10620 5116 5114 5115 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.354e-11 ps=1.17e-05 pd=1.759e-05 
+ nrs=0.08 nrd=0.14 
m10621 5074 5113 5116 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m10622 5115 5106 5074 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=1.416e-11 ps=2.04e-05 pd=1.429e-05 
+ nrs=0.12 nrd=0.11 
m10623 0 4861 5114 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m10624 5117 5114 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m10625 5103 5113 5117 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m10626 5118 4855 5103 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m10627 0 4861 5118 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m10628 5113 4855 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m10629 5119 5025 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m10630 122 5108 5119 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m10631 5120 5098 122 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10632 1 5039 5120 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m10633 5121 5100 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10634 5098 5103 5121 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m10635 5122 5101 5098 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m10636 1 5104 5122 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m10637 5100 5104 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.308e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.42 nrd=0.4 
m10638 1 5106 5105 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m10639 5123 5101 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10640 5108 5106 5123 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m10641 5124 5105 5108 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m10642 1 5103 5124 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m10643 5101 5103 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10644 5072 5104 5125 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m10645 5126 5113 5072 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m10646 1 5114 5126 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m10647 5125 5114 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m10648 1 5113 5125 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m10649 5127 5113 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m10650 1 5114 5127 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m10651 5128 5114 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m10652 5074 5113 5128 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m10653 5127 5106 5074 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m10654 1 4861 5114 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m10655 5129 5114 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.45e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m10656 5103 4855 5129 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.033e-11 ad=7.53e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.11 
m10657 5130 5113 5103 1 penh l=1.1e-06 w=7.6e-06 
+ as=7.02e-12 ad=9.35e-12 ps=1.01e-05 pd=9.97e-06 
+ nrs=0.12 nrd=0.16 
m10658 1 4861 5130 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=8.12e-12 ps=1.661e-05 pd=1.17e-05 
+ nrs=0.25 nrd=0.1 
m10659 5113 4855 1 1 penh l=1.1e-06 w=1e-05 
+ as=3.05e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.31 nrd=0.22 
m10660 1 5131 93 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m10661 5132 5025 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m10662 5131 5133 5132 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m10663 5134 5135 5131 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10664 1 5039 5134 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m10665 5025 5039 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.484e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m10666 1 5039 5025 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.484e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m10667 5039 5136 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m10668 1 5136 5039 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m10669 5135 5133 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.596e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.51 nrd=0.4 
m10670 1 4872 5137 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m10671 5138 5139 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m10672 5133 4872 5138 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m10673 5140 5137 5133 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m10674 1 4878 5140 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m10675 5139 4878 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m10676 0 5131 93 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.42e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.45 
m10677 5141 5025 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=7.37e-12 ad=1.506e-11 ps=1.097e-05 pd=1.425e-05 
+ nrs=0.13 nrd=0.26 
m10678 5131 5135 5141 0 nenh l=1.1e-06 w=6.4e-06 
+ as=8.77e-12 ad=6.21e-12 ps=9.49e-06 pd=9.23e-06 
+ nrs=0.21 nrd=0.15 
m10679 5142 5133 5131 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=7.67e-12 ps=7.3e-06 pd=8.31e-06 
+ nrs=0.15 nrd=0.24 
m10680 0 5039 5142 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m10681 5025 5039 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.254e-11 ad=1.506e-11 ps=1.09e-05 pd=1.425e-05 
+ nrs=0.22 nrd=0.26 
m10682 0 5039 5025 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.506e-11 ad=1.254e-11 ps=1.425e-05 pd=1.09e-05 
+ nrs=0.26 nrd=0.22 
m10683 5039 5136 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m10684 0 5136 5039 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m10685 5135 5133 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10686 5143 4872 5104 1 penh l=1.1e-06 w=1.44e-05 
+ as=1.224e-11 ad=4.04e-11 ps=1.61e-05 pd=3.49e-05 
+ nrs=0.06 nrd=0.19 
m10687 1 4878 5143 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.224e-11 ps=2.718e-05 pd=1.61e-05 
+ nrs=0.15 nrd=0.06 
m10688 5136 5144 1 1 penh l=1.1e-06 w=1.44e-05 
+ as=2.376e-11 ad=3.206e-11 ps=1.77e-05 pd=2.718e-05 
+ nrs=0.11 nrd=0.15 
m10689 1 5144 5136 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=2.376e-11 ps=2.718e-05 pd=1.77e-05 
+ nrs=0.15 nrd=0.11 
m10690 5144 4915 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.98e-11 ad=2.672e-11 ps=1.53e-05 pd=2.265e-05 
+ nrs=0.14 nrd=0.19 
m10691 5145 5010 5144 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.02e-11 ad=1.98e-11 ps=1.37e-05 pd=1.53e-05 
+ nrs=0.07 nrd=0.14 
m10692 1 4922 5145 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.02e-11 ps=2.265e-05 pd=1.37e-05 
+ nrs=0.19 nrd=0.07 
m10693 5106 4872 1 1 penh l=1.1e-06 w=1.28e-05 
+ as=1.264e-11 ad=2.85e-11 ps=1.53e-05 pd=2.416e-05 
+ nrs=0.08 nrd=0.17 
m10694 1 4878 5106 1 penh l=1.1e-06 w=1.28e-05 
+ as=2.85e-11 ad=1.264e-11 ps=2.416e-05 pd=1.53e-05 
+ nrs=0.17 nrd=0.08 
m10695 0 4872 5137 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.031e-11 ad=1.586e-11 ps=9.75e-06 pd=1.65e-05 
+ nrs=0.38 nrd=0.59 
m10696 5146 5139 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.32e-12 ad=1.348e-11 ps=9.63e-06 pd=1.275e-05 
+ nrs=0.14 nrd=0.29 
m10697 5133 5137 5146 0 nenh l=1.1e-06 w=5.2e-06 
+ as=8.58e-12 ad=4.84e-12 ps=8.5e-06 pd=7.37e-06 
+ nrs=0.32 nrd=0.18 
m10698 5147 4872 5133 0 nenh l=1.1e-06 w=5.2e-06 
+ as=4.56e-12 ad=8.58e-12 ps=7.37e-06 pd=8.5e-06 
+ nrs=0.17 nrd=0.32 
m10699 0 4878 5147 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.96e-12 ps=1.275e-05 pd=9.63e-06 
+ nrs=0.29 nrd=0.13 
m10700 5139 4878 0 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.031e-11 ps=1.65e-05 pd=9.75e-06 
+ nrs=0.59 nrd=0.38 
m10701 5104 4872 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=1.06e-11 ad=2.061e-11 ps=1.29e-05 pd=1.949e-05 
+ nrs=0.1 nrd=0.19 
m10702 0 4878 5104 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.061e-11 ad=1.06e-11 ps=1.949e-05 pd=1.29e-05 
+ nrs=0.19 nrd=0.1 
m10703 5136 5144 0 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.584e-11 ad=1.903e-11 ps=1.29e-05 pd=1.799e-05 
+ nrs=0.17 nrd=0.21 
m10704 0 5144 5136 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=1.584e-11 ps=1.799e-05 pd=1.29e-05 
+ nrs=0.21 nrd=0.17 
m10705 5148 4915 0 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.955e-11 ad=1.903e-11 ps=1.68e-05 pd=1.799e-05 
+ nrs=0.21 nrd=0.21 
m10706 5144 5010 5148 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.604e-11 ad=1.955e-11 ps=1.303e-05 pd=1.68e-05 
+ nrs=0.17 nrd=0.21 
m10707 5148 4922 5144 0 nenh l=1.1e-06 w=1e-05 
+ as=2.036e-11 ad=1.67e-11 ps=1.75e-05 pd=1.357e-05 
+ nrs=0.2 nrd=0.17 
m10708 5149 4872 5106 0 nenh l=1.1e-06 w=1.28e-05 
+ as=1.088e-11 ad=3.904e-11 ps=1.45e-05 pd=3.17e-05 
+ nrs=0.07 nrd=0.24 
m10709 0 4878 5149 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.088e-11 ps=2.399e-05 pd=1.45e-05 
+ nrs=0.15 nrd=0.07 
m10710 5150 5151 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=5.99e-12 ad=1.348e-11 ps=9.58e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m10711 296 5152 5150 0 nenh l=1.1e-06 w=6.4e-06 
+ as=7.52e-12 ad=5.63e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.14 
m10712 5153 5154 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10713 5152 5155 5153 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10714 5156 5157 5152 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10715 0 5158 5156 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10716 5154 5158 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10717 0 5160 5159 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m10718 5161 5155 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10719 5162 5159 5161 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10720 5163 5160 5162 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10721 0 5157 5163 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10722 5155 5157 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10723 5164 5162 296 0 nenh l=1.1e-06 w=6.4e-06 
+ as=5.63e-12 ad=7.52e-12 ps=9.02e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10724 0 5165 5164 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.99e-12 ps=1.275e-05 pd=9.58e-06 
+ nrs=0.29 nrd=0.13 
m10725 5166 5151 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m10726 296 5162 5166 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m10727 5167 5152 296 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10728 1 5165 5167 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m10729 5168 5154 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10730 5152 5157 5168 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m10731 5169 5155 5152 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m10732 1 5158 5169 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m10733 5154 5158 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10734 5170 5158 5171 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.745e-11 ps=1.429e-05 pd=2.077e-05 
+ nrs=0.11 nrd=0.13 
m10735 5172 5173 5170 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m10736 5171 5174 5172 0 nenh l=1.1e-06 w=1e-05 
+ as=1.505e-11 ad=8.5e-12 ps=1.791e-05 pd=1.17e-05 
+ nrs=0.15 nrd=0.08 
m10737 0 5174 5171 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.745e-11 ps=2.174e-05 pd=2.077e-05 
+ nrs=0.17 nrd=0.13 
m10738 5171 5173 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=1.625e-11 ad=2.141e-11 ps=1.934e-05 pd=2.024e-05 
+ nrs=0.14 nrd=0.18 
m10739 0 5173 5175 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.625e-11 ps=2.024e-05 pd=1.934e-05 
+ nrs=0.18 nrd=0.14 
m10740 5175 5174 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.745e-11 ad=2.299e-11 ps=2.077e-05 pd=2.174e-05 
+ nrs=0.13 nrd=0.17 
m10741 5176 5174 5175 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.505e-11 ps=1.17e-05 pd=1.791e-05 
+ nrs=0.08 nrd=0.15 
m10742 5177 5173 5176 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m10743 5175 5160 5177 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.745e-11 ad=1.416e-11 ps=2.077e-05 pd=1.429e-05 
+ nrs=0.13 nrd=0.11 
m10744 0 4759 5174 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m10745 5178 5174 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m10746 5157 5173 5178 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m10747 5179 4753 5157 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m10748 0 4759 5179 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m10749 5173 4753 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m10750 1 5160 5159 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m10751 5180 5155 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m10752 5162 5160 5180 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m10753 5181 5159 5162 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m10754 1 5157 5181 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m10755 5155 5157 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m10756 5170 5158 5182 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m10757 5183 5173 5170 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m10758 1 5174 5183 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m10759 5182 5174 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m10760 1 5173 5182 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m10761 5184 5173 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m10762 1 5174 5184 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m10763 5185 5174 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m10764 5177 5173 5185 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m10765 5184 5160 5177 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m10766 1 4759 5174 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m10767 5186 5174 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.45e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m10768 5157 4753 5186 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.033e-11 ad=7.53e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.11 
m10769 5187 5173 5157 1 penh l=1.1e-06 w=7.6e-06 
+ as=7.02e-12 ad=9.35e-12 ps=1.01e-05 pd=9.97e-06 
+ nrs=0.12 nrd=0.16 
m10770 1 4759 5187 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=8.12e-12 ps=1.661e-05 pd=1.17e-05 
+ nrs=0.25 nrd=0.1 
m10771 5173 4753 1 1 penh l=1.1e-06 w=1e-05 
+ as=3.05e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.31 nrd=0.22 
m10772 1 5188 267 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m10773 5189 5151 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m10774 5188 5190 5189 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m10775 5191 5192 5188 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10776 1 5165 5191 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m10777 5193 5194 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10778 5192 5195 5193 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m10779 5196 5197 5192 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m10780 1 5198 5196 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m10781 5194 5198 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10782 1 5200 5199 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m10783 5201 5197 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m10784 5190 5200 5201 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m10785 5202 5199 5190 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m10786 1 5195 5202 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m10787 5197 5195 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m10788 0 5188 267 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.031e-11 ad=1.586e-11 ps=9.75e-06 pd=1.65e-05 
+ nrs=0.38 nrd=0.59 
m10789 5203 5151 0 0 nenh l=1.1e-06 w=7.2e-06 
+ as=6.43e-12 ad=1.427e-11 ps=1.058e-05 pd=1.35e-05 
+ nrs=0.12 nrd=0.28 
m10790 5188 5192 5203 0 nenh l=1.1e-06 w=6e-06 
+ as=8.27e-12 ad=5.35e-12 ps=9.11e-06 pd=8.82e-06 
+ nrs=0.23 nrd=0.15 
m10791 5204 5190 5188 0 nenh l=1.1e-06 w=5.2e-06 
+ as=4.53e-12 ad=7.17e-12 ps=7.26e-06 pd=7.89e-06 
+ nrs=0.17 nrd=0.27 
m10792 0 5165 5204 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=5.57e-12 ps=1.2e-05 pd=8.94e-06 
+ nrs=0.31 nrd=0.14 
m10793 1 4770 5205 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=2.196e-11 ps=1.359e-05 pd=2.05e-05 
+ nrs=0.31 nrd=0.42 
m10794 5206 5207 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.55e-12 ad=1.603e-11 ps=9.05e-06 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10795 5195 4770 5206 1 penh l=1.1e-06 w=7.6e-06 
+ as=8.13e-12 ad=6.91e-12 ps=9.97e-06 pd=9.55e-06 
+ nrs=0.14 nrd=0.12 
m10796 5208 5205 5195 1 penh l=1.1e-06 w=8.4e-06 
+ as=8.56e-12 ad=8.99e-12 ps=1.088e-05 pd=1.103e-05 
+ nrs=0.12 nrd=0.13 
m10797 1 4776 5208 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=7.34e-12 ps=1.359e-05 pd=9.32e-06 
+ nrs=0.31 nrd=0.14 
m10798 5207 4776 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=2.196e-11 ad=1.603e-11 ps=2.05e-05 pd=1.359e-05 
+ nrs=0.42 nrd=0.31 
m10799 5209 5198 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.55e-11 ad=2.672e-11 ps=1.478e-05 pd=2.265e-05 
+ nrs=0.11 nrd=0.19 
m10800 5158 4770 5209 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.151e-11 ad=1.498e-11 ps=1.394e-05 pd=1.428e-05 
+ nrs=0.09 nrd=0.11 
m10801 5209 4776 5158 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.705e-11 ad=1.309e-11 ps=1.625e-05 pd=1.586e-05 
+ nrs=0.1 nrd=0.08 
m10802 5210 4776 5209 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.498e-11 ps=1.33e-05 pd=1.428e-05 
+ nrs=0.07 nrd=0.11 
m10803 1 4770 5210 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m10804 5211 4770 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m10805 5212 4776 5211 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=9.86e-12 ps=1.428e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m10806 5160 4776 5212 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.309e-11 ad=1.705e-11 ps=1.586e-05 pd=1.625e-05 
+ nrs=0.08 nrd=0.1 
m10807 5212 4770 5160 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=1.151e-11 ps=1.428e-05 pd=1.394e-05 
+ nrs=0.11 nrd=0.09 
m10808 1 5200 5212 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.55e-11 ps=2.265e-05 pd=1.478e-05 
+ nrs=0.19 nrd=0.11 
m10809 5213 5194 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10810 5192 5197 5213 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10811 5214 5195 5192 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10812 0 5198 5214 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10813 5194 5198 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10814 0 5200 5199 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m10815 5215 5197 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10816 5190 5199 5215 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10817 5216 5200 5190 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10818 0 5195 5216 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10819 5197 5195 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10820 0 4770 5205 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m10821 5217 5207 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m10822 5195 5205 5217 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m10823 5218 4770 5195 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m10824 0 4776 5218 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m10825 5207 4776 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m10826 5158 5198 5219 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.175e-11 ad=1.755e-11 ps=1.429e-05 pd=1.841e-05 
+ nrs=0.09 nrd=0.13 
m10827 5220 4770 5158 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.013e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.1 
m10828 0 4776 5220 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=8.5e-12 ps=1.874e-05 pd=1.17e-05 
+ nrs=0.2 nrd=0.08 
m10829 5219 4776 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=2.299e-11 ps=1.841e-05 pd=2.174e-05 
+ nrs=0.13 nrd=0.17 
m10830 0 4770 5219 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=1.513e-11 ps=1.874e-05 pd=1.587e-05 
+ nrs=0.2 nrd=0.15 
m10831 5221 4770 0 0 nenh l=1.1e-06 w=1e-05 
+ as=1.513e-11 ad=1.982e-11 ps=1.587e-05 pd=1.874e-05 
+ nrs=0.15 nrd=0.2 
m10832 0 4776 5221 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.755e-11 ps=2.174e-05 pd=1.841e-05 
+ nrs=0.17 nrd=0.13 
m10833 5222 4776 0 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.982e-11 ps=1.17e-05 pd=1.874e-05 
+ nrs=0.08 nrd=0.2 
m10834 5160 4770 5222 0 nenh l=1.1e-06 w=1e-05 
+ as=1.013e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.1 nrd=0.08 
m10835 5221 5200 5160 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=1.175e-11 ps=1.841e-05 pd=1.429e-05 
+ nrs=0.13 nrd=0.09 
m10836 5223 5151 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.04e-12 ad=1.348e-11 ps=9.88e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m10837 238 5224 5223 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=5.33e-12 ps=8.5e-06 pd=8.72e-06 
+ nrs=0.19 nrd=0.15 
m10838 5225 5226 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10839 5224 5227 5225 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10840 5228 5229 5224 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10841 0 5230 5228 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10842 5226 5230 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10843 0 5232 5231 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m10844 5233 5227 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10845 5234 5231 5233 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10846 5235 5232 5234 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10847 0 5229 5235 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10848 5227 5229 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10849 5236 5234 238 0 nenh l=1.1e-06 w=6e-06 
+ as=5.29e-12 ad=6.86e-12 ps=8.61e-06 pd=8.5e-06 
+ nrs=0.15 nrd=0.19 
m10850 0 5165 5236 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=5.65e-12 ps=1.2e-05 pd=9.19e-06 
+ nrs=0.31 nrd=0.14 
m10851 5198 5230 5237 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.57e-11 ps=1.429e-05 pd=2.04e-05 
+ nrs=0.11 nrd=0.12 
m10852 5238 5239 5198 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m10853 5237 5240 5238 0 nenh l=1.1e-06 w=1e-05 
+ as=1.354e-11 ad=8.5e-12 ps=1.759e-05 pd=1.17e-05 
+ nrs=0.14 nrd=0.08 
m10854 0 5240 5237 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m10855 5237 5239 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m10856 0 5239 5241 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m10857 5241 5240 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m10858 5242 5240 5241 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.354e-11 ps=1.17e-05 pd=1.759e-05 
+ nrs=0.08 nrd=0.14 
m10859 5200 5239 5242 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m10860 5241 5232 5200 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=1.416e-11 ps=2.04e-05 pd=1.429e-05 
+ nrs=0.12 nrd=0.11 
m10861 0 4793 5240 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m10862 5243 5240 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m10863 5229 5239 5243 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m10864 5244 4787 5229 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m10865 0 4793 5244 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m10866 5239 4787 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m10867 5245 5151 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m10868 238 5234 5245 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m10869 5246 5224 238 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10870 1 5165 5246 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m10871 5247 5226 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10872 5224 5229 5247 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m10873 5248 5227 5224 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m10874 1 5230 5248 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m10875 5226 5230 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.308e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.42 nrd=0.4 
m10876 1 5232 5231 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m10877 5249 5227 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10878 5234 5232 5249 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m10879 5250 5231 5234 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m10880 1 5229 5250 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m10881 5227 5229 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10882 5198 5230 5251 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m10883 5252 5239 5198 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m10884 1 5240 5252 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m10885 5251 5240 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m10886 1 5239 5251 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m10887 5253 5239 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m10888 1 5240 5253 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m10889 5254 5240 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m10890 5200 5239 5254 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m10891 5253 5232 5200 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m10892 1 4793 5240 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m10893 5255 5240 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.45e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m10894 5229 4787 5255 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.033e-11 ad=7.53e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.11 
m10895 5256 5239 5229 1 penh l=1.1e-06 w=7.6e-06 
+ as=7.02e-12 ad=9.35e-12 ps=1.01e-05 pd=9.97e-06 
+ nrs=0.12 nrd=0.16 
m10896 1 4793 5256 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=8.12e-12 ps=1.661e-05 pd=1.17e-05 
+ nrs=0.25 nrd=0.1 
m10897 5239 4787 1 1 penh l=1.1e-06 w=1e-05 
+ as=3.05e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.31 nrd=0.22 
m10898 1 5257 209 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m10899 5258 5151 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m10900 5257 5259 5258 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m10901 5260 5261 5257 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10902 1 5165 5260 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m10903 5151 5165 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.484e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m10904 1 5165 5151 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.484e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m10905 5165 5262 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m10906 1 5262 5165 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m10907 5261 5259 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.596e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.51 nrd=0.4 
m10908 1 4804 5263 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m10909 5264 5265 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m10910 5259 4804 5264 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m10911 5266 5263 5259 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m10912 1 4810 5266 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m10913 5265 4810 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m10914 0 5257 209 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.42e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.45 
m10915 5267 5151 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=7.37e-12 ad=1.506e-11 ps=1.097e-05 pd=1.425e-05 
+ nrs=0.13 nrd=0.26 
m10916 5257 5261 5267 0 nenh l=1.1e-06 w=6.4e-06 
+ as=8.77e-12 ad=6.21e-12 ps=9.49e-06 pd=9.23e-06 
+ nrs=0.21 nrd=0.15 
m10917 5268 5259 5257 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=7.67e-12 ps=7.3e-06 pd=8.31e-06 
+ nrs=0.15 nrd=0.24 
m10918 0 5165 5268 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m10919 5151 5165 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.254e-11 ad=1.506e-11 ps=1.09e-05 pd=1.425e-05 
+ nrs=0.22 nrd=0.26 
m10920 0 5165 5151 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.506e-11 ad=1.254e-11 ps=1.425e-05 pd=1.09e-05 
+ nrs=0.26 nrd=0.22 
m10921 5165 5262 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m10922 0 5262 5165 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m10923 5261 5259 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10924 5269 4804 5230 1 penh l=1.1e-06 w=1.44e-05 
+ as=1.224e-11 ad=4.04e-11 ps=1.61e-05 pd=3.49e-05 
+ nrs=0.06 nrd=0.19 
m10925 1 4810 5269 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.224e-11 ps=2.718e-05 pd=1.61e-05 
+ nrs=0.15 nrd=0.06 
m10926 5262 5270 1 1 penh l=1.1e-06 w=1.44e-05 
+ as=2.376e-11 ad=3.206e-11 ps=1.77e-05 pd=2.718e-05 
+ nrs=0.11 nrd=0.15 
m10927 1 5270 5262 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=2.376e-11 ps=2.718e-05 pd=1.77e-05 
+ nrs=0.15 nrd=0.11 
m10928 5270 5044 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.98e-11 ad=2.672e-11 ps=1.53e-05 pd=2.265e-05 
+ nrs=0.14 nrd=0.19 
m10929 5271 5136 5270 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.02e-11 ad=1.98e-11 ps=1.37e-05 pd=1.53e-05 
+ nrs=0.07 nrd=0.14 
m10930 1 5051 5271 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.02e-11 ps=2.265e-05 pd=1.37e-05 
+ nrs=0.19 nrd=0.07 
m10931 5232 4804 1 1 penh l=1.1e-06 w=1.28e-05 
+ as=1.264e-11 ad=2.85e-11 ps=1.53e-05 pd=2.416e-05 
+ nrs=0.08 nrd=0.17 
m10932 1 4810 5232 1 penh l=1.1e-06 w=1.28e-05 
+ as=2.85e-11 ad=1.264e-11 ps=2.416e-05 pd=1.53e-05 
+ nrs=0.17 nrd=0.08 
m10933 0 4804 5263 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.031e-11 ad=1.586e-11 ps=9.75e-06 pd=1.65e-05 
+ nrs=0.38 nrd=0.59 
m10934 5272 5265 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.32e-12 ad=1.348e-11 ps=9.63e-06 pd=1.275e-05 
+ nrs=0.14 nrd=0.29 
m10935 5259 5263 5272 0 nenh l=1.1e-06 w=5.2e-06 
+ as=8.58e-12 ad=4.84e-12 ps=8.5e-06 pd=7.37e-06 
+ nrs=0.32 nrd=0.18 
m10936 5273 4804 5259 0 nenh l=1.1e-06 w=5.2e-06 
+ as=4.56e-12 ad=8.58e-12 ps=7.37e-06 pd=8.5e-06 
+ nrs=0.17 nrd=0.32 
m10937 0 4810 5273 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.96e-12 ps=1.275e-05 pd=9.63e-06 
+ nrs=0.29 nrd=0.13 
m10938 5265 4810 0 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.031e-11 ps=1.65e-05 pd=9.75e-06 
+ nrs=0.59 nrd=0.38 
m10939 5230 4804 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=1.06e-11 ad=2.061e-11 ps=1.29e-05 pd=1.949e-05 
+ nrs=0.1 nrd=0.19 
m10940 0 4810 5230 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.061e-11 ad=1.06e-11 ps=1.949e-05 pd=1.29e-05 
+ nrs=0.19 nrd=0.1 
m10941 5262 5270 0 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.584e-11 ad=1.903e-11 ps=1.29e-05 pd=1.799e-05 
+ nrs=0.17 nrd=0.21 
m10942 0 5270 5262 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=1.584e-11 ps=1.799e-05 pd=1.29e-05 
+ nrs=0.21 nrd=0.17 
m10943 5274 5044 0 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.955e-11 ad=1.903e-11 ps=1.68e-05 pd=1.799e-05 
+ nrs=0.21 nrd=0.21 
m10944 5270 5136 5274 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.604e-11 ad=1.955e-11 ps=1.303e-05 pd=1.68e-05 
+ nrs=0.17 nrd=0.21 
m10945 5274 5051 5270 0 nenh l=1.1e-06 w=1e-05 
+ as=2.036e-11 ad=1.67e-11 ps=1.75e-05 pd=1.357e-05 
+ nrs=0.2 nrd=0.17 
m10946 5275 4804 5232 0 nenh l=1.1e-06 w=1.28e-05 
+ as=1.088e-11 ad=3.904e-11 ps=1.45e-05 pd=3.17e-05 
+ nrs=0.07 nrd=0.24 
m10947 0 4810 5275 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.088e-11 ps=2.399e-05 pd=1.45e-05 
+ nrs=0.15 nrd=0.07 
m10948 5276 5277 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=5.99e-12 ad=1.348e-11 ps=9.58e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m10949 412 5278 5276 0 nenh l=1.1e-06 w=6.4e-06 
+ as=7.52e-12 ad=5.63e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.14 
m10950 5279 5280 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10951 5278 5281 5279 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10952 5282 5283 5278 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10953 0 5284 5282 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10954 5280 5284 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10955 0 5286 5285 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m10956 5287 5281 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m10957 5288 5285 5287 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m10958 5289 5286 5288 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m10959 0 5283 5289 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m10960 5281 5283 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m10961 5290 5288 412 0 nenh l=1.1e-06 w=6.4e-06 
+ as=5.63e-12 ad=7.52e-12 ps=9.02e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10962 0 5291 5290 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.99e-12 ps=1.275e-05 pd=9.58e-06 
+ nrs=0.29 nrd=0.13 
m10963 5292 5277 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m10964 412 5288 5292 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m10965 5293 5278 412 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m10966 1 5291 5293 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m10967 5294 5280 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m10968 5278 5283 5294 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m10969 5295 5281 5278 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m10970 1 5284 5295 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m10971 5280 5284 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m10972 5296 5284 5297 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.745e-11 ps=1.429e-05 pd=2.077e-05 
+ nrs=0.11 nrd=0.13 
m10973 5298 5299 5296 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m10974 5297 5300 5298 0 nenh l=1.1e-06 w=1e-05 
+ as=1.505e-11 ad=8.5e-12 ps=1.791e-05 pd=1.17e-05 
+ nrs=0.15 nrd=0.08 
m10975 0 5300 5297 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.745e-11 ps=2.174e-05 pd=2.077e-05 
+ nrs=0.17 nrd=0.13 
m10976 5297 5299 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=1.625e-11 ad=2.141e-11 ps=1.934e-05 pd=2.024e-05 
+ nrs=0.14 nrd=0.18 
m10977 0 5299 5301 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.625e-11 ps=2.024e-05 pd=1.934e-05 
+ nrs=0.18 nrd=0.14 
m10978 5301 5300 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.745e-11 ad=2.299e-11 ps=2.077e-05 pd=2.174e-05 
+ nrs=0.13 nrd=0.17 
m10979 5302 5300 5301 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.505e-11 ps=1.17e-05 pd=1.791e-05 
+ nrs=0.08 nrd=0.15 
m10980 5303 5299 5302 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m10981 5301 5286 5303 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.745e-11 ad=1.416e-11 ps=2.077e-05 pd=1.429e-05 
+ nrs=0.13 nrd=0.11 
m10982 0 4691 5300 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m10983 5304 5300 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m10984 5283 5299 5304 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m10985 5305 4685 5283 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m10986 0 4691 5305 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m10987 5299 4685 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m10988 1 5286 5285 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m10989 5306 5281 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m10990 5288 5286 5306 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m10991 5307 5285 5288 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m10992 1 5283 5307 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m10993 5281 5283 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m10994 5296 5284 5308 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m10995 5309 5299 5296 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m10996 1 5300 5309 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m10997 5308 5300 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m10998 1 5299 5308 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m10999 5310 5299 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m11000 1 5300 5310 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m11001 5311 5300 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m11002 5303 5299 5311 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m11003 5310 5286 5303 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m11004 1 4691 5300 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m11005 5312 5300 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.45e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m11006 5283 4685 5312 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.033e-11 ad=7.53e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.11 
m11007 5313 5299 5283 1 penh l=1.1e-06 w=7.6e-06 
+ as=7.02e-12 ad=9.35e-12 ps=1.01e-05 pd=9.97e-06 
+ nrs=0.12 nrd=0.16 
m11008 1 4691 5313 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=8.12e-12 ps=1.661e-05 pd=1.17e-05 
+ nrs=0.25 nrd=0.1 
m11009 5299 4685 1 1 penh l=1.1e-06 w=1e-05 
+ as=3.05e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.31 nrd=0.22 
m11010 1 5314 383 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m11011 5315 5277 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m11012 5314 5316 5315 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m11013 5317 5318 5314 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m11014 1 5291 5317 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m11015 5319 5320 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m11016 5318 5321 5319 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m11017 5322 5323 5318 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m11018 1 5324 5322 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m11019 5320 5324 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m11020 1 5326 5325 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m11021 5327 5323 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m11022 5316 5326 5327 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m11023 5328 5325 5316 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m11024 1 5321 5328 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m11025 5323 5321 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m11026 0 5314 383 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.031e-11 ad=1.586e-11 ps=9.75e-06 pd=1.65e-05 
+ nrs=0.38 nrd=0.59 
m11027 5329 5277 0 0 nenh l=1.1e-06 w=7.2e-06 
+ as=6.43e-12 ad=1.427e-11 ps=1.058e-05 pd=1.35e-05 
+ nrs=0.12 nrd=0.28 
m11028 5314 5318 5329 0 nenh l=1.1e-06 w=6e-06 
+ as=8.27e-12 ad=5.35e-12 ps=9.11e-06 pd=8.82e-06 
+ nrs=0.23 nrd=0.15 
m11029 5330 5316 5314 0 nenh l=1.1e-06 w=5.2e-06 
+ as=4.53e-12 ad=7.17e-12 ps=7.26e-06 pd=7.89e-06 
+ nrs=0.17 nrd=0.27 
m11030 0 5291 5330 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=5.57e-12 ps=1.2e-05 pd=8.94e-06 
+ nrs=0.31 nrd=0.14 
m11031 1 4702 5331 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=2.196e-11 ps=1.359e-05 pd=2.05e-05 
+ nrs=0.31 nrd=0.42 
m11032 5332 5333 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.55e-12 ad=1.603e-11 ps=9.05e-06 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m11033 5321 4702 5332 1 penh l=1.1e-06 w=7.6e-06 
+ as=8.13e-12 ad=6.91e-12 ps=9.97e-06 pd=9.55e-06 
+ nrs=0.14 nrd=0.12 
m11034 5334 5331 5321 1 penh l=1.1e-06 w=8.4e-06 
+ as=8.56e-12 ad=8.99e-12 ps=1.088e-05 pd=1.103e-05 
+ nrs=0.12 nrd=0.13 
m11035 1 4708 5334 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=7.34e-12 ps=1.359e-05 pd=9.32e-06 
+ nrs=0.31 nrd=0.14 
m11036 5333 4708 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=2.196e-11 ad=1.603e-11 ps=2.05e-05 pd=1.359e-05 
+ nrs=0.42 nrd=0.31 
m11037 5335 5324 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.55e-11 ad=2.672e-11 ps=1.478e-05 pd=2.265e-05 
+ nrs=0.11 nrd=0.19 
m11038 5284 4702 5335 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.151e-11 ad=1.498e-11 ps=1.394e-05 pd=1.428e-05 
+ nrs=0.09 nrd=0.11 
m11039 5335 4708 5284 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.705e-11 ad=1.309e-11 ps=1.625e-05 pd=1.586e-05 
+ nrs=0.1 nrd=0.08 
m11040 5336 4708 5335 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.498e-11 ps=1.33e-05 pd=1.428e-05 
+ nrs=0.07 nrd=0.11 
m11041 1 4702 5336 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m11042 5337 4702 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m11043 5338 4708 5337 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=9.86e-12 ps=1.428e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m11044 5286 4708 5338 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.309e-11 ad=1.705e-11 ps=1.586e-05 pd=1.625e-05 
+ nrs=0.08 nrd=0.1 
m11045 5338 4702 5286 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=1.151e-11 ps=1.428e-05 pd=1.394e-05 
+ nrs=0.11 nrd=0.09 
m11046 1 5326 5338 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.55e-11 ps=2.265e-05 pd=1.478e-05 
+ nrs=0.19 nrd=0.11 
m11047 5339 5320 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m11048 5318 5323 5339 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m11049 5340 5321 5318 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m11050 0 5324 5340 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m11051 5320 5324 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11052 0 5326 5325 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m11053 5341 5323 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m11054 5316 5325 5341 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m11055 5342 5326 5316 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m11056 0 5321 5342 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m11057 5323 5321 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11058 0 4702 5331 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m11059 5343 5333 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m11060 5321 5331 5343 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m11061 5344 4702 5321 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m11062 0 4708 5344 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m11063 5333 4708 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m11064 5284 5324 5345 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.175e-11 ad=1.755e-11 ps=1.429e-05 pd=1.841e-05 
+ nrs=0.09 nrd=0.13 
m11065 5346 4702 5284 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.013e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.1 
m11066 0 4708 5346 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=8.5e-12 ps=1.874e-05 pd=1.17e-05 
+ nrs=0.2 nrd=0.08 
m11067 5345 4708 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=2.299e-11 ps=1.841e-05 pd=2.174e-05 
+ nrs=0.13 nrd=0.17 
m11068 0 4702 5345 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=1.513e-11 ps=1.874e-05 pd=1.587e-05 
+ nrs=0.2 nrd=0.15 
m11069 5347 4702 0 0 nenh l=1.1e-06 w=1e-05 
+ as=1.513e-11 ad=1.982e-11 ps=1.587e-05 pd=1.874e-05 
+ nrs=0.15 nrd=0.2 
m11070 0 4708 5347 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.755e-11 ps=2.174e-05 pd=1.841e-05 
+ nrs=0.17 nrd=0.13 
m11071 5348 4708 0 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.982e-11 ps=1.17e-05 pd=1.874e-05 
+ nrs=0.08 nrd=0.2 
m11072 5286 4702 5348 0 nenh l=1.1e-06 w=1e-05 
+ as=1.013e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.1 nrd=0.08 
m11073 5347 5326 5286 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=1.175e-11 ps=1.841e-05 pd=1.429e-05 
+ nrs=0.13 nrd=0.09 
m11074 5349 5277 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.04e-12 ad=1.348e-11 ps=9.88e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m11075 354 5350 5349 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=5.33e-12 ps=8.5e-06 pd=8.72e-06 
+ nrs=0.19 nrd=0.15 
m11076 5351 5352 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m11077 5350 5353 5351 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m11078 5354 5355 5350 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m11079 0 5356 5354 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m11080 5352 5356 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11081 0 5358 5357 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m11082 5359 5353 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m11083 5360 5357 5359 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m11084 5361 5358 5360 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m11085 0 5355 5361 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m11086 5353 5355 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11087 5362 5360 354 0 nenh l=1.1e-06 w=6e-06 
+ as=5.29e-12 ad=6.86e-12 ps=8.61e-06 pd=8.5e-06 
+ nrs=0.15 nrd=0.19 
m11088 0 5291 5362 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=5.65e-12 ps=1.2e-05 pd=9.19e-06 
+ nrs=0.31 nrd=0.14 
m11089 5324 5356 5363 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.57e-11 ps=1.429e-05 pd=2.04e-05 
+ nrs=0.11 nrd=0.12 
m11090 5364 5365 5324 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m11091 5363 5366 5364 0 nenh l=1.1e-06 w=1e-05 
+ as=1.354e-11 ad=8.5e-12 ps=1.759e-05 pd=1.17e-05 
+ nrs=0.14 nrd=0.08 
m11092 0 5366 5363 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m11093 5363 5365 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m11094 0 5365 5367 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m11095 5367 5366 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m11096 5368 5366 5367 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.354e-11 ps=1.17e-05 pd=1.759e-05 
+ nrs=0.08 nrd=0.14 
m11097 5326 5365 5368 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m11098 5367 5358 5326 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=1.416e-11 ps=2.04e-05 pd=1.429e-05 
+ nrs=0.12 nrd=0.11 
m11099 0 4725 5366 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m11100 5369 5366 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m11101 5355 5365 5369 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m11102 5370 4719 5355 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m11103 0 4725 5370 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m11104 5365 4719 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m11105 5371 5277 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m11106 354 5360 5371 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m11107 5372 5350 354 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m11108 1 5291 5372 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m11109 5373 5352 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m11110 5350 5355 5373 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m11111 5374 5353 5350 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m11112 1 5356 5374 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m11113 5352 5356 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.308e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.42 nrd=0.4 
m11114 1 5358 5357 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m11115 5375 5353 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m11116 5360 5358 5375 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m11117 5376 5357 5360 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m11118 1 5355 5376 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m11119 5353 5355 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m11120 5324 5356 5377 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m11121 5378 5365 5324 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m11122 1 5366 5378 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m11123 5377 5366 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m11124 1 5365 5377 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m11125 5379 5365 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m11126 1 5366 5379 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m11127 5380 5366 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m11128 5326 5365 5380 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m11129 5379 5358 5326 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m11130 1 4725 5366 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m11131 5381 5366 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.45e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m11132 5355 4719 5381 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.033e-11 ad=7.53e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.11 
m11133 5382 5365 5355 1 penh l=1.1e-06 w=7.6e-06 
+ as=7.02e-12 ad=9.35e-12 ps=1.01e-05 pd=9.97e-06 
+ nrs=0.12 nrd=0.16 
m11134 1 4725 5382 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=8.12e-12 ps=1.661e-05 pd=1.17e-05 
+ nrs=0.25 nrd=0.1 
m11135 5365 4719 1 1 penh l=1.1e-06 w=1e-05 
+ as=3.05e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.31 nrd=0.22 
m11136 1 5383 325 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m11137 5384 5277 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m11138 5383 5385 5384 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m11139 5386 5387 5383 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m11140 1 5291 5386 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m11141 5277 5291 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.484e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m11142 1 5291 5277 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.484e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m11143 5291 5388 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m11144 1 5388 5291 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m11145 5387 5385 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.596e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.51 nrd=0.4 
m11146 1 4736 5389 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m11147 5390 5391 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m11148 5385 4736 5390 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m11149 5392 5389 5385 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m11150 1 4742 5392 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m11151 5391 4742 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m11152 0 5383 325 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.42e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.45 
m11153 5393 5277 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=7.37e-12 ad=1.506e-11 ps=1.097e-05 pd=1.425e-05 
+ nrs=0.13 nrd=0.26 
m11154 5383 5387 5393 0 nenh l=1.1e-06 w=6.4e-06 
+ as=8.77e-12 ad=6.21e-12 ps=9.49e-06 pd=9.23e-06 
+ nrs=0.21 nrd=0.15 
m11155 5394 5385 5383 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=7.67e-12 ps=7.3e-06 pd=8.31e-06 
+ nrs=0.15 nrd=0.24 
m11156 0 5291 5394 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m11157 5277 5291 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.254e-11 ad=1.506e-11 ps=1.09e-05 pd=1.425e-05 
+ nrs=0.22 nrd=0.26 
m11158 0 5291 5277 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.506e-11 ad=1.254e-11 ps=1.425e-05 pd=1.09e-05 
+ nrs=0.26 nrd=0.22 
m11159 5291 5388 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m11160 0 5388 5291 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m11161 5387 5385 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11162 5395 4736 5356 1 penh l=1.1e-06 w=1.44e-05 
+ as=1.224e-11 ad=4.04e-11 ps=1.61e-05 pd=3.49e-05 
+ nrs=0.06 nrd=0.19 
m11163 1 4742 5395 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.224e-11 ps=2.718e-05 pd=1.61e-05 
+ nrs=0.15 nrd=0.06 
m11164 5388 5396 1 1 penh l=1.1e-06 w=1.44e-05 
+ as=2.376e-11 ad=3.206e-11 ps=1.77e-05 pd=2.718e-05 
+ nrs=0.11 nrd=0.15 
m11165 1 5396 5388 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=2.376e-11 ps=2.718e-05 pd=1.77e-05 
+ nrs=0.15 nrd=0.11 
m11166 5396 5170 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.98e-11 ad=2.672e-11 ps=1.53e-05 pd=2.265e-05 
+ nrs=0.14 nrd=0.19 
m11167 5397 5262 5396 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.02e-11 ad=1.98e-11 ps=1.37e-05 pd=1.53e-05 
+ nrs=0.07 nrd=0.14 
m11168 1 5177 5397 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.02e-11 ps=2.265e-05 pd=1.37e-05 
+ nrs=0.19 nrd=0.07 
m11169 5358 4736 1 1 penh l=1.1e-06 w=1.28e-05 
+ as=1.264e-11 ad=2.85e-11 ps=1.53e-05 pd=2.416e-05 
+ nrs=0.08 nrd=0.17 
m11170 1 4742 5358 1 penh l=1.1e-06 w=1.28e-05 
+ as=2.85e-11 ad=1.264e-11 ps=2.416e-05 pd=1.53e-05 
+ nrs=0.17 nrd=0.08 
m11171 0 4736 5389 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.031e-11 ad=1.586e-11 ps=9.75e-06 pd=1.65e-05 
+ nrs=0.38 nrd=0.59 
m11172 5398 5391 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.32e-12 ad=1.348e-11 ps=9.63e-06 pd=1.275e-05 
+ nrs=0.14 nrd=0.29 
m11173 5385 5389 5398 0 nenh l=1.1e-06 w=5.2e-06 
+ as=8.58e-12 ad=4.84e-12 ps=8.5e-06 pd=7.37e-06 
+ nrs=0.32 nrd=0.18 
m11174 5399 4736 5385 0 nenh l=1.1e-06 w=5.2e-06 
+ as=4.56e-12 ad=8.58e-12 ps=7.37e-06 pd=8.5e-06 
+ nrs=0.17 nrd=0.32 
m11175 0 4742 5399 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.96e-12 ps=1.275e-05 pd=9.63e-06 
+ nrs=0.29 nrd=0.13 
m11176 5391 4742 0 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.031e-11 ps=1.65e-05 pd=9.75e-06 
+ nrs=0.59 nrd=0.38 
m11177 5356 4736 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=1.06e-11 ad=2.061e-11 ps=1.29e-05 pd=1.949e-05 
+ nrs=0.1 nrd=0.19 
m11178 0 4742 5356 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.061e-11 ad=1.06e-11 ps=1.949e-05 pd=1.29e-05 
+ nrs=0.19 nrd=0.1 
m11179 5388 5396 0 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.584e-11 ad=1.903e-11 ps=1.29e-05 pd=1.799e-05 
+ nrs=0.17 nrd=0.21 
m11180 0 5396 5388 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=1.584e-11 ps=1.799e-05 pd=1.29e-05 
+ nrs=0.21 nrd=0.17 
m11181 5400 5170 0 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.955e-11 ad=1.903e-11 ps=1.68e-05 pd=1.799e-05 
+ nrs=0.21 nrd=0.21 
m11182 5396 5262 5400 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.604e-11 ad=1.955e-11 ps=1.303e-05 pd=1.68e-05 
+ nrs=0.17 nrd=0.21 
m11183 5400 5177 5396 0 nenh l=1.1e-06 w=1e-05 
+ as=2.036e-11 ad=1.67e-11 ps=1.75e-05 pd=1.357e-05 
+ nrs=0.2 nrd=0.17 
m11184 5401 4736 5358 0 nenh l=1.1e-06 w=1.28e-05 
+ as=1.088e-11 ad=3.904e-11 ps=1.45e-05 pd=3.17e-05 
+ nrs=0.07 nrd=0.24 
m11185 0 4742 5401 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.088e-11 ps=2.399e-05 pd=1.45e-05 
+ nrs=0.15 nrd=0.07 
m11186 5402 5403 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=5.99e-12 ad=1.348e-11 ps=9.58e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m11187 528 5404 5402 0 nenh l=1.1e-06 w=6.4e-06 
+ as=7.52e-12 ad=5.63e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.14 
m11188 5405 5406 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m11189 5404 5407 5405 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m11190 5408 5409 5404 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m11191 0 5410 5408 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m11192 5406 5410 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11193 0 5412 5411 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m11194 5413 5407 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m11195 5414 5411 5413 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m11196 5415 5412 5414 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m11197 0 5409 5415 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m11198 5407 5409 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11199 5416 5414 528 0 nenh l=1.1e-06 w=6.4e-06 
+ as=5.63e-12 ad=7.52e-12 ps=9.02e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m11200 0 5417 5416 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.99e-12 ps=1.275e-05 pd=9.58e-06 
+ nrs=0.29 nrd=0.13 
m11201 5418 5403 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m11202 528 5414 5418 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m11203 5419 5404 528 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m11204 1 5417 5419 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m11205 5420 5406 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m11206 5404 5409 5420 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m11207 5421 5407 5404 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m11208 1 5410 5421 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m11209 5406 5410 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m11210 5422 5410 5423 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.745e-11 ps=1.429e-05 pd=2.077e-05 
+ nrs=0.11 nrd=0.13 
m11211 5424 5425 5422 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m11212 5423 5426 5424 0 nenh l=1.1e-06 w=1e-05 
+ as=1.505e-11 ad=8.5e-12 ps=1.791e-05 pd=1.17e-05 
+ nrs=0.15 nrd=0.08 
m11213 0 5426 5423 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.745e-11 ps=2.174e-05 pd=2.077e-05 
+ nrs=0.17 nrd=0.13 
m11214 5423 5425 0 0 nenh l=1.1e-06 w=1.08e-05 
+ as=1.625e-11 ad=2.141e-11 ps=1.934e-05 pd=2.024e-05 
+ nrs=0.14 nrd=0.18 
m11215 0 5425 5427 0 nenh l=1.1e-06 w=1.08e-05 
+ as=2.141e-11 ad=1.625e-11 ps=2.024e-05 pd=1.934e-05 
+ nrs=0.18 nrd=0.14 
m11216 5427 5426 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.745e-11 ad=2.299e-11 ps=2.077e-05 pd=2.174e-05 
+ nrs=0.13 nrd=0.17 
m11217 5428 5426 5427 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.505e-11 ps=1.17e-05 pd=1.791e-05 
+ nrs=0.08 nrd=0.15 
m11218 5429 5425 5428 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m11219 5427 5412 5429 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.745e-11 ad=1.416e-11 ps=2.077e-05 pd=1.429e-05 
+ nrs=0.13 nrd=0.11 
m11220 0 4623 5426 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m11221 5430 5426 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m11222 5409 5425 5430 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m11223 5431 4617 5409 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m11224 0 4623 5431 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m11225 5425 4617 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m11226 1 5412 5411 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m11227 5432 5407 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m11228 5414 5412 5432 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m11229 5433 5411 5414 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m11230 1 5409 5433 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m11231 5407 5409 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m11232 5422 5410 5434 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m11233 5435 5425 5422 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m11234 1 5426 5435 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m11235 5434 5426 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m11236 1 5425 5434 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m11237 5436 5425 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m11238 1 5426 5436 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m11239 5437 5426 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m11240 5429 5425 5437 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m11241 5436 5412 5429 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m11242 1 4623 5426 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m11243 5438 5426 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.45e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m11244 5409 4617 5438 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.033e-11 ad=7.53e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.11 
m11245 5439 5425 5409 1 penh l=1.1e-06 w=7.6e-06 
+ as=7.02e-12 ad=9.35e-12 ps=1.01e-05 pd=9.97e-06 
+ nrs=0.12 nrd=0.16 
m11246 1 4623 5439 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=8.12e-12 ps=1.661e-05 pd=1.17e-05 
+ nrs=0.25 nrd=0.1 
m11247 5425 4617 1 1 penh l=1.1e-06 w=1e-05 
+ as=3.05e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.31 nrd=0.22 
m11248 1 5440 499 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m11249 5441 5403 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m11250 5440 5442 5441 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m11251 5443 5444 5440 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m11252 1 5417 5443 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m11253 5445 5446 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m11254 5444 5447 5445 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m11255 5448 5449 5444 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m11256 1 5450 5448 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m11257 5446 5450 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m11258 1 5452 5451 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m11259 5453 5449 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m11260 5442 5452 5453 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m11261 5454 5451 5442 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m11262 1 5447 5454 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m11263 5449 5447 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m11264 0 5440 499 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.031e-11 ad=1.586e-11 ps=9.75e-06 pd=1.65e-05 
+ nrs=0.38 nrd=0.59 
m11265 5455 5403 0 0 nenh l=1.1e-06 w=7.2e-06 
+ as=6.43e-12 ad=1.427e-11 ps=1.058e-05 pd=1.35e-05 
+ nrs=0.12 nrd=0.28 
m11266 5440 5444 5455 0 nenh l=1.1e-06 w=6e-06 
+ as=8.27e-12 ad=5.35e-12 ps=9.11e-06 pd=8.82e-06 
+ nrs=0.23 nrd=0.15 
m11267 5456 5442 5440 0 nenh l=1.1e-06 w=5.2e-06 
+ as=4.53e-12 ad=7.17e-12 ps=7.26e-06 pd=7.89e-06 
+ nrs=0.17 nrd=0.27 
m11268 0 5417 5456 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=5.57e-12 ps=1.2e-05 pd=8.94e-06 
+ nrs=0.31 nrd=0.14 
m11269 1 4634 5457 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=2.196e-11 ps=1.359e-05 pd=2.05e-05 
+ nrs=0.31 nrd=0.42 
m11270 5458 5459 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.55e-12 ad=1.603e-11 ps=9.05e-06 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m11271 5447 4634 5458 1 penh l=1.1e-06 w=7.6e-06 
+ as=8.13e-12 ad=6.91e-12 ps=9.97e-06 pd=9.55e-06 
+ nrs=0.14 nrd=0.12 
m11272 5460 5457 5447 1 penh l=1.1e-06 w=8.4e-06 
+ as=8.56e-12 ad=8.99e-12 ps=1.088e-05 pd=1.103e-05 
+ nrs=0.12 nrd=0.13 
m11273 1 4640 5460 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=7.34e-12 ps=1.359e-05 pd=9.32e-06 
+ nrs=0.31 nrd=0.14 
m11274 5459 4640 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=2.196e-11 ad=1.603e-11 ps=2.05e-05 pd=1.359e-05 
+ nrs=0.42 nrd=0.31 
m11275 5461 5450 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.55e-11 ad=2.672e-11 ps=1.478e-05 pd=2.265e-05 
+ nrs=0.11 nrd=0.19 
m11276 5410 4634 5461 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.151e-11 ad=1.498e-11 ps=1.394e-05 pd=1.428e-05 
+ nrs=0.09 nrd=0.11 
m11277 5461 4640 5410 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.705e-11 ad=1.309e-11 ps=1.625e-05 pd=1.586e-05 
+ nrs=0.1 nrd=0.08 
m11278 5462 4640 5461 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.498e-11 ps=1.33e-05 pd=1.428e-05 
+ nrs=0.07 nrd=0.11 
m11279 1 4634 5462 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m11280 5463 4634 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m11281 5464 4640 5463 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=9.86e-12 ps=1.428e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m11282 5412 4640 5464 1 penh l=1.1e-06 w=1.32e-05 
+ as=1.309e-11 ad=1.705e-11 ps=1.586e-05 pd=1.625e-05 
+ nrs=0.08 nrd=0.1 
m11283 5464 4634 5412 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.498e-11 ad=1.151e-11 ps=1.428e-05 pd=1.394e-05 
+ nrs=0.11 nrd=0.09 
m11284 1 5452 5464 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.55e-11 ps=2.265e-05 pd=1.478e-05 
+ nrs=0.19 nrd=0.11 
m11285 5465 5446 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m11286 5444 5449 5465 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m11287 5466 5447 5444 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m11288 0 5450 5466 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m11289 5446 5450 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11290 0 5452 5451 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m11291 5467 5449 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m11292 5442 5451 5467 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m11293 5468 5452 5442 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m11294 0 5447 5468 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m11295 5449 5447 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11296 0 4634 5457 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m11297 5469 5459 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m11298 5447 5457 5469 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m11299 5470 4634 5447 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m11300 0 4640 5470 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m11301 5459 4640 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m11302 5410 5450 5471 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.175e-11 ad=1.755e-11 ps=1.429e-05 pd=1.841e-05 
+ nrs=0.09 nrd=0.13 
m11303 5472 4634 5410 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.013e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.1 
m11304 0 4640 5472 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=8.5e-12 ps=1.874e-05 pd=1.17e-05 
+ nrs=0.2 nrd=0.08 
m11305 5471 4640 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=2.299e-11 ps=1.841e-05 pd=2.174e-05 
+ nrs=0.13 nrd=0.17 
m11306 0 4634 5471 0 nenh l=1.1e-06 w=1e-05 
+ as=1.982e-11 ad=1.513e-11 ps=1.874e-05 pd=1.587e-05 
+ nrs=0.2 nrd=0.15 
m11307 5473 4634 0 0 nenh l=1.1e-06 w=1e-05 
+ as=1.513e-11 ad=1.982e-11 ps=1.587e-05 pd=1.874e-05 
+ nrs=0.15 nrd=0.2 
m11308 0 4640 5473 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.755e-11 ps=2.174e-05 pd=1.841e-05 
+ nrs=0.17 nrd=0.13 
m11309 5474 4640 0 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.982e-11 ps=1.17e-05 pd=1.874e-05 
+ nrs=0.08 nrd=0.2 
m11310 5412 4634 5474 0 nenh l=1.1e-06 w=1e-05 
+ as=1.013e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.1 nrd=0.08 
m11311 5473 5452 5412 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.755e-11 ad=1.175e-11 ps=1.841e-05 pd=1.429e-05 
+ nrs=0.13 nrd=0.09 
m11312 5475 5403 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.04e-12 ad=1.348e-11 ps=9.88e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m11313 470 5476 5475 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=5.33e-12 ps=8.5e-06 pd=8.72e-06 
+ nrs=0.19 nrd=0.15 
m11314 5477 5478 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m11315 5476 5479 5477 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m11316 5480 5481 5476 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m11317 0 5482 5480 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m11318 5478 5482 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11319 0 5484 5483 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m11320 5485 5479 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m11321 5486 5483 5485 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m11322 5487 5484 5486 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m11323 0 5481 5487 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m11324 5479 5481 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11325 5488 5486 470 0 nenh l=1.1e-06 w=6e-06 
+ as=5.29e-12 ad=6.86e-12 ps=8.61e-06 pd=8.5e-06 
+ nrs=0.15 nrd=0.19 
m11326 0 5417 5488 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=5.65e-12 ps=1.2e-05 pd=9.19e-06 
+ nrs=0.31 nrd=0.14 
m11327 5450 5482 5489 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.416e-11 ad=1.57e-11 ps=1.429e-05 pd=2.04e-05 
+ nrs=0.11 nrd=0.12 
m11328 5490 5491 5450 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.22e-11 ps=1.17e-05 pd=1.231e-05 
+ nrs=0.08 nrd=0.12 
m11329 5489 5492 5490 0 nenh l=1.1e-06 w=1e-05 
+ as=1.354e-11 ad=8.5e-12 ps=1.759e-05 pd=1.17e-05 
+ nrs=0.14 nrd=0.08 
m11330 0 5492 5489 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m11331 5489 5491 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m11332 0 5491 5493 0 nenh l=1.1e-06 w=1.16e-05 
+ as=2.299e-11 ad=1.57e-11 ps=2.174e-05 pd=2.04e-05 
+ nrs=0.17 nrd=0.12 
m11333 5493 5492 0 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=2.299e-11 ps=2.04e-05 pd=2.174e-05 
+ nrs=0.12 nrd=0.17 
m11334 5494 5492 5493 0 nenh l=1.1e-06 w=1e-05 
+ as=8.5e-12 ad=1.354e-11 ps=1.17e-05 pd=1.759e-05 
+ nrs=0.08 nrd=0.14 
m11335 5452 5491 5494 0 nenh l=1.1e-06 w=1e-05 
+ as=1.22e-11 ad=8.5e-12 ps=1.231e-05 pd=1.17e-05 
+ nrs=0.12 nrd=0.08 
m11336 5493 5484 5452 0 nenh l=1.1e-06 w=1.16e-05 
+ as=1.57e-11 ad=1.416e-11 ps=2.04e-05 pd=1.429e-05 
+ nrs=0.12 nrd=0.11 
m11337 0 4657 5492 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m11338 5495 5492 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m11339 5481 5491 5495 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m11340 5496 4651 5481 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m11341 0 4657 5496 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m11342 5491 4651 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m11343 5497 5403 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m11344 470 5486 5497 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m11345 5498 5476 470 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m11346 1 5417 5498 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m11347 5499 5478 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m11348 5476 5481 5499 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m11349 5500 5479 5476 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m11350 1 5482 5500 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m11351 5478 5482 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.308e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.42 nrd=0.4 
m11352 1 5484 5483 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m11353 5501 5479 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m11354 5486 5484 5501 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m11355 5502 5483 5486 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m11356 1 5481 5502 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m11357 5479 5481 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m11358 5450 5482 5503 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.569e-11 ad=1.453e-11 ps=1.515e-05 pd=1.849e-05 
+ nrs=0.11 nrd=0.1 
m11359 5504 5491 5450 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=1.517e-11 ps=1.33e-05 pd=1.465e-05 
+ nrs=0.07 nrd=0.11 
m11360 1 5492 5504 1 penh l=1.1e-06 w=1.16e-05 
+ as=2.583e-11 ad=9.86e-12 ps=2.19e-05 pd=1.33e-05 
+ nrs=0.19 nrd=0.07 
m11361 5503 5492 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m11362 1 5491 5503 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m11363 5505 5491 1 1 penh l=1.1e-06 w=1.24e-05 
+ as=1.501e-11 ad=2.761e-11 ps=1.911e-05 pd=2.341e-05 
+ nrs=0.1 nrd=0.18 
m11364 1 5492 5505 1 penh l=1.1e-06 w=1.24e-05 
+ as=2.761e-11 ad=1.501e-11 ps=2.341e-05 pd=1.911e-05 
+ nrs=0.18 nrd=0.1 
m11365 5506 5492 1 1 penh l=1.1e-06 w=1.16e-05 
+ as=9.86e-12 ad=2.583e-11 ps=1.33e-05 pd=2.19e-05 
+ nrs=0.07 nrd=0.19 
m11366 5452 5491 5506 1 penh l=1.1e-06 w=1.16e-05 
+ as=1.517e-11 ad=9.86e-12 ps=1.465e-05 pd=1.33e-05 
+ nrs=0.11 nrd=0.07 
m11367 5505 5484 5452 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.453e-11 ad=1.569e-11 ps=1.849e-05 pd=1.515e-05 
+ nrs=0.1 nrd=0.11 
m11368 1 4657 5492 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m11369 5507 5492 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.45e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m11370 5481 4651 5507 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.033e-11 ad=7.53e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.11 
m11371 5508 5491 5481 1 penh l=1.1e-06 w=7.6e-06 
+ as=7.02e-12 ad=9.35e-12 ps=1.01e-05 pd=9.97e-06 
+ nrs=0.12 nrd=0.16 
m11372 1 4657 5508 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=8.12e-12 ps=1.661e-05 pd=1.17e-05 
+ nrs=0.25 nrd=0.1 
m11373 5491 4651 1 1 penh l=1.1e-06 w=1e-05 
+ as=3.05e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.31 nrd=0.22 
m11374 1 5509 441 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m11375 5510 5403 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m11376 5509 5511 5510 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m11377 5512 5513 5509 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m11378 1 5417 5512 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m11379 5403 5417 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.484e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m11380 1 5417 5403 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.484e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m11381 5417 5514 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m11382 1 5514 5417 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m11383 5513 5511 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.596e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.51 nrd=0.4 
m11384 1 4668 5515 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m11385 5516 5517 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m11386 5511 4668 5516 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m11387 5518 5515 5511 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m11388 1 4674 5518 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m11389 5517 4674 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m11390 0 5509 441 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.42e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.45 
m11391 5519 5403 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=7.37e-12 ad=1.506e-11 ps=1.097e-05 pd=1.425e-05 
+ nrs=0.13 nrd=0.26 
m11392 5509 5513 5519 0 nenh l=1.1e-06 w=6.4e-06 
+ as=8.77e-12 ad=6.21e-12 ps=9.49e-06 pd=9.23e-06 
+ nrs=0.21 nrd=0.15 
m11393 5520 5511 5509 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=7.67e-12 ps=7.3e-06 pd=8.31e-06 
+ nrs=0.15 nrd=0.24 
m11394 0 5417 5520 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m11395 5403 5417 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.254e-11 ad=1.506e-11 ps=1.09e-05 pd=1.425e-05 
+ nrs=0.22 nrd=0.26 
m11396 0 5417 5403 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.506e-11 ad=1.254e-11 ps=1.425e-05 pd=1.09e-05 
+ nrs=0.26 nrd=0.22 
m11397 5417 5514 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m11398 0 5514 5417 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m11399 5513 5511 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11400 5521 4668 5482 1 penh l=1.1e-06 w=1.44e-05 
+ as=1.224e-11 ad=4.04e-11 ps=1.61e-05 pd=3.49e-05 
+ nrs=0.06 nrd=0.19 
m11401 1 4674 5521 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.224e-11 ps=2.718e-05 pd=1.61e-05 
+ nrs=0.15 nrd=0.06 
m11402 5514 5522 1 1 penh l=1.1e-06 w=1.44e-05 
+ as=2.376e-11 ad=3.206e-11 ps=1.77e-05 pd=2.718e-05 
+ nrs=0.11 nrd=0.15 
m11403 1 5522 5514 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=2.376e-11 ps=2.718e-05 pd=1.77e-05 
+ nrs=0.15 nrd=0.11 
m11404 5522 5296 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.98e-11 ad=2.672e-11 ps=1.53e-05 pd=2.265e-05 
+ nrs=0.14 nrd=0.19 
m11405 5523 5388 5522 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.02e-11 ad=1.98e-11 ps=1.37e-05 pd=1.53e-05 
+ nrs=0.07 nrd=0.14 
m11406 1 5303 5523 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.02e-11 ps=2.265e-05 pd=1.37e-05 
+ nrs=0.19 nrd=0.07 
m11407 5484 4668 1 1 penh l=1.1e-06 w=1.28e-05 
+ as=1.264e-11 ad=2.85e-11 ps=1.53e-05 pd=2.416e-05 
+ nrs=0.08 nrd=0.17 
m11408 1 4674 5484 1 penh l=1.1e-06 w=1.28e-05 
+ as=2.85e-11 ad=1.264e-11 ps=2.416e-05 pd=1.53e-05 
+ nrs=0.17 nrd=0.08 
m11409 0 4668 5515 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.031e-11 ad=1.586e-11 ps=9.75e-06 pd=1.65e-05 
+ nrs=0.38 nrd=0.59 
m11410 5524 5517 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.32e-12 ad=1.348e-11 ps=9.63e-06 pd=1.275e-05 
+ nrs=0.14 nrd=0.29 
m11411 5511 5515 5524 0 nenh l=1.1e-06 w=5.2e-06 
+ as=8.58e-12 ad=4.84e-12 ps=8.5e-06 pd=7.37e-06 
+ nrs=0.32 nrd=0.18 
m11412 5525 4668 5511 0 nenh l=1.1e-06 w=5.2e-06 
+ as=4.56e-12 ad=8.58e-12 ps=7.37e-06 pd=8.5e-06 
+ nrs=0.17 nrd=0.32 
m11413 0 4674 5525 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.96e-12 ps=1.275e-05 pd=9.63e-06 
+ nrs=0.29 nrd=0.13 
m11414 5517 4674 0 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.031e-11 ps=1.65e-05 pd=9.75e-06 
+ nrs=0.59 nrd=0.38 
m11415 5482 4668 0 0 nenh l=1.1e-06 w=1.04e-05 
+ as=1.06e-11 ad=2.061e-11 ps=1.29e-05 pd=1.949e-05 
+ nrs=0.1 nrd=0.19 
m11416 0 4674 5482 0 nenh l=1.1e-06 w=1.04e-05 
+ as=2.061e-11 ad=1.06e-11 ps=1.949e-05 pd=1.29e-05 
+ nrs=0.19 nrd=0.1 
m11417 5514 5522 0 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.584e-11 ad=1.903e-11 ps=1.29e-05 pd=1.799e-05 
+ nrs=0.17 nrd=0.21 
m11418 0 5522 5514 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.903e-11 ad=1.584e-11 ps=1.799e-05 pd=1.29e-05 
+ nrs=0.21 nrd=0.17 
m11419 5526 5296 0 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.955e-11 ad=1.903e-11 ps=1.68e-05 pd=1.799e-05 
+ nrs=0.21 nrd=0.21 
m11420 5522 5388 5526 0 nenh l=1.1e-06 w=9.6e-06 
+ as=1.604e-11 ad=1.955e-11 ps=1.303e-05 pd=1.68e-05 
+ nrs=0.17 nrd=0.21 
m11421 5526 5303 5522 0 nenh l=1.1e-06 w=1e-05 
+ as=2.036e-11 ad=1.67e-11 ps=1.75e-05 pd=1.357e-05 
+ nrs=0.2 nrd=0.17 
m11422 5527 4668 5484 0 nenh l=1.1e-06 w=1.28e-05 
+ as=1.088e-11 ad=3.904e-11 ps=1.45e-05 pd=3.17e-05 
+ nrs=0.07 nrd=0.24 
m11423 0 4674 5527 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.088e-11 ps=2.399e-05 pd=1.45e-05 
+ nrs=0.15 nrd=0.07 
m11424 5528 5529 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.04e-12 ad=1.348e-11 ps=9.88e-06 pd=1.275e-05 
+ nrs=0.13 nrd=0.29 
m11425 584 5530 5528 0 nenh l=1.1e-06 w=6e-06 
+ as=6.86e-12 ad=5.33e-12 ps=8.5e-06 pd=8.72e-06 
+ nrs=0.19 nrd=0.15 
m11426 5531 5532 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m11427 5530 5533 5531 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m11428 5534 5535 5530 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m11429 0 5536 5534 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m11430 5532 5536 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11431 0 5538 5537 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m11432 5539 5533 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=5.55e-12 ps=4.5e-06 pd=5.25e-06 
+ nrs=0.3 nrd=0.71 
m11433 5540 5537 5539 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=2.38e-12 ps=6.1e-06 pd=4.5e-06 
+ nrs=0.59 nrd=0.3 
m11434 5541 5538 5540 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.38e-12 ad=4.62e-12 ps=4.5e-06 pd=6.1e-06 
+ nrs=0.3 nrd=0.59 
m11435 0 5535 5541 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=2.38e-12 ps=5.25e-06 pd=4.5e-06 
+ nrs=0.71 nrd=0.3 
m11436 5533 5535 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11437 5542 5540 584 0 nenh l=1.1e-06 w=6e-06 
+ as=5.29e-12 ad=6.86e-12 ps=8.61e-06 pd=8.5e-06 
+ nrs=0.15 nrd=0.19 
m11438 0 5543 5542 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=5.65e-12 ps=1.2e-05 pd=9.19e-06 
+ nrs=0.31 nrd=0.14 
m11439 0 4589 5544 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.708e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.54 
m11440 5545 5544 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.11e-11 ps=7.3e-06 pd=1.05e-05 
+ nrs=0.15 nrd=0.35 
m11441 5535 5546 5545 0 nenh l=1.1e-06 w=5.6e-06 
+ as=9.24e-12 ad=4.76e-12 ps=8.9e-06 pd=7.3e-06 
+ nrs=0.29 nrd=0.15 
m11442 5547 4569 5535 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=9.24e-12 ps=7.3e-06 pd=8.9e-06 
+ nrs=0.15 nrd=0.29 
m11443 0 4589 5547 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m11444 5546 4569 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.11e-11 ps=1.73e-05 pd=1.05e-05 
+ nrs=0.54 nrd=0.35 
m11445 5548 5529 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m11446 584 5540 5548 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m11447 5549 5530 584 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m11448 1 5543 5549 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m11449 5550 5532 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.77e-12 ad=1.603e-11 ps=1.015e-05 pd=1.359e-05 
+ nrs=0.13 nrd=0.31 
m11450 5530 5535 5550 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.65e-12 ps=8.34e-06 pd=8.45e-06 
+ nrs=0.19 nrd=0.16 
m11451 5551 5533 5530 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.6e-12 ad=7.65e-12 ps=9.81e-06 pd=9.46e-06 
+ nrs=0.14 nrd=0.17 
m11452 1 5536 5551 1 penh l=1.1e-06 w=7.2e-06 
+ as=1.603e-11 ad=6.98e-12 ps=1.359e-05 pd=1.039e-05 
+ nrs=0.31 nrd=0.13 
m11453 5532 5536 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.308e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.42 nrd=0.4 
m11454 1 5538 5537 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m11455 5552 5533 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.88e-12 ad=1.247e-11 ps=7.43e-06 pd=1.057e-05 
+ nrs=0.16 nrd=0.4 
m11456 5540 5538 5552 1 penh l=1.1e-06 w=6e-06 
+ as=6.75e-12 ad=5.22e-12 ps=8.34e-06 pd=7.97e-06 
+ nrs=0.19 nrd=0.15 
m11457 5553 5537 5540 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.17e-12 ad=7.65e-12 ps=9.32e-06 pd=9.46e-06 
+ nrs=0.13 nrd=0.17 
m11458 1 5535 5553 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=5.09e-12 ps=1.057e-05 pd=7.68e-06 
+ nrs=0.4 nrd=0.16 
m11459 5533 5535 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.708e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.54 nrd=0.4 
m11460 1 4589 5544 1 penh l=1.1e-06 w=1e-05 
+ as=2.227e-11 ad=3.05e-11 ps=1.888e-05 pd=2.61e-05 
+ nrs=0.22 nrd=0.31 
m11461 5554 5544 1 1 penh l=1.1e-06 w=7.2e-06 
+ as=6.45e-12 ad=1.603e-11 ps=9.32e-06 pd=1.359e-05 
+ nrs=0.12 nrd=0.31 
m11462 5535 4569 5554 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.033e-11 ad=7.53e-12 ps=1.103e-05 pd=1.088e-05 
+ nrs=0.15 nrd=0.11 
m11463 5555 5546 5535 1 penh l=1.1e-06 w=7.6e-06 
+ as=7.02e-12 ad=9.35e-12 ps=1.01e-05 pd=9.97e-06 
+ nrs=0.12 nrd=0.16 
m11464 1 4589 5555 1 penh l=1.1e-06 w=8.8e-06 
+ as=1.959e-11 ad=8.12e-12 ps=1.661e-05 pd=1.17e-05 
+ nrs=0.25 nrd=0.1 
m11465 5546 4569 1 1 penh l=1.1e-06 w=1e-05 
+ as=3.05e-11 ad=2.227e-11 ps=2.61e-05 pd=1.888e-05 
+ nrs=0.31 nrd=0.22 
m11466 1 5556 556 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.708e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.54 
m11467 5557 5529 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6.4e-12 ad=1.514e-11 ps=9.58e-06 pd=1.284e-05 
+ nrs=0.14 nrd=0.33 
m11468 5556 5558 5557 1 penh l=1.1e-06 w=6.4e-06 
+ as=7.2e-12 ad=6.02e-12 ps=8.9e-06 pd=9.02e-06 
+ nrs=0.18 nrd=0.15 
m11469 5559 5560 5556 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.7e-12 ad=7.2e-12 ps=8.64e-06 pd=8.9e-06 
+ nrs=0.14 nrd=0.18 
m11470 1 5543 5559 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=4.98e-12 ps=1.057e-05 pd=7.56e-06 
+ nrs=0.4 nrd=0.16 
m11471 5529 5543 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.484e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m11472 1 5543 5529 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.484e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m11473 5543 5561 1 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.42e-11 ad=2.672e-11 ps=1.45e-05 pd=2.265e-05 
+ nrs=0.1 nrd=0.19 
m11474 1 5561 5543 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.42e-11 ps=2.265e-05 pd=1.45e-05 
+ nrs=0.19 nrd=0.1 
m11475 5560 5558 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.596e-11 ad=1.247e-11 ps=1.73e-05 pd=1.057e-05 
+ nrs=0.51 nrd=0.4 
m11476 1 4600 5562 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.158e-11 ad=1.586e-11 ps=9.82e-06 pd=1.65e-05 
+ nrs=0.43 nrd=0.59 
m11477 5563 5564 1 1 penh l=1.1e-06 w=6.8e-06 
+ as=6e-12 ad=1.514e-11 ps=9.76e-06 pd=1.284e-05 
+ nrs=0.13 nrd=0.33 
m11478 5558 4600 5563 1 penh l=1.1e-06 w=5.6e-06 
+ as=6.4e-12 ad=4.94e-12 ps=7.93e-06 pd=8.04e-06 
+ nrs=0.2 nrd=0.16 
m11479 5565 5562 5558 1 penh l=1.1e-06 w=6.4e-06 
+ as=5.71e-12 ad=7.32e-12 ps=9.41e-06 pd=9.07e-06 
+ nrs=0.14 nrd=0.18 
m11480 1 4606 5565 1 penh l=1.1e-06 w=6.8e-06 
+ as=1.514e-11 ad=6.07e-12 ps=1.284e-05 pd=9.99e-06 
+ nrs=0.33 nrd=0.13 
m11481 5564 4606 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.59 nrd=0.43 
m11482 0 5556 556 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=1.42e-11 ps=1.05e-05 pd=1.73e-05 
+ nrs=0.35 nrd=0.45 
m11483 5566 5529 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=7.37e-12 ad=1.506e-11 ps=1.097e-05 pd=1.425e-05 
+ nrs=0.13 nrd=0.26 
m11484 5556 5560 5566 0 nenh l=1.1e-06 w=6.4e-06 
+ as=8.77e-12 ad=6.21e-12 ps=9.49e-06 pd=9.23e-06 
+ nrs=0.21 nrd=0.15 
m11485 5567 5558 5556 0 nenh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=7.67e-12 ps=7.3e-06 pd=8.31e-06 
+ nrs=0.15 nrd=0.24 
m11486 0 5543 5567 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.11e-11 ad=4.76e-12 ps=1.05e-05 pd=7.3e-06 
+ nrs=0.35 nrd=0.15 
m11487 5529 5543 0 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.254e-11 ad=1.506e-11 ps=1.09e-05 pd=1.425e-05 
+ nrs=0.22 nrd=0.26 
m11488 0 5543 5529 0 nenh l=1.1e-06 w=7.6e-06 
+ as=1.506e-11 ad=1.254e-11 ps=1.425e-05 pd=1.09e-05 
+ nrs=0.26 nrd=0.22 
m11489 5543 5561 0 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.386e-11 ad=1.665e-11 ps=1.17e-05 pd=1.575e-05 
+ nrs=0.2 nrd=0.24 
m11490 0 5561 5543 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.665e-11 ad=1.386e-11 ps=1.575e-05 pd=1.17e-05 
+ nrs=0.24 nrd=0.2 
m11491 5560 5558 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.54e-12 ad=5.55e-12 ps=1.17e-05 pd=5.25e-06 
+ nrs=1.09 nrd=0.71 
m11492 5568 4600 5536 1 penh l=1.1e-06 w=1.28e-05 
+ as=1.088e-11 ad=3.68e-11 ps=1.45e-05 pd=3.17e-05 
+ nrs=0.07 nrd=0.22 
m11493 1 4606 5568 1 penh l=1.1e-06 w=1.28e-05 
+ as=2.85e-11 ad=1.088e-11 ps=2.416e-05 pd=1.45e-05 
+ nrs=0.17 nrd=0.07 
m11494 5561 5569 1 1 penh l=1.1e-06 w=1.28e-05 
+ as=2.112e-11 ad=2.85e-11 ps=1.61e-05 pd=2.416e-05 
+ nrs=0.13 nrd=0.17 
m11495 1 5569 5561 1 penh l=1.1e-06 w=1.28e-05 
+ as=2.85e-11 ad=2.112e-11 ps=2.416e-05 pd=1.61e-05 
+ nrs=0.17 nrd=0.13 
m11496 5569 5422 1 1 penh l=1.1e-06 w=1.04e-05 
+ as=1.716e-11 ad=2.316e-11 ps=1.37e-05 pd=1.963e-05 
+ nrs=0.16 nrd=0.21 
m11497 5570 5514 5569 1 penh l=1.1e-06 w=1.04e-05 
+ as=8.84e-12 ad=1.716e-11 ps=1.21e-05 pd=1.37e-05 
+ nrs=0.08 nrd=0.16 
m11498 1 5429 5570 1 penh l=1.1e-06 w=1.04e-05 
+ as=2.316e-11 ad=8.84e-12 ps=1.963e-05 pd=1.21e-05 
+ nrs=0.21 nrd=0.08 
m11499 5538 4600 1 1 penh l=1.1e-06 w=1.12e-05 
+ as=1.128e-11 ad=2.494e-11 ps=1.37e-05 pd=2.114e-05 
+ nrs=0.09 nrd=0.2 
m11500 1 4606 5538 1 penh l=1.1e-06 w=1.12e-05 
+ as=2.494e-11 ad=1.128e-11 ps=2.114e-05 pd=1.37e-05 
+ nrs=0.2 nrd=0.09 
m11501 0 4600 5562 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.031e-11 ad=1.586e-11 ps=9.75e-06 pd=1.65e-05 
+ nrs=0.38 nrd=0.59 
m11502 5571 5564 0 0 nenh l=1.1e-06 w=6.8e-06 
+ as=6.32e-12 ad=1.348e-11 ps=9.63e-06 pd=1.275e-05 
+ nrs=0.14 nrd=0.29 
m11503 5558 5562 5571 0 nenh l=1.1e-06 w=5.2e-06 
+ as=8.58e-12 ad=4.84e-12 ps=8.5e-06 pd=7.37e-06 
+ nrs=0.32 nrd=0.18 
m11504 5572 4600 5558 0 nenh l=1.1e-06 w=5.2e-06 
+ as=4.56e-12 ad=8.58e-12 ps=7.37e-06 pd=8.5e-06 
+ nrs=0.17 nrd=0.32 
m11505 0 4606 5572 0 nenh l=1.1e-06 w=6.8e-06 
+ as=1.348e-11 ad=5.96e-12 ps=1.275e-05 pd=9.63e-06 
+ nrs=0.29 nrd=0.13 
m11506 5564 4606 0 0 nenh l=1.1e-06 w=5.2e-06 
+ as=1.586e-11 ad=1.031e-11 ps=1.65e-05 pd=9.75e-06 
+ nrs=0.59 nrd=0.38 
m11507 5536 4600 0 0 nenh l=1.1e-06 w=8.8e-06 
+ as=9.24e-12 ad=1.744e-11 ps=1.13e-05 pd=1.65e-05 
+ nrs=0.12 nrd=0.23 
m11508 0 4606 5536 0 nenh l=1.1e-06 w=8.8e-06 
+ as=1.744e-11 ad=9.24e-12 ps=1.65e-05 pd=1.13e-05 
+ nrs=0.23 nrd=0.12 
m11509 5561 5569 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.32e-11 ad=1.586e-11 ps=1.13e-05 pd=1.5e-05 
+ nrs=0.21 nrd=0.25 
m11510 0 5569 5561 0 nenh l=1.1e-06 w=8e-06 
+ as=1.586e-11 ad=1.32e-11 ps=1.5e-05 pd=1.13e-05 
+ nrs=0.25 nrd=0.21 
m11511 5573 5422 0 0 nenh l=1.1e-06 w=8e-06 
+ as=1.616e-11 ad=1.586e-11 ps=1.466e-05 pd=1.5e-05 
+ nrs=0.25 nrd=0.25 
m11512 5569 5514 5573 0 nenh l=1.1e-06 w=8e-06 
+ as=1.34e-11 ad=1.616e-11 ps=1.141e-05 pd=1.466e-05 
+ nrs=0.21 nrd=0.25 
m11513 5573 5429 5569 0 nenh l=1.1e-06 w=8.4e-06 
+ as=1.697e-11 ad=1.406e-11 ps=1.539e-05 pd=1.199e-05 
+ nrs=0.24 nrd=0.2 
m11514 5574 4600 5538 0 nenh l=1.1e-06 w=1.12e-05 
+ as=9.52e-12 ad=3.416e-11 ps=1.29e-05 pd=2.85e-05 
+ nrs=0.08 nrd=0.27 
m11515 0 4606 5574 0 nenh l=1.1e-06 w=1.12e-05 
+ as=2.22e-11 ad=9.52e-12 ps=2.099e-05 pd=1.29e-05 
+ nrs=0.18 nrd=0.08 
m11516 0 5575 4923 0 nenh l=1.1e-06 w=1.44e-05 
+ as=2.854e-11 ad=3.144e-11 ps=2.699e-05 pd=3.25e-05 
+ nrs=0.14 nrd=0.15 
m11517 5576 5577 0 0 nenh l=1.1e-06 w=1.52e-05 
+ as=2.083e-11 ad=3.013e-11 ps=2.27e-05 pd=2.849e-05 
+ nrs=0.09 nrd=0.13 
m11518 0 4514 5576 0 nenh l=1.1e-06 w=1.52e-05 
+ as=3.013e-11 ad=2.083e-11 ps=2.849e-05 pd=2.27e-05 
+ nrs=0.13 nrd=0.09 
m11519 5578 5577 0 0 nenh l=1.1e-06 w=1.64e-05 
+ as=1.415e-11 ad=3.25e-11 ps=1.928e-05 pd=3.074e-05 
+ nrs=0.05 nrd=0.12 
m11520 5575 4514 5578 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.423e-11 ad=1.243e-11 ps=1.795e-05 pd=1.692e-05 
+ nrs=0.07 nrd=0.06 
m11521 5576 4520 5575 0 nenh l=1.1e-06 w=1.4e-05 
+ as=1.919e-11 ad=1.383e-11 ps=2.091e-05 pd=1.745e-05 
+ nrs=0.1 nrd=0.07 
m11522 5579 4520 0 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.352e-11 ad=2.854e-11 ps=1.61e-05 pd=2.699e-05 
+ nrs=0.07 nrd=0.14 
m11523 5580 5575 5579 0 nenh l=1.1e-06 w=1.44e-05 
+ as=1.449e-11 ad=1.352e-11 ps=1.785e-05 pd=1.61e-05 
+ nrs=0.07 nrd=0.07 
m11524 5581 4514 5580 0 nenh l=1.1e-06 w=1.48e-05 
+ as=1.27e-11 ad=1.489e-11 ps=1.701e-05 pd=1.835e-05 
+ nrs=0.06 nrd=0.07 
m11525 5582 4520 5581 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.372e-11 ad=1.372e-11 ps=1.822e-05 pd=1.839e-05 
+ nrs=0.05 nrd=0.05 
m11526 0 5577 5582 0 nenh l=1.1e-06 w=1.72e-05 
+ as=3.409e-11 ad=1.474e-11 ps=3.224e-05 pd=1.958e-05 
+ nrs=0.12 nrd=0.05 
m11527 5579 4514 0 0 nenh l=1.1e-06 w=1.6e-05 
+ as=1.502e-11 ad=3.171e-11 ps=1.789e-05 pd=2.999e-05 
+ nrs=0.06 nrd=0.12 
m11528 0 5577 5579 0 nenh l=1.1e-06 w=1.28e-05 
+ as=2.537e-11 ad=1.202e-11 ps=2.399e-05 pd=1.431e-05 
+ nrs=0.15 nrd=0.07 
m11529 1 5575 4923 1 penh l=1.1e-06 w=1.8e-05 
+ as=4.008e-11 ad=3.314e-11 ps=3.398e-05 pd=3.89e-05 
+ nrs=0.12 nrd=0.1 
m11530 4950 5580 0 0 nenh l=1.1e-06 w=2.24e-05 
+ as=3.312e-11 ad=4.44e-11 ps=4.45e-05 pd=4.199e-05 
+ nrs=0.07 nrd=0.09 
m11531 5583 5577 1 1 penh l=1.1e-06 w=1.8e-05 
+ as=1.542e-11 ad=4.008e-11 ps=2.038e-05 pd=3.398e-05 
+ nrs=0.05 nrd=0.12 
m11532 5584 4514 5583 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.692e-11 ad=1.44e-11 ps=1.967e-05 pd=1.902e-05 
+ nrs=0.06 nrd=0.05 
m11533 5575 5577 5584 1 penh l=1.1e-06 w=1.68e-05 
+ as=1.615e-11 ad=1.692e-11 ps=1.96e-05 pd=1.967e-05 
+ nrs=0.06 nrd=0.06 
m11534 5584 4514 5575 1 penh l=1.1e-06 w=1.56e-05 
+ as=1.571e-11 ad=1.499e-11 ps=1.827e-05 pd=1.82e-05 
+ nrs=0.06 nrd=0.06 
m11535 1 4520 5584 1 penh l=1.1e-06 w=1.4e-05 
+ as=3.117e-11 ad=1.41e-11 ps=2.643e-05 pd=1.639e-05 
+ nrs=0.16 nrd=0.07 
m11536 1 5585 4954 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.247e-11 ad=1.484e-11 ps=1.057e-05 pd=1.73e-05 
+ nrs=0.4 nrd=0.47 
m11537 5586 4582 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=4.76e-12 ad=1.247e-11 ps=7.3e-06 pd=1.057e-05 
+ nrs=0.15 nrd=0.4 
m11538 5585 4563 5586 1 penh l=1.1e-06 w=5.6e-06 
+ as=1.372e-11 ad=4.76e-12 ps=1.73e-05 pd=7.3e-06 
+ nrs=0.44 nrd=0.15 
m11539 1 5587 5577 1 penh l=1.1e-06 w=8.4e-06 
+ as=1.87e-11 ad=1.89e-11 ps=1.586e-05 pd=2.29e-05 
+ nrs=0.27 nrd=0.27 
m11540 5580 5575 5588 1 penh l=1.1e-06 w=1.2e-05 
+ as=1.447e-11 ad=1.386e-11 ps=1.722e-05 pd=1.719e-05 
+ nrs=0.1 nrd=0.1 
m11541 5589 4514 5580 1 penh l=1.1e-06 w=1.88e-05 
+ as=1.621e-11 ad=2.267e-11 ps=2.153e-05 pd=2.698e-05 
+ nrs=0.05 nrd=0.06 
m11542 5590 4520 5589 1 penh l=1.1e-06 w=2.12e-05 
+ as=1.814e-11 ad=1.827e-11 ps=2.344e-05 pd=2.427e-05 
+ nrs=0.04 nrd=0.04 
m11543 5588 5577 5590 1 penh l=1.1e-06 w=2.24e-05 
+ as=2.588e-11 ad=1.916e-11 ps=3.21e-05 pd=2.476e-05 
+ nrs=0.05 nrd=0.04 
m11544 1 4514 5588 1 penh l=1.1e-06 w=1.44e-05 
+ as=3.206e-11 ad=1.664e-11 ps=2.718e-05 pd=2.063e-05 
+ nrs=0.15 nrd=0.08 
m11545 5588 5577 1 1 penh l=1.1e-06 w=1.52e-05 
+ as=1.756e-11 ad=3.384e-11 ps=2.178e-05 pd=2.869e-05 
+ nrs=0.08 nrd=0.15 
m11546 1 4520 5588 1 penh l=1.1e-06 w=1.2e-05 
+ as=2.672e-11 ad=1.386e-11 ps=2.265e-05 pd=1.719e-05 
+ nrs=0.19 nrd=0.1 
m11547 5587 5591 1 1 penh l=1.1e-06 w=5.2e-06 
+ as=1.202e-11 ad=1.158e-11 ps=1.65e-05 pd=9.82e-06 
+ nrs=0.44 nrd=0.43 
m11548 4950 5580 1 1 penh l=1.1e-06 w=2.2e-05 
+ as=3.446e-11 ad=4.898e-11 ps=4.69e-05 pd=4.153e-05 
+ nrs=0.07 nrd=0.1 
m11549 0 5585 4954 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=8.54e-12 ps=5.25e-06 pd=1.17e-05 
+ nrs=0.71 nrd=1.09 
m11550 5585 4582 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=4.62e-12 ad=5.55e-12 ps=6.1e-06 pd=5.25e-06 
+ nrs=0.59 nrd=0.71 
m11551 0 4563 5585 0 nenh l=1.1e-06 w=2.8e-06 
+ as=5.55e-12 ad=4.62e-12 ps=5.25e-06 pd=6.1e-06 
+ nrs=0.71 nrd=0.59 
m11552 0 5587 5577 0 nenh l=1.1e-06 w=6.4e-06 
+ as=1.268e-11 ad=1.52e-11 ps=1.2e-05 pd=1.89e-05 
+ nrs=0.31 nrd=0.37 
m11553 0 5591 5587 0 nenh l=1.1e-06 w=6e-06 
+ as=1.189e-11 ad=1.446e-11 ps=1.125e-05 pd=1.81e-05 
+ nrs=0.33 nrd=0.4 
m11554 0 4567 5591 0 nenh l=1.1e-06 w=3.2e-06 
+ as=6.34e-12 ad=6.09e-12 ps=6e-06 pd=7.29e-06 
+ nrs=0.62 nrd=0.6 
m11555 5591 4582 1 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.098e-11 ps=8.2e-06 pd=1.406e-05 
+ nrs=0.53 nrd=0.85 
m11556 0 4571 5591 0 nenh l=1.1e-06 w=3.6e-06 
+ as=7.14e-12 ad=6.86e-12 ps=6.75e-06 pd=8.2e-06 
+ nrs=0.55 nrd=0.53 
m11557 5591 4580 858 0 nenh l=1.1e-06 w=3.6e-06 
+ as=6.86e-12 ad=1.036e-11 ps=8.2e-06 pd=1.246e-05 
+ nrs=0.53 nrd=0.8 
m11558 852 4563 5591 0 nenh l=1.1e-06 w=3.6e-06 
+ as=1.003e-11 ad=6.86e-12 ps=1.202e-05 pd=8.2e-06 
+ nrs=0.77 nrd=0.53 
c0 4571 0 3.14973e-13
c1 5585 0 7.46e-15
c2 5588 0 1.984e-15
c3 5584 0 8.1e-16
c4 5538 0 3.7244e-14
c5 5573 0 7.58e-16
c6 5536 0 2.3203e-14
c7 5562 0 1.354e-14
c8 5564 0 1.4292e-14
c9 5558 0 2.7971e-14
c10 5560 0 1.8387e-14
c11 5546 0 1.2507e-14
c12 5544 0 1.2867e-14
c13 5537 0 1.2546e-14
c14 5533 0 2.061e-14
c15 5532 0 1.346e-14
c16 5540 0 2.019e-14
c17 5530 0 1.5093e-14
c18 5515 0 1.354e-14
c19 5517 0 1.4292e-14
c20 5511 0 2.7971e-14
c21 5513 0 1.8387e-14
c22 5505 0 1.356e-15
c23 5503 0 1.31e-15
c24 5483 0 1.2892e-14
c25 5479 0 2.1812e-14
c26 5478 0 1.346e-14
c27 5486 0 2.0361e-14
c28 5476 0 1.5093e-14
c29 5451 0 1.4445e-14
c30 5449 0 2.3269e-14
c31 5446 0 1.4818e-14
c32 5442 0 2.5005e-14
c33 5444 0 1.4174e-14
c34 5440 0 1.2715e-14
c35 5464 0 5.74e-16
c36 5461 0 5.74e-16
c37 5436 0 1.356e-15
c38 5434 0 1.31e-15
c39 5411 0 1.292e-14
c40 5407 0 2.2234e-14
c41 5406 0 1.3439e-14
c42 5414 0 2.0225e-14
c43 5404 0 1.2854e-14
c44 5389 0 1.354e-14
c45 5391 0 1.4292e-14
c46 5385 0 2.7971e-14
c47 5387 0 1.8387e-14
c48 5379 0 1.356e-15
c49 5377 0 1.31e-15
c50 5357 0 1.2892e-14
c51 5353 0 2.1812e-14
c52 5352 0 1.346e-14
c53 5360 0 2.0361e-14
c54 5350 0 1.5093e-14
c55 5325 0 1.4445e-14
c56 5323 0 2.3269e-14
c57 5320 0 1.4818e-14
c58 5316 0 2.5005e-14
c59 5318 0 1.4174e-14
c60 5314 0 1.2715e-14
c61 5338 0 5.74e-16
c62 5335 0 5.74e-16
c63 5310 0 1.356e-15
c64 5308 0 1.31e-15
c65 5285 0 1.292e-14
c66 5281 0 2.2234e-14
c67 5280 0 1.3439e-14
c68 5288 0 2.0225e-14
c69 5278 0 1.2854e-14
c70 5263 0 1.354e-14
c71 5265 0 1.4292e-14
c72 5259 0 2.7971e-14
c73 5261 0 1.8387e-14
c74 5253 0 1.356e-15
c75 5251 0 1.31e-15
c76 5231 0 1.2892e-14
c77 5227 0 2.1812e-14
c78 5226 0 1.346e-14
c79 5234 0 2.0361e-14
c80 5224 0 1.5093e-14
c81 5199 0 1.4445e-14
c82 5197 0 2.3269e-14
c83 5194 0 1.4818e-14
c84 5190 0 2.5005e-14
c85 5192 0 1.4174e-14
c86 5188 0 1.2715e-14
c87 5212 0 5.74e-16
c88 5209 0 5.74e-16
c89 5184 0 1.356e-15
c90 5182 0 1.31e-15
c91 5159 0 1.292e-14
c92 5155 0 2.2234e-14
c93 5154 0 1.3439e-14
c94 5162 0 2.0225e-14
c95 5152 0 1.2854e-14
c96 5137 0 1.354e-14
c97 5139 0 1.4292e-14
c98 5133 0 2.7971e-14
c99 5135 0 1.8387e-14
c100 5127 0 1.356e-15
c101 5125 0 1.31e-15
c102 5105 0 1.2892e-14
c103 5101 0 2.1812e-14
c104 5100 0 1.346e-14
c105 5108 0 2.0361e-14
c106 5098 0 1.4841e-14
c107 5073 0 1.4445e-14
c108 5071 0 2.3269e-14
c109 5068 0 1.4818e-14
c110 5064 0 2.4782e-14
c111 5066 0 1.4031e-14
c112 5062 0 1.2661e-14
c113 5086 0 5.74e-16
c114 5083 0 5.74e-16
c115 5058 0 1.356e-15
c116 5056 0 1.31e-15
c117 5033 0 1.292e-14
c118 5029 0 2.2234e-14
c119 5028 0 1.3439e-14
c120 5036 0 2.0225e-14
c121 5026 0 1.2854e-14
c122 4549 0 2.7482e-14
c123 4980 0 3.9197e-14
c124 5018 0 1.1959e-14
c125 5022 0 7.58e-16
c126 5011 0 1.2441e-14
c127 5013 0 1.2627e-14
c128 4978 0 2.8569e-14
c129 5007 0 2.8206e-14
c130 5009 0 1.8429e-14
c131 5005 0 1.3439e-14
c132 4991 0 3.5449e-14
c133 4992 0 2.7179e-14
c134 4977 0 3.7753e-14
c135 5001 0 1.356e-15
c136 4999 0 1.31e-15
c137 4979 0 1.2712e-14
c138 4975 0 2.233e-14
c139 4974 0 1.348e-14
c140 4982 0 2.1059e-14
c141 4972 0 1.4886e-14
c142 4905 0 3.795e-14
c143 4949 0 1.4239e-14
c144 4952 0 1.5303e-14
c145 4903 0 2.8534e-14
c146 4941 0 3.1837e-14
c147 4945 0 1.4719e-14
c148 4943 0 2.349e-14
c149 4940 0 1.4618e-14
c150 4936 0 2.374e-14
c151 4938 0 1.4447e-14
c152 4934 0 1.3211e-14
c153 4960 0 5.74e-16
c154 4957 0 5.74e-16
c155 4918 0 3.5676e-14
c156 4919 0 2.6686e-14
c157 4902 0 3.8301e-14
c158 4930 0 1.356e-15
c159 4928 0 1.31e-15
c160 4904 0 1.3057e-14
c161 4900 0 2.3069e-14
c162 4899 0 1.3038e-14
c163 4907 0 2.151e-14
c164 4897 0 1.3101e-14
c165 4894 0 1.1019e-14
c166 4893 0 1.0554e-14
c167 4890 0 2.606e-15
c168 4888 0 1.225e-15
c169 4877 0 1.0881e-14
c170 4876 0 1.0232e-14
c171 4873 0 2.606e-15
c172 4871 0 1.225e-15
c173 4860 0 1.1019e-14
c174 4859 0 1.0488e-14
c175 4856 0 2.606e-15
c176 4854 0 1.225e-15
c177 4843 0 1.1019e-14
c178 4842 0 1.0488e-14
c179 4839 0 2.606e-15
c180 4837 0 1.225e-15
c181 4826 0 1.0818e-14
c182 4825 0 1.0309e-14
c183 4822 0 2.606e-15
c184 4820 0 1.225e-15
c185 4809 0 1.1019e-14
c186 4808 0 1.0327e-14
c187 4805 0 2.606e-15
c188 4803 0 1.225e-15
c189 4792 0 1.1019e-14
c190 4791 0 1.0488e-14
c191 4788 0 2.606e-15
c192 4786 0 1.225e-15
c193 4775 0 1.1019e-14
c194 4774 0 1.0488e-14
c195 4771 0 2.606e-15
c196 4769 0 1.225e-15
c197 4758 0 1.0839e-14
c198 4757 0 1.0488e-14
c199 4754 0 2.606e-15
c200 4752 0 1.225e-15
c201 4741 0 1.1019e-14
c202 4740 0 1.0488e-14
c203 4737 0 2.606e-15
c204 4735 0 1.225e-15
c205 4724 0 1.1019e-14
c206 4723 0 1.0488e-14
c207 4720 0 2.606e-15
c208 4718 0 1.225e-15
c209 4707 0 1.086e-14
c210 4706 0 1.0341e-14
c211 4703 0 2.606e-15
c212 4701 0 1.225e-15
c213 4690 0 1.1019e-14
c214 4689 0 1.0296e-14
c215 4686 0 2.606e-15
c216 4684 0 1.225e-15
c217 4673 0 1.1019e-14
c218 4672 0 1.0488e-14
c219 4669 0 2.606e-15
c220 4667 0 1.225e-15
c221 4656 0 1.1019e-14
c222 4655 0 1.0488e-14
c223 4652 0 2.606e-15
c224 4650 0 1.225e-15
c225 4639 0 1.0797e-14
c226 4638 0 1.0245e-14
c227 4635 0 2.606e-15
c228 4633 0 1.225e-15
c229 4622 0 1.1019e-14
c230 4621 0 1.0488e-14
c231 4618 0 2.606e-15
c232 4616 0 1.225e-15
c233 4605 0 1.1033e-14
c234 4604 0 1.0488e-14
c235 4601 0 2.606e-15
c236 4599 0 1.225e-15
c237 4577 0 1.0817e-14
c238 4570 0 1.3624e-14
c239 4559 0 2.2032e-14
c240 4558 0 9.475e-15
c241 4550 0 7.46e-15
c242 4553 0 1.984e-15
c243 4548 0 8.1e-16
c244 4536 0 1.1818e-14
c245 4535 0 1.0591e-14
c246 4532 0 2.606e-15
c247 4530 0 1.225e-15
c248 4519 0 1.1818e-14
c249 4518 0 1.0591e-14
c250 4515 0 2.606e-15
c251 4513 0 1.225e-15
c252 4502 0 1.1818e-14
c253 4501 0 1.0591e-14
c254 4498 0 2.606e-15
c255 4496 0 1.225e-15
c256 4485 0 1.1818e-14
c257 4484 0 1.0591e-14
c258 4481 0 2.606e-15
c259 4479 0 1.225e-15
c260 4468 0 1.1818e-14
c261 4467 0 1.0591e-14
c262 4464 0 2.606e-15
c263 4462 0 1.225e-15
c264 4451 0 1.1818e-14
c265 4450 0 1.0591e-14
c266 4447 0 2.606e-15
c267 4445 0 1.225e-15
c268 4434 0 1.1818e-14
c269 4433 0 1.0591e-14
c270 4430 0 2.606e-15
c271 4428 0 1.225e-15
c272 4417 0 1.1818e-14
c273 4416 0 1.0591e-14
c274 4413 0 2.606e-15
c275 4411 0 1.225e-15
c276 4400 0 1.1818e-14
c277 4399 0 1.0591e-14
c278 4396 0 2.606e-15
c279 4394 0 1.225e-15
c280 4383 0 1.1818e-14
c281 4382 0 1.0591e-14
c282 4379 0 2.606e-15
c283 4377 0 1.225e-15
c284 4366 0 1.1818e-14
c285 4365 0 1.0591e-14
c286 4362 0 2.606e-15
c287 4360 0 1.225e-15
c288 4349 0 1.1818e-14
c289 4348 0 1.0591e-14
c290 4345 0 2.606e-15
c291 4343 0 1.225e-15
c292 4332 0 1.1818e-14
c293 4331 0 1.0591e-14
c294 4328 0 2.606e-15
c295 4326 0 1.225e-15
c296 4315 0 1.1818e-14
c297 4314 0 1.0591e-14
c298 4311 0 2.606e-15
c299 4309 0 1.225e-15
c300 4298 0 1.1818e-14
c301 4297 0 1.0591e-14
c302 4294 0 2.606e-15
c303 4292 0 1.225e-15
c304 4281 0 1.1818e-14
c305 4280 0 1.0591e-14
c306 4277 0 2.606e-15
c307 4275 0 1.225e-15
c308 4264 0 1.1818e-14
c309 4263 0 1.0591e-14
c310 4260 0 2.606e-15
c311 4258 0 1.225e-15
c312 4247 0 1.1818e-14
c313 4246 0 1.0591e-14
c314 4243 0 2.606e-15
c315 4241 0 1.225e-15
c316 4225 0 1.3665e-14
c317 4217 0 2.2391e-14
c318 4226 0 1.5034e-14
c319 4223 0 8.428e-15
c320 4218 0 1.5318e-14
c321 4204 0 1.4918e-14
c322 4207 0 1.3549e-14
c323 4199 0 2.2275e-14
c324 4205 0 8.372e-15
c325 4200 0 1.5255e-14
c326 4190 0 1.3665e-14
c327 4182 0 2.2391e-14
c328 4191 0 1.5034e-14
c329 4188 0 8.428e-15
c330 4183 0 1.5318e-14
c331 4171 0 1.4918e-14
c332 4174 0 1.3549e-14
c333 4166 0 2.2275e-14
c334 4172 0 8.372e-15
c335 4167 0 1.5255e-14
c336 4158 0 1.3665e-14
c337 4150 0 2.2391e-14
c338 4159 0 1.5034e-14
c339 4156 0 8.428e-15
c340 4151 0 1.5318e-14
c341 4139 0 1.4918e-14
c342 4142 0 1.3549e-14
c343 4134 0 2.2275e-14
c344 4140 0 8.372e-15
c345 4135 0 1.5255e-14
c346 4126 0 1.3665e-14
c347 4118 0 2.2391e-14
c348 4127 0 1.5034e-14
c349 4124 0 8.428e-15
c350 4119 0 1.5318e-14
c351 4107 0 1.4918e-14
c352 4110 0 1.3549e-14
c353 4102 0 2.2275e-14
c354 4108 0 8.372e-15
c355 4103 0 1.5255e-14
c356 4094 0 1.3665e-14
c357 4086 0 2.2391e-14
c358 4095 0 1.5034e-14
c359 4092 0 8.428e-15
c360 4087 0 1.5318e-14
c361 4075 0 1.4918e-14
c362 4078 0 1.3549e-14
c363 4070 0 2.2275e-14
c364 4076 0 8.372e-15
c365 4071 0 1.5255e-14
c366 4062 0 1.3665e-14
c367 4054 0 2.2391e-14
c368 4063 0 1.5034e-14
c369 4060 0 8.428e-15
c370 4055 0 1.5318e-14
c371 4043 0 1.4918e-14
c372 4046 0 1.3549e-14
c373 4038 0 2.2275e-14
c374 4044 0 8.372e-15
c375 4039 0 1.5255e-14
c376 4030 0 1.3665e-14
c377 4022 0 2.2391e-14
c378 4031 0 1.5034e-14
c379 4028 0 8.428e-15
c380 4023 0 1.5318e-14
c381 4011 0 1.4918e-14
c382 4014 0 1.3549e-14
c383 4006 0 2.2275e-14
c384 4012 0 8.372e-15
c385 4007 0 1.5255e-14
c386 3998 0 1.3665e-14
c387 3990 0 2.2391e-14
c388 3999 0 1.5034e-14
c389 3996 0 8.428e-15
c390 3991 0 1.5318e-14
c391 3979 0 1.4918e-14
c392 3982 0 1.3549e-14
c393 3974 0 2.2275e-14
c394 3980 0 8.372e-15
c395 3975 0 1.5255e-14
c396 3966 0 1.3578e-14
c397 3958 0 2.2391e-14
c398 3967 0 1.5034e-14
c399 3964 0 8.428e-15
c400 3959 0 1.5318e-14
c401 3947 0 1.4918e-14
c402 3950 0 1.3549e-14
c403 3942 0 2.2275e-14
c404 3948 0 8.372e-15
c405 3943 0 1.5255e-14
c406 3934 0 1.3665e-14
c407 3926 0 2.2391e-14
c408 3935 0 1.5034e-14
c409 3932 0 8.428e-15
c410 3927 0 1.5318e-14
c411 3914 0 1.4918e-14
c412 3917 0 1.3549e-14
c413 3909 0 2.2275e-14
c414 3915 0 8.372e-15
c415 3910 0 1.5255e-14
c416 3895 0 1.0292e-14
c417 3875 0 1.4941e-14
c418 3872 0 2.0685e-14
c419 3871 0 8.578e-15
c420 3863 0 7.46e-15
c421 3866 0 1.984e-15
c422 3862 0 8.1e-16
c423 3840 0 1.3582e-14
c424 3842 0 1.4338e-14
c425 3836 0 2.8059e-14
c426 3838 0 1.8475e-14
c427 3806 0 3.7591e-14
c428 3830 0 1.356e-15
c429 3828 0 1.31e-15
c430 3808 0 1.2712e-14
c431 3804 0 2.233e-14
c432 3803 0 1.348e-14
c433 3811 0 2.1059e-14
c434 3801 0 1.4886e-14
c435 3780 0 1.2701e-14
c436 3783 0 1.3522e-14
c437 3770 0 3.2684e-14
c438 3774 0 1.4719e-14
c439 3772 0 2.349e-14
c440 3769 0 1.4906e-14
c441 3765 0 2.3688e-14
c442 3767 0 1.4226e-14
c443 3763 0 1.2709e-14
c444 3789 0 5.74e-16
c445 3786 0 5.74e-16
c446 3731 0 3.782e-14
c447 3759 0 1.356e-15
c448 3757 0 1.31e-15
c449 3733 0 1.3057e-14
c450 3729 0 2.2866e-14
c451 3728 0 1.3061e-14
c452 3736 0 2.0899e-14
c453 3726 0 1.3115e-14
c454 3723 0 1.1818e-14
c455 3722 0 1.0591e-14
c456 3719 0 2.606e-15
c457 3717 0 1.225e-15
c458 3706 0 1.1818e-14
c459 3705 0 1.0591e-14
c460 3702 0 2.606e-15
c461 3700 0 1.225e-15
c462 3689 0 1.1818e-14
c463 3688 0 1.0591e-14
c464 3685 0 2.606e-15
c465 3683 0 1.225e-15
c466 3672 0 1.1818e-14
c467 3671 0 1.0591e-14
c468 3668 0 2.606e-15
c469 3666 0 1.225e-15
c470 3655 0 1.1818e-14
c471 3654 0 1.0591e-14
c472 3651 0 2.606e-15
c473 3649 0 1.225e-15
c474 3638 0 1.1818e-14
c475 3637 0 1.0591e-14
c476 3634 0 2.606e-15
c477 3632 0 1.225e-15
c478 3621 0 1.1818e-14
c479 3620 0 1.0591e-14
c480 3617 0 2.606e-15
c481 3615 0 1.225e-15
c482 3604 0 1.1818e-14
c483 3603 0 1.0591e-14
c484 3600 0 2.606e-15
c485 3598 0 1.225e-15
c486 3587 0 1.1818e-14
c487 3586 0 1.0591e-14
c488 3583 0 2.606e-15
c489 3581 0 1.225e-15
c490 3570 0 1.1818e-14
c491 3569 0 1.0591e-14
c492 3566 0 2.606e-15
c493 3564 0 1.225e-15
c494 3553 0 1.1818e-14
c495 3552 0 1.0591e-14
c496 3549 0 2.606e-15
c497 3547 0 1.225e-15
c498 3536 0 1.1818e-14
c499 3535 0 1.0591e-14
c500 3532 0 2.606e-15
c501 3530 0 1.225e-15
c502 3519 0 1.1818e-14
c503 3518 0 1.0591e-14
c504 3515 0 2.606e-15
c505 3513 0 1.225e-15
c506 3502 0 1.1818e-14
c507 3501 0 1.0591e-14
c508 3498 0 2.606e-15
c509 3496 0 1.225e-15
c510 3485 0 1.1818e-14
c511 3484 0 1.0591e-14
c512 3481 0 2.606e-15
c513 3479 0 1.225e-15
c514 3468 0 1.1818e-14
c515 3467 0 1.0591e-14
c516 3464 0 2.606e-15
c517 3462 0 1.225e-15
c518 3451 0 1.1818e-14
c519 3450 0 1.0591e-14
c520 3447 0 2.606e-15
c521 3445 0 1.225e-15
c522 3434 0 1.1818e-14
c523 3433 0 1.0591e-14
c524 3430 0 2.606e-15
c525 3428 0 1.225e-15
c526 3406 0 1.0292e-14
c527 3386 0 1.5028e-14
c528 3383 0 2.0685e-14
c529 3382 0 8.578e-15
c530 3374 0 7.46e-15
c531 3377 0 1.984e-15
c532 3372 0 8.1e-16
c533 3360 0 1.1818e-14
c534 3359 0 1.0591e-14
c535 3356 0 2.606e-15
c536 3354 0 1.225e-15
c537 3343 0 1.1818e-14
c538 3342 0 1.0591e-14
c539 3339 0 2.606e-15
c540 3337 0 1.225e-15
c541 3326 0 1.1818e-14
c542 3325 0 1.0591e-14
c543 3322 0 2.606e-15
c544 3320 0 1.225e-15
c545 3309 0 1.1818e-14
c546 3308 0 1.0591e-14
c547 3305 0 2.606e-15
c548 3303 0 1.225e-15
c549 3292 0 1.1818e-14
c550 3291 0 1.0591e-14
c551 3288 0 2.606e-15
c552 3286 0 1.225e-15
c553 3275 0 1.1818e-14
c554 3274 0 1.0591e-14
c555 3271 0 2.606e-15
c556 3269 0 1.225e-15
c557 3258 0 1.1818e-14
c558 3257 0 1.0591e-14
c559 3254 0 2.606e-15
c560 3252 0 1.225e-15
c561 3241 0 1.1818e-14
c562 3240 0 1.0591e-14
c563 3237 0 2.606e-15
c564 3235 0 1.225e-15
c565 3224 0 1.1818e-14
c566 3223 0 1.0591e-14
c567 3220 0 2.606e-15
c568 3218 0 1.225e-15
c569 3207 0 1.1818e-14
c570 3206 0 1.0591e-14
c571 3203 0 2.606e-15
c572 3201 0 1.225e-15
c573 3190 0 1.1818e-14
c574 3189 0 1.0591e-14
c575 3186 0 2.606e-15
c576 3184 0 1.225e-15
c577 3173 0 1.1818e-14
c578 3172 0 1.0591e-14
c579 3169 0 2.606e-15
c580 3167 0 1.225e-15
c581 3156 0 1.1818e-14
c582 3155 0 1.0591e-14
c583 3152 0 2.606e-15
c584 3150 0 1.225e-15
c585 3139 0 1.1818e-14
c586 3138 0 1.0591e-14
c587 3135 0 2.606e-15
c588 3133 0 1.225e-15
c589 3122 0 1.1818e-14
c590 3121 0 1.0591e-14
c591 3118 0 2.606e-15
c592 3116 0 1.225e-15
c593 3105 0 1.1818e-14
c594 3104 0 1.0591e-14
c595 3101 0 2.606e-15
c596 3099 0 1.225e-15
c597 3088 0 1.1818e-14
c598 3087 0 1.0591e-14
c599 3084 0 2.606e-15
c600 3082 0 1.225e-15
c601 3071 0 1.1818e-14
c602 3070 0 1.0591e-14
c603 3067 0 2.606e-15
c604 3065 0 1.225e-15
c605 3043 0 1.0292e-14
c606 3023 0 1.5028e-14
c607 3020 0 2.0685e-14
c608 3019 0 8.578e-15
c609 3011 0 7.46e-15
c610 3014 0 1.984e-15
c611 3010 0 8.1e-16
c612 2988 0 1.3582e-14
c613 2990 0 1.4338e-14
c614 2984 0 2.8059e-14
c615 2986 0 1.8475e-14
c616 2954 0 3.7591e-14
c617 2978 0 1.356e-15
c618 2976 0 1.31e-15
c619 2956 0 1.2712e-14
c620 2952 0 2.233e-14
c621 2951 0 1.348e-14
c622 2959 0 2.1059e-14
c623 2949 0 1.4886e-14
c624 2928 0 1.2701e-14
c625 2931 0 1.3522e-14
c626 2918 0 3.2684e-14
c627 2922 0 1.4719e-14
c628 2920 0 2.349e-14
c629 2917 0 1.4906e-14
c630 2913 0 2.3688e-14
c631 2915 0 1.4226e-14
c632 2911 0 1.2709e-14
c633 2937 0 5.74e-16
c634 2934 0 5.74e-16
c635 2879 0 3.782e-14
c636 2907 0 1.356e-15
c637 2905 0 1.31e-15
c638 2881 0 1.3057e-14
c639 2877 0 2.2866e-14
c640 2876 0 1.3061e-14
c641 2884 0 2.0899e-14
c642 2874 0 1.3115e-14
c643 2871 0 1.1818e-14
c644 2870 0 1.0591e-14
c645 2867 0 2.606e-15
c646 2865 0 1.225e-15
c647 2854 0 1.1818e-14
c648 2853 0 1.0591e-14
c649 2850 0 2.606e-15
c650 2848 0 1.225e-15
c651 2837 0 1.1818e-14
c652 2836 0 1.0591e-14
c653 2833 0 2.606e-15
c654 2831 0 1.225e-15
c655 2820 0 1.1818e-14
c656 2819 0 1.0591e-14
c657 2816 0 2.606e-15
c658 2814 0 1.225e-15
c659 2803 0 1.1818e-14
c660 2802 0 1.0591e-14
c661 2799 0 2.606e-15
c662 2797 0 1.225e-15
c663 2786 0 1.1818e-14
c664 2785 0 1.0591e-14
c665 2782 0 2.606e-15
c666 2780 0 1.225e-15
c667 2769 0 1.1818e-14
c668 2768 0 1.0591e-14
c669 2765 0 2.606e-15
c670 2763 0 1.225e-15
c671 2752 0 1.1818e-14
c672 2751 0 1.0591e-14
c673 2748 0 2.606e-15
c674 2746 0 1.225e-15
c675 2735 0 1.1818e-14
c676 2734 0 1.0591e-14
c677 2731 0 2.606e-15
c678 2729 0 1.225e-15
c679 2718 0 1.1818e-14
c680 2717 0 1.0591e-14
c681 2714 0 2.606e-15
c682 2712 0 1.225e-15
c683 2701 0 1.1818e-14
c684 2700 0 1.0591e-14
c685 2697 0 2.606e-15
c686 2695 0 1.225e-15
c687 2684 0 1.1818e-14
c688 2683 0 1.0591e-14
c689 2680 0 2.606e-15
c690 2678 0 1.225e-15
c691 2667 0 1.1818e-14
c692 2666 0 1.0591e-14
c693 2663 0 2.606e-15
c694 2661 0 1.225e-15
c695 2650 0 1.1818e-14
c696 2649 0 1.0591e-14
c697 2646 0 2.606e-15
c698 2644 0 1.225e-15
c699 2633 0 1.1818e-14
c700 2632 0 1.0591e-14
c701 2629 0 2.606e-15
c702 2627 0 1.225e-15
c703 2616 0 1.1818e-14
c704 2615 0 1.0591e-14
c705 2612 0 2.606e-15
c706 2610 0 1.225e-15
c707 2599 0 1.1818e-14
c708 2598 0 1.0591e-14
c709 2595 0 2.606e-15
c710 2593 0 1.225e-15
c711 2582 0 1.1818e-14
c712 2581 0 1.0591e-14
c713 2578 0 2.606e-15
c714 2576 0 1.225e-15
c715 2554 0 1.0292e-14
c716 2534 0 1.4933e-14
c717 2531 0 2.0685e-14
c718 2530 0 8.578e-15
c719 2522 0 7.46e-15
c720 2525 0 1.984e-15
c721 2520 0 8.1e-16
c722 2508 0 1.1818e-14
c723 2507 0 1.0591e-14
c724 2504 0 2.606e-15
c725 2502 0 1.225e-15
c726 2491 0 1.1818e-14
c727 2490 0 1.0591e-14
c728 2487 0 2.606e-15
c729 2485 0 1.225e-15
c730 2474 0 1.1818e-14
c731 2473 0 1.0591e-14
c732 2470 0 2.606e-15
c733 2468 0 1.225e-15
c734 2457 0 1.1818e-14
c735 2456 0 1.0591e-14
c736 2453 0 2.606e-15
c737 2451 0 1.225e-15
c738 2440 0 1.1818e-14
c739 2439 0 1.0591e-14
c740 2436 0 2.606e-15
c741 2434 0 1.225e-15
c742 2423 0 1.1818e-14
c743 2422 0 1.0591e-14
c744 2419 0 2.606e-15
c745 2417 0 1.225e-15
c746 2406 0 1.1818e-14
c747 2405 0 1.0591e-14
c748 2402 0 2.606e-15
c749 2400 0 1.225e-15
c750 2389 0 1.1818e-14
c751 2388 0 1.0591e-14
c752 2385 0 2.606e-15
c753 2383 0 1.225e-15
c754 2372 0 1.1818e-14
c755 2371 0 1.0591e-14
c756 2368 0 2.606e-15
c757 2366 0 1.225e-15
c758 2355 0 1.1818e-14
c759 2354 0 1.0591e-14
c760 2351 0 2.606e-15
c761 2349 0 1.225e-15
c762 2338 0 1.1818e-14
c763 2337 0 1.0591e-14
c764 2334 0 2.606e-15
c765 2332 0 1.225e-15
c766 2321 0 1.1818e-14
c767 2320 0 1.0591e-14
c768 2317 0 2.606e-15
c769 2315 0 1.225e-15
c770 2304 0 1.1818e-14
c771 2303 0 1.0591e-14
c772 2300 0 2.606e-15
c773 2298 0 1.225e-15
c774 2287 0 1.1818e-14
c775 2286 0 1.0591e-14
c776 2283 0 2.606e-15
c777 2281 0 1.225e-15
c778 2270 0 1.1818e-14
c779 2269 0 1.0591e-14
c780 2266 0 2.606e-15
c781 2264 0 1.225e-15
c782 2253 0 1.1818e-14
c783 2252 0 1.0591e-14
c784 2249 0 2.606e-15
c785 2247 0 1.225e-15
c786 2236 0 1.1818e-14
c787 2235 0 1.0591e-14
c788 2232 0 2.606e-15
c789 2230 0 1.225e-15
c790 2219 0 1.1818e-14
c791 2218 0 1.0591e-14
c792 2215 0 2.606e-15
c793 2213 0 1.225e-15
c794 2191 0 1.0292e-14
c795 2171 0 1.4931e-14
c796 2168 0 2.0685e-14
c797 2167 0 8.578e-15
c798 2159 0 7.46e-15
c799 2162 0 1.984e-15
c800 2158 0 8.1e-16
c801 2137 0 1.3582e-14
c802 2139 0 1.4338e-14
c803 2133 0 2.8059e-14
c804 2135 0 1.8475e-14
c805 2103 0 3.7591e-14
c806 2127 0 1.356e-15
c807 2125 0 1.31e-15
c808 2105 0 1.2712e-14
c809 2101 0 2.233e-14
c810 2100 0 1.348e-14
c811 2108 0 2.1059e-14
c812 2098 0 1.4886e-14
c813 2077 0 1.2701e-14
c814 2080 0 1.3522e-14
c815 2067 0 3.2684e-14
c816 2071 0 1.4719e-14
c817 2069 0 2.349e-14
c818 2066 0 1.4906e-14
c819 2062 0 2.3688e-14
c820 2064 0 1.4226e-14
c821 2060 0 1.2709e-14
c822 2086 0 5.74e-16
c823 2083 0 5.74e-16
c824 2028 0 3.782e-14
c825 2056 0 1.356e-15
c826 2054 0 1.31e-15
c827 2030 0 1.3057e-14
c828 2026 0 2.2866e-14
c829 2025 0 1.3061e-14
c830 2033 0 2.0899e-14
c831 2023 0 1.3115e-14
c832 2020 0 1.1818e-14
c833 2019 0 1.0591e-14
c834 2016 0 2.606e-15
c835 2014 0 1.225e-15
c836 2003 0 1.1818e-14
c837 2002 0 1.0591e-14
c838 1999 0 2.606e-15
c839 1997 0 1.225e-15
c840 1986 0 1.1818e-14
c841 1985 0 1.0591e-14
c842 1982 0 2.606e-15
c843 1980 0 1.225e-15
c844 1969 0 1.1818e-14
c845 1968 0 1.0591e-14
c846 1965 0 2.606e-15
c847 1963 0 1.225e-15
c848 1952 0 1.1818e-14
c849 1951 0 1.0591e-14
c850 1948 0 2.606e-15
c851 1946 0 1.225e-15
c852 1935 0 1.1818e-14
c853 1934 0 1.0591e-14
c854 1931 0 2.606e-15
c855 1929 0 1.225e-15
c856 1918 0 1.1818e-14
c857 1917 0 1.0591e-14
c858 1914 0 2.606e-15
c859 1912 0 1.225e-15
c860 1901 0 1.1818e-14
c861 1900 0 1.0591e-14
c862 1897 0 2.606e-15
c863 1895 0 1.225e-15
c864 1884 0 1.1818e-14
c865 1883 0 1.0591e-14
c866 1880 0 2.606e-15
c867 1878 0 1.225e-15
c868 1867 0 1.1818e-14
c869 1866 0 1.0591e-14
c870 1863 0 2.606e-15
c871 1861 0 1.225e-15
c872 1850 0 1.1818e-14
c873 1849 0 1.0591e-14
c874 1846 0 2.606e-15
c875 1844 0 1.225e-15
c876 1833 0 1.1818e-14
c877 1832 0 1.0591e-14
c878 1829 0 2.606e-15
c879 1827 0 1.225e-15
c880 1816 0 1.1818e-14
c881 1815 0 1.0591e-14
c882 1812 0 2.606e-15
c883 1810 0 1.225e-15
c884 1799 0 1.1818e-14
c885 1798 0 1.0591e-14
c886 1795 0 2.606e-15
c887 1793 0 1.225e-15
c888 1782 0 1.1818e-14
c889 1781 0 1.0591e-14
c890 1778 0 2.606e-15
c891 1776 0 1.225e-15
c892 1765 0 1.1818e-14
c893 1764 0 1.0591e-14
c894 1761 0 2.606e-15
c895 1759 0 1.225e-15
c896 1748 0 1.1818e-14
c897 1747 0 1.0591e-14
c898 1744 0 2.606e-15
c899 1742 0 1.225e-15
c900 1731 0 1.1818e-14
c901 1730 0 1.0591e-14
c902 1727 0 2.606e-15
c903 1725 0 1.225e-15
c904 1703 0 1.0292e-14
c905 1683 0 1.5028e-14
c906 1680 0 2.0685e-14
c907 1679 0 8.578e-15
c908 1671 0 7.46e-15
c909 1674 0 1.984e-15
c910 1669 0 8.1e-16
c911 1657 0 1.1818e-14
c912 1656 0 1.0591e-14
c913 1653 0 2.606e-15
c914 1651 0 1.225e-15
c915 1640 0 1.1818e-14
c916 1639 0 1.0591e-14
c917 1636 0 2.606e-15
c918 1634 0 1.225e-15
c919 1623 0 1.1818e-14
c920 1622 0 1.0591e-14
c921 1619 0 2.606e-15
c922 1617 0 1.225e-15
c923 1606 0 1.1818e-14
c924 1605 0 1.0591e-14
c925 1602 0 2.606e-15
c926 1600 0 1.225e-15
c927 1589 0 1.1818e-14
c928 1588 0 1.0591e-14
c929 1585 0 2.606e-15
c930 1583 0 1.225e-15
c931 1572 0 1.1818e-14
c932 1571 0 1.0591e-14
c933 1568 0 2.606e-15
c934 1566 0 1.225e-15
c935 1555 0 1.1818e-14
c936 1554 0 1.0591e-14
c937 1551 0 2.606e-15
c938 1549 0 1.225e-15
c939 1538 0 1.1818e-14
c940 1537 0 1.0591e-14
c941 1534 0 2.606e-15
c942 1532 0 1.225e-15
c943 1521 0 1.1818e-14
c944 1520 0 1.0591e-14
c945 1517 0 2.606e-15
c946 1515 0 1.225e-15
c947 1504 0 1.1818e-14
c948 1503 0 1.0591e-14
c949 1500 0 2.606e-15
c950 1498 0 1.225e-15
c951 1487 0 1.1818e-14
c952 1486 0 1.0591e-14
c953 1483 0 2.606e-15
c954 1481 0 1.225e-15
c955 1470 0 1.1818e-14
c956 1469 0 1.0591e-14
c957 1466 0 2.606e-15
c958 1464 0 1.225e-15
c959 1453 0 1.1818e-14
c960 1452 0 1.0591e-14
c961 1449 0 2.606e-15
c962 1447 0 1.225e-15
c963 1436 0 1.1818e-14
c964 1435 0 1.0591e-14
c965 1432 0 2.606e-15
c966 1430 0 1.225e-15
c967 1419 0 1.1818e-14
c968 1418 0 1.0591e-14
c969 1415 0 2.606e-15
c970 1413 0 1.225e-15
c971 1402 0 1.1818e-14
c972 1401 0 1.0591e-14
c973 1398 0 2.606e-15
c974 1396 0 1.225e-15
c975 1385 0 1.1818e-14
c976 1384 0 1.0591e-14
c977 1381 0 2.606e-15
c978 1379 0 1.225e-15
c979 1368 0 1.1818e-14
c980 1367 0 1.0591e-14
c981 1364 0 2.606e-15
c982 1362 0 1.225e-15
c983 1340 0 1.0292e-14
c984 1320 0 1.5758e-14
c985 1317 0 2.0685e-14
c986 1316 0 8.578e-15
c987 1299 0 1.7549e-14
c988 1307 0 1.4789e-14
c989 1309 0 1.1292e-14
c990 1306 0 1.2538e-14
c991 1305 0 7.123e-15
c992 1300 0 1.363e-14
c993 1294 0 1.0389e-14
c994 1297 0 1.1329e-14
c995 1293 0 1.2827e-14
c996 1276 0 1.2618e-14
c997 1278 0 1.3929e-14
c998 1275 0 1.553e-14
c999 1269 0 1.3865e-14
c1000 1272 0 1.3888e-14
c1001 1273 0 1.5379e-14
c1002 1268 0 1.3555e-14
c1003 1284 0 5.74e-16
c1004 1280 0 5.74e-16
c1005 1248 0 2.4453e-14
c1006 1264 0 1.356e-15
c1007 1262 0 1.31e-15
c1008 1242 0 1.3284e-14
c1009 1245 0 1.3911e-14
c1010 1246 0 1.3864e-14
c1011 920 0 3.23309e-13
c1012 1240 0 7.494e-15
c1013 919 0 3.08903e-13
c1014 1232 0 7.432e-15
c1015 1216 0 1.026e-14
c1016 1201 0 9.835e-15
c1017 1186 0 9.929e-15
c1018 1171 0 1.026e-14
c1019 1156 0 1.026e-14
c1020 1141 0 9.853e-15
c1021 1126 0 9.832e-15
c1022 1111 0 1.026e-14
c1023 1096 0 1.026e-14
c1024 1081 0 9.961e-15
c1025 1066 0 1.026e-14
c1026 1051 0 1.026e-14
c1027 1036 0 9.917e-15
c1028 1021 0 9.864e-15
c1029 1006 0 1.026e-14
c1030 991 0 1.026e-14
c1031 976 0 9.993e-15
c1032 961 0 1.0728e-14
c1033 944 0 1.1544e-14
c1034 942 0 1.2613e-14
c1035 941 0 9.788e-15
c1036 933 0 1.2004e-14
c1037 936 0 8.994e-15
c1038 918 0 1.7198e-14
c1039 932 0 7.109e-15
c1040 882 0 1.4477e-14
c1041 879 0 1.7796e-14
c1042 878 0 1.0263e-14
c1043 872 0 9.788e-15
c1044 863 0 1.2004e-14
c1045 866 0 8.672e-15
c1046 856 0 9.788e-15
c1047 847 0 1.2004e-14
c1048 850 0 8.672e-15
c1049 841 0 9.788e-15
c1050 832 0 1.2004e-14
c1051 835 0 8.672e-15
c1052 826 0 9.788e-15
c1053 817 0 1.2004e-14
c1054 820 0 8.672e-15
c1055 811 0 9.788e-15
c1056 802 0 1.2004e-14
c1057 805 0 8.672e-15
c1058 796 0 9.788e-15
c1059 787 0 1.2004e-14
c1060 790 0 8.672e-15
c1061 781 0 9.788e-15
c1062 772 0 1.2004e-14
c1063 775 0 8.672e-15
c1064 766 0 9.788e-15
c1065 757 0 1.2004e-14
c1066 760 0 8.672e-15
c1067 751 0 9.788e-15
c1068 742 0 1.2004e-14
c1069 745 0 8.672e-15
c1070 736 0 9.788e-15
c1071 727 0 1.2004e-14
c1072 730 0 8.672e-15
c1073 721 0 9.788e-15
c1074 712 0 1.2004e-14
c1075 715 0 8.672e-15
c1076 706 0 9.788e-15
c1077 697 0 1.2004e-14
c1078 700 0 8.672e-15
c1079 691 0 9.788e-15
c1080 682 0 1.2004e-14
c1081 685 0 8.672e-15
c1082 676 0 9.788e-15
c1083 667 0 1.2004e-14
c1084 670 0 8.672e-15
c1085 661 0 9.788e-15
c1086 652 0 1.2004e-14
c1087 655 0 8.672e-15
c1088 646 0 9.788e-15
c1089 637 0 1.2004e-14
c1090 640 0 8.672e-15
c1091 631 0 9.788e-15
c1092 622 0 1.2004e-14
c1093 625 0 8.672e-15
c1094 616 0 9.788e-15
c1095 607 0 1.2004e-14
c1096 610 0 8.672e-15
c1097 600 0 9.788e-15
c1098 589 0 1.2004e-14
c1099 593 0 8.672e-15
c1100 581 0 1.1803e-14
c1101 580 0 9.0767e-14
c1102 577 0 2.0151e-14
c1103 576 0 1.4594e-14
c1104 553 0 1.1803e-14
c1105 552 0 9.0767e-14
c1106 549 0 2.0151e-14
c1107 548 0 1.4594e-14
c1108 524 0 1.1803e-14
c1109 523 0 9.0767e-14
c1110 520 0 2.0151e-14
c1111 519 0 1.4594e-14
c1112 495 0 1.1803e-14
c1113 494 0 9.0767e-14
c1114 491 0 2.0151e-14
c1115 490 0 1.4594e-14
c1116 466 0 1.1803e-14
c1117 465 0 9.0767e-14
c1118 462 0 2.0151e-14
c1119 461 0 1.4594e-14
c1120 437 0 1.1803e-14
c1121 436 0 9.0325e-14
c1122 433 0 2.0151e-14
c1123 432 0 1.4594e-14
c1124 408 0 1.1803e-14
c1125 407 0 9.0767e-14
c1126 404 0 2.0151e-14
c1127 403 0 1.4594e-14
c1128 379 0 1.1803e-14
c1129 378 0 9.0767e-14
c1130 375 0 2.0151e-14
c1131 374 0 1.4594e-14
c1132 350 0 1.1803e-14
c1133 349 0 9.0767e-14
c1134 346 0 2.0151e-14
c1135 345 0 1.4594e-14
c1136 321 0 1.1803e-14
c1137 320 0 9.0546e-14
c1138 317 0 2.0151e-14
c1139 316 0 1.4594e-14
c1140 292 0 1.1803e-14
c1141 291 0 9.0767e-14
c1142 288 0 2.0151e-14
c1143 287 0 1.4594e-14
c1144 263 0 1.1803e-14
c1145 262 0 9.0767e-14
c1146 259 0 2.0151e-14
c1147 258 0 1.4594e-14
c1148 234 0 1.1803e-14
c1149 233 0 9.0767e-14
c1150 230 0 2.0151e-14
c1151 229 0 1.4594e-14
c1152 205 0 1.1803e-14
c1153 204 0 9.0767e-14
c1154 201 0 2.0151e-14
c1155 200 0 1.4594e-14
c1156 176 0 1.1803e-14
c1157 175 0 9.0767e-14
c1158 172 0 2.0151e-14
c1159 171 0 1.4594e-14
c1160 147 0 1.1803e-14
c1161 146 0 9.0325e-14
c1162 143 0 2.0151e-14
c1163 142 0 1.4594e-14
c1164 118 0 1.1803e-14
c1165 117 0 9.0767e-14
c1166 114 0 2.0151e-14
c1167 113 0 1.4594e-14
c1168 89 0 1.1803e-14
c1169 88 0 9.0767e-14
c1170 85 0 2.0151e-14
c1171 84 0 1.4594e-14
c1172 60 0 1.1803e-14
c1173 59 0 9.0767e-14
c1174 56 0 2.0151e-14
c1175 55 0 1.4594e-14
c1176 28 0 1.1803e-14
c1177 27 0 9.0767e-14
c1178 22 0 2.0151e-14
c1179 21 0 1.4594e-14
c1180 2730 777 1.58e-16
c1181 2747 762 3.79e-16
c1182 2713 3235 1.96e-16
c1183 2719 3230 1.96e-16
c1184 3162 677 1.9e-16
c1185 2057 2056 1.6e-16
c1186 2067 1 6.62e-16
c1187 612 1715 1.58e-16
c1188 601 2215 7.68e-16
c1189 602 1682 1.58e-16
c1190 349 570 1.88e-16
c1191 909 1007 4.35e-16
c1192 907 1006 1.88e-16
c1193 890 999 1.58e-16
c1194 4305 662 1.84e-16
c1195 2824 2435 2.386e-15
c1196 2807 2452 1.58e-16
c1197 4567 4847 1.58e-16
c1198 3243 1 1.716e-15
c1199 1788 662 5.03e-16
c1200 2351 707 3.64e-16
c1201 3619 1 1.056e-15
c1202 1969 812 7.38e-16
c1203 1583 1574 3.46e-16
c1204 4639 632 1.23e-16
c1205 4642 4643 2.48e-16
c1206 4647 4646 2.83e-16
c1207 4650 4259 1.96e-16
c1208 3150 2628 1.96e-16
c1209 2194 842 4.46e-16
c1210 4752 1 8.43e-16
c1211 4971 526 2.51e-16
c1212 2713 752 1.58e-16
c1213 2165 2161 1.96e-16
c1214 747 1516 3.79e-16
c1215 277 291 1.58e-16
c1216 1 148 4.92e-16
c1217 15 137 4.88e-16
c1218 9 117 5.8e-16
c1219 288 274 3.84e-16
c1220 3679 3678 1.6e-16
c1221 3293 3674 3.92e-16
c1222 687 2671 1.58e-16
c1223 2461 1 5.808e-15
c1224 596 725 5.28e-16
c1225 657 3117 3.79e-16
c1226 601 2567 1.339e-15
c1227 2463 0 3.466e-15
c1228 136 0 7.3842e-14
c1229 2265 2260 1.642e-15
c1230 1508 737 1.58e-16
c1231 1076 732 3.79e-16
c1232 5530 5543 1.96e-16
c1233 4810 381 1.88e-16
c1234 2545 2469 5.5e-16
c1235 2849 2844 1.642e-15
c1236 1573 807 1.58e-16
c1237 1345 1041 1.58e-16
c1238 1343 1031 5.5e-16
c1239 1331 1486 1.58e-16
c1240 767 1 3.1284e-14
c1241 3718 3713 1.642e-15
c1242 1830 1829 1.6e-16
c1243 1822 1820 2.15e-16
c1244 642 1694 7.99e-16
c1245 4175 19 3.84e-16
c1246 4184 0 2.0707e-14
c1247 4926 4907 6.67e-16
c1248 1755 1756 5.65e-16
c1249 762 1113 1.58e-16
c1250 4463 4435 2.64e-16
c1251 4830 4836 7.25e-16
c1252 5010 265 1.88e-16
c1253 3048 3224 3.92e-16
c1254 1641 1690 1.58e-16
c1255 1196 0 7.482e-14
c1256 3589 3592 6.44e-16
c1257 4733 4730 3.01e-16
c1258 50 54 1.372e-15
c1259 27 5 1.325e-15
c1260 31 34 4.6e-16
c1261 4563 4276 5.88e-16
c1262 4571 4282 1.58e-16
c1263 1913 2430 2.38e-15
c1264 3773 3809 1.58e-16
c1265 4387 732 1.58e-16
c1266 883 1113 3.54e-16
c1267 894 1134 1.58e-16
c1268 5353 5357 5.6e-16
c1269 1465 722 1.58e-16
c1270 392 88 1.88e-16
c1271 3036 3035 6.97e-16
c1272 3037 3033 1.71e-16
c1273 911 921 3.45e-16
c1274 3983 19 3.84e-16
c1275 3992 0 2.0707e-14
c1276 1643 1644 2.48e-16
c1277 1046 1 5.821e-15
c1278 3590 3592 2.03e-16
c1279 4327 4711 1.36e-15
c1280 4720 4714 1.6e-16
c1281 2856 852 1.58e-16
c1282 1794 1783 1.58e-16
c1283 822 1619 2.65e-16
c1284 2186 1698 3.84e-16
c1285 0 588 2.87e-16
c1286 19 577 3.84e-16
c1287 3876 777 3.15e-16
c1288 5175 0 2.156e-15
c1289 2282 1 5.97e-15
c1290 1104 1111 2.27e-16
c1291 894 931 1.58e-16
c1292 222 15 6.58e-16
c1293 4283 647 1.339e-15
c1294 5352 5350 5.48e-16
c1295 4855 294 1.88e-16
c1296 2172 2004 1.58e-16
c1297 2178 1998 5.88e-16
c1298 4741 722 1.23e-16
c1299 1579 797 1.84e-16
c1300 1331 722 3.15e-16
c1301 1388 966 2.48e-16
c1302 1327 1161 1.58e-16
c1303 2594 3112 2.38e-15
c1304 747 749 5.59e-16
c1305 4353 1 5.808e-15
c1306 4355 0 3.466e-15
c1307 3554 747 5.73e-16
c1308 2899 2895 1.64e-16
c1309 3489 672 1.58e-16
c1310 3492 647 1.58e-16
c1311 4891 1 9.25e-16
c1312 1 322 4.92e-16
c1313 9 304 6.48e-16
c1314 4810 4816 5.87e-16
c1315 2004 2512 1.361e-15
c1316 1998 2182 5.5e-16
c1317 2417 1 8.43e-16
c1318 1008 1021 1.58e-16
c1319 762 26 1.58e-16
c1320 5530 526 3.54e-16
c1321 5526 0 1.376e-15
c1322 3009 1 5.01e-16
c1323 1226 1225 2.07e-16
c1324 1061 1059 1.931e-15
c1325 3886 732 7.99e-16
c1326 3898 722 4.46e-16
c1327 642 997 1.58e-16
c1328 632 982 6.38e-16
c1329 2048 0 1.8423e-14
c1330 2541 2390 1.58e-16
c1331 4267 4269 2.03e-16
c1332 3174 0 3.583e-14
c1333 3690 4523 7.84e-16
c1334 1095 1 3.06e-16
c1335 3048 3160 1.58e-16
c1336 608 607 1.96e-16
c1337 3207 722 7.38e-16
c1338 3409 3502 3.92e-16
c1339 465 447 1.58e-16
c1340 5337 1 3.36e-16
c1341 3713 858 1.84e-16
c1342 5296 5286 1.58e-16
c1343 4878 91 1.88e-16
c1344 1163 1164 1.213e-15
c1345 3385 3418 1.418e-15
c1346 4249 4251 1.862e-15
c1347 3429 3384 2.64e-16
c1348 3898 4502 3.92e-16
c1349 3769 1 2.53e-16
c1350 601 4232 1.339e-15
c1351 2668 3177 7.84e-16
c1352 3474 3089 1.96e-16
c1353 3479 3083 1.96e-16
c1354 1979 1 6.15e-16
c1355 482 494 1.58e-16
c1356 490 491 6.4e-16
c1357 5126 1 3.36e-16
c1358 3030 852 4.03e-16
c1359 3387 3259 1.58e-16
c1360 2776 2390 5.66e-16
c1361 392 390 1.88e-16
c1362 99 102 1.099e-15
c1363 4719 381 1.88e-16
c1364 601 3441 1.58e-16
c1365 1557 782 1.339e-15
c1366 3882 3469 1.58e-16
c1367 1727 1318 1.96e-16
c1368 922 920 4.274e-15
c1369 919 921 4.694e-15
c1370 1331 1121 5.5e-16
c1371 856 19 1.96e-16
c1372 996 0 3.7129e-14
c1373 4412 3571 1.136e-15
c1374 84 19 3.45e-16
c1375 368 364 1.58e-16
c1376 3292 782 1.58e-16
c1377 3048 702 3.58e-16
c1378 2223 2221 1.862e-15
c1379 3321 2804 1.136e-15
c1380 2072 2080 3.54e-16
c1381 238 207 1.88e-16
c1382 4657 4663 5.87e-16
c1383 4567 4774 1.58e-16
c1384 4580 4378 5.5e-16
c1385 4582 4384 1.58e-16
c1386 5238 5237 1.6e-16
c1387 2570 0 6.62e-16
c1388 596 635 5.28e-16
c1389 3736 3732 1.96e-16
c1390 3385 3872 1.58e-16
c1391 4039 4036 1.58e-16
c1392 3142 0 2.93e-15
c1393 2214 2209 1.642e-15
c1394 375 19 8.4e-16
c1395 378 25 5.71e-16
c1396 5482 5478 5.7e-16
c1397 5422 5435 9.34e-16
c1398 1760 647 3.15e-16
c1399 2671 2683 2.32e-16
c1400 919 1069 1.58e-16
c1401 3510 0 6.72e-16
c1402 2952 2954 1.133e-15
c1403 1202 0 1.0183e-14
c1404 3048 2804 1.58e-16
c1405 3046 2798 5.5e-16
c1406 3248 3245 5.5e-16
c1407 1767 0 1.6491e-14
c1408 4666 1 6.42e-16
c1409 4395 4774 1.58e-16
c1410 4463 0 6.9337e-14
c1411 3409 3438 1.58e-16
c1412 2559 868 3.58e-16
c1413 2107 2108 5.07e-16
c1414 2082 2070 5.37e-16
c1415 233 455 1.88e-16
c1416 5190 5195 3.54e-16
c1417 566 565 1.079e-15
c1418 3542 3543 1.6e-16
c1419 3538 3157 3.92e-16
c1420 3960 857 3.1e-16
c1421 2398 2395 3.01e-16
c1422 2394 2391 6.44e-16
c1423 2167 1 1.96e-16
c1424 88 276 1.88e-16
c1425 5452 5492 4.39e-16
c1426 890 852 4.14e-16
c1427 3855 3411 3.25e-16
c1428 602 3069 4.81e-16
c1429 2967 0 1.65e-16
c1430 919 717 3.15e-16
c1431 971 975 2.03e-16
c1432 1321 1372 1.58e-16
c1433 4135 4132 1.58e-16
c1434 1833 677 1.58e-16
c1435 1455 1016 1.532e-15
c1436 3673 4505 2.48e-16
c1437 2535 2751 1.58e-16
c1438 2557 2739 1.58e-16
c1439 4070 37 1.88e-16
c1440 4400 3565 1.96e-16
c1441 3248 3255 6.73e-16
c1442 3024 2645 5.5e-16
c1443 3046 2628 5.5e-16
c1444 3179 702 2.72e-16
c1445 2106 1211 1.12e-15
c1446 4466 1 1.056e-15
c1447 4626 0 3.4653e-14
c1448 4693 4692 2.03e-16
c1449 1562 0 1.4092e-14
c1450 3538 717 1.58e-16
c1451 5232 0 3.974e-14
c1452 4982 4974 3.54e-16
c1453 3385 3386 3.36e-16
c1454 3034 837 7.99e-16
c1455 642 2541 4.03e-16
c1456 777 1684 3.15e-16
c1457 909 702 3.15e-16
c1458 5046 0 1.65e-16
c1459 2217 2215 1.6e-16
c1460 1682 2171 1.62e-16
c1461 5591 4531 1.58e-16
c1462 2724 0 3.466e-15
c1463 1070 707 5.74e-16
c1464 858 864 1.078e-15
c1465 1343 807 3.15e-16
c1466 4094 3918 6.32e-16
c1467 4623 5426 3.92e-16
c1468 3301 0 8e-16
c1469 601 3046 4.46e-16
c1470 2628 2623 1.642e-15
c1471 3886 3429 5.5e-16
c1472 3859 0 6.72e-16
c1473 1603 1602 1.6e-16
c1474 1595 1593 2.15e-16
c1475 1343 1538 3.92e-16
c1476 811 19 1.96e-16
c1477 1694 1815 1.58e-16
c1478 1392 1 2.054e-15
c1479 3080 3077 3.01e-16
c1480 3076 3073 6.44e-16
c1481 1394 0 8e-16
c1482 1875 1873 1.6e-16
c1483 1870 1869 2.03e-16
c1484 4979 4978 3.54e-16
c1485 2195 2189 1.988e-15
c1486 2196 1 2.222e-15
c1487 1067 717 2.68e-16
c1488 852 859 1.065e-15
c1489 3219 3617 4.36e-16
c1490 617 2603 1.832e-15
c1491 2004 0 3.7647e-14
c1492 2031 2045 2.217e-15
c1493 4606 4610 1.81e-16
c1494 5437 1 3.36e-16
c1495 4922 31 3.84e-16
c1496 4759 0 3.13327e-13
c1497 2477 1970 2.48e-16
c1498 2172 1732 1.58e-16
c1499 2178 1726 5.88e-16
c1500 1706 722 4.46e-16
c1501 1694 732 7.99e-16
c1502 3496 1 8.43e-16
c1503 4488 3650 4.97e-16
c1504 1162 0 1.8851e-14
c1505 3219 3610 4.11e-16
c1506 2662 677 3.15e-16
c1507 2334 1 1.868e-15
c1508 1 483 9.8e-16
c1509 459 19 3.2e-16
c1510 0 488 6.224e-15
c1511 3225 767 1.75e-16
c1512 2542 2186 2.035e-15
c1513 2324 0 2.93e-15
c1514 2182 1726 5.5e-16
c1515 862 850 7.23e-16
c1516 853 854 1.6e-16
c1517 91 1 3.36e-15
c1518 3497 3492 1.642e-15
c1519 4770 5195 1.152e-15
c1520 1443 677 1.84e-16
c1521 883 1187 3.92e-16
c1522 890 1186 1.88e-16
c1523 601 907 4.8e-16
c1524 4043 1 6.66e-16
c1525 4472 4484 2.32e-16
c1526 3341 3339 1.6e-16
c1527 2545 2305 1.58e-16
c1528 3034 3088 4.63e-16
c1529 657 1769 1.58e-16
c1530 3613 3610 3.01e-16
c1531 4743 4746 6.67e-16
c1532 1708 1956 1.58e-16
c1533 822 1331 7.99e-16
c1534 30 178 3.84e-16
c1535 5032 5031 3.92e-16
c1536 601 1682 3.15e-16
c1537 627 1715 5.73e-16
c1538 4940 1 1.23e-16
c1539 2678 1 8.43e-16
c1540 894 1022 3.92e-16
c1541 909 1021 1.88e-16
c1542 883 1014 1.58e-16
c1543 4322 672 1.58e-16
c1544 4922 5149 2.24e-16
c1545 4878 5106 1.279e-15
c1546 4567 4864 1.58e-16
c1547 1321 767 4.48e-16
c1548 4024 25 7.01e-16
c1549 1845 707 3.15e-16
c1550 1331 1677 6.18e-16
c1551 4746 4744 2.03e-16
c1552 766 19 1.96e-16
c1553 3126 3138 2.32e-16
c1554 1362 1 8.43e-16
c1555 3898 822 3.15e-16
c1556 1351 0 3.22e-16
c1557 4557 4558 1.76e-16
c1558 1488 1 4.41e-15
c1559 4769 1 8.43e-16
c1560 1872 0 6.62e-16
c1561 3409 3168 5.5e-16
c1562 3857 852 2.42e-16
c1563 5590 1 8e-16
c1564 2758 2367 4.11e-16
c1565 2481 1 2.054e-15
c1566 2483 0 8e-16
c1567 1528 737 1.58e-16
c1568 2817 2810 6.73e-16
c1569 2532 0 4.4158e-14
c1570 1321 1046 5.5e-16
c1571 1331 1491 1.58e-16
c1572 4218 1 4.45e-16
c1573 1998 852 1.13e-15
c1574 1134 1 2.972e-15
c1575 1135 0 6.29e-16
c1576 4452 4463 1.58e-16
c1577 3316 3315 1.6e-16
c1578 2271 1 4.41e-15
c1579 3797 3796 1.6e-16
c1580 4563 4293 5.88e-16
c1581 5081 91 3.54e-16
c1582 4793 207 1.88e-16
c1583 5440 439 3.54e-16
c1584 165 0 9.3149e-14
c1585 149 33 1.88e-16
c1586 2835 1 1.056e-15
c1587 3401 1 8.822e-15
c1588 2806 2424 2.48e-16
c1589 1882 722 4.81e-16
c1590 1500 1056 1.96e-16
c1591 1501 1494 6.73e-16
c1592 3047 3041 1.988e-15
c1593 632 1391 5.03e-16
c1594 2882 2929 2.851e-15
c1595 2931 2928 4.87e-16
c1596 2946 2933 3.92e-16
c1597 931 1 4.632e-15
c1598 4837 4828 3.46e-16
c1599 945 0 8.475e-15
c1600 4344 4711 1.58e-16
c1601 3030 3020 3.54e-16
c1602 3046 3023 1.58e-16
c1603 822 1166 3.79e-16
c1604 447 450 1.099e-15
c1605 433 436 3.54e-16
c1606 3900 792 3.58e-16
c1607 1326 886 7.67e-16
c1608 4899 4900 6.09e-16
c1609 1098 737 1.58e-16
c1610 401 1 2.87e-16
c1611 2636 2638 2.03e-16
c1612 395 0 9.795e-15
c1613 4770 0 3.91995e-13
c1614 4657 33 1.88e-16
c1615 4069 4070 3.15e-16
c1616 642 3429 1.58e-16
c1617 3211 0 3.3874e-14
c1618 146 223 1.88e-16
c1619 3974 19 7.04e-16
c1620 4369 3537 2.48e-16
c1621 2577 2572 1.642e-15
c1622 2321 702 2.4e-16
c1623 1343 1176 1.58e-16
c1624 924 0 1.1387e-14
c1625 4373 1 2.054e-15
c1626 2775 782 5.03e-16
c1627 187 194 7.76e-16
c1628 4375 0 8e-16
c1629 1253 0 3.5494e-14
c1630 5281 352 9.68e-16
c1631 5291 5316 3.54e-16
c1632 1 28 1.456e-15
c1633 17 0 1.4803e-14
c1634 3411 827 3.15e-16
c1635 3387 868 3.15e-16
c1636 4827 4830 6.02e-16
c1637 5267 5151 1.52e-16
c1638 5253 5232 1.96e-16
c1639 1028 1029 1.213e-15
c1640 3019 1 1.96e-16
c1641 1218 883 1.96e-16
c1642 59 421 1.88e-16
c1643 3900 737 3.15e-16
c1644 4855 62 7.67e-16
c1645 2559 0 3.396e-13
c1646 2557 2407 1.58e-16
c1647 920 1115 3.92e-16
c1648 921 1114 2.54e-16
c1649 3701 4535 1.58e-16
c1650 2557 3017 4.22e-16
c1651 617 1369 2.33e-16
c1652 1109 1 3.06e-16
c1653 4879 4503 4.51e-16
c1654 4891 4890 1.6e-16
c1655 3030 2668 1.58e-16
c1656 2135 2133 1.167e-15
c1657 15 571 4.88e-16
c1658 3191 3574 7.84e-16
c1659 2412 1896 4.11e-16
c1660 1732 0 3.6368e-14
c1661 816 805 7.23e-16
c1662 5286 0 3.8102e-14
c1663 70 0 9.795e-15
c1664 53 19 3.2e-16
c1665 3370 2899 1.96e-16
c1666 3842 2892 2.12e-16
c1667 3537 722 1.75e-16
c1668 4793 5229 6.5e-16
c1669 921 926 2.712e-15
c1670 3562 0 8e-16
c1671 1850 717 2.4e-16
c1672 3876 4519 3.92e-16
c1673 3007 3006 1.6e-16
c1674 722 26 7.12e-16
c1675 4143 19 3.84e-16
c1676 3886 4332 4.63e-16
c1677 4440 3599 4.11e-16
c1678 2679 3189 1.58e-16
c1679 2541 732 4.03e-16
c1680 1618 1985 1.58e-16
c1681 1690 1884 1.96e-16
c1682 612 1731 2.4e-16
c1683 509 515 1.372e-15
c1684 505 504 6.67e-16
c1685 2225 0 3.466e-15
c1686 1988 1 1.716e-15
c1687 5106 1 3.914e-15
c1688 2322 2323 1.35e-16
c1689 5025 0 5.736e-14
c1690 3411 3276 1.58e-16
c1691 1087 1088 7.46e-16
c1692 890 882 1.58e-16
c1693 883 904 1.58e-16
c1694 70 69 6.67e-16
c1695 2584 0 1.6491e-14
c1696 4567 4580 4.369e-15
c1697 5587 4563 6.89e-16
c1698 4657 5492 3.92e-16
c1699 4640 5452 7.84e-16
c1700 627 3455 1.58e-16
c1701 617 3441 1.84e-16
c1702 2557 2773 1.58e-16
c1703 1131 1132 8.58e-16
c1704 2559 2203 1.58e-16
c1705 2557 2170 5.5e-16
c1706 2545 2598 1.58e-16
c1707 675 1 1.65e-16
c1708 3180 3179 1.6e-16
c1709 1904 1905 2.48e-16
c1710 822 1706 3.15e-16
c1711 4864 4863 2.48e-16
c1712 4867 4868 2.83e-16
c1713 5165 178 4.02e-16
c1714 3397 3100 5.5e-16
c1715 2585 0 2.93e-15
c1716 1 567 4.22e-16
c1717 3411 812 3.15e-16
c1718 4567 4791 1.58e-16
c1719 4580 4395 5.5e-16
c1720 4582 4401 1.58e-16
c1721 5503 1 7.49e-16
c1722 2493 1987 3.92e-16
c1723 2497 2498 1.6e-16
c1724 3031 2549 2.035e-15
c1725 1343 1572 3.92e-16
c1726 2015 2508 1.96e-16
c1727 612 3411 3.58e-16
c1728 3185 747 1.58e-16
c1729 2955 2954 5.88e-16
c1730 3360 2849 1.96e-16
c1731 3024 2815 5.5e-16
c1732 3625 3632 1.96e-16
c1733 4683 1 6.42e-16
c1734 4412 4774 1.58e-16
c1735 4401 4782 5.66e-16
c1736 4788 4779 3.92e-16
c1737 2679 717 1.813e-15
c1738 2072 2071 6.26e-16
c1739 480 479 7.08e-16
c1740 427 436 1.58e-16
c1741 15 187 5.8e-16
c1742 306 303 2.142e-15
c1743 0 197 1.4803e-14
c1744 5490 0 1.65e-16
c1745 5131 5133 1.609e-15
c1746 5039 5135 9.36e-16
c1747 3770 3767 1.732e-15
c1748 3765 3792 5.87e-16
c1749 3935 3926 1.96e-16
c1750 1474 702 1.58e-16
c1751 596 837 1.96e-16
c1752 612 2533 1.813e-15
c1753 2308 2320 2.32e-16
c1754 4233 3384 2.48e-16
c1755 4355 707 5.03e-16
c1756 2674 2681 6.73e-16
c1757 1345 1389 1.58e-16
c1758 3091 3093 2.03e-16
c1759 2584 2203 3.92e-16
c1760 3876 4455 1.58e-16
c1761 3900 4467 5.42e-16
c1762 3030 2538 1.96e-16
c1763 851 1 5.57e-16
c1764 4112 0 1.18545e-13
c1765 2070 2067 9.58e-16
c1766 4482 1 9.28e-16
c1767 4643 0 3.485e-14
c1768 2557 692 4.46e-16
c1769 2545 702 7.99e-16
c1770 1971 1982 1.96e-16
c1771 3151 3539 4.97e-16
c1772 4582 4570 2.14e-16
c1773 5105 5103 5.25e-16
c1774 3174 707 2.33e-16
c1775 632 2535 4.48e-16
c1776 792 1708 3.58e-16
c1777 894 717 8.34e-16
c1778 111 117 1.58e-16
c1779 5257 149 3.54e-16
c1780 2765 762 2.65e-16
c1781 2744 0 8e-16
c1782 2203 2585 2.48e-16
c1783 2531 1 2.346e-15
c1784 602 3426 1.09e-16
c1785 3317 0 6.72e-16
c1786 3136 1 9.28e-16
c1787 617 3046 4.46e-16
c1788 2178 792 4.03e-16
c1789 378 9 5.8e-16
c1790 4532 842 3.64e-16
c1791 2781 792 3.79e-16
c1792 1862 732 3.79e-16
c1793 824 25 1.13e-15
c1794 828 19 1.58e-16
c1795 1410 0 6.72e-16
c1796 3055 3438 7.84e-16
c1797 1499 1867 1.96e-16
c1798 190 194 1.58e-16
c1799 368 262 1.88e-16
c1800 2849 868 3.79e-16
c1801 3262 767 1.832e-15
c1802 1681 2205 2.48e-16
c1803 1752 1 5.808e-15
c1804 5590 4950 1.6e-16
c1805 2782 2384 4.36e-16
c1806 3123 1 4.41e-15
c1807 4022 4024 3.54e-16
c1808 4623 4625 4.93e-16
c1809 2182 792 7.99e-16
c1810 2841 2853 2.32e-16
c1811 2918 1 6.62e-16
c1812 919 842 3.15e-16
c1813 920 1173 1.58e-16
c1814 3669 1 9.28e-16
c1815 1973 827 1.58e-16
c1816 1708 737 3.15e-16
c1817 2731 737 7.68e-16
c1818 2178 737 3.15e-16
c1819 1741 1 6.15e-16
c1820 3411 3406 1.58e-16
c1821 1828 1 5.97e-15
c1822 2065 2064 8.03e-16
c1823 1652 2007 1.58e-16
c1824 5240 1 2.424e-15
c1825 3885 3883 3.67e-16
c1826 1511 1508 5.5e-16
c1827 4577 4578 1.796e-15
c1828 657 996 4e-16
c1829 3472 0 3.3691e-14
c1830 2770 1 4.41e-15
c1831 617 907 4.8e-16
c1832 3886 3588 1.58e-16
c1833 4677 4299 7.84e-16
c1834 2418 812 1.58e-16
c1835 2430 797 1.84e-16
c1836 2182 737 3.15e-16
c1837 1784 1397 1.532e-15
c1838 1790 1789 5.65e-16
c1839 4595 1 2.378e-15
c1840 1690 1590 1.58e-16
c1841 4594 0 3.466e-15
c1842 3509 3506 5.5e-16
c1843 5254 1 3.36e-16
c1844 2387 2385 1.6e-16
c1845 627 2249 2.65e-16
c1846 617 1682 1.58e-16
c1847 4993 4991 3.92e-16
c1848 4977 4537 6.29e-16
c1849 910 2532 3.75e-16
c1850 2286 1777 1.58e-16
c1851 1142 767 1.58e-16
c1852 894 1036 1.58e-16
c1853 907 1008 3.54e-16
c1854 277 276 1.079e-15
c1855 161 175 1.58e-16
c1856 2659 2656 3.01e-16
c1857 2655 2652 6.44e-16
c1858 657 655 3.327e-15
c1859 4567 4881 1.58e-16
c1860 2136 2036 6.72e-16
c1861 1322 1326 1.988e-15
c1862 3894 1 1.002e-15
c1863 4389 4390 1.6e-16
c1864 4385 3554 3.92e-16
c1865 5558 5562 1.202e-15
c1866 657 1767 1.58e-16
c1867 3387 0 3.17834e-13
c1868 4659 4660 2.48e-16
c1869 4664 4663 2.83e-16
c1870 4667 4276 1.96e-16
c1871 3565 0 6.9481e-14
c1872 5383 265 3.54e-16
c1873 5009 4896 1.58e-16
c1874 2987 2923 1.58e-16
c1875 1897 1 1.868e-15
c1876 749 750 1.6e-16
c1877 4786 1 8.43e-16
c1878 2174 2173 6.67e-16
c1879 1887 0 2.93e-15
c1880 3387 3586 1.58e-16
c1881 5294 5278 7.48e-16
c1882 5170 5182 3.18e-16
c1883 1044 692 1.58e-16
c1884 687 3117 1.58e-16
c1885 3786 3732 1.191e-15
c1886 4100 4104 3.84e-16
c1887 4044 3918 2.87e-16
c1888 1309 1239 8.9e-16
c1889 1299 1295 1.96e-16
c1890 910 945 6.76e-16
c1891 3156 2645 1.96e-16
c1892 1973 812 1.832e-15
c1893 1601 807 2.22e-16
c1894 2529 3020 4.65e-16
c1895 1835 1846 1.96e-16
c1896 1769 1768 2.48e-16
c1897 1705 1 2.94e-16
c1898 792 1132 1.58e-16
c1899 4748 0 1.4233e-14
c1900 1697 0 6.35e-16
c1901 4563 4310 5.88e-16
c1902 4571 4316 1.58e-16
c1903 822 26 1.58e-16
c1904 2453 1936 1.96e-16
c1905 2454 2447 6.73e-16
c1906 0 183 2.87e-16
c1907 5529 5543 5.12e-16
c1908 2178 2190 6.67e-16
c1909 3834 3844 1.98e-16
c1910 3016 2486 1.23e-16
c1911 2851 1 9.28e-16
c1912 1001 662 3.15e-16
c1913 911 925 7.25e-16
c1914 528 524 6.38e-16
c1915 149 147 6.01e-16
c1916 632 1411 1.09e-16
c1917 967 1 3.54e-16
c1918 4015 1 5.284e-15
c1919 4462 4455 1.96e-16
c1920 3616 4464 4.36e-16
c1921 3312 2798 4.97e-16
c1922 2408 782 1.339e-15
c1923 4005 0 1.5061e-14
c1924 4007 19 3.45e-16
c1925 964 0 9.347e-15
c1926 4546 4547 3.01e-16
c1927 4344 4728 1.36e-15
c1928 4737 4731 1.6e-16
c1929 3390 3038 7.84e-16
c1930 3126 662 1.58e-16
c1931 1694 1550 5.5e-16
c1932 1514 1 6.15e-16
c1933 21 5 1.108e-15
c1934 4215 0 5.525e-14
c1935 1938 1940 2.03e-16
c1936 5057 5056 1.6e-16
c1937 5028 5031 3.54e-16
c1938 5049 5048 3.92e-16
c1939 272 1 4.22e-16
c1940 910 2559 5.03e-16
c1941 1117 752 1.58e-16
c1942 1098 1104 1.58e-16
c1943 4304 647 1.9e-16
c1944 2640 0 1.4092e-14
c1945 4204 3918 8.1e-16
c1946 1146 797 2.33e-16
c1947 3411 747 3.58e-16
c1948 2611 2600 1.58e-16
c1949 1311 1 5.5e-16
c1950 1920 1922 1.862e-15
c1951 1533 1539 1.418e-15
c1952 647 638 1.078e-15
c1953 5010 5011 3.54e-16
c1954 4582 4299 1.58e-16
c1955 3048 3046 4.506e-15
c1956 602 2173 5.18e-16
c1957 592 682 1.96e-16
c1958 239 30 6.83e-16
c1959 4719 4333 1.179e-15
c1960 2333 2339 1.418e-15
c1961 1389 1401 2.32e-16
c1962 4055 857 6.23e-16
c1963 3734 3781 2.851e-15
c1964 3209 0 1.6491e-14
c1965 3639 807 1.58e-16
c1966 2535 2424 1.58e-16
c1967 3707 4543 8.31e-16
c1968 2684 692 7.38e-16
c1969 3046 2685 1.58e-16
c1970 1181 1 5.821e-15
c1971 4711 1 4.832e-15
c1972 19 316 3.45e-16
c1973 136 565 1.88e-16
c1974 3202 3557 1.58e-16
c1975 3672 812 7.38e-16
c1976 5529 526 3.54e-16
c1977 4861 439 1.88e-16
c1978 2413 0 1.4092e-14
c1979 1177 1158 1.546e-15
c1980 3702 827 3.64e-16
c1981 4279 4277 1.6e-16
c1982 2237 2620 7.84e-16
c1983 3578 0 6.72e-16
c1984 1481 1472 3.46e-16
c1985 2541 3003 3.16e-16
c1986 3024 762 3.15e-16
c1987 2879 2895 2.062e-15
c1988 3693 1 5.808e-15
c1989 1539 1540 1.35e-16
c1990 3203 3197 1.6e-16
c1991 2679 3194 2.386e-15
c1992 2696 3177 1.58e-16
c1993 2854 827 1.58e-16
c1994 1618 1990 1.58e-16
c1995 1706 1901 3.92e-16
c1996 453 452 6.67e-16
c1997 465 455 1.88e-16
c1998 3577 3576 1.6e-16
c1999 3491 3100 4.11e-16
c2000 2245 0 8e-16
c2001 4855 5113 9.98e-16
c2002 6 13 3.84e-16
c2003 3387 3287 5.5e-16
c2004 4855 4850 1.536e-15
c2005 2786 2418 1.96e-16
c2006 919 925 3.92e-16
c2007 4657 526 1.88e-16
c2008 2849 0 7.0008e-14
c2009 3886 4331 1.58e-16
c2010 3599 4434 1.96e-16
c2011 1319 1315 1.58e-16
c2012 3928 25 7.01e-16
c2013 4589 64 1.88e-16
c2014 2535 2214 5.5e-16
c2015 2545 2603 1.58e-16
c2016 1181 1622 1.58e-16
c2017 685 1 3.79e-16
c2018 1690 1883 1.58e-16
c2019 921 1 9.72e-16
c2020 1706 1703 1.58e-16
c2021 1684 1704 3.92e-16
c2022 5114 0 2.9101e-14
c2023 3024 3359 1.58e-16
c2024 3046 3347 1.58e-16
c2025 3279 807 1.58e-16
c2026 2249 2251 1.6e-16
c2027 3409 3655 3.92e-16
c2028 2103 2130 9.6e-16
c2029 4065 4062 1.76e-16
c2030 4567 4808 1.58e-16
c2031 4580 4412 5.5e-16
c2032 4582 4418 1.58e-16
c2033 5239 5237 3.92e-16
c2034 4872 323 1.88e-16
c2035 1327 702 4.03e-16
c2036 91 94 4.6e-16
c2037 3322 822 2.65e-16
c2038 2178 2303 1.58e-16
c2039 3616 782 3.15e-16
c2040 1252 1250 1.6e-16
c2041 4346 4339 6.73e-16
c2042 4345 3503 1.96e-16
c2043 1321 1589 3.92e-16
c2044 627 3411 3.58e-16
c2045 3157 1 4.41e-15
c2046 2691 2688 5.5e-16
c2047 1541 1542 2.48e-16
c2048 1802 1804 2.03e-16
c2049 762 883 3.15e-16
c2050 4571 797 1.33e-16
c2051 4865 4862 6.67e-16
c2052 3048 2832 5.5e-16
c2053 4700 1 6.42e-16
c2054 4412 4791 1.58e-16
c2055 2103 2105 3.73e-16
c2056 2117 2119 3.92e-16
c2057 1 336 4.22e-16
c2058 523 516 3.54e-16
c2059 0 323 1.21052e-13
c2060 3555 3168 1.532e-15
c2061 762 2401 2.22e-16
c2062 2182 2303 1.58e-16
c2063 2172 1760 5.5e-16
c2064 894 1235 3.54e-16
c2065 909 907 4.754e-15
c2066 1234 890 5.49e-16
c2067 627 2533 1.58e-16
c2068 4375 707 1.09e-16
c2069 2288 2299 1.58e-16
c2070 2015 2507 1.58e-16
c2071 1327 981 1.58e-16
c2072 59 47 1.58e-16
c2073 717 1 4.1542e-14
c2074 595 1364 2.65e-16
c2075 602 880 2.33e-16
c2076 1196 1192 3.78e-16
c2077 3900 4472 1.58e-16
c2078 2659 662 1.09e-16
c2079 2461 837 1.58e-16
c2080 747 1097 2.68e-16
c2081 1058 0 1.4198e-14
c2082 3046 3139 3.92e-16
c2083 4782 4781 1.6e-16
c2084 2101 2105 5.6e-16
c2085 4495 1 6.15e-16
c2086 4660 0 3.4756e-14
c2087 2559 707 3.15e-16
c2088 602 1704 1.58e-16
c2089 5104 5103 3.92e-16
c2090 5106 5127 1.96e-16
c2091 1885 2393 7.84e-16
c2092 4954 4905 2.45e-16
c2093 5301 0 2.156e-15
c2094 4938 4936 5.66e-16
c2095 657 2559 3.58e-16
c2096 2311 2318 6.73e-16
c2097 2760 0 6.72e-16
c2098 2579 1 9.28e-16
c2099 2541 2175 1.96e-16
c2100 3731 3747 2.062e-15
c2101 612 3440 2.72e-16
c2102 3149 1 6.15e-16
c2103 1355 1362 1.96e-16
c2104 3565 4404 2.386e-15
c2105 4413 4407 1.6e-16
c2106 3701 842 3.15e-16
c2107 4640 5410 2.69e-16
c2108 2379 737 1.58e-16
c2109 1608 1619 1.96e-16
c2110 4486 4487 1.35e-16
c2111 3066 3450 1.58e-16
c2112 3562 707 1.09e-16
c2113 4977 4946 1.58e-16
c2114 5048 0 2.8602e-14
c2115 792 1922 1.58e-16
c2116 3409 3620 1.58e-16
c2117 5286 5285 5.25e-16
c2118 5010 381 1.88e-16
c2119 2550 0 6.35e-16
c2120 4640 4647 1.81e-16
c2121 4668 439 1.88e-16
c2122 2178 1919 1.58e-16
c2123 1331 672 7.99e-16
c2124 1357 877 4.11e-16
c2125 2541 2553 6.67e-16
c2126 643 1 1.65e-16
c2127 3682 1 6.15e-16
c2128 1993 827 1.58e-16
c2129 1990 868 1.58e-16
c2130 1321 1554 1.58e-16
c2131 1343 1542 1.58e-16
c2132 4223 4230 7.81e-16
c2133 2566 3075 7.84e-16
c2134 1880 1871 3.92e-16
c2135 1488 1874 5.66e-16
c2136 1499 1866 1.58e-16
c2137 632 2242 5.03e-16
c2138 4097 1 2.3688e-14
c2139 4283 0 1.6491e-14
c2140 3350 3356 1.6e-16
c2141 3347 2832 2.386e-15
c2142 2849 3330 1.58e-16
c2143 2172 752 4.48e-16
c2144 1750 1 1.716e-15
c2145 4841 1 1.013e-15
c2146 3620 3621 9.1e-16
c2147 3411 3021 1.58e-16
c2148 2370 1 1.056e-15
c2149 4725 4726 9.93e-16
c2150 2478 2490 2.32e-16
c2151 2182 1919 1.58e-16
c2152 0 430 6.224e-15
c2153 3636 767 4.81e-16
c2154 3781 3344 1.958e-15
c2155 3876 647 4.48e-16
c2156 3898 672 3.15e-16
c2157 894 842 3.15e-16
c2158 890 1173 3.54e-16
c2159 909 1194 1.58e-16
c2160 919 1023 1.58e-16
c2161 4217 4216 3.15e-16
c2162 5399 5170 1.33e-16
c2163 911 3411 3.45e-16
c2164 910 3387 5.22e-16
c2165 3492 0 1.4092e-14
c2166 1436 1016 1.96e-16
c2167 4492 4489 5.5e-16
c2168 3345 2838 3.92e-16
c2169 2452 797 1.58e-16
c2170 2633 647 7.38e-16
c2171 1032 0 6.29e-16
c2172 4612 1 2.378e-15
c2173 1706 1607 1.58e-16
c2174 4611 0 3.466e-15
c2175 1961 1958 3.01e-16
c2176 1957 1954 6.44e-16
c2177 25 494 5.71e-16
c2178 0 484 1.79784e-13
c2179 3911 3909 3.54e-16
c2180 5091 5069 6.67e-16
c2181 93 31 1.58e-16
c2182 911 2533 1.88e-16
c2183 602 3025 5.18e-16
c2184 2291 1777 2.386e-15
c2185 96 0 2.87e-16
c2186 2569 2581 2.32e-16
c2187 1801 677 1.339e-15
c2188 1421 986 1.532e-15
c2189 1427 1426 5.65e-16
c2190 1328 1326 8.67e-16
c2191 4040 37 5.71e-16
c2192 2541 2701 1.96e-16
c2193 1249 1250 3.18e-16
c2194 794 1 7.18e-16
c2195 3409 792 3.15e-16
c2196 3146 3143 5.5e-16
c2197 3419 3018 1.532e-15
c2198 3425 3424 5.65e-16
c2199 3397 3038 1.58e-16
c2200 2270 1760 1.96e-16
c2201 1516 1 5.97e-15
c2202 1987 1 4.41e-15
c2203 777 1903 1.58e-16
c2204 1038 1052 1.96e-16
c2205 88 570 1.88e-16
c2206 2496 0 6.62e-16
c2207 4063 3918 8.1e-16
c2208 2831 2824 1.96e-16
c2209 687 677 3.28e-16
c2210 2577 0 6.894e-14
c2211 3005 2492 2.91e-16
c2212 392 391 1.88e-16
c2213 4298 3463 1.96e-16
c2214 4244 1 9.28e-16
c2215 4197 4568 3.84e-16
c2216 1358 0 1.4092e-14
c2217 1148 1 4.59e-16
c2218 3410 3394 3.54e-16
c2219 1145 0 1.0077e-14
c2220 4217 26 4.48e-16
c2221 3333 3334 5.65e-16
c2222 1781 1414 1.58e-16
c2223 4765 0 1.4233e-14
c2224 1712 0 1.23e-16
c2225 1 369 1.607e-15
c2226 3409 737 4.46e-16
c2227 4872 265 1.88e-16
c2228 1947 1936 1.58e-16
c2229 3825 3806 7.95e-16
c2230 2864 1 6.15e-16
c2231 747 2339 5.73e-16
c2232 1197 827 4.98e-16
c2233 1193 842 1.58e-16
c2234 5410 5472 6.67e-16
c2235 921 1010 1.96e-16
c2236 542 291 1.88e-16
c2237 1773 1771 1.6e-16
c2238 1768 1767 2.03e-16
c2239 4849 4463 4.11e-16
c2240 4854 4845 3.46e-16
c2241 3146 662 1.58e-16
c2242 2033 2026 8.3e-16
c2243 1523 1 1.716e-15
c2244 0 265 1.21158e-13
c2245 1760 0 6.9481e-14
c2246 2085 1 3.36e-16
c2247 2356 2367 1.58e-16
c2248 2196 2200 1.6e-16
c2249 407 421 1.88e-16
c2250 64 354 1.88e-16
c2251 2653 2265 4.97e-16
c2252 1324 898 7.84e-16
c2253 1039 1040 7.51e-16
c2254 1136 812 1.58e-16
c2255 1293 1297 4.52e-16
c2256 1635 842 3.15e-16
c2257 1321 1181 5.5e-16
c2258 1331 1644 1.58e-16
c2259 749 1 7.18e-16
c2260 1575 1577 2.03e-16
c2261 3506 3117 2.386e-15
c2262 3554 1 4.41e-15
c2263 455 450 1.88e-16
c2264 4388 0 6.62e-16
c2265 3515 672 2.65e-16
c2266 4902 4918 2.072e-15
c2267 3397 3552 1.58e-16
c2268 4982 526 1.038e-15
c2269 404 25 7.06e-16
c2270 400 19 8.82e-16
c2271 284 274 8.86e-16
c2272 281 291 1.88e-16
c2273 657 3472 1.58e-16
c2274 5044 5265 2.12e-16
c2275 1772 647 1.84e-16
c2276 902 929 5.8e-16
c2277 4006 3918 2.48e-16
c2278 5540 5537 1.958e-15
c2279 5514 5517 3.54e-16
c2280 4702 5326 1.53e-15
c2281 1273 1269 2.45e-15
c2282 1076 1072 3.78e-16
c2283 4370 4382 2.32e-16
c2284 2559 2441 1.58e-16
c2285 1557 1559 1.862e-15
c2286 1106 1116 1.418e-15
c2287 1690 1352 1.58e-16
c2288 1825 1822 3.01e-16
c2289 1821 1818 6.44e-16
c2290 1290 0 1.65e-16
c2291 4917 4916 1.6e-16
c2292 3024 2702 1.58e-16
c2293 3030 2696 5.88e-16
c2294 1676 1 8e-16
c2295 4728 1 4.832e-15
c2296 1641 2154 8.31e-16
c2297 1 43 1.073e-15
c2298 12 5 5.8e-16
c2299 4844 4845 9.93e-16
c2300 0 44 1.024e-14
c2301 41 40 6.67e-16
c2302 27 37 1.88e-16
c2303 3387 707 4.48e-16
c2304 2435 0 6.9484e-14
c2305 2434 2425 3.46e-16
c2306 826 824 5.88e-16
c2307 5324 0 4.0816e-14
c2308 1001 999 1.931e-15
c2309 146 305 1.88e-16
c2310 657 3387 3.15e-16
c2311 3565 707 1.58e-16
c2312 4398 722 4.81e-16
c2313 1706 672 3.15e-16
c2314 1684 647 4.48e-16
c2315 911 878 1.81e-16
c2316 2248 2603 1.58e-16
c2317 3380 1 9.43e-16
c2318 3026 3025 6.67e-16
c2319 1487 1486 9.1e-16
c2320 3839 3747 1.772e-15
c2321 2196 837 3.58e-16
c2322 4165 0 1.5061e-14
c2323 4167 19 3.45e-16
c2324 752 0 2.80197e-13
c2325 3048 777 3.58e-16
c2326 2882 2907 1.96e-16
c2327 1735 1744 3.92e-16
c2328 1738 1352 5.66e-16
c2329 1363 1730 1.58e-16
c2330 937 1 6.2e-16
c2331 2144 1667 5.5e-16
c2332 4713 4327 4.11e-16
c2333 4718 4709 3.46e-16
c2334 1 584 7.348e-15
c2335 2261 0 6.72e-16
c2336 3338 3854 4.78e-16
c2337 3344 3853 3.92e-16
c2338 5262 207 1.58e-16
c2339 632 3101 7.68e-16
c2340 165 565 1.88e-16
c2341 4810 5265 1.628e-15
c2342 5326 5284 3.41e-16
c2343 2799 2407 1.96e-16
c2344 2237 2618 3.92e-16
c2345 2623 2622 1.6e-16
c2346 592 866 6.34e-16
c2347 1854 717 1.58e-16
c2348 3194 1 5.808e-15
c2349 1136 1140 2.03e-16
c2350 3886 4336 1.58e-16
c2351 3876 3497 5.5e-16
c2352 4668 5482 2.037e-15
c2353 2719 747 1.58e-16
c2354 2559 2231 5.5e-16
c2355 704 1 7.18e-16
c2356 3942 25 3.84e-16
c2357 3197 3198 5.65e-16
c2358 1181 1627 1.58e-16
c2359 1706 1900 1.58e-16
c2360 1690 1888 1.58e-16
c2361 3116 3107 3.46e-16
c2362 3100 3485 1.96e-16
c2363 792 922 3.15e-16
c2364 4881 4880 2.48e-16
c2365 3299 807 1.58e-16
c2366 3024 722 4.48e-16
c2367 1990 0 3.3874e-14
c2368 3270 3637 1.58e-16
c2369 3259 3645 5.66e-16
c2370 3651 3642 3.92e-16
c2371 812 805 5.58e-16
c2372 9 306 4.88e-16
c2373 3748 3734 2.217e-15
c2374 4218 857 6.23e-16
c2375 4567 4825 1.58e-16
c2376 4580 4429 5.5e-16
c2377 4582 4435 1.58e-16
c2378 642 3453 1.58e-16
c2379 2704 2322 2.48e-16
c2380 1321 717 3.15e-16
c2381 881 1381 4.36e-16
c2382 1379 1372 1.96e-16
c2383 5509 0 1.1948e-14
c2384 2815 822 3.79e-16
c2385 2194 2320 1.58e-16
c2386 2178 2308 1.58e-16
c2387 2136 1 4.67e-15
c2388 684 1 5.57e-16
c2389 3514 3503 1.58e-16
c2390 3566 1 1.868e-15
c2391 2594 3105 1.96e-16
c2392 1694 1683 1.58e-16
c2393 1235 1 4.42e-16
c2394 1222 0 2.2077e-14
c2395 2458 842 1.75e-16
c2396 911 2177 1.58e-16
c2397 777 909 3.15e-16
c2398 3277 807 1.58e-16
c2399 3393 3501 1.58e-16
c2400 4429 4791 1.58e-16
c2401 4418 4799 5.66e-16
c2402 4805 4796 3.92e-16
c2403 3192 732 1.58e-16
c2404 657 2640 1.58e-16
c2405 2151 2078 9.61e-16
c2406 3642 797 1.58e-16
c2407 4571 4604 1.58e-16
c2408 5491 0 3.4847e-14
c2409 4793 497 1.88e-16
c2410 2182 2308 1.58e-16
c2411 1715 1 4.41e-15
c2412 879 878 5.89e-16
c2413 895 896 6.73e-16
c2414 2328 2325 5.5e-16
c2415 922 737 5.14e-16
c2416 921 1068 1.58e-16
c2417 4250 3385 4.97e-16
c2418 2688 2695 1.96e-16
c2419 1663 858 1.58e-16
c2420 601 880 1.75e-16
c2421 852 25 1.58e-16
c2422 3882 3656 1.58e-16
c2423 2855 3367 8.31e-16
c2424 2481 837 1.58e-16
c2425 1431 1403 2.64e-16
c2426 3919 1 5.649e-15
c2427 612 4247 2.4e-16
c2428 3271 3272 1.6e-16
c2429 3262 3264 2.15e-16
c2430 3024 3156 3.92e-16
c2431 4504 1 1.716e-15
c2432 4677 0 3.4686e-14
c2433 1997 1601 1.96e-16
c2434 1992 1607 1.96e-16
c2435 480 494 1.58e-16
c2436 305 320 1.88e-16
c2437 3253 2736 1.136e-15
c2438 1149 807 1.58e-16
c2439 883 722 6.45e-16
c2440 909 1082 4.35e-16
c2441 907 1081 1.88e-16
c2442 890 1074 1.58e-16
c2443 4234 4246 2.32e-16
c2444 4776 5212 1.96e-16
c2445 3397 3253 5.5e-16
c2446 5320 5319 2.67e-16
c2447 5262 5229 1.58e-16
c2448 1068 1069 1.21e-16
c2449 595 593 3.327e-15
c2450 2838 1 4.41e-15
c2451 1818 702 1.58e-16
c2452 1657 842 1.58e-16
c2453 642 592 5.8e-16
c2454 3348 0 6.62e-16
c2455 397 395 1.257e-15
c2456 398 407 1.58e-16
c2457 361 403 9.5e-16
c2458 3914 1 6.66e-16
c2459 4542 852 2.42e-16
c2460 1720 1716 1.96e-16
c2461 3819 0 1.65e-16
c2462 1432 1 1.868e-15
c2463 4567 3890 1.58e-16
c2464 92 1 4.92e-16
c2465 4196 4581 1.846e-15
c2466 1422 0 2.93e-15
c2467 3464 3458 1.6e-16
c2468 3066 3455 2.386e-15
c2469 3083 3438 1.58e-16
c2470 2310 1794 4.11e-16
c2471 1682 2222 4.97e-16
c2472 792 1942 1.58e-16
c2473 1068 717 1.58e-16
c2474 2549 0 8.0911e-14
c2475 238 209 3.75e-16
c2476 4657 4665 1.81e-16
c2477 612 3434 2.4e-16
c2478 2194 1936 1.58e-16
c2479 1345 677 3.15e-16
c2480 2861 2858 5.5e-16
c2481 392 0 1.08834e-13
c2482 2559 2552 3.54e-16
c2483 3691 1 1.716e-15
c2484 4326 4317 3.46e-16
c2485 1777 647 3.15e-16
c2486 1091 1521 1.96e-16
c2487 842 1 3.1284e-14
c2488 2577 3087 1.58e-16
c2489 1499 1871 1.58e-16
c2490 632 2262 1.09e-16
c2491 1776 1 8.43e-16
c2492 4858 1 1.013e-15
c2493 5188 5192 1.088e-15
c2494 3387 3022 5.5e-16
c2495 5051 1 1.113e-15
c2496 883 1188 3.54e-16
c2497 894 1209 1.58e-16
c2498 5506 5505 1.6e-16
c2499 2933 0 3.0577e-14
c2500 2666 2667 9.1e-16
c2501 1936 812 1.75e-16
c2502 4629 1 2.378e-15
c2503 4764 4767 3.01e-16
c2504 3024 3121 1.58e-16
c2505 3046 3109 1.58e-16
c2506 1563 0 6.72e-16
c2507 4628 0 3.466e-15
c2508 777 1106 1.813e-15
c2509 762 1121 4.21e-16
c2510 335 341 1.372e-15
c2511 5151 0 5.7679e-14
c2512 3514 662 1.58e-16
c2513 894 1023 3.54e-16
c2514 1331 797 3.15e-16
c2515 1335 1338 2.109e-15
c2516 3882 4434 1.96e-16
c2517 2557 2718 3.92e-16
c2518 672 26 1.58e-16
c2519 1598 1595 3.01e-16
c2520 1594 1591 6.44e-16
c2521 4676 4677 2.48e-16
c2522 4681 4680 2.83e-16
c2523 4684 4293 1.96e-16
c2524 4999 4992 3.92e-16
c2525 4944 4978 1.24e-16
c2526 4972 4910 3.54e-16
c2527 2289 1777 1.532e-15
c2528 3393 3202 5.88e-16
c2529 2525 1 1.601e-15
c2530 1058 707 1.58e-16
c2531 4776 1 2.552e-14
c2532 4582 0 3.3892e-13
c2533 4736 497 1.88e-16
c2534 2513 0 6.78e-16
c2535 3886 807 7.99e-16
c2536 3898 797 4.46e-16
c2537 4489 827 1.58e-16
c2538 1091 752 3.15e-16
c2539 1101 1104 1.58e-16
c2540 3900 4234 1.58e-16
c2541 1331 1086 1.58e-16
c2542 3625 0 3.3874e-14
c2543 4257 1 6.15e-16
c2544 3056 2529 1.532e-15
c2545 3062 3061 5.65e-16
c2546 1861 1465 1.96e-16
c2547 1856 1471 1.96e-16
c2548 1170 1 3.06e-16
c2549 1902 1903 1.35e-16
c2550 4782 0 1.4233e-14
c2551 5288 5280 3.54e-16
c2552 9 494 5.8e-16
c2553 245 246 5.8e-16
c2554 5160 5157 7.84e-16
c2555 1947 2470 4.36e-16
c2556 2468 2461 1.96e-16
c2557 1436 662 7.38e-16
c2558 1215 842 6.48e-16
c2559 121 1 4.92e-16
c2560 4404 752 1.58e-16
c2561 920 1024 1.58e-16
c2562 3455 1 5.808e-15
c2563 1327 1326 3.15e-16
c2564 3457 0 3.466e-15
c2565 4039 1 6.03e-16
c2566 3876 4400 3.92e-16
c2567 4474 4472 2.15e-16
c2568 4482 4481 1.6e-16
c2569 1397 1765 1.96e-16
c2570 1567 1562 1.642e-15
c2571 0 168 1.4803e-14
c2572 3361 3821 5.71e-16
c2573 2196 2206 1.58e-16
c2574 2031 0 3.7984e-14
c2575 632 648 1.621e-15
c2576 170 166 1.372e-15
c2577 161 159 1.58e-16
c2578 2739 2356 7.84e-16
c2579 1621 812 4.81e-16
c2580 1166 797 3.57e-16
c2581 657 4283 1.58e-16
c2582 3882 4399 1.58e-16
c2583 4467 4468 9.1e-16
c2584 3024 822 3.15e-16
c2585 2887 2874 5.78e-16
c2586 2535 2666 1.58e-16
c2587 2557 2654 1.58e-16
c2588 3901 1 2.86e-16
c2589 2153 852 2.42e-16
c2590 632 1765 7.38e-16
c2591 1196 1345 5.5e-16
c2592 1671 1661 1.65e-16
c2593 3883 0 4.1004e-14
c2594 1338 1 7.228e-15
c2595 3136 3135 1.6e-16
c2596 3128 3126 2.15e-16
c2597 1950 1948 1.6e-16
c2598 5010 5001 7.01e-16
c2599 3506 677 1.58e-16
c2600 4402 762 1.58e-16
c2601 1981 1590 1.136e-15
c2602 5277 5291 5.12e-16
c2603 5390 5385 9.94e-16
c2604 3397 3557 1.58e-16
c2605 276 0 7.7571e-14
c2606 657 3492 1.58e-16
c2607 3338 858 3.15e-16
c2608 1409 1406 5.5e-16
c2609 2172 2372 3.92e-16
c2610 944 943 1.39e-15
c2611 3667 807 2.22e-16
c2612 4489 812 1.832e-15
c2613 3067 1 1.868e-15
c2614 2809 2805 1.96e-16
c2615 1270 1276 3.54e-16
c2616 3057 0 2.93e-15
c2617 919 1144 1.58e-16
c2618 1958 812 5.03e-16
c2619 3611 762 1.58e-16
c2620 1314 0 2.94e-16
c2621 4201 1 5.1e-16
c2622 1448 0 6.9481e-14
c2623 596 700 2.45e-16
c2624 9 246 6.48e-16
c2625 5064 91 3.15e-16
c2626 602 2572 1.58e-16
c2627 2440 2439 9.1e-16
c2628 157 1 4.59e-16
c2629 1016 993 6.54e-16
c2630 143 19 8.4e-16
c2631 139 0 1.4803e-14
c2632 4287 4288 1.6e-16
c2633 4283 3452 3.92e-16
c2634 5410 5407 3.54e-16
c2635 1493 1489 1.96e-16
c2636 3886 4556 6.18e-16
c2637 822 883 3.15e-16
c2638 2545 2820 4.63e-16
c2639 2194 662 4.46e-16
c2640 1735 1363 1.58e-16
c2641 2016 1624 1.96e-16
c2642 2017 2010 6.73e-16
c2643 3304 807 2.22e-16
c2644 4571 632 1.33e-16
c2645 5162 5157 3.73e-16
c2646 2196 1851 1.58e-16
c2647 335 349 1.58e-16
c2648 3591 737 1.832e-15
c2649 642 2594 1.813e-15
c2650 592 732 5.8e-16
c2651 5388 5291 6.72e-16
c2652 4753 1 2.111e-14
c2653 1115 737 1.58e-16
c2654 4623 0 3.49986e-13
c2655 3214 1 2.054e-15
c2656 3900 3514 5.5e-16
c2657 1733 1744 1.96e-16
c2658 925 1 2.48e-16
c2659 891 0 4.0542e-14
c2660 2078 858 1.58e-16
c2661 2645 672 3.79e-16
c2662 2628 647 3.15e-16
c2663 1684 1917 1.58e-16
c2664 1706 1905 1.58e-16
c2665 2181 1698 5.8e-16
c2666 2195 1687 3.54e-16
c2667 1694 1730 1.58e-16
c2668 747 1508 1.58e-16
c2669 1254 1 2.36e-15
c2670 5029 5026 1.075e-15
c2671 2351 1834 1.96e-16
c2672 2352 2345 6.73e-16
c2673 3723 852 2.4e-16
c2674 2790 2418 1.58e-16
c2675 2626 1 6.15e-16
c2676 3270 3642 1.58e-16
c2677 6 27 3.84e-16
c2678 13 0 4.2131e-14
c2679 4166 3918 2.48e-16
c2680 4567 4842 1.58e-16
c2681 4580 4446 5.5e-16
c2682 4582 4452 1.58e-16
c2683 2172 2337 1.58e-16
c2684 2194 2325 1.58e-16
c2685 4453 797 1.339e-15
c2686 4702 5284 1.925e-15
c2687 4360 4353 1.96e-16
c2688 3514 4362 4.36e-16
c2689 1706 797 4.46e-16
c2690 1694 807 7.99e-16
c2691 3185 1 5.97e-15
c2692 2545 777 7.99e-16
c2693 1265 1 3.36e-16
c2694 657 1760 1.813e-15
c2695 1256 0 1.65e-16
c2696 4150 1 7.08e-16
c2697 3364 3367 5.5e-16
c2698 3034 2855 1.58e-16
c2699 4429 4808 1.58e-16
c2700 3288 3279 3.92e-16
c2701 2770 3282 5.66e-16
c2702 2702 722 2.33e-16
c2703 2134 2036 3.87e-16
c2704 2103 2104 5.88e-16
c2705 3651 3640 1.96e-16
c2706 5165 5234 3.54e-16
c2707 1014 672 1.58e-16
c2708 812 804 1.74e-16
c2709 2249 1 1.868e-15
c2710 0 516 1.4803e-14
c2711 3662 797 1.58e-16
c2712 4015 857 1.88e-16
c2713 4897 64 1.049e-15
c2714 72 1 1.073e-15
c2715 3967 3964 4.41e-16
c2716 5388 5303 8.28e-16
c2717 3840 3370 2.241e-15
c2718 1345 996 1.58e-16
c2719 1343 986 5.5e-16
c2720 1331 1435 1.58e-16
c2721 4156 4159 4.41e-16
c2722 612 1381 2.65e-16
c2723 3747 1 2.269e-15
c2724 3898 3673 1.58e-16
c2725 2470 827 7.68e-16
c2726 1814 1812 1.6e-16
c2727 4132 19 3.84e-16
c2728 3955 1 6.78e-16
c2729 2545 2785 1.58e-16
c2730 4799 4798 1.6e-16
c2731 3196 722 5.03e-16
c2732 2106 2108 1.001e-15
c2733 2104 2101 5.5e-16
c2734 1151 0 7.4292e-14
c2735 4694 0 3.485e-14
c2736 1766 1767 1.35e-16
c2737 526 524 6.01e-16
c2738 513 509 1.58e-16
c2739 291 565 1.88e-16
c2740 3640 797 1.339e-15
c2741 523 570 1.88e-16
c2742 5131 1 1.88e-16
c2743 2325 2332 1.96e-16
c2744 3710 868 1.58e-16
c2745 2782 1 1.868e-15
c2746 2695 2686 3.46e-16
c2747 687 2559 3.58e-16
c2748 894 1097 3.92e-16
c2749 909 1096 1.88e-16
c2750 883 1089 1.58e-16
c2751 2772 0 2.93e-15
c2752 47 42 1.482e-15
c2753 4150 4151 1.58e-16
c2754 1454 692 2.33e-16
c2755 1321 842 4.48e-16
c2756 392 281 1.88e-16
c2757 3839 3739 6.72e-16
c2758 602 4237 1.58e-16
c2759 3264 3260 1.96e-16
c2760 3175 3176 2.03e-16
c2761 602 1720 1.9e-16
c2762 1634 1166 1.96e-16
c2763 1629 1176 1.96e-16
c2764 1694 1471 1.58e-16
c2765 5029 120 9.68e-16
c2766 5092 0 1.23e-16
c2767 1081 1082 1.238e-15
c2768 1072 732 1.58e-16
c2769 596 845 5.28e-16
c2770 2499 2497 1.6e-16
c2771 2494 2493 2.03e-16
c2772 2172 1953 1.58e-16
c2773 2178 1947 5.88e-16
c2774 3900 827 3.15e-16
c2775 3876 868 3.15e-16
c2776 4332 4331 9.1e-16
c2777 1327 1116 1.58e-16
c2778 4302 1 5.808e-15
c2779 3101 3095 1.6e-16
c2780 2577 3092 2.386e-15
c2781 1499 1891 2.38e-15
c2782 1209 1 2.972e-15
c2783 1210 0 6.29e-16
c2784 4304 0 3.466e-15
c2785 5198 178 1.58e-16
c2786 3281 782 1.9e-16
c2787 456 460 1.372e-15
c2788 458 459 1.58e-16
c2789 427 425 1.58e-16
c2790 1 198 2.87e-16
c2791 390 433 1.88e-16
c2792 4651 4646 1.536e-15
c2793 3411 3066 5.5e-16
c2794 2182 1947 5.5e-16
c2795 2374 1 1.716e-15
c2796 0 193 1.5723e-14
c2797 3918 3915 2.87e-16
c2798 5471 0 1.963e-15
c2799 1485 692 4.81e-16
c2800 397 291 1.88e-16
c2801 5296 381 1.96e-16
c2802 2777 2776 5.65e-16
c2803 638 0 1.1593e-14
c2804 1091 1520 1.58e-16
c2805 1023 1 1.56e-15
c2806 4116 1 6.78e-16
c2807 2470 812 3.64e-16
c2808 1806 1414 2.38e-15
c2809 1698 1691 7.37e-16
c2810 4646 1 2.378e-15
c2811 1684 1618 5.5e-16
c2812 1694 2007 1.58e-16
c2813 594 593 6.67e-16
c2814 4742 4746 1.81e-16
c2815 642 2265 2.22e-16
c2816 4645 0 3.466e-15
c2817 1969 1584 1.96e-16
c2818 37 433 5.71e-16
c2819 3723 3409 3.92e-16
c2820 4563 4566 1.96e-16
c2821 5118 5103 7.95e-16
c2822 2303 2304 9.1e-16
c2823 107 117 1.88e-16
c2824 3893 3885 1.606e-15
c2825 4339 692 1.84e-16
c2826 1128 782 1.58e-16
c2827 1822 677 1.9e-16
c2828 1627 842 1.58e-16
c2829 1181 837 3.79e-16
c2830 1440 1016 1.58e-16
c2831 3898 4451 3.92e-16
c2832 2535 2735 3.92e-16
c2833 677 19 1.676e-15
c2834 1573 1956 7.84e-16
c2835 158 163 1.482e-15
c2836 4438 792 1.58e-16
c2837 3437 3438 2.48e-16
c2838 1667 0 5.5851e-14
c2839 1928 1 6.15e-16
c2840 777 1924 2.72e-16
c2841 842 873 1.621e-15
c2842 868 872 2.19e-16
c2843 3693 837 1.58e-16
c2844 5300 5297 3.92e-16
c2845 4827 236 1.88e-16
c2846 4922 4902 1.58e-16
c2847 3900 812 3.15e-16
c2848 4506 868 1.58e-16
c2849 4509 827 1.58e-16
c2850 2851 2850 1.6e-16
c2851 2843 2841 2.15e-16
c2852 3882 3418 1.58e-16
c2853 920 1190 3.92e-16
c2854 921 1189 2.54e-16
c2855 3645 0 1.4092e-14
c2856 952 0 3.7285e-14
c2857 1184 1 3.06e-16
c2858 612 3900 3.58e-16
c2859 4266 1 1.716e-15
c2860 3030 3274 1.58e-16
c2861 4799 0 1.4233e-14
c2862 3393 3390 1.123e-15
c2863 3397 3386 1.58e-16
c2864 3514 3486 2.64e-16
c2865 3110 0 6.62e-16
c2866 921 837 3.15e-16
c2867 1026 1033 7.95e-16
c2868 3463 4302 2.386e-15
c2869 4311 4305 1.6e-16
c2870 4424 752 1.58e-16
c2871 3475 1 2.054e-15
c2872 1907 752 1.9e-16
c2873 1506 1517 1.96e-16
c2874 3477 0 8e-16
c2875 4060 1 4.64e-16
c2876 4679 4299 1.96e-16
c2877 2923 2922 6.26e-16
c2878 2921 2931 1.58e-16
c2879 797 26 7.12e-16
c2880 3034 2583 1.58e-16
c2881 1716 0 1.6491e-14
c2882 2541 807 4.03e-16
c2883 1 382 4.92e-16
c2884 421 252 1.88e-16
c2885 3504 3515 1.96e-16
c2886 4564 0 4.0997e-14
c2887 0 355 1.4515e-14
c2888 281 276 1.88e-16
c2889 4317 677 1.339e-15
c2890 3898 3875 1.58e-16
c2891 3882 3872 3.54e-16
c2892 1166 1164 1.931e-15
c2893 1386 1772 5.66e-16
c2894 2730 0 6.9481e-14
c2895 2559 2683 5.42e-16
c2896 2535 2671 1.58e-16
c2897 992 0 1.0183e-14
c2898 3411 1 2.222e-15
c2899 4386 4385 2.03e-16
c2900 4391 4389 1.6e-16
c2901 3877 0 1.4835e-14
c2902 4415 1 1.056e-15
c2903 1525 0 3.3688e-14
c2904 30 267 3.84e-16
c2905 565 484 1.88e-16
c2906 49 247 1.88e-16
c2907 3526 677 1.58e-16
c2908 762 1901 2.4e-16
c2909 3656 3657 1.35e-16
c2910 4563 4859 1.58e-16
c2911 5170 5171 3.18e-16
c2912 2737 2356 3.92e-16
c2913 1403 662 1.75e-16
c2914 3250 0 8e-16
c2915 2533 1 5.277e-15
c2916 757 1 5.62e-16
c2917 1684 868 3.15e-16
c2918 1708 827 3.15e-16
c2919 1978 812 1.09e-16
c2920 1587 1585 1.6e-16
c2921 528 1 5.848e-15
c2922 1684 1386 1.58e-16
c2923 1690 1380 5.88e-16
c2924 2705 717 1.58e-16
c2925 2178 827 3.15e-16
c2926 1833 1448 1.96e-16
c2927 3048 2713 5.5e-16
c2928 2165 1690 2e-16
c2929 275 274 5.8e-16
c2930 1 117 4.22e-16
c2931 3304 3671 1.58e-16
c2932 3202 3208 1.418e-15
c2933 3589 3591 1.862e-15
c2934 4750 0 8e-16
c2935 3219 3191 2.64e-16
c2936 601 2572 1.84e-16
c2937 5136 5058 1.58e-16
c2938 5051 5059 9.34e-16
c2939 4922 323 1.88e-16
c2940 2441 2435 1.418e-15
c2941 1953 0 3.5724e-14
c2942 2424 2452 2.64e-16
c2943 2446 2442 1.96e-16
c2944 752 745 5.58e-16
c2945 1292 1291 1.6e-16
c2946 1289 1231 3.92e-16
c2947 687 3387 3.15e-16
c2948 506 513 7.76e-16
c2949 146 129 1.325e-15
c2950 2182 827 3.15e-16
c2951 1437 1820 7.84e-16
c2952 3710 0 3.3749e-14
c2953 4004 1 2.259e-15
c2954 4184 19 7.35e-16
c2955 2423 767 1.58e-16
c2956 1755 1363 2.38e-15
c2957 2713 2685 2.64e-16
c2958 1673 0 1.1956e-14
c2959 3591 3590 2.48e-16
c2960 4730 4344 4.11e-16
c2961 4735 4726 3.46e-16
c2962 2557 767 4.46e-16
c2963 777 1327 4.03e-16
c2964 37 21 1.88e-16
c2965 5054 5036 6.67e-16
c2966 3804 3807 5.5e-16
c2967 2333 2731 4.36e-16
c2968 5324 5355 1.58e-16
c2969 2866 858 3.15e-16
c2970 2805 0 1.6491e-14
c2971 4175 4168 1.88e-16
c2972 1471 732 5.73e-16
c2973 2172 2528 3.54e-16
c2974 2194 2178 4.274e-15
c2975 2920 2917 3.54e-16
c2976 2882 2937 1.141e-15
c2977 2545 2819 1.58e-16
c2978 3306 3305 1.6e-16
c2979 2545 2254 1.58e-16
c2980 3785 0 3.0577e-14
c2981 3992 19 7.35e-16
c2982 3211 3210 2.48e-16
c2983 1653 1191 1.96e-16
c2984 1654 1647 6.73e-16
c2985 3876 0 3.12587e-13
c2986 1921 1533 4.97e-16
c2987 1694 1735 1.58e-16
c2988 747 1528 1.58e-16
c2989 1489 0 1.6491e-14
c2990 37 580 1.88e-16
c2991 5010 4549 5.8e-16
c2992 1845 1834 1.58e-16
c2993 4889 4881 5.87e-16
c2994 2635 1 1.716e-15
c2995 883 962 3.92e-16
c2996 890 961 1.58e-16
c2997 215 1 4.59e-16
c2998 4288 647 1.84e-16
c2999 5355 5350 1.493e-15
c3000 5366 5367 3.92e-16
c3001 4827 5031 6.58e-16
c3002 221 0 9.795e-15
c3003 3270 3662 2.38e-15
c3004 3855 852 2.8e-16
c3005 2194 2182 4.369e-15
c3006 2178 2524 6.89e-16
c3007 632 3474 1.9e-16
c3008 3218 1 8.43e-16
c3009 1399 1398 1.6e-16
c3010 1391 1389 2.15e-16
c3011 2172 2342 1.58e-16
c3012 2557 2282 5.5e-16
c3013 2541 2265 5.88e-16
c3014 712 1 5.62e-16
c3015 1794 692 1.58e-16
c3016 1708 812 3.15e-16
c3017 1448 1443 1.642e-15
c3018 3520 0 3.6368e-14
c3019 2178 812 3.15e-16
c3020 612 1708 3.58e-16
c3021 3134 677 3.15e-16
c3022 2781 812 1.58e-16
c3023 2256 1743 4.97e-16
c3024 4446 4808 1.58e-16
c3025 4435 4816 5.66e-16
c3026 4822 4813 3.92e-16
c3027 2696 737 1.58e-16
c3028 1670 2104 3.65e-16
c3029 1 304 1.073e-15
c3030 2418 1 5.97e-15
c3031 1008 647 1.58e-16
c3032 2414 0 6.72e-16
c3033 612 2178 4.03e-16
c3034 602 2172 3.46e-16
c3035 3397 692 3.15e-16
c3036 5535 526 5.5e-16
c3037 3006 1 1.871e-15
c3038 777 1896 1.813e-15
c3039 1913 762 2.22e-16
c3040 1491 722 1.58e-16
c3041 1061 717 3.79e-16
c3042 1226 1222 5.5e-16
c3043 5406 5407 3.54e-16
c3044 3005 0 3.792e-15
c3045 2705 2707 2.15e-16
c3046 2736 2737 1.35e-16
c3047 1473 1475 2.03e-16
c3048 601 1383 4.81e-16
c3049 1964 827 3.15e-16
c3050 2182 812 3.15e-16
c3051 747 1098 1.58e-16
c3052 3288 3277 1.96e-16
c3053 3216 722 1.09e-16
c3054 1862 1471 1.136e-15
c3055 3572 3573 2.03e-16
c3056 612 2182 7.99e-16
c3057 812 1172 1.58e-16
c3058 894 1111 1.58e-16
c3059 907 1083 3.54e-16
c3060 4254 4251 5.5e-16
c3061 3379 1 8e-16
c3062 2771 792 1.58e-16
c3063 1448 707 1.58e-16
c3064 1455 1457 1.862e-15
c3065 878 1 5.1e-16
c3066 601 4237 1.84e-16
c3067 612 4251 1.58e-16
c3068 1879 752 3.15e-16
c3069 2679 3173 1.96e-16
c3070 601 1720 5.03e-16
c3071 1450 1 9.28e-16
c3072 1777 1386 1.136e-15
c3073 4506 0 3.3724e-14
c3074 478 484 3.84e-16
c3075 556 584 3.75e-16
c3076 3900 747 3.58e-16
c3077 5074 1 1.021e-15
c3078 2332 2323 3.46e-16
c3079 1973 1 5.808e-15
c3080 1975 0 3.466e-15
c3081 3393 3654 1.58e-16
c3082 1089 722 8.3e-16
c3083 5321 5316 3.54e-16
c3084 2797 2401 1.96e-16
c3085 5200 5221 1.96e-16
c3086 1998 2491 1.96e-16
c3087 2194 1964 5.5e-16
c3088 389 390 1.482e-15
c3089 4047 4054 2.45e-16
c3090 4872 381 1.88e-16
c3091 1562 782 1.84e-16
c3092 921 1238 2.45e-16
c3093 3911 37 5.71e-16
c3094 4338 4334 1.96e-16
c3095 5509 5513 8.88e-16
c3096 2287 662 7.38e-16
c3097 1343 1131 1.58e-16
c3098 632 1331 3.15e-16
c3099 3030 3343 1.96e-16
c3100 1 325 5.798e-15
c3101 216 218 1.88e-16
c3102 4759 4760 9.93e-16
c3103 3385 3895 2.79e-16
c3104 4036 4037 7.45e-16
c3105 4044 4046 2.239e-15
c3106 3520 3521 1.35e-16
c3107 381 0 1.21533e-13
c3108 2172 1777 5.5e-16
c3109 1222 1224 7.46e-16
c3110 1046 1044 1.931e-15
c3111 3882 692 3.15e-16
c3112 5482 5481 3.92e-16
c3113 5509 5519 1.98e-16
c3114 5422 5426 2.95e-16
c3115 1533 767 3.15e-16
c3116 1091 1525 1.58e-16
c3117 632 3898 4.46e-16
c3118 3874 4577 2.79e-16
c3119 4118 1 7.08e-16
c3120 3684 4501 1.58e-16
c3121 2979 2923 9.34e-16
c3122 2976 2969 3.92e-16
c3123 2954 2981 9.6e-16
c3124 1964 812 3.15e-16
c3125 1057 1 3.54e-16
c3126 1054 0 9.602e-15
c3127 4663 1 2.378e-15
c3128 3190 707 7.38e-16
c3129 3030 2617 1.58e-16
c3130 2120 2119 1.6e-16
c3131 2098 2100 3.54e-16
c3132 1772 0 1.4092e-14
c3133 3168 3535 1.58e-16
c3134 3157 3543 5.66e-16
c3135 3549 3540 3.92e-16
c3136 2177 1 6.056e-15
c3137 4662 0 3.466e-15
c3138 4922 265 1.88e-16
c3139 2392 2393 2.48e-16
c3140 5325 323 3.54e-16
c3141 2174 0 5.96e-16
c3142 146 450 1.88e-16
c3143 3397 3393 4.431e-15
c3144 2873 323 1.707e-15
c3145 4132 4133 7.45e-16
c3146 4140 4142 2.239e-15
c3147 1460 1016 2.38e-15
c3148 2559 2752 3.92e-16
c3149 3839 2892 4.35e-16
c3150 3739 1 4.083e-15
c3151 4088 26 1.075e-15
c3152 3725 0 5.5809e-14
c3153 4693 4694 2.48e-16
c3154 4698 4697 2.83e-16
c3155 4701 4310 1.96e-16
c3156 2662 3155 1.58e-16
c3157 1584 1968 1.58e-16
c3158 1706 1816 3.92e-16
c3159 117 363 1.88e-16
c3160 5074 5081 3.54e-16
c3161 4977 4979 3.73e-16
c3162 3366 858 1.58e-16
c3163 1684 0 3.09567e-13
c3164 1937 1 1.716e-15
c3165 3411 3225 1.58e-16
c3166 4776 410 1.88e-16
c3167 2528 0 2.0654e-14
c3168 3599 3208 1.136e-15
c3169 1540 767 1.339e-15
c3170 3898 3435 1.58e-16
c3171 1146 1593 7.84e-16
c3172 622 1 5.62e-16
c3173 627 3900 3.58e-16
c3174 4292 1 8.43e-16
c3175 1873 1482 4.11e-16
c3176 194 247 1.88e-16
c3177 3046 3291 1.58e-16
c3178 3030 3279 1.58e-16
c3179 3024 672 3.15e-16
c3180 3048 647 3.15e-16
c3181 4816 0 1.4233e-14
c3182 4606 4607 9.93e-16
c3183 4878 33 1.88e-16
c3184 2339 1 4.41e-15
c3185 2488 2487 1.6e-16
c3186 2480 2478 2.15e-16
c3187 2196 2423 3.92e-16
c3188 2342 0 3.3692e-14
c3189 3919 857 1.88e-16
c3190 1743 647 1.58e-16
c3191 919 1040 3.92e-16
c3192 922 1039 2.54e-16
c3193 910 3877 7.06e-16
c3194 3493 0 6.72e-16
c3195 4487 4498 1.96e-16
c3196 2440 807 2.4e-16
c3197 3351 3349 1.6e-16
c3198 3346 3345 2.03e-16
c3199 4751 4745 7.25e-16
c3200 4361 4367 9.42e-16
c3201 3387 3388 1.487e-15
c3202 245 256 2.45e-16
c3203 131 117 1.88e-16
c3204 233 368 1.88e-16
c3205 602 0 3.02143e-13
c3206 26 491 1.03e-15
c3207 0 502 2.87e-16
c3208 19 488 3.2e-16
c3209 5066 5064 8.35e-16
c3210 89 1 1.456e-15
c3211 3910 3907 1.58e-16
c3212 1440 662 1.832e-15
c3213 64 439 1.88e-16
c3214 919 662 3.15e-16
c3215 881 882 5.43e-16
c3216 3886 3884 5.93e-16
c3217 1343 1341 1.96e-16
c3218 1327 1340 1.58e-16
c3219 2579 2578 1.6e-16
c3220 1176 1178 7.72e-16
c3221 657 4304 2.72e-16
c3222 3876 4404 1.58e-16
c3223 3900 4416 5.42e-16
c3224 2559 2688 1.58e-16
c3225 795 1 1.65e-16
c3226 4040 0 2.0592e-14
c3227 4431 1 9.28e-16
c3228 3141 3152 1.96e-16
c3229 320 450 1.88e-16
c3230 5034 5047 1.138e-15
c3231 672 678 1.097e-15
c3232 2119 0 2.078e-15
c3233 244 246 2.84e-16
c3234 2270 1777 1.96e-16
c3235 747 1708 3.58e-16
c3236 883 672 3.15e-16
c3237 909 647 3.15e-16
c3238 2807 822 1.58e-16
c3239 2549 2552 2.109e-15
c3240 4563 4876 1.58e-16
c3241 2675 0 6.72e-16
c3242 2178 747 4.03e-16
c3243 4007 4008 6.4e-16
c3244 3103 1 1.056e-15
c3245 3896 0 1.2366e-14
c3246 4298 3480 1.96e-16
c3247 1321 1504 3.92e-16
c3248 777 779 5.59e-16
c3249 392 397 1.88e-16
c3250 1708 1403 1.58e-16
c3251 1706 1397 5.5e-16
c3252 1359 0 6.72e-16
c3253 3702 1 1.868e-15
c3254 3406 3407 1.736e-15
c3255 2194 852 3.15e-16
c3256 1769 1781 2.32e-16
c3257 3387 3570 3.92e-16
c3258 3676 3304 1.58e-16
c3259 3293 827 1.75e-16
c3260 5177 1 1.113e-15
c3261 2182 747 7.99e-16
c3262 2172 2376 1.58e-16
c3263 2194 2168 1.58e-16
c3264 2172 2171 1.58e-16
c3265 146 137 1.58e-16
c3266 3801 3803 3.54e-16
c3267 4318 3486 2.48e-16
c3268 5442 5449 8.94e-16
c3269 5444 5447 1.342e-15
c3270 2541 2486 5.88e-16
c3271 2954 2503 9.63e-16
c3272 1690 692 3.15e-16
c3273 1327 1503 1.58e-16
c3274 1397 966 1.136e-15
c3275 2248 2254 1.418e-15
c3276 910 3876 5.22e-16
c3277 911 3900 3.45e-16
c3278 1448 1832 1.58e-16
c3279 632 1706 4.46e-16
c3280 1133 0 1.4198e-14
c3281 3508 3123 1.96e-16
c3282 3313 3322 3.92e-16
c3283 3316 2804 5.66e-16
c3284 2815 3308 1.58e-16
c3285 2559 782 3.15e-16
c3286 2285 1 1.056e-15
c3287 792 1343 3.15e-16
c3288 117 310 1.88e-16
c3289 5451 439 3.54e-16
c3290 1777 0 6.909e-14
c3291 842 837 2.77e-16
c3292 920 963 1.58e-16
c3293 4753 410 1.88e-16
c3294 2557 2271 1.58e-16
c3295 2637 2636 2.48e-16
c3296 2649 2282 1.58e-16
c3297 1880 732 2.65e-16
c3298 3029 3027 1.041e-15
c3299 632 966 1.75e-16
c3300 2719 1 4.41e-15
c3301 632 4281 7.38e-16
c3302 2545 2824 1.58e-16
c3303 1759 1363 1.96e-16
c3304 945 19 1.58e-16
c3305 3396 3027 1.176e-15
c3306 3048 3031 3.62e-16
c3307 3046 3038 4.63e-16
c3308 1196 1191 1.58e-16
c3309 3139 647 1.58e-16
c3310 1690 1539 1.58e-16
c3311 429 419 8.86e-16
c3312 1845 2368 4.36e-16
c3313 2366 2359 1.96e-16
c3314 2056 1 7.51e-16
c3315 4531 4894 1.96e-16
c3316 4900 4902 1.134e-15
c3317 2257 2256 2.48e-16
c3318 883 976 1.88e-16
c3319 907 969 1.58e-16
c3320 226 216 8.86e-16
c3321 426 9 5.8e-16
c3322 2634 2635 1.35e-16
c3323 4651 33 1.88e-16
c3324 2911 2913 6.91e-16
c3325 1343 737 4.46e-16
c3326 4372 4370 2.15e-16
c3327 4380 4379 1.6e-16
c3328 4474 812 5.03e-16
c3329 2336 692 4.81e-16
c3330 3215 3213 1.6e-16
c3331 3210 3209 2.03e-16
c3332 3597 1 6.15e-16
c3333 1558 1106 4.97e-16
c3334 1251 1 5.398e-15
c3335 2305 692 2.33e-16
c3336 1431 1 5.97e-15
c3337 627 1708 3.58e-16
c3338 4898 4897 5.87e-16
c3339 3324 812 4.81e-16
c3340 2815 797 1.58e-16
c3341 4446 4825 1.58e-16
c3342 1 33 2.2651e-14
c3343 8 5 2.142e-15
c3344 17 19 8.82e-16
c3345 3387 3506 1.58e-16
c3346 3411 3518 5.42e-16
c3347 3276 3661 1.96e-16
c3348 3270 3666 1.96e-16
c3349 3409 827 4.46e-16
c3350 5257 5259 1.609e-15
c3351 5165 5261 9.36e-16
c3352 1027 662 1.58e-16
c3353 677 1037 1.58e-16
c3354 632 3468 7.38e-16
c3355 627 2178 4.03e-16
c3356 601 2172 4.48e-16
c3357 3293 812 2.33e-16
c3358 4039 857 6.23e-16
c3359 3951 943 2.566e-15
c3360 2426 2428 2.03e-16
c3361 5530 5531 5.87e-16
c3362 3026 0 5.96e-16
c3363 919 1098 1.58e-16
c3364 1550 807 1.58e-16
c3365 1761 1369 1.96e-16
c3366 4609 4621 2.62e-16
c3367 3751 3731 1.69e-16
c3368 4164 1 2.259e-15
c3369 4344 3503 1.136e-15
c3370 3886 4523 1.58e-16
c3371 3876 3684 5.5e-16
c3372 2673 692 5.03e-16
c3373 1107 0 6.29e-16
c3374 4156 25 1.88e-16
c3375 4816 4815 1.6e-16
c3376 4429 4811 1.443e-15
c3377 2291 1783 7.84e-16
c3378 627 2182 7.99e-16
c3379 1 573 1.44e-16
c3380 310 304 3.84e-16
c3381 117 339 1.88e-16
c3382 3661 812 5.03e-16
c3383 2408 2410 1.862e-15
c3384 1896 1902 1.418e-15
c3385 0 570 2.14091e-13
c3386 2342 2344 2.15e-16
c3387 59 5 1.88e-16
c3388 3866 3338 4.69e-16
c3389 4872 5139 5.5e-16
c3390 2800 1 9.28e-16
c3391 2707 2703 1.96e-16
c3392 1865 707 4.81e-16
c3393 1482 692 1.58e-16
c3394 3010 3003 2.15e-16
c3395 627 4251 1.58e-16
c3396 3599 3605 1.418e-15
c3397 4436 4438 1.862e-15
c3398 687 1829 2.65e-16
c3399 2850 842 7.68e-16
c3400 2843 827 1.9e-16
c3401 1694 1499 5.5e-16
c3402 1463 1 6.15e-16
c3403 1993 1 2.054e-15
c3404 1995 0 8e-16
c3405 564 570 3.84e-16
c3406 3393 3659 1.58e-16
c3407 3409 3276 1.58e-16
c3408 5039 31 7.46e-16
c3409 890 905 3.92e-16
c3410 909 915 1.13e-16
c3411 592 847 1.96e-16
c3412 2589 0 1.4092e-14
c3413 4580 5591 4.22e-16
c3414 64 238 1.88e-16
c3415 617 984 8.3e-16
c3416 1223 1 7.34e-16
c3417 2758 767 5.03e-16
c3418 1914 1522 1.96e-16
c3419 1915 1908 6.73e-16
c3420 1694 1695 1.027e-15
c3421 1220 0 1.0077e-14
c3422 1947 1942 1.642e-15
c3423 2158 2078 3.2e-16
c3424 13 565 1.88e-16
c3425 3409 812 4.46e-16
c3426 5492 1 2.424e-15
c3427 5200 5197 7.46e-16
c3428 4793 468 1.88e-16
c3429 2504 2495 3.92e-16
c3430 1987 2498 5.66e-16
c3431 993 999 1.58e-16
c3432 797 787 6.38e-16
c3433 2178 2287 1.96e-16
c3434 1056 1058 7.72e-16
c3435 3876 707 4.48e-16
c3436 2535 2373 1.58e-16
c3437 921 1085 1.96e-16
c3438 612 3409 3.15e-16
c3439 657 3876 3.15e-16
c3440 3684 4506 1.58e-16
c3441 2957 2968 1.138e-15
c3442 911 1708 3.45e-16
c3443 910 1684 5.22e-16
c3444 3089 3090 1.35e-16
c3445 1136 1 5.821e-15
c3446 4680 1 2.378e-15
c3447 657 2633 2.4e-16
c3448 465 459 1.58e-16
c3449 426 419 7.76e-16
c3450 423 424 6.67e-16
c3451 4679 0 3.466e-15
c3452 314 303 2.45e-16
c3453 19 197 8.82e-16
c3454 3168 3540 1.58e-16
c3455 2376 0 3.3588e-14
c3456 911 2178 7.6e-16
c3457 3785 3775 7.84e-16
c3458 4827 178 1.88e-16
c3459 2182 2287 4.63e-16
c3460 107 479 1.88e-16
c3461 3520 707 1.75e-16
c3462 1147 1149 7.84e-16
c3463 4236 4234 2.15e-16
c3464 4244 4243 1.6e-16
c3465 2595 2586 3.92e-16
c3466 2203 2589 5.66e-16
c3467 1439 1011 2.48e-16
c3468 850 1 3.79e-16
c3469 3910 1 4.45e-16
c3470 1982 1976 1.6e-16
c3471 1584 1973 2.386e-15
c3472 1601 1956 1.58e-16
c3473 1684 1833 3.92e-16
c3474 1016 1 5.821e-15
c3475 632 26 7.12e-16
c3476 5127 5074 3.18e-16
c3477 5125 5113 1.96e-16
c3478 911 2182 3.45e-16
c3479 5420 5404 7.48e-16
c3480 107 189 1.88e-16
c3481 592 802 1.96e-16
c3482 2586 2588 2.15e-16
c3483 4150 857 1.88e-16
c3484 361 15 5.8e-16
c3485 378 1 4.22e-16
c3486 5580 5581 1.6e-16
c3487 4520 5579 2.91e-16
c3488 595 3018 1.655e-15
c3489 602 3430 3.64e-16
c3490 2798 0 6.9481e-14
c3491 2856 2867 1.96e-16
c3492 2617 2618 1.35e-16
c3493 3882 3446 5.88e-16
c3494 3876 3452 1.58e-16
c3495 4318 4320 2.03e-16
c3496 2557 2531 1.58e-16
c3497 2535 2534 1.58e-16
c3498 2257 647 1.58e-16
c3499 1151 1605 1.58e-16
c3500 3066 3434 1.96e-16
c3501 602 910 4.07e-16
c3502 181 180 3.84e-16
c3503 3024 3308 1.58e-16
c3504 3046 3296 1.58e-16
c3505 2206 2208 2.15e-16
c3506 4833 0 1.4233e-14
c3507 2095 2078 1.96e-16
c3508 2080 2082 7.3e-16
c3509 3387 782 4.48e-16
c3510 5193 5192 8.03e-16
c3511 2628 0 6.8998e-14
c3512 922 827 5.14e-16
c3513 4430 767 7.68e-16
c3514 5486 5479 9.81e-16
c3515 4787 5239 9.98e-16
c3516 4861 149 1.88e-16
c3517 3073 3074 2.03e-16
c3518 1532 1076 1.96e-16
c3519 1527 1086 1.96e-16
c3520 1315 1316 1.76e-16
c3521 4268 0 3.3724e-14
c3522 1737 0 3.466e-15
c3523 4378 4367 1.58e-16
c3524 3409 3406 1.58e-16
c3525 3160 692 1.58e-16
c3526 2074 2069 3.07e-16
c3527 601 0 2.79469e-13
c3528 4708 4714 5.87e-16
c3529 2196 2422 5.42e-16
c3530 3525 3140 1.96e-16
c3531 5529 497 5.11e-16
c3532 5257 1 1.88e-16
c3533 747 2379 1.58e-16
c3534 1879 2372 1.96e-16
c3535 2340 0 1.6491e-14
c3536 910 3896 1.58e-16
c3537 4568 3890 1.018e-15
c3538 2857 2469 4.97e-16
c3539 2654 2652 1.862e-15
c3540 1327 880 1.58e-16
c3541 4327 3486 1.136e-15
c3542 3900 4421 1.58e-16
c3543 2622 647 5.03e-16
c3544 1397 1789 2.38e-15
c3545 642 920 3.15e-16
c3546 805 1 3.79e-16
c3547 2892 1 1.113e-15
c3548 3030 3105 1.96e-16
c3549 4444 1 6.15e-16
c3550 2803 797 7.38e-16
c3551 2545 647 3.15e-16
c3552 1684 1798 1.58e-16
c3553 2384 2379 1.642e-15
c3554 4440 777 2.72e-16
c3555 3532 692 7.68e-16
c3556 3024 797 4.48e-16
c3557 2274 2272 1.862e-15
c3558 1766 1760 1.418e-15
c3559 894 662 3.15e-16
c3560 275 273 2.84e-16
c3561 3712 868 2.72e-16
c3562 2827 822 1.58e-16
c3563 3397 3208 1.58e-16
c3564 4563 4893 1.58e-16
c3565 4736 468 1.88e-16
c3566 2567 2571 1.96e-16
c3567 2511 1 4.03e-16
c3568 4124 4127 4.41e-16
c3569 4657 497 1.88e-16
c3570 3263 0 6.62e-16
c3571 3565 4382 1.58e-16
c3572 3554 4390 5.66e-16
c3573 4396 4387 3.92e-16
c3574 5536 5561 1.58e-16
c3575 2545 2492 1.58e-16
c3576 3628 1 2.054e-15
c3577 3893 0 5.4943e-14
c3578 1345 1521 3.92e-16
c3579 3634 777 2.65e-16
c3580 4980 4978 5.88e-16
c3581 4549 3744 6.11e-16
c3582 3839 3751 1.02e-15
c3583 3245 752 1.832e-15
c3584 3034 2736 1.58e-16
c3585 762 1905 1.58e-16
c3586 1 479 3.0375e-14
c3587 3411 3587 3.92e-16
c3588 4582 4480 5.5e-16
c3589 4861 4866 5.53e-16
c3590 5262 5174 1.237e-15
c3591 692 702 3.28e-16
c3592 601 2203 2.33e-16
c3593 595 2214 2.22e-16
c3594 461 19 3.45e-16
c3595 4046 3918 6.32e-16
c3596 4878 526 1.88e-16
c3597 1236 596 2.9e-16
c3598 4793 64 1.88e-16
c3599 922 812 5.14e-16
c3600 921 1143 1.58e-16
c3601 602 884 5.47e-16
c3602 1684 707 4.48e-16
c3603 542 27 1.88e-16
c3604 3627 777 2.72e-16
c3605 1846 1840 1.6e-16
c3606 1448 1837 2.386e-15
c3607 1465 1820 1.58e-16
c3608 657 1684 3.15e-16
c3609 4030 1 6.76e-16
c3610 4473 4470 6.44e-16
c3611 4477 4474 3.01e-16
c3612 612 922 3.15e-16
c3613 3313 2815 1.58e-16
c3614 2301 1 9.28e-16
c3615 1694 1952 4.63e-16
c3616 1 189 1.1938e-14
c3617 100 37 1.88e-16
c3618 4567 4707 3.92e-16
c3619 3617 752 3.64e-16
c3620 381 441 1.58e-16
c3621 3808 3811 1.931e-15
c3622 3003 2486 1.885e-15
c3623 2749 2748 1.6e-16
c3624 883 797 6.45e-16
c3625 909 1157 4.35e-16
c3626 907 1156 1.88e-16
c3627 890 1149 1.58e-16
c3628 2663 1 1.868e-15
c3629 3327 3713 5.66e-16
c3630 1871 737 1.58e-16
c3631 1499 732 3.79e-16
c3632 632 1415 3.64e-16
c3633 4606 5561 5.5e-16
c3634 4589 5538 4.06e-16
c3635 3744 3734 1.58e-16
c3636 4024 1 5.1e-16
c3637 3311 3322 1.96e-16
c3638 2401 797 1.58e-16
c3639 2413 782 1.84e-16
c3640 4005 19 9.67e-16
c3641 2342 707 1.832e-15
c3642 1196 1674 4.69e-16
c3643 1659 1664 2.029e-15
c3644 1508 1 5.808e-15
c3645 4546 4543 8.32e-16
c3646 1706 1556 1.58e-16
c3647 3131 3128 3.01e-16
c3648 762 1086 5.73e-16
c3649 1510 0 3.466e-15
c3650 3610 752 1.9e-16
c3651 5056 5048 3.92e-16
c3652 3390 3398 3.84e-16
c3653 890 963 3.54e-16
c3654 909 984 1.58e-16
c3655 3469 647 2.33e-16
c3656 282 0 1.0822e-14
c3657 281 27 1.88e-16
c3658 3685 3293 1.96e-16
c3659 1345 752 3.15e-16
c3660 1404 1415 1.96e-16
c3661 4494 812 1.09e-16
c3662 2541 2650 1.96e-16
c3663 941 25 7.64e-16
c3664 3409 747 3.15e-16
c3665 1295 1 8.135e-15
c3666 1925 1922 5.5e-16
c3667 1848 1 1.056e-15
c3668 4904 4907 2.208e-15
c3669 4452 4833 5.66e-16
c3670 4839 4830 3.92e-16
c3671 229 19 3.45e-16
c3672 3411 3523 1.58e-16
c3673 3397 3536 4.63e-16
c3674 5543 1 2.102e-15
c3675 1936 1 4.41e-15
c3676 2445 0 6.62e-16
c3677 617 2172 4.48e-16
c3678 147 1 1.456e-15
c3679 657 1006 1.35e-16
c3680 146 26 8.41e-16
c3681 140 0 6.224e-15
c3682 4284 4283 2.03e-16
c3683 4289 4287 1.6e-16
c3684 3122 2628 1.96e-16
c3685 1380 1369 1.58e-16
c3686 3604 762 2.4e-16
c3687 4550 4540 1.65e-16
c3688 3701 3900 5.5e-16
c3689 4606 4617 4.67e-16
c3690 4623 4634 4.67e-16
c3691 4640 4651 4.67e-16
c3692 4657 4668 4.67e-16
c3693 2693 692 1.09e-16
c3694 2498 842 1.58e-16
c3695 2787 3298 1.96e-16
c3696 3660 3657 6.44e-16
c3697 3664 3661 3.01e-16
c3698 4333 0 3.6274e-14
c3699 2009 2005 1.96e-16
c3700 1642 0 1.6491e-14
c3701 19 291 3.84e-16
c3702 891 901 1.008e-15
c3703 3393 702 4.03e-16
c3704 3681 812 1.09e-16
c3705 3972 3974 4.33e-16
c3706 4708 439 1.88e-16
c3707 378 363 1.88e-16
c3708 1179 1186 2.27e-16
c3709 894 1098 3.54e-16
c3710 986 963 6.54e-16
c3711 238 234 6.38e-16
c3712 4640 1 1.262e-14
c3713 2792 792 2.72e-16
c3714 1485 1483 1.6e-16
c3715 908 1 2.508e-15
c3716 3984 1 1.4213e-14
c3717 627 4271 1.58e-16
c3718 3882 4349 1.96e-16
c3719 2391 767 1.339e-15
c3720 687 1448 3.79e-16
c3721 1731 1319 1.96e-16
c3722 3696 0 1.4092e-14
c3723 3109 647 1.58e-16
c3724 2860 868 2.72e-16
c3725 2289 1783 3.92e-16
c3726 1472 1 1.716e-15
c3727 3100 3106 1.418e-15
c3728 3487 3489 1.862e-15
c3729 204 186 1.58e-16
c3730 4915 236 1.88e-16
c3731 4915 4928 3.18e-16
c3732 2322 2350 2.64e-16
c3733 2344 2340 1.96e-16
c3734 1103 737 3.57e-16
c3735 1083 1096 1.58e-16
c3736 4 1 4.59e-16
c3737 4651 526 1.88e-16
c3738 886 0 8.2827e-14
c3739 4736 64 1.88e-16
c3740 2541 2615 1.58e-16
c3741 1321 1136 5.5e-16
c3742 1331 1593 1.58e-16
c3743 3484 3117 1.58e-16
c3744 3503 1 4.41e-15
c3745 657 1777 3.79e-16
c3746 1690 1691 1.239e-15
c3747 4337 0 6.62e-16
c3748 3481 647 7.68e-16
c3749 3048 3360 3.92e-16
c3750 911 2168 1.88e-16
c3751 3253 3638 1.96e-16
c3752 2072 2117 1.817e-15
c3753 1012 1014 7.84e-16
c3754 1 526 3.36e-15
c3755 9 513 5.8e-16
c3756 3411 837 3.58e-16
c3757 4702 4316 1.179e-15
c3758 5229 5226 3.54e-16
c3759 1998 2495 1.58e-16
c3760 94 89 1.059e-15
c3761 4004 857 1.88e-16
c3762 2194 2304 3.92e-16
c3763 75 1 4.22e-16
c3764 5525 5296 1.33e-16
c3765 920 1099 1.58e-16
c3766 627 3409 3.15e-16
c3767 1551 1101 1.96e-16
c3768 1552 1545 6.73e-16
c3769 1321 1016 5.5e-16
c3770 1343 1001 5.5e-16
c3771 4590 3873 3.92e-16
c3772 4602 4601 1.6e-16
c3773 2048 2518 1.96e-16
c3774 2136 2521 1.96e-16
c3775 2667 677 7.38e-16
c3776 612 971 4.21e-16
c3777 4866 4486 1.96e-16
c3778 1621 1 1.056e-15
c3779 3393 3485 1.96e-16
c3780 3387 3134 5.5e-16
c3781 4697 1 2.378e-15
c3782 2117 2125 1.96e-16
c3783 4696 0 3.466e-15
c3784 4776 4780 1.81e-16
c3785 5226 5227 3.54e-16
c3786 511 513 1.257e-15
c3787 26 320 8.41e-16
c3788 3168 3560 2.38e-15
c3789 4759 352 1.88e-16
c3790 149 209 1.58e-16
c3791 5044 120 1.58e-16
c3792 920 732 3.15e-16
c3793 3321 868 1.813e-15
c3794 4379 707 3.64e-16
c3795 5303 5283 1.58e-16
c3796 4776 5160 2.45e-16
c3797 2687 2689 2.03e-16
c3798 3524 0 6.62e-16
c3799 2769 777 2.4e-16
c3800 2214 2586 1.58e-16
c3801 1653 858 7.68e-16
c3802 78 72 3.84e-16
c3803 2985 2887 3.87e-16
c3804 3712 0 3.466e-15
c3805 3739 410 3.39e-16
c3806 4124 25 1.88e-16
c3807 4420 3588 2.48e-16
c3808 5026 180 1.188e-15
c3809 4489 1 5.808e-15
c3810 2557 717 3.15e-16
c3811 1708 1850 3.92e-16
c3812 4491 0 3.466e-15
c3813 3393 3869 2e-16
c3814 4685 4299 1.179e-15
c3815 4970 4969 1.6e-16
c3816 4943 4941 1.471e-15
c3817 3048 868 3.58e-16
c3818 2232 2223 3.92e-16
c3819 1715 2226 5.66e-16
c3820 1726 2218 1.58e-16
c3821 612 3055 1.58e-16
c3822 601 3430 7.68e-16
c3823 602 3022 1.58e-16
c3824 3143 1 5.808e-15
c3825 1561 767 1.9e-16
c3826 4634 5471 1.96e-16
c3827 3839 3807 1.58e-16
c3828 3145 0 3.466e-15
c3829 1315 1680 4.65e-16
c3830 919 1219 1.58e-16
c3831 2559 2166 1.58e-16
c3832 2277 647 1.58e-16
c3833 2274 672 1.58e-16
c3834 1619 1613 1.6e-16
c3835 1151 1610 2.386e-15
c3836 1166 1593 1.58e-16
c3837 601 972 4.98e-16
c3838 1684 1832 1.58e-16
c3839 1706 1820 1.58e-16
c3840 2752 752 7.38e-16
c3841 1895 1886 3.46e-16
c3842 484 262 1.88e-16
c3843 747 922 3.15e-16
c3844 3048 3325 5.42e-16
c3845 3024 3313 1.58e-16
c3846 1939 0 3.3874e-14
c3847 3236 3620 1.58e-16
c3848 2544 0 1.5577e-14
c3849 448 456 2.218e-15
c3850 1 206 4.92e-16
c3851 4567 4367 1.58e-16
c3852 4821 439 1.88e-16
c3853 642 3030 4.03e-16
c3854 1327 647 3.15e-16
c3855 877 880 1.606e-15
c3856 3599 767 3.15e-16
c3857 5513 381 3.54e-16
c3858 919 852 3.15e-16
c3859 3497 3469 2.64e-16
c3860 3678 0 3.466e-15
c3861 4226 4225 5.5e-16
c3862 1331 1385 4.63e-16
c3863 2577 3071 1.96e-16
c3864 4288 0 1.4092e-14
c3865 4508 3673 1.96e-16
c3866 4513 3667 1.96e-16
c3867 2248 647 3.15e-16
c3868 2208 2204 1.96e-16
c3869 1757 0 8e-16
c3870 4395 4367 2.64e-16
c3871 4768 4762 7.25e-16
c3872 4378 4384 9.42e-16
c3873 3409 3021 1.58e-16
c3874 3393 3421 1.58e-16
c3875 3180 692 1.58e-16
c3876 642 2620 1.58e-16
c3877 632 2606 1.84e-16
c3878 2080 2067 8.07e-16
c3879 2031 2029 1.96e-16
c3880 1635 1624 1.58e-16
c3881 1 442 5.62e-16
c3882 617 0 2.80251e-13
c3883 4725 4728 6.02e-16
c3884 2196 2427 1.58e-16
c3885 19 430 3.2e-16
c3886 777 2367 1.58e-16
c3887 2172 1743 5.5e-16
c3888 3781 3867 4.06e-16
c3889 909 868 3.15e-16
c3890 592 807 5.8e-16
c3891 1145 782 5.74e-16
c3892 957 959 6.13e-16
c3893 911 3409 9.54e-16
c3894 662 1 3.1284e-14
c3895 1442 1001 4.11e-16
c3896 1181 1177 3.78e-16
c3897 4310 4305 1.642e-15
c3898 3882 3605 1.58e-16
c3899 2642 647 1.09e-16
c3900 2444 807 1.58e-16
c3901 3279 792 1.58e-16
c3902 1008 0 4.6535e-14
c3903 824 1 7.18e-16
c3904 120 180 3.45e-16
c3905 2535 677 4.48e-16
c3906 1955 1956 2.48e-16
c3907 3521 3524 6.44e-16
c3908 5069 5081 8.45e-16
c3909 5032 5034 1.96e-16
c3910 1257 1 1.113e-15
c3911 3542 702 2.72e-16
c3912 3151 692 3.15e-16
c3913 5358 265 1.58e-16
c3914 3347 868 1.58e-16
c3915 2768 2384 1.58e-16
c3916 2706 0 6.62e-16
c3917 1806 677 1.84e-16
c3918 986 1426 2.38e-15
c3919 642 890 3.35e-16
c3920 3278 0 2.93e-15
c3921 3107 1 1.716e-15
c3922 1338 1330 1.606e-15
c3923 2846 2843 3.01e-16
c3924 2842 2839 6.44e-16
c3925 2350 737 3.15e-16
c3926 2545 2316 5.5e-16
c3927 2362 722 1.58e-16
c3928 804 1 5.57e-16
c3929 1381 1 1.868e-15
c3930 3253 777 3.79e-16
c3931 3236 792 1.58e-16
c3932 1371 0 2.93e-15
c3933 4434 777 2.4e-16
c3934 3018 3424 2.38e-15
c3935 4903 4907 1.96e-16
c3936 1903 0 1.6491e-14
c3937 4582 4497 5.5e-16
c3938 3397 3398 1.027e-15
c3939 617 2203 1.75e-16
c3940 2325 1 5.808e-15
c3941 4118 857 1.88e-16
c3942 4759 294 1.88e-16
c3943 4770 352 1.88e-16
c3944 2194 1885 1.58e-16
c3945 4674 5517 1.628e-15
c3946 2559 2503 3.92e-16
c3947 2518 2004 1.958e-15
c3948 781 25 7.64e-16
c3949 389 391 2.84e-16
c3950 379 383 6.38e-16
c3951 3480 4302 1.58e-16
c3952 3142 3144 2.03e-16
c3953 1973 837 1.58e-16
c3954 1345 1520 5.42e-16
c3955 1321 1508 1.58e-16
c3956 1504 1061 1.96e-16
c3957 627 922 3.15e-16
c3958 4059 1 6.78e-16
c3959 3333 2815 2.38e-15
c3960 1725 1 8.43e-16
c3961 3700 3304 1.96e-16
c3962 1714 0 3.22e-16
c3963 4581 1 2.471e-15
c3964 3370 3378 4.06e-16
c3965 2314 1 6.15e-16
c3966 479 310 1.88e-16
c3967 5158 5169 1.37e-16
c3968 0 360 9.795e-15
c3969 3236 737 1.58e-16
c3970 4417 737 1.58e-16
c3971 4691 5300 3.92e-16
c3972 2858 1 5.808e-15
c3973 1173 827 1.58e-16
c3974 894 1172 3.92e-16
c3975 909 1171 1.88e-16
c3976 883 1164 1.58e-16
c3977 2860 0 3.466e-15
c3978 922 993 1.58e-16
c3979 281 282 6.96e-16
c3980 5358 5324 1.58e-16
c3981 2657 2265 2.38e-15
c3982 1891 737 1.58e-16
c3983 642 986 3.79e-16
c3984 3731 3726 1.078e-15
c3985 3256 1 1.056e-15
c3986 2435 782 1.58e-16
c3987 1771 1380 4.11e-16
c3988 4463 4856 1.914e-15
c3989 2719 3227 2.48e-16
c3990 3024 3070 1.58e-16
c3991 3046 3058 1.58e-16
c3992 3021 3020 3.54e-16
c3993 1528 1 2.054e-15
c3994 1530 0 8e-16
c3995 4915 4905 1.58e-16
c3996 657 2628 3.79e-16
c3997 5286 352 7.46e-16
c3998 911 3020 1.88e-16
c3999 883 978 3.54e-16
c4000 894 999 1.58e-16
c4001 596 936 2.85e-16
c4002 412 413 3.84e-16
c4003 3463 662 1.58e-16
c4004 2833 2435 4.36e-16
c4005 3755 3736 6.67e-16
c4006 2967 2966 1.6e-16
c4007 632 4285 1.832e-15
c4008 1304 1270 7.53e-16
c4009 1297 1218 7.01e-16
c4010 1327 1656 1.58e-16
c4011 759 1 5.57e-16
c4012 632 1754 5.03e-16
c4013 2801 782 4.81e-16
c4014 1322 0 1.4835e-14
c4015 3751 1 5.21e-16
c4016 1760 2253 1.96e-16
c4017 1864 1 9.28e-16
c4018 3393 3151 5.88e-16
c4019 3287 3678 4.11e-16
c4020 687 2680 2.65e-16
c4021 2470 1 1.868e-15
c4022 427 0 1.0822e-14
c4023 1 135 9.8e-16
c4024 410 33 2.84e-16
c4025 4079 4088 3.84e-16
c4026 2460 0 2.93e-15
c4027 5051 5050 1.062e-15
c4028 1517 737 7.68e-16
c4029 1331 898 1.58e-16
c4030 1275 1278 7.27e-16
c4031 1284 1226 1.96e-16
c4032 5535 5555 9.6e-16
c4033 5548 5529 5.82e-16
c4034 5514 5522 3.258e-15
c4035 4922 381 1.88e-16
c4036 736 25 7.64e-16
c4037 1562 1559 5.5e-16
c4038 1331 1041 1.58e-16
c4039 4626 4638 2.62e-16
c4040 506 517 2.45e-16
c4041 4190 1 6.76e-16
c4042 2493 852 1.58e-16
c4043 1819 1820 2.48e-16
c4044 1098 1 1.56e-15
c4045 3321 0 6.9481e-14
c4046 3034 3224 4.63e-16
c4047 1661 1 6.636e-15
c4048 4833 4832 1.6e-16
c4049 4446 4828 1.443e-15
c4050 1635 1708 5.5e-16
c4051 2159 2151 1.65e-16
c4052 4350 0 3.5736e-14
c4053 5232 5275 1.617e-15
c4054 31 30 3.84e-16
c4055 45 49 1.58e-16
c4056 479 339 1.88e-16
c4057 5291 1 4.669e-15
c4058 2438 2436 1.6e-16
c4059 3480 3475 1.642e-15
c4060 5046 5045 1.6e-16
c4061 3361 3370 1.37e-16
c4062 2814 1 8.43e-16
c4063 1173 812 1.58e-16
c4064 4396 732 2.65e-16
c4065 910 886 1.977e-15
c4066 4171 4172 4.41e-16
c4067 5375 5353 1.74e-16
c4068 5360 5352 3.54e-16
c4069 3382 1 1.96e-16
c4070 627 633 1.097e-15
c4071 3048 0 3.44963e-13
c4072 2929 2900 1.37e-16
c4073 911 922 1.251e-15
c4074 752 19 1.676e-15
c4075 3998 1 6.76e-16
c4076 4165 19 9.67e-16
c4077 3898 4366 3.92e-16
c4078 3301 3298 3.01e-16
c4079 3297 3294 6.44e-16
c4080 3734 0 3.8149e-14
c4081 1646 1642 1.96e-16
c4082 3900 1 2.222e-15
c4083 4718 4711 1.96e-16
c4084 4327 4720 1.914e-15
c4085 3034 3032 5.93e-16
c4086 1498 1 8.43e-16
c4087 3707 0 3.7647e-14
c4088 1743 0 6.9481e-14
c4089 1624 1 4.41e-15
c4090 26 577 1.03e-15
c4091 3857 3860 1.6e-16
c4092 5183 1 3.36e-16
c4093 5010 4991 1.58e-16
c4094 5171 0 2.156e-15
c4095 2008 0 6.62e-16
c4096 1103 1104 1.213e-15
c4097 4167 4168 6.4e-16
c4098 4770 294 1.88e-16
c4099 4668 5388 1.96e-16
c4100 1121 797 1.58e-16
c4101 1394 1391 3.01e-16
c4102 1390 1387 6.44e-16
c4103 3882 4348 1.58e-16
c4104 2685 0 3.519e-14
c4105 3951 37 1.88e-16
c4106 2557 2632 1.58e-16
c4107 2541 2620 1.58e-16
c4108 1345 1151 5.5e-16
c4109 714 1 5.57e-16
c4110 3120 3118 1.6e-16
c4111 3489 3117 1.58e-16
c4112 4362 1 1.868e-15
c4113 204 252 1.88e-16
c4114 450 368 1.88e-16
c4115 4352 0 2.93e-15
c4116 564 580 3.84e-16
c4117 3100 647 3.15e-16
c4118 3030 732 4.03e-16
c4119 2899 2879 1.69e-16
c4120 2892 2896 3.01e-16
c4121 1025 647 1.58e-16
c4122 1 306 1.65e-15
c4123 4810 4429 5.2e-16
c4124 5492 410 7.62e-16
c4125 5303 1 1.113e-15
c4126 2525 2515 7.29e-16
c4127 2510 2512 2.861e-15
c4128 2172 2321 3.92e-16
c4129 3179 0 3.466e-15
c4130 1061 1057 3.78e-16
c4131 2957 0 4.0391e-14
c4132 687 3876 3.15e-16
c4133 3591 747 1.58e-16
c4134 4533 4526 6.73e-16
c4135 4532 3690 1.96e-16
c4136 627 971 3.79e-16
c4137 909 0 3.3925e-13
c4138 3034 3160 1.58e-16
c4139 1637 1 9.28e-16
c4140 4793 4795 4.93e-16
c4141 0 541 1.5723e-14
c4142 33 556 6.83e-16
c4143 37 552 1.88e-16
c4144 27 565 1.88e-16
c4145 4582 4605 3.92e-16
c4146 5425 468 9.42e-16
c4147 3706 3338 1.96e-16
c4148 3951 3959 3.45e-16
c4149 1162 1163 7.46e-16
c4150 392 262 1.88e-16
c4151 3702 837 2.65e-16
c4152 4249 4260 1.96e-16
c4153 3548 692 1.58e-16
c4154 2015 2196 3.92e-16
c4155 2214 2606 2.38e-15
c4156 3539 0 2.93e-15
c4157 2518 2990 5.5e-16
c4158 1196 858 3.15e-16
c4159 1206 1209 1.58e-16
c4160 3347 0 3.3749e-14
c4161 3928 1 5.1e-16
c4162 1721 1727 1.6e-16
c4163 1718 1315 2.386e-15
c4164 4509 1 2.054e-15
c4165 3186 2668 1.96e-16
c4166 3187 3180 6.73e-16
c4167 5144 5010 1.37e-15
c4168 911 2538 1.58e-16
c4169 884 886 1.013e-15
c4170 717 719 5.59e-16
c4171 3471 3089 2.48e-16
c4172 4511 0 8e-16
c4173 2207 0 6.62e-16
c4174 565 570 1.88e-16
c4175 3168 732 1.58e-16
c4176 2324 2326 2.03e-16
c4177 890 732 3.35e-16
c4178 5116 0 1.65e-16
c4179 1726 2223 1.58e-16
c4180 1440 1452 2.32e-16
c4181 4047 4055 3.45e-16
c4182 601 3022 3.15e-16
c4183 627 3055 5.73e-16
c4184 1121 1125 2.03e-16
c4185 3900 3463 5.5e-16
c4186 3701 852 1.13e-15
c4187 3143 2634 7.84e-16
c4188 2883 2884 5.87e-16
c4189 2815 2424 1.136e-15
c4190 1716 1318 3.92e-16
c4191 919 922 4.274e-15
c4192 3911 0 2.0592e-14
c4193 2294 672 1.58e-16
c4194 1708 1849 5.42e-16
c4195 1684 1837 1.58e-16
c4196 1901 1900 9.1e-16
c4197 4941 4946 7.46e-16
c4198 1794 1800 1.418e-15
c4199 3048 3330 1.58e-16
c4200 3046 692 4.46e-16
c4201 3034 702 7.99e-16
c4202 2232 2221 1.96e-16
c4203 596 820 2.45e-16
c4204 3253 3608 1.58e-16
c4205 4164 857 1.88e-16
c4206 4657 4276 5.2e-16
c4207 4567 4384 1.58e-16
c4208 632 3024 4.48e-16
c4209 2299 2294 1.642e-15
c4210 1321 662 4.48e-16
c4211 881 1320 1.62e-16
c4212 396 15 6.58e-16
c4213 4674 5514 5.5e-16
c4214 2172 2257 1.58e-16
c4215 389 0 9.795e-15
c4216 375 26 1.03e-15
c4217 397 27 1.88e-16
c4218 4804 5051 1.96e-16
c4219 4330 4328 1.6e-16
c4220 2272 672 1.58e-16
c4221 3517 1 1.056e-15
c4222 3698 0 8e-16
c4223 2288 2671 7.84e-16
c4224 646 25 7.64e-16
c4225 4119 1 4.45e-16
c4226 3034 2804 1.58e-16
c4227 3254 3248 1.6e-16
c4228 2730 3245 2.386e-15
c4229 1773 0 6.72e-16
c4230 4395 4384 1.58e-16
c4231 3175 717 1.58e-16
c4232 2557 842 4.46e-16
c4233 2545 868 7.99e-16
c4234 552 548 1.58e-16
c4235 3542 3151 4.11e-16
c4236 3625 782 1.58e-16
c4237 762 1868 5.73e-16
c4238 5505 5491 1.96e-16
c4239 5481 5452 1.58e-16
c4240 1026 702 5.73e-16
c4241 894 852 8.34e-16
c4242 595 3060 2.72e-16
c4243 612 3056 1.58e-16
c4244 4349 702 2.4e-16
c4245 1345 952 1.58e-16
c4246 1343 881 5.5e-16
c4247 2798 2793 1.642e-15
c4248 2634 662 2.33e-16
c4249 4070 19 7.04e-16
c4250 4085 0 1.5176e-14
c4251 1691 1693 3.67e-16
c4252 2736 3243 3.92e-16
c4253 3248 3247 1.6e-16
c4254 3048 3122 3.92e-16
c4255 2071 2067 3.54e-16
c4256 1106 0 7.4135e-14
c4257 1708 1 2.222e-15
c4258 5074 5064 1.021e-15
c4259 5072 5093 1.96e-16
c4260 1879 2376 1.58e-16
c4261 1641 0 3.7647e-14
c4262 4944 4977 1.58e-16
c4263 4982 4981 5.07e-16
c4264 2731 1 1.868e-15
c4265 907 692 4.8e-16
c4266 883 1052 3.92e-16
c4267 890 1051 1.88e-16
c4268 2721 0 2.93e-15
c4269 2178 1 2.824e-15
c4270 2781 1 5.97e-15
c4271 632 883 6.45e-16
c4272 1555 752 1.58e-16
c4273 3807 1 4.651e-15
c4274 2756 2768 2.32e-16
c4275 3344 0 3.7647e-14
c4276 1592 1593 2.48e-16
c4277 2807 797 1.832e-15
c4278 2722 737 1.58e-16
c4279 175 252 1.88e-16
c4280 3536 702 2.4e-16
c4281 3345 852 1.58e-16
c4282 642 1726 1.58e-16
c4283 2736 767 1.75e-16
c4284 2186 2179 7.37e-16
c4285 2182 1 4.57e-15
c4286 596 775 2.45e-16
c4287 3606 3219 1.532e-15
c4288 617 2612 3.64e-16
c4289 601 2231 1.58e-16
c4290 2510 0 1.7608e-14
c4291 3397 767 3.15e-16
c4292 3722 3393 1.58e-16
c4293 4844 0 3.00416e-13
c4294 2483 2480 3.01e-16
c4295 2479 2476 6.44e-16
c4296 2905 1 7.49e-16
c4297 1993 837 1.58e-16
c4298 1345 1525 1.58e-16
c4299 3486 1 4.41e-15
c4300 4251 1 5.808e-15
c4301 2529 3061 2.38e-15
c4302 687 1684 3.15e-16
c4303 4253 0 3.466e-15
c4304 3030 3258 1.96e-16
c4305 1 494 4.22e-16
c4306 120 123 4.6e-16
c4307 276 262 1.88e-16
c4308 3219 3607 4.97e-16
c4309 3881 3401 9.72e-16
c4310 2652 2271 3.92e-16
c4311 627 2605 2.72e-16
c4312 2323 1 1.716e-15
c4313 857 850 4.19e-16
c4314 0 485 1.0822e-14
c4315 3910 857 6.23e-16
c4316 4708 5345 3.92e-16
c4317 2754 2765 1.96e-16
c4318 1445 662 1.09e-16
c4319 1217 842 1.58e-16
c4320 894 1186 1.58e-16
c4321 907 1158 3.54e-16
c4322 3072 0 3.6368e-14
c4323 910 1322 7.06e-16
c4324 999 1 2.972e-15
c4325 4037 1 7.71e-16
c4326 3639 4472 7.84e-16
c4327 3337 2815 1.96e-16
c4328 3332 2821 1.96e-16
c4329 1000 0 6.29e-16
c4330 3048 3087 5.42e-16
c4331 3024 3075 1.58e-16
c4332 3022 3023 3.36e-16
c4333 1684 1567 5.5e-16
c4334 1694 1956 1.58e-16
c4335 1567 1935 1.96e-16
c4336 19 168 8.82e-16
c4337 3820 3821 1.353e-15
c4338 5158 1 1.0125e-14
c4339 5062 5065 1.98e-16
c4340 1119 767 1.58e-16
c4341 165 166 6.96e-16
c4342 4690 677 1.23e-16
c4343 2559 2667 3.92e-16
c4344 1635 852 1.13e-15
c4345 1673 1345 6.7e-16
c4346 632 1774 1.09e-16
c4347 2617 3126 7.84e-16
c4348 1706 1414 5.5e-16
c4349 1328 0 4.1004e-14
c4350 3390 3401 4.097e-15
c4351 1877 1 6.15e-16
c4352 1964 1 5.97e-15
c4353 2172 1783 1.58e-16
c4354 1038 677 1.58e-16
c4355 596 730 2.45e-16
c4356 3858 852 1.58e-16
c4357 5584 1 8.43e-16
c4358 2755 2367 4.97e-16
c4359 5422 0 2.148e-14
c4360 3882 767 3.15e-16
c4361 910 3048 5.03e-16
c4362 2809 2810 1.6e-16
c4363 1076 737 3.15e-16
c4364 1086 1089 1.58e-16
c4365 657 1008 1.58e-16
c4366 1573 812 1.75e-16
c4367 4222 1 6.78e-16
c4368 2004 858 3.69e-16
c4369 1325 0 6.78e-16
c4370 1132 1 3.54e-16
c4371 1129 0 9.602e-15
c4372 4209 0 1.68557e-13
c4373 1764 1765 9.1e-16
c4374 4915 178 1.88e-16
c4375 2035 2023 1.74e-16
c4376 1 246 1.073e-15
c4377 136 305 1.88e-16
c4378 4878 207 1.88e-16
c4379 3785 3732 2.45e-16
c4380 2257 0 3.357e-14
c4381 1419 647 7.38e-16
c4382 1173 1179 1.58e-16
c4383 161 0 1.051e-14
c4384 139 19 8.82e-16
c4385 142 37 1.88e-16
c4386 3452 4288 5.66e-16
c4387 4294 4285 3.92e-16
c4388 4387 737 1.58e-16
c4389 920 980 3.92e-16
c4390 921 979 2.54e-16
c4391 542 541 3.84e-16
c4392 1489 1056 3.92e-16
c4393 1493 1494 1.6e-16
c4394 2880 2933 2.45e-16
c4395 2947 2946 1.6e-16
c4396 959 1 3.06e-16
c4397 2412 767 1.9e-16
c4398 3211 3223 2.32e-16
c4399 3886 792 7.99e-16
c4400 447 455 1.58e-16
c4401 5155 236 9.68e-16
c4402 239 236 4.6e-16
c4403 4076 4070 1.96e-16
c4404 4685 0 4.14862e-13
c4405 2725 2339 5.66e-16
c4406 1151 782 3.57e-16
c4407 4259 4254 1.642e-15
c4408 3882 4353 1.58e-16
c4409 3898 4365 1.58e-16
c4410 910 909 5.33e-16
c4411 3974 26 4.48e-16
c4412 4371 4368 6.44e-16
c4413 4375 4372 3.01e-16
c4414 1474 0 3.3846e-14
c4415 1283 1 3.36e-16
c4416 3531 1 5.97e-15
c4417 687 1777 1.58e-16
c4418 5010 4957 8.95e-16
c4419 2622 0 3.466e-15
c4420 1027 1028 7.46e-16
c4421 12 0 1.5723e-14
c4422 792 2390 5.73e-16
c4423 3886 737 3.15e-16
c4424 4458 797 1.84e-16
c4425 3199 0 8e-16
c4426 1254 1248 1.473e-15
c4427 632 1002 4.98e-16
c4428 2545 0 3.3139e-13
c4429 919 1115 3.92e-16
c4430 922 1114 2.54e-16
c4431 1941 797 5.03e-16
c4432 1343 1436 3.92e-16
c4433 4607 4231 3.92e-16
c4434 4619 4618 1.6e-16
c4435 1684 1318 1.58e-16
c4436 1690 1315 1.58e-16
c4437 3572 0 1.6491e-14
c4438 2559 2535 4.383e-15
c4439 3701 3690 1.58e-16
c4440 1431 1799 1.96e-16
c4441 4883 4503 1.96e-16
c4442 3048 2662 5.5e-16
c4443 2117 2106 1.138e-15
c4444 2022 2135 1.58e-16
c4445 4810 4817 1.81e-16
c4446 1 562 4.59e-16
c4447 19 516 8.82e-16
c4448 37 520 5.71e-16
c4449 306 310 1.58e-16
c4450 3584 3577 6.73e-16
c4451 3583 3191 1.96e-16
c4452 4024 857 3.1e-16
c4453 4582 4622 3.92e-16
c4454 2409 1896 4.97e-16
c4455 79 1 1.607e-15
c4456 3783 3770 8.07e-16
c4457 3370 3842 5.5e-16
c4458 3355 3387 3.92e-16
c4459 5344 0 1.23e-16
c4460 617 3092 1.832e-15
c4461 68 0 2.87e-16
c4462 59 37 1.88e-16
c4463 922 926 3.54e-16
c4464 3005 3001 1.96e-16
c4465 2299 672 2.22e-16
c4466 4134 37 1.88e-16
c4467 3942 1 7.44e-16
c4468 4437 3599 4.97e-16
c4469 3274 2764 1.58e-16
c4470 2679 2668 1.58e-16
c4471 1618 1590 2.64e-16
c4472 509 508 1.079e-15
c4473 30 326 6.83e-16
c4474 4571 4592 1.58e-16
c4475 911 2540 1.58e-16
c4476 2196 1794 5.5e-16
c4477 2222 0 2.93e-15
c4478 3202 717 2.22e-16
c4479 3574 722 1.832e-15
c4480 3446 3441 1.642e-15
c4481 596 702 1.96e-16
c4482 5426 5423 3.92e-16
c4483 2699 2697 1.6e-16
c4484 1726 2243 2.38e-15
c4485 5286 5347 1.6e-16
c4486 2773 777 1.58e-16
c4487 2214 2610 1.96e-16
c4488 2220 2605 1.96e-16
c4489 894 882 1.58e-16
c4490 2990 2988 3.92e-16
c4491 1657 852 2.4e-16
c4492 1327 868 4.03e-16
c4493 1343 827 4.46e-16
c4494 627 3464 2.65e-16
c4495 617 3022 1.58e-16
c4496 612 3083 2.22e-16
c4497 1367 881 1.58e-16
c4498 1131 1138 7.95e-16
c4499 3839 3821 1.58e-16
c4500 4421 4433 2.32e-16
c4501 5585 4582 1.96e-16
c4502 4657 5481 6.5e-16
c4503 3313 822 1.58e-16
c4504 2696 747 1.58e-16
c4505 2545 2203 1.58e-16
c4506 2662 3179 4.11e-16
c4507 595 1727 2.65e-16
c4508 602 1318 2.33e-16
c4509 1708 1854 1.58e-16
c4510 1907 1903 1.96e-16
c4511 3048 707 3.15e-16
c4512 3393 3638 1.96e-16
c4513 5330 5314 7.38e-16
c4514 797 789 1.74e-16
c4515 4567 4401 1.58e-16
c4516 5025 62 6.86e-16
c4517 657 3048 3.58e-16
c4518 2497 1981 4.11e-16
c4519 3948 3956 6.67e-16
c4520 3954 3944 6.67e-16
c4521 2785 2773 2.32e-16
c4522 2276 662 5.03e-16
c4523 1690 767 3.15e-16
c4524 1211 842 3.57e-16
c4525 3533 1 9.28e-16
c4526 3270 822 1.58e-16
c4527 852 1 3.6821e-14
c4528 2957 2952 7.46e-16
c4529 657 1743 1.58e-16
c4530 1208 0 1.4198e-14
c4531 3469 0 3.5926e-14
c4532 1607 1608 1.35e-16
c4533 4412 4384 2.64e-16
c4534 4785 4779 7.25e-16
c4535 4395 4401 9.42e-16
c4536 2685 707 2.33e-16
c4537 2559 858 3.15e-16
c4538 1783 0 3.6368e-14
c4539 1 207 3.36e-15
c4540 3628 3629 5.65e-16
c4541 3236 3623 1.532e-15
c4542 4563 4758 1.96e-16
c4543 4742 4748 5.87e-16
c4544 3409 3066 5.5e-16
c4545 2379 1 2.054e-15
c4546 0 212 2.87e-16
c4547 526 556 1.88e-16
c4548 3645 782 1.58e-16
c4549 5025 5039 5.12e-16
c4550 5138 5133 9.94e-16
c4551 2381 0 8e-16
c4552 2168 1 2.346e-15
c4553 3734 3775 2.45e-16
c4554 3770 3772 1.462e-15
c4555 3918 3917 6.32e-16
c4556 3932 3935 4.41e-16
c4557 1483 702 2.65e-16
c4558 4235 4232 6.44e-16
c4559 4239 4236 3.01e-16
c4560 2288 2669 3.92e-16
c4561 2674 2673 1.6e-16
c4562 1331 1389 1.58e-16
c4563 3886 4467 1.58e-16
c4564 3898 3616 5.5e-16
c4565 3900 3622 1.58e-16
c4566 822 1164 1.58e-16
c4567 3179 707 5.03e-16
c4568 1690 2019 1.58e-16
c4569 599 598 1.6e-16
c4570 3167 3158 3.46e-16
c4571 3151 3536 1.96e-16
c4572 4567 4570 1.58e-16
c4573 350 349 7.03e-16
c4574 792 1694 7.99e-16
c4575 106 117 3.84e-16
c4576 110 100 8.86e-16
c4577 5296 5297 3.18e-16
c4578 909 707 3.15e-16
c4579 883 1066 1.88e-16
c4580 907 1059 1.58e-16
c4581 5177 5160 1.92e-16
c4582 2584 2587 6.44e-16
c4583 3324 1 1.056e-15
c4584 1437 677 2.33e-16
c4585 1343 812 4.46e-16
c4586 657 909 3.15e-16
c4587 4028 4030 2.254e-15
c4588 4107 3918 8.1e-16
c4589 832 1 5.62e-16
c4590 3293 1 4.41e-15
c4591 1417 1 1.056e-15
c4592 612 1343 3.15e-16
c4593 602 1345 3.15e-16
c4594 2742 737 1.58e-16
c4595 181 176 1.059e-15
c4596 175 169 1.58e-16
c4597 3447 3055 1.96e-16
c4598 3448 3441 6.73e-16
c4599 1922 1 5.808e-15
c4600 1924 0 3.466e-15
c4601 3271 767 3.64e-16
c4602 777 1539 1.58e-16
c4603 5584 4950 3.2e-16
c4604 2771 2384 1.532e-15
c4605 2585 2587 2.03e-16
c4606 617 2231 3.15e-16
c4607 2172 1896 5.5e-16
c4608 602 3388 5.18e-16
c4609 4707 692 1.23e-16
c4610 5417 5442 3.54e-16
c4611 3109 0 3.3691e-14
c4612 919 1173 1.58e-16
c4613 602 933 2.322e-15
c4614 1982 827 7.68e-16
c4615 1694 737 3.15e-16
c4616 1701 1335 5.8e-16
c4617 4271 1 2.054e-15
c4618 2720 737 1.339e-15
c4619 1182 0 6.29e-16
c4620 4273 0 8e-16
c4621 3046 3275 3.92e-16
c4622 4850 4463 2.196e-15
c4623 4708 4716 1.81e-16
c4624 4580 4711 1.58e-16
c4625 4571 4723 1.58e-16
c4626 2349 1 8.43e-16
c4627 1468 677 4.81e-16
c4628 5450 5459 1.58e-16
c4629 5452 5451 5.01e-16
c4630 2843 2458 1.96e-16
c4631 2541 2322 1.58e-16
c4632 1522 752 2.33e-16
c4633 1517 1511 1.6e-16
c4634 1061 1508 2.386e-15
c4635 2923 2946 1.96e-16
c4636 3650 4484 1.58e-16
c4637 4686 4299 1.96e-16
c4638 1913 797 1.58e-16
c4639 1793 1784 3.46e-16
c4640 3870 1 5.663e-15
c4641 3048 3092 1.58e-16
c4642 1708 1584 5.5e-16
c4643 1101 1 4.044e-15
c4644 1543 0 6.62e-16
c4645 3515 3509 1.6e-16
c4646 677 667 6.38e-16
c4647 687 2628 1.58e-16
c4648 2383 1862 1.96e-16
c4649 2378 1868 1.96e-16
c4650 5490 5489 1.6e-16
c4651 1766 1777 1.58e-16
c4652 165 158 7.76e-16
c4653 174 172 7.1e-16
c4654 146 194 1.88e-16
c4655 3715 842 1.09e-16
c4656 4322 677 1.84e-16
c4657 5391 5385 6.23e-16
c4658 2673 2282 4.11e-16
c4659 1113 1127 1.96e-16
c4660 3900 3904 1.6e-16
c4661 3882 3895 1.58e-16
c4662 4514 1 5.46e-15
c4663 4657 468 1.88e-16
c4664 5560 5558 1.167e-15
c4665 4389 3548 4.11e-16
c4666 3409 1 4.77e-16
c4667 2322 732 5.73e-16
c4668 3393 777 4.03e-16
c4669 1567 1934 1.58e-16
c4670 5009 5005 9.73e-16
c4671 1886 1 1.716e-15
c4672 418 426 1.58e-16
c4673 3387 3191 1.58e-16
c4674 1042 692 6.38e-16
c4675 4580 4860 3.92e-16
c4676 2552 2544 1.606e-15
c4677 3876 782 4.48e-16
c4678 4489 837 1.58e-16
c4679 5560 5556 8.88e-16
c4680 3073 0 1.6491e-14
c4681 921 1160 1.96e-16
c4682 1982 812 3.64e-16
c4683 4643 4655 2.62e-16
c4684 538 0 1.051e-14
c4685 4367 4368 1.35e-16
c4686 1701 1 7.228e-15
c4687 3046 3240 1.58e-16
c4688 3030 3228 1.58e-16
c4689 637 638 1.96e-16
c4690 4896 33 3.222e-15
c4691 4361 0 6.9337e-14
c4692 1692 0 4.64e-16
c4693 100 0 4.6653e-14
c4694 3594 3591 5.5e-16
c4695 5277 412 3.54e-16
c4696 4742 323 1.88e-16
c4697 2442 1936 3.92e-16
c4698 2446 2447 1.6e-16
c4699 3882 3401 3.15e-16
c4700 5566 5556 1.98e-16
c4701 2277 0 1.4092e-14
c4702 3803 3806 3.54e-16
c4703 3838 3739 9.36e-16
c4704 78 479 1.88e-16
c4705 3010 2486 1.96e-16
c4706 2744 2741 3.01e-16
c4707 2740 2737 6.44e-16
c4708 1114 1115 7.51e-16
c4709 506 508 1.88e-16
c4710 151 149 3.84e-16
c4711 143 129 3.84e-16
c4712 4186 4184 7.1e-16
c4713 3038 3031 7.37e-16
c4714 4459 4458 5.65e-16
c4715 4453 3616 1.532e-15
c4716 2541 2837 1.96e-16
c4717 3309 2798 1.96e-16
c4718 4559 1 3.882e-15
c4719 4735 4728 1.96e-16
c4720 4344 4737 1.914e-15
c4721 3135 662 7.68e-16
c4722 1327 0 3.57642e-13
c4723 22 5 3.84e-16
c4724 5045 5048 3.92e-16
c4725 165 305 1.88e-16
c4726 280 15 6.58e-16
c4727 78 189 1.88e-16
c4728 5379 5366 3.92e-16
c4729 4844 5083 1.96e-16
c4730 4855 236 1.88e-16
c4731 2810 0 1.4092e-14
c4732 910 2545 5.03e-16
c4733 2248 0 6.9484e-14
c4734 632 4270 5.03e-16
c4735 3898 4370 1.58e-16
c4736 3876 4382 1.58e-16
c4737 2559 2637 1.58e-16
c4738 939 0 7.868e-15
c4739 3030 3027 1.123e-15
c4740 1211 1254 6.35e-16
c4741 4723 4724 8.22e-16
c4742 4565 0 4.64e-16
c4743 1920 1931 1.96e-16
c4744 1690 1747 1.58e-16
c4745 1494 0 1.4092e-14
c4746 1270 1 4.17e-16
c4747 5010 4546 7.76e-16
c4748 4567 4299 1.58e-16
c4749 5010 120 1.88e-16
c4750 3034 3046 4.369e-15
c4751 3376 3030 6.89e-16
c4752 224 1 1.607e-15
c4753 2642 0 8e-16
c4754 596 695 5.28e-16
c4755 632 3089 2.33e-16
c4756 3387 858 4.48e-16
c4757 2048 2028 1.69e-16
c4758 966 1389 7.84e-16
c4759 926 927 6.52e-16
c4760 179 1 4.92e-16
c4761 146 15 5.8e-16
c4762 3994 3992 7.1e-16
c4763 3215 0 6.72e-16
c4764 3020 1 2.346e-15
c4765 1236 921 1.17e-16
c4766 1800 702 5.73e-16
c4767 2541 792 4.03e-16
c4768 1321 1453 3.92e-16
c4769 4538 4543 2.029e-15
c4770 3701 4553 4.69e-16
c4771 2491 827 1.58e-16
c4772 573 563 5.32e-16
c4773 4720 1 1.749e-15
c4774 1651 1 8.43e-16
c4775 1 296 5.798e-15
c4776 4827 4835 1.81e-16
c4777 4712 0 7.67e-16
c4778 0 309 1.5723e-14
c4779 4582 4639 3.92e-16
c4780 5410 468 4.44e-16
c4781 5161 5162 5.87e-16
c4782 1896 0 6.9124e-14
c4783 3702 3704 1.6e-16
c4784 2790 2802 2.32e-16
c4785 5324 294 1.58e-16
c4786 3310 827 2.33e-16
c4787 4270 3435 1.96e-16
c4788 4275 3429 1.96e-16
c4789 5407 5409 1.441e-15
c4790 5427 5425 3.92e-16
c4791 2557 2418 5.5e-16
c4792 2629 2237 1.96e-16
c4793 2630 2623 6.73e-16
c4794 149 64 1.88e-16
c4795 2905 2896 3.92e-16
c4796 2406 752 1.58e-16
c4797 882 1 2.97e-15
c4798 4571 677 1.33e-16
c4799 3279 2764 2.386e-15
c4800 2781 3262 1.58e-16
c4801 2679 3203 4.36e-16
c4802 3185 3576 4.11e-16
c4803 901 886 5.71e-16
c4804 3690 1 4.41e-15
c4805 2541 737 3.15e-16
c4806 747 1343 3.15e-16
c4807 37 549 5.71e-16
c4808 4571 4609 1.58e-16
c4809 4582 4621 1.58e-16
c4810 193 195 1.58e-16
c4811 5350 294 3.54e-16
c4812 8 6 1.58e-16
c4813 3397 3688 1.58e-16
c4814 1454 717 5.73e-16
c4815 1321 852 3.15e-16
c4816 1460 1457 5.5e-16
c4817 3726 3727 5.87e-16
c4818 4159 3918 8.1e-16
c4819 617 3466 4.81e-16
c4820 627 3083 3.79e-16
c4821 2668 1 4.41e-15
c4822 2194 2491 3.92e-16
c4823 2879 2877 1.082e-15
c4824 2895 2897 3.92e-16
c4825 4657 64 1.88e-16
c4826 887 0 6.78e-16
c4827 872 19 1.96e-16
c4828 601 1318 1.75e-16
c4829 1690 1488 1.58e-16
c4830 922 1 5.66e-16
c4831 565 580 1.88e-16
c4832 494 487 3.54e-16
c4833 3472 3484 2.32e-16
c4834 3397 3123 1.58e-16
c4835 2336 2334 1.6e-16
c4836 657 2257 1.58e-16
c4837 1590 0 3.5724e-14
c4838 5103 0 3.6193e-14
c4839 1726 2247 1.96e-16
c4840 1732 2242 1.96e-16
c4841 737 732 2.77e-16
c4842 2608 2605 3.01e-16
c4843 2604 2601 6.44e-16
c4844 4567 4418 1.58e-16
c4845 4787 323 1.88e-16
c4846 4056 4054 3.54e-16
c4847 5524 5511 8.94e-16
c4848 5521 5482 1.738e-15
c4849 2921 1 1.021e-15
c4850 4338 4339 1.6e-16
c4851 4334 3503 3.92e-16
c4852 2296 662 1.09e-16
c4853 2020 858 7.38e-16
c4854 1684 782 4.48e-16
c4855 1211 1209 1.931e-15
c4856 3546 1 6.15e-16
c4857 1935 782 7.38e-16
c4858 1544 1540 1.96e-16
c4859 4593 4590 6.67e-16
c4860 2955 2957 5.88e-16
c4861 3034 2832 5.5e-16
c4862 4412 4401 1.58e-16
c4863 2118 2115 3.92e-16
c4864 2072 2120 1.062e-15
c4865 15 320 5.8e-16
c4866 3387 3484 1.58e-16
c4867 4759 4762 6.02e-16
c4868 4563 4775 1.96e-16
c4869 5238 5198 1.062e-15
c4870 5114 62 7.62e-16
c4871 3564 3555 3.46e-16
c4872 4038 4043 1.96e-16
c4873 2216 1 9.28e-16
c4874 520 523 3.54e-16
c4875 0 335 1.051e-14
c4876 1474 707 1.58e-16
c4877 1046 702 3.79e-16
c4878 1224 909 3.08e-16
c4879 5484 5491 1.138e-15
c4880 601 3077 1.9e-16
c4881 2871 2503 1.96e-16
c4882 2015 1987 2.64e-16
c4883 1143 1144 1.21e-16
c4884 2923 2968 1.817e-15
c4885 3720 1 9.28e-16
c4886 3886 4472 1.58e-16
c4887 3876 3633 5.5e-16
c4888 2282 702 1.58e-16
c4889 4395 4781 4.11e-16
c4890 3199 707 1.09e-16
c4891 2108 2100 3.54e-16
c4892 2545 707 3.15e-16
c4893 548 549 6.4e-16
c4894 4742 265 5.88e-16
c4895 5131 5132 1.08e-15
c4896 5106 5105 5.68e-16
c4897 2402 1885 1.96e-16
c4898 2403 2396 6.73e-16
c4899 5297 0 2.156e-15
c4900 5085 1 3.36e-16
c4901 2311 2310 1.6e-16
c4902 2187 0 6.35e-16
c4903 3877 3878 6.67e-16
c4904 4353 702 1.58e-16
c4905 602 3071 1.58e-16
c4906 2767 1 1.056e-15
c4907 657 2545 7.99e-16
c4908 4134 4139 1.96e-16
c4909 4514 4950 9.7e-16
c4910 5308 5299 1.96e-16
c4911 5283 5313 9.6e-16
c4912 3340 1 9.28e-16
c4913 392 223 1.88e-16
c4914 3821 1 2.397e-15
c4915 3839 3847 3.422e-15
c4916 4411 4404 1.96e-16
c4917 3565 4413 4.36e-16
c4918 1862 737 3.15e-16
c4919 627 1343 3.15e-16
c4920 601 1345 3.15e-16
c4921 642 25 1.58e-16
c4922 1887 1889 2.03e-16
c4923 371 378 3.54e-16
c4924 3066 3055 1.58e-16
c4925 2849 858 3.15e-16
c4926 1942 1 2.054e-15
c4927 1944 0 8e-16
c4928 3393 3608 1.58e-16
c4929 3409 3225 1.58e-16
c4930 2538 1 8.766e-15
c4931 5284 5281 3.54e-16
c4932 5440 1 1.88e-16
c4933 3327 3338 1.58e-16
c4934 4108 3918 2.87e-16
c4935 3900 837 3.58e-16
c4936 1545 767 1.84e-16
c4937 1354 877 4.97e-16
c4938 1601 827 3.15e-16
c4939 1321 1101 1.58e-16
c4940 1327 1091 5.88e-16
c4941 612 961 1.35e-16
c4942 4564 4583 1.94e-16
c4943 3084 2566 1.96e-16
c4944 3085 3078 6.73e-16
c4945 1869 1871 1.862e-15
c4946 1482 1488 1.418e-15
c4947 1499 1471 2.64e-16
c4948 4289 0 6.72e-16
c4949 3347 3354 1.96e-16
c4950 3024 3292 3.92e-16
c4951 2082 2083 1.96e-16
c4952 9 451 4.88e-16
c4953 1 429 1.44e-16
c4954 538 542 1.58e-16
c4955 4606 4609 6.02e-16
c4956 4617 4231 1.179e-15
c4957 4580 4728 1.58e-16
c4958 4571 4740 1.58e-16
c4959 4725 4730 5.53e-16
c4960 4725 33 1.88e-16
c4961 1970 2478 7.84e-16
c4962 963 977 1.96e-16
c4963 3781 3862 3.2e-16
c4964 3928 857 3.1e-16
c4965 5112 5111 1.6e-16
c4966 2935 1 3.36e-16
c4967 894 1173 3.54e-16
c4968 1031 1029 1.931e-15
c4969 2557 2339 1.58e-16
c4970 3100 0 6.9481e-14
c4971 3667 4472 1.58e-16
c4972 3650 4489 2.386e-15
c4973 4498 4492 1.6e-16
c4974 2455 797 4.81e-16
c4975 1028 1 4.59e-16
c4976 3349 2832 4.11e-16
c4977 1025 0 1.0077e-14
c4978 3874 1 5.611e-15
c4979 4748 4745 5.5e-16
c4980 3890 3401 3.84e-16
c4981 2143 1 3.36e-16
c4982 602 19 1.676e-15
c4983 0 476 9.795e-15
c4984 3907 3908 7.55e-16
c4985 3915 3917 2.239e-15
c4986 5064 5069 3.54e-16
c4987 2072 0 4.4394e-14
c4988 1133 782 1.58e-16
c4989 3882 3894 6.67e-16
c4990 4208 4218 3.45e-16
c4991 2169 2569 7.84e-16
c4992 1799 662 7.38e-16
c4993 1430 1421 3.46e-16
c4994 657 3469 1.58e-16
c4995 4044 25 1.88e-16
c4996 4040 19 7.35e-16
c4997 3152 3146 1.6e-16
c4998 1567 1939 1.58e-16
c4999 971 1 5.821e-15
c5000 3428 3419 3.46e-16
c5001 3343 827 1.58e-16
c5002 1912 1 8.43e-16
c5003 2501 1 6.15e-16
c5004 4580 4877 3.92e-16
c5005 4119 857 6.23e-16
c5006 964 965 9.71e-16
c5007 4016 4014 1.76e-16
c5008 4509 837 1.58e-16
c5009 2828 2827 5.65e-16
c5010 920 1174 1.58e-16
c5011 1601 812 3.15e-16
c5012 1136 1571 1.58e-16
c5013 779 0 7.709e-15
c5014 397 389 1.58e-16
c5015 910 1327 7.97e-16
c5016 911 1343 9.54e-16
c5017 877 0 4.7451e-14
c5018 4214 4566 5.8e-16
c5019 4223 26 4.58e-16
c5020 827 843 1.621e-15
c5021 4378 0 6.9337e-14
c5022 4787 265 1.88e-16
c5023 822 2424 5.73e-16
c5024 953 931 1.546e-15
c5025 3693 3397 1.58e-16
c5026 3801 3811 8.28e-16
c5027 1190 827 5.74e-16
c5028 920 807 3.15e-16
c5029 129 136 7.76e-16
c5030 910 939 5.59e-16
c5031 2640 2637 5.5e-16
c5032 922 1010 3.92e-16
c5033 3886 3887 1.027e-15
c5034 3055 1 4.41e-15
c5035 642 1001 4.21e-16
c5036 3439 0 6.62e-16
c5037 2557 2854 3.92e-16
c5038 1 256 2.87e-16
c5039 657 3109 1.58e-16
c5040 1423 647 1.832e-15
c5041 407 390 1.138e-15
c5042 408 412 6.38e-16
c5043 276 223 1.88e-16
c5044 3480 662 3.15e-16
c5045 2807 2424 7.84e-16
c5046 2650 2265 1.96e-16
c5047 2640 2647 6.73e-16
c5048 632 4290 1.09e-16
c5049 2541 2836 1.58e-16
c5050 2196 702 3.58e-16
c5051 1301 1293 6.67e-16
c5052 3030 3029 3.15e-16
c5053 762 766 2.19e-16
c5054 4393 1 6.15e-16
c5055 1706 1764 1.58e-16
c5056 1690 1752 1.58e-16
c5057 437 442 1.059e-15
c5058 3515 3117 4.36e-16
c5059 262 570 1.88e-16
c5060 4928 4919 3.92e-16
c5061 4902 4933 6.67e-16
c5062 2260 2267 6.73e-16
c5063 426 1 2.6688e-14
c5064 229 233 1.58e-16
c5065 416 0 2.87e-16
c5066 1 118 1.456e-15
c5067 407 37 1.88e-16
c5068 3397 3157 1.58e-16
c5069 4804 33 1.88e-16
c5070 1380 647 1.58e-16
c5071 3639 812 1.75e-16
c5072 5552 5540 6.67e-16
c5073 5530 5532 5.48e-16
c5074 1268 1273 3.54e-16
c5075 3537 4370 7.84e-16
c5076 2334 702 2.65e-16
c5077 1708 837 3.58e-16
c5078 3591 1 5.808e-15
c5079 2545 2441 1.58e-16
c5080 1952 807 2.4e-16
c5081 1557 1568 1.96e-16
c5082 1345 1470 3.92e-16
c5083 734 0 7.709e-15
c5084 4624 4248 3.92e-16
c5085 4636 4635 1.6e-16
c5086 1708 1319 5.5e-16
c5087 617 1402 1.58e-16
c5088 3719 1 1.868e-15
c5089 2178 837 4.03e-16
c5090 4889 4884 1.977e-15
c5091 4737 1 1.749e-15
c5092 4896 526 1.395e-15
c5093 1635 2162 4.69e-16
c5094 2149 2154 2.029e-15
c5095 747 1871 1.58e-16
c5096 1818 0 1.6491e-14
c5097 1669 1 1.106e-15
c5098 3409 3518 1.58e-16
c5099 4571 4463 5.5e-16
c5100 4844 4849 5.53e-16
c5101 4729 0 7.67e-16
c5102 27 19 3.84e-16
c5103 3397 717 7.99e-16
c5104 4582 4656 3.92e-16
c5105 1345 886 3.54e-16
c5106 1251 1248 1.96e-16
c5107 3039 0 6.35e-16
c5108 1190 812 1.58e-16
c5109 1001 997 3.78e-16
c5110 2535 2435 5.5e-16
c5111 2717 2333 1.58e-16
c5112 1321 1452 1.58e-16
c5113 1343 1440 1.58e-16
c5114 3839 3759 1.58e-16
c5115 3882 4535 1.58e-16
c5116 2182 837 7.99e-16
c5117 1431 1803 1.58e-16
c5118 3034 777 7.99e-16
c5119 1735 1733 1.862e-15
c5120 1083 0 4.6723e-14
c5121 927 1 1.503e-15
c5122 2104 1667 2.037e-15
c5123 4553 1 1.601e-15
c5124 2535 752 4.48e-16
c5125 2015 842 1.58e-16
c5126 2268 1 1.056e-15
c5127 291 305 1.88e-16
c5128 4571 4626 1.58e-16
c5129 4582 4638 1.58e-16
c5130 2413 2410 5.5e-16
c5131 0 569 1.5723e-14
c5132 5367 0 2.078e-15
c5133 2342 1834 7.84e-16
c5134 48 50 1.58e-16
c5135 42 37 1.88e-16
c5136 3862 3853 7.53e-16
c5137 4872 5144 5.5e-16
c5138 632 3090 1.339e-15
c5139 2237 1 4.41e-15
c5140 4173 4172 7.81e-16
c5141 5326 5323 7.46e-16
c5142 2788 2407 3.92e-16
c5143 2231 2622 4.11e-16
c5144 1863 717 2.65e-16
c5145 2172 2508 3.92e-16
c5146 3203 1 1.868e-15
c5147 4441 4438 5.5e-16
c5148 2880 2884 1.96e-16
c5149 732 25 1.58e-16
c5150 3277 2764 1.532e-15
c5151 2545 2231 5.5e-16
c5152 3937 37 1.88e-16
c5153 3951 0 2.069e-14
c5154 3192 3201 3.46e-16
c5155 612 1744 2.65e-16
c5156 1457 1 5.808e-15
c5157 1706 1505 1.58e-16
c5158 601 4605 1.23e-16
c5159 1459 0 3.466e-15
c5160 657 2277 1.58e-16
c5161 5144 0 1.5838e-14
c5162 5137 31 3.54e-16
c5163 909 901 3.54e-16
c5164 3253 3259 1.418e-15
c5165 4567 4435 1.58e-16
c5166 5478 410 3.54e-16
c5167 5511 1 1.81e-16
c5168 3270 3242 2.64e-16
c5169 2520 2510 7.53e-16
c5170 2514 1998 3.92e-16
c5171 1008 1009 1.21e-16
c5172 687 3048 3.58e-16
c5173 1327 707 3.15e-16
c5174 1370 881 1.532e-15
c5175 1376 1375 5.65e-16
c5176 3967 3958 1.96e-16
c5177 2541 2599 1.96e-16
c5178 2319 677 4.81e-16
c5179 657 1327 4.03e-16
c5180 3555 1 1.716e-15
c5181 1234 1 1.842e-15
c5182 4525 4521 1.96e-16
c5183 2892 2893 3.18e-16
c5184 2288 677 2.33e-16
c5185 2798 782 1.58e-16
c5186 2245 2242 3.01e-16
c5187 2241 2238 6.44e-16
c5188 4429 4401 2.64e-16
c5189 4802 4796 7.25e-16
c5190 4412 4418 9.42e-16
c5191 3387 3489 1.58e-16
c5192 3411 3501 5.42e-16
c5193 3393 3106 1.58e-16
c5194 4563 4792 1.96e-16
c5195 5165 5190 3.54e-16
c5196 657 2248 1.813e-15
c5197 1885 1 4.41e-15
c5198 647 998 1.58e-16
c5199 2394 0 6.62e-16
c5200 3651 797 7.68e-16
c5201 3944 3951 1.88e-16
c5202 5406 468 3.54e-16
c5203 4878 497 1.88e-16
c5204 1494 707 1.58e-16
c5205 3882 717 4.03e-16
c5206 617 3077 5.03e-16
c5207 2691 2692 5.65e-16
c5208 922 1068 1.58e-16
c5209 4247 3385 1.96e-16
c5210 3350 1 2.054e-15
c5211 3900 3650 5.5e-16
c5212 1964 837 1.813e-15
c5213 2849 3377 4.69e-16
c5214 3362 3367 2.029e-15
c5215 3815 410 9.36e-16
c5216 3262 3261 2.48e-16
c5217 1591 0 1.6491e-14
c5218 1989 1607 2.48e-16
c5219 887 884 5.6e-16
c5220 319 317 7.1e-16
c5221 136 450 1.88e-16
c5222 5104 5106 1.96e-16
c5223 3559 722 5.03e-16
c5224 2186 0 8.0614e-14
c5225 601 3071 7.38e-16
c5226 2870 2503 1.58e-16
c5227 1156 1157 1.238e-15
c5228 1147 807 1.58e-16
c5229 883 1053 3.54e-16
c5230 894 1074 1.58e-16
c5231 966 968 7.72e-16
c5232 3384 4234 7.84e-16
c5233 3353 1 6.15e-16
c5234 1465 677 1.58e-16
c5235 1647 868 1.58e-16
c5236 1450 1449 1.6e-16
c5237 1442 1440 2.15e-16
c5238 687 909 3.15e-16
c5239 411 408 6.67e-16
c5240 107 108 6.96e-16
c5241 3908 1 7.71e-16
c5242 4104 37 5.71e-16
c5243 3882 4298 1.96e-16
c5244 3900 3480 5.5e-16
c5245 1722 1720 1.6e-16
c5246 1717 1716 2.03e-16
c5247 4783 4781 1.6e-16
c5248 1421 1 1.716e-15
c5249 617 1345 3.15e-16
c5250 5114 5113 1.559e-15
c5251 352 355 4.6e-16
c5252 3066 3464 4.36e-16
c5253 3462 3455 1.96e-16
c5254 2307 1794 4.97e-16
c5255 2540 1 6.056e-15
c5256 1682 2219 1.96e-16
c5257 792 1550 1.813e-15
c5258 2555 0 1.2366e-14
c5259 4127 3918 8.1e-16
c5260 5577 5584 2.15e-16
c5261 2867 2861 1.6e-16
c5262 1331 677 3.15e-16
c5263 2559 2558 1.866e-15
c5264 602 923 1.58e-16
c5265 644 0 7.709e-15
c5266 2577 2566 1.58e-16
c5267 1173 1 1.56e-15
c5268 2741 752 5.03e-16
c5269 1667 1674 3.96e-16
c5270 3048 3309 3.92e-16
c5271 5202 5197 3.07e-16
c5272 3397 3450 1.58e-16
c5273 1981 2461 1.58e-16
c5274 3942 857 1.88e-16
c5275 1222 858 1.58e-16
c5276 1203 1216 1.58e-16
c5277 3898 677 4.46e-16
c5278 5450 5503 3.18e-16
c5279 2947 0 1.65e-16
c5280 1321 971 5.5e-16
c5281 1343 957 5.5e-16
c5282 4093 1 6.78e-16
c5283 3024 2600 1.58e-16
c5284 3030 2594 5.88e-16
c5285 1352 0 3.5936e-14
c5286 1570 1 1.056e-15
c5287 4242 1 6.275e-15
c5288 233 484 1.88e-16
c5289 601 19 1.676e-15
c5290 2345 0 1.4092e-14
c5291 2162 1 1.601e-15
c5292 5491 5489 3.92e-16
c5293 2152 0 6.78e-16
c5294 160 107 1.88e-16
c5295 2969 2970 3.92e-16
c5296 910 877 1.58e-16
c5297 1335 1344 1.846e-15
c5298 3847 1 1.672e-15
c5299 4054 37 1.88e-16
c5300 4063 25 4.68e-16
c5301 4400 4399 9.1e-16
c5302 792 799 1.6e-16
c5303 4438 1 5.808e-15
c5304 2812 797 1.09e-16
c5305 1708 1799 3.92e-16
c5306 3605 777 1.58e-16
c5307 4440 0 3.466e-15
c5308 4905 4919 2.208e-15
c5309 4977 4980 7.84e-16
c5310 3030 807 4.03e-16
c5311 3411 3202 5.5e-16
c5312 2866 3024 3.92e-16
c5313 852 857 1.58e-16
c5314 4787 4782 1.536e-15
c5315 4580 4894 3.92e-16
c5316 4861 1 4.1966e-14
c5317 2572 2571 1.6e-16
c5318 4567 0 3.27017e-13
c5319 4651 497 1.88e-16
c5320 4498 827 7.68e-16
c5321 1101 1102 8.58e-16
c5322 3886 4234 1.58e-16
c5323 3876 3381 3.54e-16
c5324 1136 1576 1.58e-16
c5325 4660 4672 2.62e-16
c5326 3146 3147 5.65e-16
c5327 3065 3056 3.46e-16
c5328 1853 1471 2.48e-16
c5329 4546 3744 4.72e-16
c5330 3342 3343 9.1e-16
c5331 3048 3245 1.58e-16
c5332 1888 0 3.372e-14
c5333 1 471 5.62e-16
c5334 421 117 1.88e-16
c5335 3409 3587 3.92e-16
c5336 4395 0 6.9337e-14
c5337 1 497 3.36e-15
c5338 245 248 2.142e-15
c5339 136 137 6.96e-16
c5340 448 37 1.88e-16
c5341 5136 5093 3.1e-16
c5342 4855 178 1.88e-16
c5343 4725 526 1.88e-16
c5344 2459 1947 1.532e-15
c5345 2465 2464 5.65e-16
c5346 2194 2218 1.58e-16
c5347 2178 2206 1.58e-16
c5348 108 1 1.607e-15
c5349 4413 752 7.68e-16
c5350 1690 717 4.03e-16
c5351 919 1024 1.58e-16
c5352 3627 0 3.466e-15
c5353 4205 4213 6.67e-16
c5354 4211 4201 7.1e-16
c5355 3464 1 1.868e-15
c5356 3454 0 2.93e-15
c5357 4471 4472 2.48e-16
c5358 2535 2871 3.92e-16
c5359 4033 0 6.113e-14
c5360 4766 0 6.72e-16
c5361 236 267 1.88e-16
c5362 0 181 1.4515e-14
c5363 747 2350 1.813e-15
c5364 2182 2206 1.58e-16
c5365 3739 3837 3.87e-16
c5366 3811 3826 6.67e-16
c5367 890 807 3.35e-16
c5368 146 247 1.88e-16
c5369 4188 4190 2.254e-15
c5370 3882 3554 1.58e-16
c5371 4600 5429 1.96e-16
c5372 2557 2853 1.58e-16
c5373 2541 2841 1.58e-16
c5374 3248 762 1.58e-16
c5375 969 0 2.7176e-14
c5376 3897 1 2.94e-16
c5377 4006 25 3.84e-16
c5378 1206 1661 1.361e-15
c5379 1196 1331 5.5e-16
c5380 4740 4741 8.22e-16
c5381 1946 1550 1.96e-16
c5382 1941 1556 1.96e-16
c5383 1684 1781 1.58e-16
c5384 1706 1769 1.58e-16
c5385 1071 0 3.7577e-14
c5386 1344 1 2.471e-15
c5387 5048 5047 1.334e-15
c5388 662 653 1.078e-15
c5389 602 2209 1.58e-16
c5390 3508 662 1.9e-16
c5391 3515 677 7.68e-16
c5392 3046 767 4.46e-16
c5393 293 1 4.92e-16
c5394 5393 5383 1.98e-16
c5395 4844 5095 3.92e-16
c5396 4827 5034 5.87e-16
c5397 642 640 3.327e-15
c5398 287 37 1.88e-16
c5399 5569 1 9.22e-16
c5400 2866 3359 1.58e-16
c5401 2655 0 6.62e-16
c5402 1055 677 1.58e-16
c5403 657 3100 1.813e-15
c5404 1397 672 1.58e-16
c5405 1797 647 4.81e-16
c5406 1415 1409 1.6e-16
c5407 3056 1 1.716e-15
c5408 1270 1269 6.84e-16
c5409 4498 812 3.64e-16
c5410 4821 149 1.88e-16
c5411 2811 2809 1.6e-16
c5412 2806 2805 2.03e-16
c5413 3548 4353 1.58e-16
c5414 1828 702 3.79e-16
c5415 3124 3123 1.35e-16
c5416 3236 747 2.22e-16
c5417 3219 762 1.813e-15
c5418 5417 528 1.76e-16
c5419 4213 1 6.78e-16
c5420 2305 717 5.73e-16
c5421 777 596 1.96e-16
c5422 3228 737 1.832e-15
c5423 747 1891 1.58e-16
c5424 3409 3523 1.58e-16
c5425 602 2166 1.58e-16
c5426 612 2169 5.73e-16
c5427 2260 1 2.054e-15
c5428 902 898 9.02e-16
c5429 937 936 6.67e-16
c5430 9 248 4.88e-16
c5431 3293 837 5.73e-16
c5432 3734 3732 1.96e-16
c5433 3996 3998 2.254e-15
c5434 4582 4673 3.92e-16
c5435 5062 91 3.54e-16
c5436 2178 1851 1.58e-16
c5437 1511 732 1.58e-16
c5438 160 1 1.5821e-14
c5439 143 26 1.03e-15
c5440 140 19 3.2e-16
c5441 3038 0 8.1163e-14
c5442 3480 3486 1.418e-15
c5443 2559 2452 5.5e-16
c5444 2725 2731 1.6e-16
c5445 2722 2333 2.386e-15
c5446 1016 1019 6.13e-16
c5447 4287 3446 4.11e-16
c5448 1706 677 4.46e-16
c5449 1345 1469 5.42e-16
c5450 1321 1457 1.58e-16
c5451 1495 1493 1.6e-16
c5452 1490 1489 2.03e-16
c5453 542 552 3.75e-16
c5454 4552 3900 6.7e-16
c5455 2697 692 3.64e-16
c5456 2922 2918 3.54e-16
c5457 3221 3220 1.6e-16
c5458 1647 0 1.4092e-14
c5459 4531 3690 1.136e-15
c5460 2871 858 7.38e-16
c5461 2005 1624 3.92e-16
c5462 2009 2010 1.6e-16
c5463 37 274 1.88e-16
c5464 4571 4643 1.58e-16
c5465 4582 4655 1.58e-16
c5466 5488 470 8.44e-16
c5467 5178 5157 1.6e-16
c5468 2182 1851 1.58e-16
c5469 447 446 6.67e-16
c5470 335 332 2.142e-15
c5471 3600 737 3.64e-16
c5472 2354 1845 1.58e-16
c5473 1186 837 1.35e-16
c5474 907 767 4.8e-16
c5475 883 1127 3.92e-16
c5476 890 1126 1.88e-16
c5477 223 221 1.257e-15
c5478 4668 1 1.8371e-14
c5479 2620 2265 1.58e-16
c5480 1482 717 3.79e-16
c5481 2696 1 5.97e-15
c5482 3886 3514 5.5e-16
c5483 2396 767 1.84e-16
c5484 3918 25 9.168e-15
c5485 2311 692 1.84e-16
c5486 3206 3207 9.1e-16
c5487 601 1746 4.81e-16
c5488 612 1363 3.79e-16
c5489 1477 1 2.054e-15
c5490 3718 4536 1.96e-16
c5491 1684 1522 1.58e-16
c5492 1690 1516 5.88e-16
c5493 822 1593 1.58e-16
c5494 2177 1698 9.72e-16
c5495 1479 0 8e-16
c5496 3492 3489 5.5e-16
c5497 3593 737 1.9e-16
c5498 4915 4919 2.95e-16
c5499 3276 3277 1.35e-16
c5500 2340 1834 3.92e-16
c5501 2344 2345 1.6e-16
c5502 5108 122 1.345e-15
c5503 3299 812 1.84e-16
c5504 8 0 1.051e-14
c5505 3397 842 3.15e-16
c5506 4567 4452 1.58e-16
c5507 4804 526 1.88e-16
c5508 2172 2507 1.58e-16
c5509 2194 2495 1.58e-16
c5510 3013 1 1.052e-15
c5511 4357 4356 5.65e-16
c5512 4351 3514 1.532e-15
c5513 2557 2616 3.92e-16
c5514 1327 1605 1.58e-16
c5515 703 1 1.65e-16
c5516 3581 1 8.43e-16
c5517 4610 4607 6.67e-16
c5518 4156 1 4.64e-16
c5519 1813 1 9.28e-16
c5520 4486 1 4.442e-15
c5521 4429 4418 1.58e-16
c5522 4863 0 2.93e-15
c5523 1 513 3.4063e-14
c5524 3409 837 3.15e-16
c5525 4563 4809 1.96e-16
c5526 5239 5198 1.817e-15
c5527 2196 1981 5.5e-16
c5528 1021 1022 1.238e-15
c5529 1020 647 6.48e-16
c5530 1012 672 1.58e-16
c5531 807 813 1.097e-15
c5532 3270 797 3.15e-16
c5533 2994 1 3.36e-16
c5534 1261 1245 1.79e-16
c5535 1246 1242 2.092e-15
c5536 642 991 1.35e-16
c5537 56 58 7.1e-16
c5538 617 3097 1.09e-16
c5539 2923 0 4.4655e-14
c5540 1939 782 1.832e-15
c5541 1331 996 1.58e-16
c5542 3873 4592 7.84e-16
c5543 3759 1 7.51e-16
c5544 2469 842 3.15e-16
c5545 2676 677 1.09e-16
c5546 2459 827 1.339e-15
c5547 1074 1 2.972e-15
c5548 4873 4486 1.96e-16
c5549 1075 0 6.29e-16
c5550 4412 4798 4.11e-16
c5551 4794 4803 3.46e-16
c5552 910 2555 1.58e-16
c5553 30 323 3.84e-16
c5554 3393 647 3.15e-16
c5555 2328 2329 5.65e-16
c5556 2771 1 1.716e-15
c5557 687 2545 7.99e-16
c5558 1164 797 8.3e-16
c5559 3385 4246 1.58e-16
c5560 5343 5321 6.67e-16
c5561 78 79 6.96e-16
c5562 2982 2986 9.07e-16
c5563 4514 5577 1.91e-15
c5564 1367 957 1.58e-16
c5565 3724 468 8.6e-16
c5566 612 3384 5.73e-16
c5567 602 3381 1.58e-16
c5568 4423 4421 2.15e-16
c5569 4431 4430 1.6e-16
c5570 3266 3264 1.6e-16
c5571 3261 3260 2.03e-16
c5572 1626 1176 2.48e-16
c5573 2843 837 2.72e-16
c5574 3656 0 3.5724e-14
c5575 1573 1 4.41e-15
c5576 165 450 1.88e-16
c5577 1957 0 6.62e-16
c5578 3387 3637 1.58e-16
c5579 2884 352 1.098e-15
c5580 392 233 1.88e-16
c5581 3710 3355 1.58e-16
c5582 4047 4039 9.33e-16
c5583 3886 827 3.15e-16
c5584 3882 842 3.15e-16
c5585 4536 858 7.38e-16
c5586 1116 767 2.33e-16
c5587 4416 4417 9.1e-16
c5588 2557 2581 1.58e-16
c5589 2541 2569 1.58e-16
c5590 2010 842 1.58e-16
c5591 1345 1106 5.5e-16
c5592 612 963 1.58e-16
c5593 601 923 1.58e-16
c5594 2577 3101 4.36e-16
c5595 3099 3092 1.96e-16
c5596 1207 1 3.54e-16
c5597 366 361 1.482e-15
c5598 4311 1 1.868e-15
c5599 2761 752 1.09e-16
c5600 1899 1897 1.6e-16
c5601 4301 0 2.93e-15
c5602 5001 4946 3.18e-16
c5603 4990 4989 1.6e-16
c5604 1204 0 9.602e-15
c5605 5234 178 3.54e-16
c5606 1930 1539 1.136e-15
c5607 88 252 1.88e-16
c5608 3397 3455 1.58e-16
c5609 466 469 6.67e-16
c5610 461 465 1.58e-16
c5611 448 453 1.482e-15
c5612 1 209 5.798e-15
c5613 4742 4750 1.81e-16
c5614 4582 4745 1.58e-16
c5615 5207 5195 8.45e-16
c5616 5160 5158 1.96e-16
c5617 3765 3770 3.54e-16
c5618 5469 0 1.23e-16
c5619 5484 381 1.58e-16
c5620 2780 2771 3.46e-16
c5621 4103 1 6.03e-16
c5622 1049 1 3.06e-16
c5623 2747 3241 1.96e-16
c5624 1586 1 9.28e-16
c5625 538 544 1.372e-15
c5626 4259 1 6.275e-15
c5627 4765 4762 5.5e-16
c5628 617 19 1.676e-15
c5629 0 444 2.87e-16
c5630 19 433 8.4e-16
c5631 3638 767 1.58e-16
c5632 4563 4214 3.15e-16
c5633 2367 0 6.9484e-14
c5634 921 702 3.15e-16
c5635 99 100 1.482e-15
c5636 3497 692 1.58e-16
c5637 3507 0 6.62e-16
c5638 1636 842 7.68e-16
c5639 1629 827 1.9e-16
c5640 1011 1001 1.418e-15
c5641 3296 0 3.3633e-14
c5642 834 1 5.57e-16
c5643 677 26 7.12e-16
c5644 687 1783 5.73e-16
c5645 2557 662 4.46e-16
c5646 1965 1573 1.96e-16
c5647 1966 1959 6.73e-16
c5648 3523 3522 2.48e-16
c5649 5081 5079 3.92e-16
c5650 3616 762 2.22e-16
c5651 3440 3436 1.96e-16
c5652 617 2253 1.58e-16
c5653 2106 0 4.014e-14
c5654 175 171 1.58e-16
c5655 158 168 8.86e-16
c5656 3157 702 1.58e-16
c5657 102 49 1.88e-16
c5658 2765 2373 1.96e-16
c5659 3747 3757 1.96e-16
c5660 1803 662 1.832e-15
c5661 3588 3589 1.35e-16
c5662 3112 1 2.054e-15
c5663 3886 812 3.15e-16
c5664 3667 827 3.15e-16
c5665 2840 2841 2.48e-16
c5666 3900 3385 5.5e-16
c5667 3114 0 8e-16
c5668 1257 1248 1.97e-16
c5669 919 1190 3.92e-16
c5670 922 1189 2.54e-16
c5671 3253 0 6.9178e-14
c5672 612 3886 7.99e-16
c5673 2735 722 1.58e-16
c5674 253 252 6.96e-16
c5675 1760 2283 4.36e-16
c5676 4469 4846 2.48e-16
c5677 3030 2753 1.58e-16
c5678 3140 3141 1.35e-16
c5679 2179 2181 3.67e-16
c5680 1908 0 1.4092e-14
c5681 4412 0 6.8929e-14
c5682 4589 4596 1.81e-16
c5683 4674 5522 5.5e-16
c5684 4708 5388 1.596e-15
c5685 2172 2235 1.58e-16
c5686 2194 2223 1.58e-16
c5687 3582 752 3.15e-16
c5688 5450 5442 3.54e-16
c5689 922 837 3.15e-16
c5690 4309 4302 1.96e-16
c5691 3463 4311 4.36e-16
c5692 3083 1 5.97e-15
c5693 657 1419 2.4e-16
c5694 1345 1328 3.62e-16
c5695 1343 1335 4.63e-16
c5696 1785 1787 2.03e-16
c5697 3151 3123 2.64e-16
c5698 3237 3228 3.92e-16
c5699 2719 3231 5.66e-16
c5700 2730 3223 1.58e-16
c5701 1722 0 6.72e-16
c5702 4783 0 6.72e-16
c5703 3163 677 1.58e-16
c5704 2044 2049 7.46e-16
c5705 1690 1969 1.96e-16
c5706 3304 827 3.15e-16
c5707 4585 0 1.23e-16
c5708 5158 5162 1.96e-16
c5709 0 362 1.5696e-14
c5710 5423 0 2.156e-15
c5711 2310 0 3.466e-15
c5712 2196 1682 5.5e-16
c5713 677 669 1.74e-16
c5714 3819 3773 1.062e-15
c5715 3818 3820 3.92e-16
c5716 3823 3822 1.6e-16
c5717 5207 0 1.5617e-14
c5718 3900 3899 1.866e-15
c5719 4315 662 7.38e-16
c5720 2722 747 1.58e-16
c5721 3667 3276 1.136e-15
c5722 2535 2870 1.58e-16
c5723 2557 2858 1.58e-16
c5724 1166 1162 3.78e-16
c5725 1380 1386 1.418e-15
c5726 2559 2288 1.58e-16
c5727 2545 2683 1.58e-16
c5728 3701 3310 1.136e-15
c5729 3228 3230 2.15e-16
c5730 3048 3071 3.92e-16
c5731 30 265 3.84e-16
c5732 3219 2702 1.136e-15
c5733 612 2223 1.58e-16
c5734 601 2209 1.84e-16
c5735 3048 782 3.15e-16
c5736 276 233 1.88e-16
c5737 3397 3185 5.5e-16
c5738 4563 4469 1.58e-16
c5739 4872 120 1.88e-16
c5740 4022 3918 2.48e-16
c5741 3082 1 8.43e-16
c5742 1281 1299 9.23e-16
c5743 3667 812 3.15e-16
c5744 3243 777 1.58e-16
c5745 2345 707 1.58e-16
c5746 1690 842 3.15e-16
c5747 1694 827 3.15e-16
c5748 1667 858 1.58e-16
c5749 1343 1657 3.92e-16
c5750 3392 3027 7.67e-16
c5751 3235 3226 3.46e-16
c5752 1583 1121 1.96e-16
c5753 1578 1131 1.96e-16
c5754 1320 1 2.259e-15
c5755 4641 4265 3.92e-16
c5756 4653 4652 1.6e-16
c5757 792 592 5.8e-16
c5758 4546 0 5.5523e-14
c5759 4756 1 1.013e-15
c5760 4984 526 9.02e-16
c5761 3034 2713 5.5e-16
c5762 277 274 2.142e-15
c5763 3676 3674 1.862e-15
c5764 3304 3276 2.64e-16
c5765 3589 3600 1.96e-16
c5766 601 2166 1.58e-16
c5767 120 0 1.21326e-13
c5768 4582 4690 3.92e-16
c5769 2448 2446 1.6e-16
c5770 2443 2442 2.03e-16
c5771 1275 1226 1.154e-15
c5772 1290 1289 1.6e-16
c5773 4742 381 1.88e-16
c5774 617 2611 1.58e-16
c5775 3615 1 8.43e-16
c5776 1956 807 1.58e-16
c5777 1345 1474 1.58e-16
c5778 1386 1387 1.35e-16
c5779 2316 692 3.15e-16
c5780 1829 1437 1.96e-16
c5781 1830 1823 6.73e-16
c5782 542 59 1.88e-16
c5783 4193 0 1.46378e-13
c5784 4019 1 6.78e-16
c5785 4184 26 1.075e-15
c5786 1343 1 4.77e-16
c5787 777 767 3.28e-16
c5788 4463 4813 2e-16
c5789 3226 752 1.339e-15
c5790 2161 1708 6.7e-16
c5791 1664 0 1.3715e-14
c5792 3589 3593 1.96e-16
c5793 642 2194 3.15e-16
c5794 19 21 3.45e-16
c5795 37 22 5.71e-16
c5796 3304 812 3.15e-16
c5797 4571 4660 1.58e-16
c5798 4582 4672 1.58e-16
c5799 2435 2430 1.642e-15
c5800 3219 722 1.58e-16
c5801 3830 3809 1.96e-16
c5802 632 3111 1.9e-16
c5803 2720 2333 1.532e-15
c5804 909 782 3.15e-16
c5805 883 1141 1.88e-16
c5806 907 1134 1.58e-16
c5807 2811 0 6.72e-16
c5808 2648 1 1.056e-15
c5809 5360 5355 5.63e-16
c5810 5324 5378 9.34e-16
c5811 3389 0 5.96e-16
c5812 2920 2915 7.25e-16
c5813 941 1 4.03e-16
c5814 3783 1 1.3e-16
c5815 4166 25 3.84e-16
c5816 4001 0 4.3997e-14
c5817 3992 26 1.075e-15
c5818 1642 1191 3.92e-16
c5819 1646 1647 1.6e-16
c5820 3718 3876 3.92e-16
c5821 2645 677 3.15e-16
c5822 627 1363 1.813e-15
c5823 822 1613 1.58e-16
c5824 1495 0 6.72e-16
c5825 617 4622 1.23e-16
c5826 1918 1533 1.96e-16
c5827 747 1076 1.813e-15
c5828 19 580 3.84e-16
c5829 5174 1 2.386e-15
c5830 5010 5009 3.54e-16
c5831 5160 207 1.58e-16
c5832 752 1112 1.58e-16
c5833 894 961 5.9e-16
c5834 907 931 1.58e-16
c5835 216 9 5.8e-16
c5836 3446 647 1.58e-16
c5837 5366 5363 3.92e-16
c5838 5326 5368 1.017e-15
c5839 223 27 1.88e-16
c5840 3670 3668 1.6e-16
c5841 2136 2046 1.58e-16
c5842 1131 807 5.73e-16
c5843 1388 1389 2.48e-16
c5844 59 281 1.88e-16
c5845 3960 37 5.71e-16
c5846 2535 2633 3.92e-16
c5847 1694 812 3.15e-16
c5848 1343 1622 1.58e-16
c5849 1327 1610 1.58e-16
c5850 367 15 6.58e-16
c5851 687 1327 4.03e-16
c5852 1752 1369 7.84e-16
c5853 2784 767 4.81e-16
c5854 562 563 1.482e-15
c5855 4387 747 1.58e-16
c5856 4503 1 3.97e-15
c5857 2253 1743 1.96e-16
c5858 612 1694 7.99e-16
c5859 4143 3404 2.697e-15
c5860 4446 4418 2.64e-16
c5861 4429 4435 9.42e-16
c5862 4880 0 2.972e-15
c5863 1 314 2.87e-16
c5864 13 305 1.88e-16
c5865 4563 4826 1.96e-16
c5866 2421 1 1.056e-15
c5867 3016 1 8e-16
c5868 1500 722 7.68e-16
c5869 4702 5338 1.96e-16
c5870 2800 2799 1.6e-16
c5871 2792 2790 2.15e-16
c5872 2705 2704 2.48e-16
c5873 676 25 7.64e-16
c5874 3557 0 3.3874e-14
c5875 2476 868 1.58e-16
c5876 627 1370 1.58e-16
c5877 3030 3172 1.58e-16
c5878 3655 807 2.4e-16
c5879 911 2169 1.88e-16
c5880 3959 3960 6.4e-16
c5881 3710 858 1.58e-16
c5882 3429 4234 1.58e-16
c5883 3385 4251 2.386e-15
c5884 4260 4254 1.6e-16
c5885 3372 1 1.106e-15
c5886 1206 852 4e-16
c5887 1455 1466 1.96e-16
c5888 3772 1 1.23e-16
c5889 601 3381 1.58e-16
c5890 612 4260 2.65e-16
c5891 3900 4315 3.92e-16
c5892 2764 3258 1.96e-16
c5893 1533 1528 1.642e-15
c5894 4800 4798 1.6e-16
c5895 1990 2002 2.32e-16
c5896 475 476 6.67e-16
c5897 274 317 1.88e-16
c5898 465 484 1.88e-16
c5899 3474 3472 2.15e-16
c5900 3482 3481 1.6e-16
c5901 3886 747 7.99e-16
c5902 1982 1 1.868e-15
c5903 478 476 2.84e-16
c5904 482 477 1.482e-15
c5905 495 494 7.03e-16
c5906 1972 0 2.93e-15
c5907 3387 3642 1.58e-16
c5908 3411 3654 5.42e-16
c5909 3393 3259 1.58e-16
c5910 1087 722 1.58e-16
c5911 1068 1074 1.58e-16
c5912 391 407 3.84e-16
c5913 99 98 6.67e-16
c5914 378 421 1.88e-16
c5915 4055 4056 6.4e-16
c5916 3876 858 4.48e-16
c5917 4787 381 1.88e-16
c5918 2874 2876 8.88e-16
c5919 2898 2897 1.6e-16
c5920 1106 782 1.58e-16
c5921 3882 4302 1.58e-16
c5922 3898 4314 1.58e-16
c5923 1240 921 2.48e-16
c5924 922 1238 4.42e-16
c5925 3915 25 1.88e-16
c5926 3911 19 7.35e-16
c5927 4335 4334 2.03e-16
c5928 4340 4338 1.6e-16
c5929 5509 5403 6.31e-16
c5930 2005 852 1.58e-16
c5931 1431 1420 1.58e-16
c5932 627 963 1.05e-15
c5933 822 828 1.097e-15
c5934 1423 0 3.3581e-14
c5935 3467 3468 9.1e-16
c5936 2571 0 3.466e-15
c5937 4039 4038 1.58e-16
c5938 4759 4764 5.53e-16
c5939 4582 4762 1.58e-16
c5940 5100 62 3.54e-16
c5941 762 2373 1.58e-16
c5942 387 0 2.87e-16
c5943 3041 2549 5.8e-16
c5944 5484 5479 7.46e-16
c5945 5429 5437 9.34e-16
c5946 5514 5436 1.58e-16
c5947 5509 5510 1.08e-15
c5948 3148 0 8e-16
c5949 1222 1203 1.091e-15
c5950 1046 1042 3.78e-16
c5951 1327 1402 1.96e-16
c5952 3684 3656 2.64e-16
c5953 4124 1 4.64e-16
c5954 3048 2611 5.5e-16
c5955 1380 0 6.9481e-14
c5956 4276 1 6.275e-15
c5957 3005 858 1.58e-16
c5958 2541 827 3.15e-16
c5959 5199 5195 3.54e-16
c5960 792 1578 2.72e-16
c5961 552 565 1.88e-16
c5962 3151 3157 1.418e-15
c5963 3538 3540 1.862e-15
c5964 5039 5100 6.38e-16
c5965 3168 3140 2.64e-16
c5966 2390 2384 1.418e-15
c5967 2373 2401 2.64e-16
c5968 2395 2391 1.96e-16
c5969 702 704 5.59e-16
c5970 2165 0 2.0654e-14
c5971 3397 3411 4.274e-15
c5972 595 2532 1.58e-16
c5973 146 455 1.88e-16
c5974 4364 692 4.81e-16
c5975 2739 0 3.3598e-14
c5976 3731 3752 4.41e-16
c5977 4135 4134 1.58e-16
c5978 4506 4505 2.48e-16
c5979 3316 0 1.4092e-14
c5980 2545 2752 4.63e-16
c5981 3839 3370 7.46e-16
c5982 4085 19 9.67e-16
c5983 2094 2093 1.6e-16
c5984 1257 1211 1.45e-16
c5985 1584 1573 1.58e-16
c5986 291 450 1.88e-16
c5987 3151 717 1.58e-16
c5988 5058 1 7.87e-16
c5989 4861 410 1.88e-16
c5990 1623 827 7.38e-16
c5991 3294 0 1.6491e-14
c5992 2178 2423 1.96e-16
c5993 1106 1110 2.03e-16
c5994 911 3384 1.88e-16
c5995 2541 2333 5.88e-16
c5996 1602 1146 1.96e-16
c5997 1603 1596 6.73e-16
c5998 4677 4689 2.62e-16
c5999 1708 1803 1.58e-16
c6000 3077 3073 1.96e-16
c6001 1387 0 1.6491e-14
c6002 627 3886 7.99e-16
c6003 4196 4566 4.17e-16
c6004 1870 1482 4.97e-16
c6005 3046 2770 1.58e-16
c6006 3034 647 3.15e-16
c6007 3219 3611 2.38e-15
c6008 4429 0 6.8914e-14
c6009 4606 4611 5.53e-16
c6010 4691 0 3.31498e-13
c6011 2477 2478 2.48e-16
c6012 2182 2423 4.63e-16
c6013 2196 777 3.58e-16
c6014 2172 2240 1.58e-16
c6015 2895 1 2.269e-15
c6016 626 1 5.57e-16
c6017 3500 1 1.056e-15
c6018 2333 732 1.813e-15
c6019 1854 1866 2.32e-16
c6020 3418 0 3.5936e-14
c6021 2424 797 2.33e-16
c6022 2194 732 3.15e-16
c6023 4571 752 1.33e-16
c6024 4747 4748 1.6e-16
c6025 4743 4361 1.443e-15
c6026 4800 0 6.72e-16
c6027 2541 812 3.15e-16
c6028 2031 2028 7.84e-16
c6029 767 758 1.078e-15
c6030 245 255 8.86e-16
c6031 470 33 1.88e-16
c6032 3608 767 1.58e-16
c6033 2552 2186 5.8e-16
c6034 5062 5066 1.151e-15
c6035 2330 0 8e-16
c6036 1652 1 1.387e-15
c6037 4770 5219 1.96e-16
c6038 2765 2759 1.6e-16
c6039 1449 662 3.64e-16
c6040 612 2541 4.03e-16
c6041 595 2559 3.15e-16
c6042 602 2535 3.46e-16
c6043 1766 2277 5.66e-16
c6044 4201 4208 1.88e-16
c6045 1343 1317 1.58e-16
c6046 1321 1320 1.58e-16
c6047 598 25 1.13e-15
c6048 2742 747 1.58e-16
c6049 2685 2686 1.35e-16
c6050 1422 1424 2.03e-16
c6051 3886 4416 1.58e-16
c6052 3898 3565 5.5e-16
c6053 3900 3571 1.58e-16
c6054 3650 4468 1.96e-16
c6055 2545 2688 1.58e-16
c6056 998 0 1.4198e-14
c6057 4361 4744 4.97e-16
c6058 1690 1968 1.58e-16
c6059 320 455 1.88e-16
c6060 5068 5070 3.25e-16
c6061 5034 5031 7.84e-16
c6062 2126 1 3.36e-16
c6063 3420 3422 2.03e-16
c6064 627 2223 1.58e-16
c6065 2116 0 1.65e-16
c6066 251 250 2.84e-16
c6067 2682 1 1.056e-15
c6068 747 1694 7.99e-16
c6069 907 1022 3.92e-16
c6070 2720 747 1.58e-16
c6071 2549 2558 1.846e-15
c6072 72 71 5.8e-16
c6073 4111 4104 1.88e-16
c6074 1623 812 1.58e-16
c6075 1538 737 1.58e-16
c6076 4736 5356 2.037e-15
c6077 1684 858 4.48e-16
c6078 1321 1343 4.078e-15
c6079 1345 1327 4.312e-15
c6080 781 1 4.03e-16
c6081 632 1778 3.64e-16
c6082 361 375 3.84e-16
c6083 1366 1 1.056e-15
c6084 1694 1403 1.58e-16
c6085 3310 1 4.41e-15
c6086 2528 858 3.15e-16
c6087 3396 3392 5.8e-16
c6088 1871 1 5.808e-15
c6089 1873 0 3.466e-15
c6090 4773 1 1.013e-15
c6091 762 1505 5.73e-16
c6092 2476 0 1.6491e-14
c6093 5582 0 8e-16
c6094 1947 2440 1.96e-16
c6095 2194 1862 5.5e-16
c6096 2816 2807 3.92e-16
c6097 3058 0 3.3643e-14
c6098 4298 4297 9.1e-16
c6099 1327 1056 1.58e-16
c6100 911 3886 3.45e-16
c6101 2515 852 1.58e-16
c6102 1448 1437 1.58e-16
c6103 1211 1661 1.58e-16
c6104 3313 3311 1.862e-15
c6105 2815 2787 2.64e-16
c6106 2172 692 4.48e-16
c6107 4830 4463 1.58e-16
c6108 2545 782 3.15e-16
c6109 1 263 1.456e-15
c6110 4674 4678 1.81e-16
c6111 4571 4677 1.58e-16
c6112 4582 4689 1.58e-16
c6113 556 497 1.66e-16
c6114 1428 647 1.09e-16
c6115 1173 837 1.05e-15
c6116 827 1178 1.58e-16
c6117 919 963 1.58e-16
c6118 4668 410 1.88e-16
c6119 2254 2282 2.64e-16
c6120 1500 1491 3.92e-16
c6121 1056 1494 5.66e-16
c6122 543 541 1.58e-16
c6123 3031 3033 3.67e-16
c6124 2933 2929 1.583e-15
c6125 3633 4450 1.58e-16
c6126 1902 767 2.33e-16
c6127 956 0 6.29e-16
c6128 3046 3044 1.96e-16
c6129 3030 3043 1.58e-16
c6130 3048 3051 1.6e-16
c6131 1708 1533 5.5e-16
c6132 2357 1845 1.532e-15
c6133 2363 2362 5.65e-16
c6134 4992 1 3.66e-16
c6135 422 9 4.88e-16
c6136 412 1 4.848e-15
c6137 221 233 1.58e-16
c6138 1324 886 1.96e-16
c6139 909 923 3.54e-16
c6140 4569 33 1.88e-16
c6141 4838 0 3.50269e-13
c6142 4182 3918 2.48e-16
c6143 3976 25 7.01e-16
c6144 4369 4370 2.48e-16
c6145 1321 1639 1.58e-16
c6146 1343 1627 1.58e-16
c6147 736 1 4.03e-16
c6148 1555 1106 1.96e-16
c6149 4627 4624 6.67e-16
c6150 1690 1731 1.96e-16
c6151 4368 0 1.6491e-14
c6152 5194 207 6.67e-16
c6153 5162 296 1.345e-15
c6154 1827 1 8.43e-16
c6155 627 1694 7.99e-16
c6156 3276 3658 2.48e-16
c6157 4446 4435 1.58e-16
c6158 2437 1 9.28e-16
c6159 2150 1635 4.78e-16
c6160 596 670 2.45e-16
c6161 1 50 1.607e-15
c6162 3393 868 4.03e-16
c6163 4563 4843 1.96e-16
c6164 5151 5165 5.12e-16
c6165 5264 5259 9.94e-16
c6166 41 0 9.795e-15
c6167 2407 0 3.6368e-14
c6168 3548 3157 1.136e-15
c6169 3990 3918 2.48e-16
c6170 642 993 1.58e-16
c6171 632 978 1.58e-16
c6172 3017 0 2.0654e-14
c6173 698 0 1.1435e-14
c6174 2838 2839 1.35e-16
c6175 1556 797 1.75e-16
c6176 1750 1369 3.92e-16
c6177 3577 0 1.4092e-14
c6178 4231 4609 7.84e-16
c6179 4179 1 6.78e-16
c6180 1103 1 4.59e-16
c6181 4891 4884 6.73e-16
c6182 4890 4503 1.96e-16
c6183 1100 0 1.0077e-14
c6184 3046 3189 1.58e-16
c6185 3030 3177 1.58e-16
c6186 4429 4815 4.11e-16
c6187 2133 2139 6.23e-16
c6188 5232 5198 1.58e-16
c6189 292 296 6.38e-16
c6190 2408 2419 1.96e-16
c6191 2240 0 3.3692e-14
c6192 2342 2341 2.48e-16
c6193 1178 812 3.57e-16
c6194 1158 1171 1.58e-16
c6195 42 0 4.5547e-14
c6196 55 5 9.5e-16
c6197 3548 717 3.79e-16
c6198 4370 722 1.58e-16
c6199 2709 2707 1.6e-16
c6200 2704 2703 2.03e-16
c6201 2541 2786 1.96e-16
c6202 3957 1 7.19e-16
c6203 612 3429 3.79e-16
c6204 601 4262 4.81e-16
c6205 4436 4447 1.96e-16
c6206 3948 26 4.58e-16
c6207 3937 0 2.299e-14
c6208 2839 842 1.339e-15
c6209 1601 1 5.97e-15
c6210 3411 3659 1.58e-16
c6211 3397 3672 4.63e-16
c6212 2773 0 3.3717e-14
c6213 1087 1089 7.84e-16
c6214 894 905 3.92e-16
c6215 596 861 5.28e-16
c6216 3710 3717 1.96e-16
c6217 2170 0 6.9778e-14
c6218 3616 3611 1.642e-15
c6219 1587 782 4.81e-16
c6220 4582 4571 4.763e-15
c6221 4651 5481 9.43e-16
c6222 2559 2586 1.58e-16
c6223 617 982 1.58e-16
c6224 3514 4332 1.96e-16
c6225 1627 1639 2.32e-16
c6226 4329 1 9.28e-16
c6227 1903 1522 3.92e-16
c6228 1907 1908 1.6e-16
c6229 3046 717 3.15e-16
c6230 5291 5288 1.96e-16
c6231 890 893 1.96e-16
c6232 3625 3637 2.32e-16
c6233 2591 0 8e-16
c6234 4582 4779 1.58e-16
c6235 4878 468 1.88e-16
c6236 4804 207 1.88e-16
c6237 2493 2495 1.862e-15
c6238 1981 1987 1.418e-15
c6239 3937 3944 3.84e-16
c6240 3948 3947 4.41e-16
c6241 3164 0 6.72e-16
c6242 922 1085 3.92e-16
c6243 595 3387 1.511e-15
c6244 2541 747 4.03e-16
c6245 1924 782 5.03e-16
c6246 3104 3105 9.1e-16
c6247 687 1459 2.72e-16
c6248 3363 2849 4.78e-16
c6249 3030 2821 1.58e-16
c6250 911 1694 3.45e-16
c6251 2866 2475 1.136e-15
c6252 1600 1 8.43e-16
c6253 4293 1 6.275e-15
c6254 4782 4779 5.5e-16
c6255 3387 3468 3.92e-16
c6256 2557 852 3.15e-16
c6257 2072 2029 2.15e-16
c6258 422 419 2.142e-15
c6259 5198 5190 3.54e-16
c6260 302 303 1.482e-15
c6261 2196 2286 5.42e-16
c6262 3706 3387 3.92e-16
c6263 3785 3773 5.37e-16
c6264 59 565 1.88e-16
c6265 4233 4234 2.48e-16
c6266 2541 2384 5.88e-16
c6267 2299 2666 1.58e-16
c6268 1327 1401 1.58e-16
c6269 2584 2586 1.862e-15
c6270 2170 2203 1.418e-15
c6271 1445 1442 3.01e-16
c6272 1441 1438 6.44e-16
c6273 4104 0 2.0592e-14
c6274 692 0 2.80135e-13
c6275 2070 2093 1.96e-16
c6276 1706 2020 3.92e-16
c6277 3171 3169 1.6e-16
c6278 3639 1 4.41e-15
c6279 1584 1982 4.36e-16
c6280 1980 1973 1.96e-16
c6281 792 1572 2.4e-16
c6282 4580 4578 1.96e-16
c6283 4563 4577 1.58e-16
c6284 702 709 1.6e-16
c6285 4473 0 6.62e-16
c6286 3185 702 2.22e-16
c6287 3557 707 1.832e-15
c6288 3696 3703 6.73e-16
c6289 4949 4950 2.423e-15
c6290 4941 4944 9.58e-16
c6291 907 717 3.15e-16
c6292 71 117 1.88e-16
c6293 4838 4452 1.179e-15
c6294 2759 762 1.58e-16
c6295 2737 0 1.6491e-14
c6296 2586 2585 2.48e-16
c6297 596 815 5.28e-16
c6298 1640 868 2.4e-16
c6299 2617 1 4.41e-15
c6300 2194 2440 3.92e-16
c6301 411 1 4.92e-16
c6302 4526 842 1.58e-16
c6303 4514 5576 4.78e-16
c6304 1249 1243 1.58e-16
c6305 602 965 1.58e-16
c6306 646 1 4.03e-16
c6307 2266 647 7.68e-16
c6308 1151 1146 1.58e-16
c6309 2301 2300 1.6e-16
c6310 3024 2787 1.58e-16
c6311 3024 677 4.48e-16
c6312 2206 2205 2.48e-16
c6313 1539 0 3.6368e-14
c6314 2776 2384 2.38e-15
c6315 4446 0 6.9337e-14
c6316 2031 2095 1.6e-16
c6317 2178 2422 1.58e-16
c6318 4419 767 1.339e-15
c6319 1220 858 5.74e-16
c6320 3164 3162 1.6e-16
c6321 3660 0 6.62e-16
c6322 1524 1086 2.48e-16
c6323 1321 1367 1.58e-16
c6324 1343 1355 1.58e-16
c6325 397 59 1.88e-16
c6326 1158 0 4.6723e-14
c6327 4080 1 2.8425e-14
c6328 1744 1 1.868e-15
c6329 4817 0 6.72e-16
c6330 3169 692 7.68e-16
c6331 1734 0 2.93e-15
c6332 4708 4327 5.2e-16
c6333 4582 4724 3.92e-16
c6334 3411 3415 1.6e-16
c6335 2350 1 5.97e-15
c6336 642 2220 5.73e-16
c6337 2196 1902 1.58e-16
c6338 2182 2422 1.58e-16
c6339 747 1862 1.813e-15
c6340 2346 0 6.72e-16
c6341 2150 1 4.03e-16
c6342 5452 5473 1.96e-16
c6343 4770 5198 3.54e-16
c6344 1217 852 2.68e-16
c6345 627 2541 4.03e-16
c6346 601 2535 4.48e-16
c6347 910 3872 1.58e-16
c6348 2854 2469 1.96e-16
c6349 2663 2652 1.96e-16
c6350 1345 877 1.58e-16
c6351 657 1423 1.58e-16
c6352 3279 1 5.808e-15
c6353 642 919 3.15e-16
c6354 807 25 1.58e-16
c6355 3886 4421 1.58e-16
c6356 3876 3582 5.5e-16
c6357 1919 807 5.73e-16
c6358 1797 1795 1.6e-16
c6359 3370 1 5.051e-15
c6360 4055 37 1.88e-16
c6361 2753 792 5.73e-16
c6362 3162 692 5.03e-16
c6363 1706 1985 1.58e-16
c6364 1690 1973 1.58e-16
c6365 30 355 6.83e-16
c6366 198 204 1.58e-16
c6367 197 187 8.86e-16
c6368 3521 692 1.339e-15
c6369 627 2243 1.58e-16
c6370 157 175 1.58e-16
c6371 2698 1 9.28e-16
c6372 883 677 6.45e-16
c6373 909 1037 4.35e-16
c6374 907 1036 1.88e-16
c6375 890 1029 1.58e-16
c6376 4319 662 1.832e-15
c6377 2656 2652 1.96e-16
c6378 5587 1 8.88e-16
c6379 4651 468 1.88e-16
c6380 2567 2568 2.03e-16
c6381 2136 2133 7.46e-16
c6382 3268 1 6.15e-16
c6383 1327 782 3.15e-16
c6384 1322 1324 1.578e-15
c6385 1337 1330 7.06e-16
c6386 3565 3537 2.64e-16
c6387 3548 3554 1.418e-15
c6388 4385 4387 1.862e-15
c6389 3264 777 2.72e-16
c6390 2351 722 7.68e-16
c6391 657 1380 1.58e-16
c6392 632 1397 3.15e-16
c6393 542 407 1.88e-16
c6394 3236 1 5.97e-15
c6395 3393 0 3.63418e-13
c6396 3167 2645 1.96e-16
c6397 1331 1521 4.63e-16
c6398 4658 4282 3.92e-16
c6399 4670 4669 1.6e-16
c6400 3057 3059 2.03e-16
c6401 5372 354 5.93e-16
c6402 3339 842 7.68e-16
c6403 3332 827 1.9e-16
c6404 627 2221 1.58e-16
c6405 1891 1 2.054e-15
c6406 1893 0 8e-16
c6407 3393 3586 1.58e-16
c6408 4790 1 1.013e-15
c6409 3254 752 3.64e-16
c6410 762 1914 2.65e-16
c6411 1 468 3.36e-15
c6412 4104 4102 3.54e-16
c6413 4567 4480 5.5e-16
c6414 5287 5288 5.87e-16
c6415 5177 5184 3.18e-16
c6416 5170 5157 1.58e-16
c6417 448 0 4.512e-14
c6418 4103 857 6.23e-16
c6419 911 3383 1.88e-16
c6420 1295 1236 1.066e-15
c6421 5536 5568 1.738e-15
c6422 4878 64 1.88e-16
c6423 3078 0 1.4092e-14
c6424 922 1143 1.58e-16
c6425 1448 1846 4.36e-16
c6426 1844 1837 1.96e-16
c6427 3410 3404 1.988e-15
c6428 3024 3241 3.92e-16
c6429 3247 752 1.9e-16
c6430 1685 0 1.4835e-14
c6431 100 19 3.84e-16
c6432 4691 4693 4.93e-16
c6433 4571 4694 1.58e-16
c6434 4582 4706 1.58e-16
c6435 2453 2444 3.92e-16
c6436 1936 2447 5.66e-16
c6437 1947 2439 1.58e-16
c6438 0 186 9.795e-15
c6439 3803 3739 2.249e-15
c6440 3806 3811 3.73e-16
c6441 1420 662 2.33e-16
c6442 883 1128 3.54e-16
c6443 894 1149 1.58e-16
c6444 2842 0 6.62e-16
c6445 1880 737 7.68e-16
c6446 147 152 1.059e-15
c6447 139 129 8.86e-16
c6448 4600 5558 1.383e-15
c6449 3616 4458 2.38e-15
c6450 1896 782 1.58e-16
c6451 4546 4555 1.6e-16
c6452 1517 1 1.868e-15
c6453 1507 0 2.93e-15
c6454 4568 0 1.1567e-14
c6455 5059 5058 1.6e-16
c6456 279 1 3.6e-16
c6457 911 2541 7.6e-16
c6458 894 963 3.54e-16
c6459 2136 2083 9.01e-16
c6460 1414 672 1.813e-15
c6461 1593 797 1.832e-15
c6462 1331 752 3.15e-16
c6463 632 3435 1.75e-16
c6464 3241 762 2.4e-16
c6465 2611 3109 1.58e-16
c6466 1306 1 2.4e-16
c6467 1931 1925 1.6e-16
c6468 1533 1922 2.386e-15
c6469 1706 1748 3.92e-16
c6470 4531 4503 2.64e-16
c6471 3046 3380 4.22e-16
c6472 4446 4452 9.42e-16
c6473 4889 0 4.5906e-14
c6474 2450 1 6.15e-16
c6475 242 0 2.87e-16
c6476 792 2429 2.72e-16
c6477 151 1 4.848e-15
c6478 3898 752 4.46e-16
c6479 4472 807 1.58e-16
c6480 657 998 1.58e-16
c6481 4036 2175 2.573e-15
c6482 3701 3886 5.5e-16
c6483 3707 4540 1.361e-15
c6484 1981 842 3.15e-16
c6485 2497 868 2.72e-16
c6486 617 1391 1.9e-16
c6487 2787 3295 2.48e-16
c6488 3024 3206 1.58e-16
c6489 3046 3194 1.58e-16
c6490 4709 0 1.6462e-14
c6491 2011 2009 1.6e-16
c6492 2006 2005 2.03e-16
c6493 1648 0 6.72e-16
c6494 0 274 4.3729e-14
c6495 26 291 8.41e-16
c6496 27 305 1.88e-16
c6497 233 570 1.88e-16
c6498 3411 702 3.58e-16
c6499 5152 5154 5.62e-16
c6500 5176 5175 1.6e-16
c6501 4793 439 1.88e-16
c6502 910 2170 3.45e-16
c6503 2196 2355 3.92e-16
c6504 891 916 2.82e-16
c6505 1178 1179 1.213e-15
c6506 986 989 6.13e-16
c6507 361 368 7.76e-16
c6508 5434 5425 1.96e-16
c6509 5409 5439 9.6e-16
c6510 2333 2701 1.96e-16
c6511 160 78 1.88e-16
c6512 1481 1031 1.96e-16
c6513 1476 1041 1.96e-16
c6514 642 957 1.58e-16
c6515 627 3429 1.813e-15
c6516 2896 2895 1.334e-15
c6517 4817 4815 1.6e-16
c6518 3118 647 7.68e-16
c6519 3487 3498 1.96e-16
c6520 2238 0 1.6491e-14
c6521 2346 2344 1.6e-16
c6522 2341 2340 2.03e-16
c6523 13 14 6.96e-16
c6524 7 1 8.75e-16
c6525 3393 3287 5.88e-16
c6526 4569 526 3.92e-16
c6527 3367 0 1.3715e-14
c6528 1396 957 1.96e-16
c6529 3900 4319 1.58e-16
c6530 4651 64 1.88e-16
c6531 2541 2220 1.58e-16
c6532 899 0 6.35e-16
c6533 682 1 5.62e-16
c6534 4342 1 6.15e-16
c6535 4429 4424 1.642e-15
c6536 1708 1698 5.5e-16
c6537 3089 3117 2.64e-16
c6538 777 921 3.15e-16
c6539 3470 647 1.339e-15
c6540 3034 3360 4.63e-16
c6541 3292 797 7.38e-16
c6542 3185 3180 1.642e-15
c6543 2178 1698 3.15e-16
c6544 1658 1652 9.59e-16
c6545 2103 2118 1.739e-15
c6546 1 517 2.87e-16
c6547 4582 4796 1.58e-16
c6548 5229 5224 1.493e-15
c6549 5240 5241 3.92e-16
c6550 102 103 1.079e-15
c6551 64 1 2.4201e-14
c6552 2866 3809 1.12e-15
c6553 1244 1246 5.87e-16
c6554 3514 4331 1.58e-16
c6555 3503 4339 5.66e-16
c6556 4345 4336 3.92e-16
c6557 2300 662 3.64e-16
c6558 1211 852 3.15e-16
c6559 919 1099 1.58e-16
c6560 3540 1 5.808e-15
c6561 1944 782 1.09e-16
c6562 1540 1101 3.92e-16
c6563 1544 1545 1.6e-16
c6564 1345 1419 3.92e-16
c6565 4594 3873 1.96e-16
c6566 3542 0 3.466e-15
c6567 2957 2518 1.794e-15
c6568 2995 2136 1.389e-15
c6569 3752 1 8.09e-16
c6570 3046 2838 1.58e-16
c6571 4863 4480 4.97e-16
c6572 4866 4862 1.96e-16
c6573 4310 1 6.275e-15
c6574 3262 3274 2.32e-16
c6575 2182 1698 1.58e-16
c6576 229 187 9.5e-16
c6577 3411 3485 3.92e-16
c6578 592 640 6.34e-16
c6579 5224 5227 1.18e-15
c6580 0 328 2.87e-16
c6581 3568 3566 1.6e-16
c6582 4563 4196 9.51e-16
c6583 4844 352 1.88e-16
c6584 2196 2291 1.58e-16
c6585 2220 2221 1.35e-16
c6586 381 30 3.84e-16
c6587 907 1235 5.04e-16
c6588 601 2566 2.33e-16
c6589 595 2577 2.22e-16
c6590 919 732 3.15e-16
c6591 4838 5083 1.96e-16
c6592 2671 2299 1.58e-16
c6593 1343 1418 1.58e-16
c6594 1327 1406 1.58e-16
c6595 1319 1320 3.36e-16
c6596 59 60 7.03e-16
c6597 1833 692 7.38e-16
c6598 1642 858 1.339e-15
c6599 595 1358 1.58e-16
c6600 3882 4484 1.58e-16
c6601 1355 1367 2.32e-16
c6602 4422 4419 6.44e-16
c6603 4426 4423 3.01e-16
c6604 2557 2768 1.58e-16
c6605 2541 2756 1.58e-16
c6606 2389 737 1.58e-16
c6607 1059 0 2.7376e-14
c6608 5038 180 7.97e-16
c6609 2070 2126 9.34e-16
c6610 4498 1 1.868e-15
c6611 1694 1850 4.63e-16
c6612 707 698 1.078e-15
c6613 4488 0 2.93e-15
c6614 4970 4905 6.67e-16
c6615 3046 842 4.46e-16
c6616 3034 868 7.99e-16
c6617 2308 2317 3.92e-16
c6618 2311 1800 5.66e-16
c6619 1811 2303 1.58e-16
c6620 2181 0 1.5577e-14
c6621 3411 3869 3.54e-16
c6622 3393 3863 1.96e-16
c6623 3429 3021 1.136e-15
c6624 1682 1715 1.418e-15
c6625 1726 1681 2.64e-16
c6626 2888 352 9.43e-16
c6627 2169 1 4.044e-15
c6628 1343 837 3.15e-16
c6629 601 3419 1.339e-15
c6630 3152 1 1.868e-15
c6631 2172 2457 3.92e-16
c6632 4521 852 1.58e-16
c6633 4640 5412 2.45e-16
c6634 2645 2640 1.642e-15
c6635 2545 2166 3.54e-16
c6636 601 965 6.31e-16
c6637 1151 1619 4.36e-16
c6638 1617 1610 1.96e-16
c6639 1327 1555 1.96e-16
c6640 4694 4706 2.62e-16
c6641 1684 1437 1.58e-16
c6642 1690 1431 5.88e-16
c6643 367 361 5.8e-16
c6644 2855 852 1.58e-16
c6645 3034 3325 1.58e-16
c6646 2561 1 2.86e-16
c6647 3236 3225 1.58e-16
c6648 4110 3918 6.32e-16
c6649 4736 439 1.88e-16
c6650 4922 120 1.88e-16
c6651 2194 2439 1.58e-16
c6652 2178 2427 1.58e-16
c6653 1353 1364 1.96e-16
c6654 5403 381 5.11e-16
c6655 2772 2774 2.03e-16
c6656 2003 842 7.38e-16
c6657 1706 752 4.46e-16
c6658 3675 0 2.93e-15
c6659 4223 4217 1.96e-16
c6660 1345 1384 5.42e-16
c6661 1874 1871 5.5e-16
c6662 4094 1 6.76e-16
c6663 3446 0 6.9481e-14
c6664 1363 1 5.97e-15
c6665 2210 2208 1.6e-16
c6666 2205 2204 2.03e-16
c6667 4764 4765 1.6e-16
c6668 4760 4378 1.443e-15
c6669 4834 0 6.72e-16
c6670 2662 692 3.15e-16
c6671 2036 2023 5.78e-16
c6672 537 536 1.88e-16
c6673 1 451 1.65e-15
c6674 13 450 1.88e-16
c6675 4582 4741 3.92e-16
c6676 3397 3434 4.63e-16
c6677 3411 3421 1.58e-16
c6678 642 2629 2.65e-16
c6679 632 2214 1.58e-16
c6680 2182 2427 1.58e-16
c6681 0 449 1.5696e-14
c6682 3919 3909 1.88e-16
c6683 907 842 4.8e-16
c6684 883 1202 3.92e-16
c6685 890 1201 1.88e-16
c6686 2722 1 5.808e-15
c6687 617 2535 4.48e-16
c6688 5400 5396 1.243e-15
c6689 910 3393 7.97e-16
c6690 3299 1 2.054e-15
c6691 1439 1001 4.97e-16
c6692 3900 3599 5.5e-16
c6693 2832 2838 1.418e-15
c6694 2282 647 1.58e-16
c6695 2453 807 2.65e-16
c6696 3288 792 2.65e-16
c6697 1685 1689 1.988e-15
c6698 1684 2002 1.58e-16
c6699 1706 1990 1.58e-16
c6700 1958 1954 1.96e-16
c6701 3909 3914 1.96e-16
c6702 5025 5077 1.39e-16
c6703 186 188 2.84e-16
c6704 5391 265 3.54e-16
c6705 3712 858 5.03e-16
c6706 2853 2469 1.58e-16
c6707 2711 1 6.15e-16
c6708 3277 1 1.716e-15
c6709 1808 662 1.09e-16
c6710 1434 1432 1.6e-16
c6711 2887 2913 3.54e-16
c6712 642 894 8.34e-16
c6713 1338 1326 3.225e-15
c6714 1328 1324 2.074e-15
c6715 3882 4247 1.96e-16
c6716 1845 722 3.15e-16
c6717 2361 732 2.72e-16
c6718 3653 1 1.056e-15
c6719 910 1685 7.06e-16
c6720 1370 1 1.716e-15
c6721 266 263 6.67e-16
c6722 3432 3430 1.6e-16
c6723 3022 3386 1.62e-16
c6724 2832 842 3.15e-16
c6725 3349 868 2.72e-16
c6726 1909 0 6.72e-16
c6727 4807 1 1.013e-15
c6728 2747 752 3.15e-16
c6729 2495 1 5.808e-15
c6730 777 1516 1.58e-16
c6731 1057 702 1.58e-16
c6732 4567 4497 5.5e-16
c6733 4685 352 7.45e-16
c6734 4844 294 1.88e-16
c6735 2497 0 3.466e-15
c6736 2458 2459 1.35e-16
c6737 2015 1624 1.136e-15
c6738 2545 2503 3.92e-16
c6739 2518 2510 5.95e-16
c6740 1345 1071 1.58e-16
c6741 1343 1061 5.5e-16
c6742 1331 1520 1.58e-16
c6743 3384 1 4.044e-15
c6744 1149 1 2.972e-15
c6745 1150 0 6.29e-16
c6746 4219 25 7.01e-16
c6747 4235 0 6.62e-16
c6748 1691 0 4.1004e-14
c6749 1 359 4.22e-16
c6750 5010 91 1.88e-16
c6751 1947 2444 1.58e-16
c6752 955 961 2.32e-16
c6753 4319 3486 7.84e-16
c6754 5173 236 9.42e-16
c6755 2867 1 1.868e-15
c6756 1194 842 1.58e-16
c6757 5447 5457 1.462e-15
c6758 5358 5360 1.001e-15
c6759 5356 5353 3.54e-16
c6760 2857 0 2.93e-15
c6761 3898 3883 1.632e-15
c6762 1499 737 3.15e-16
c6763 4218 37 1.88e-16
c6764 2438 782 4.81e-16
c6765 1930 767 1.58e-16
c6766 1708 1420 1.58e-16
c6767 1768 1380 4.97e-16
c6768 963 1 1.56e-15
c6769 3156 677 7.38e-16
c6770 3024 2532 1.58e-16
c6771 3030 2529 1.58e-16
c6772 2026 2030 5.6e-16
c6773 1076 1 5.821e-15
c6774 0 252 1.10918e-13
c6775 2196 2179 3.62e-16
c6776 4537 4991 7.46e-16
c6777 401 390 2.45e-16
c6778 410 412 1.96e-16
c6779 5358 5367 1.96e-16
c6780 2822 2435 1.532e-15
c6781 1113 752 1.58e-16
c6782 632 4294 3.64e-16
c6783 4758 737 1.23e-16
c6784 3227 3229 2.03e-16
c6785 1327 1191 1.58e-16
c6786 4644 4641 6.67e-16
c6787 1332 1 3.009e-15
c6788 4387 1 5.808e-15
c6789 687 2310 2.72e-16
c6790 1684 1765 3.92e-16
c6791 4389 0 3.466e-15
c6792 1333 0 5.86e-16
c6793 3509 672 1.58e-16
c6794 4549 3718 1.96e-16
c6795 4889 4918 9.36e-16
c6796 3411 3151 5.5e-16
c6797 3287 3675 4.97e-16
c6798 2459 1 1.716e-15
c6799 1050 677 6.48e-16
c6800 281 274 7.76e-16
c6801 9 130 6.48e-16
c6802 1 122 4.848e-15
c6803 4736 4731 1.536e-15
c6804 3900 3390 3.54e-16
c6805 5532 5535 3.54e-16
c6806 1506 737 1.339e-15
c6807 1272 1275 6.21e-16
c6808 1967 797 4.81e-16
c6809 1568 1562 1.6e-16
c6810 1106 1559 2.386e-15
c6811 4248 4626 7.84e-16
c6812 3208 0 3.6368e-14
c6813 1291 0 2.285e-15
c6814 1124 1 3.06e-16
c6815 1822 1818 1.96e-16
c6816 4181 0 1.5176e-14
c6817 3048 3223 5.42e-16
c6818 3024 3211 1.58e-16
c6819 1823 0 1.4092e-14
c6820 4446 4832 4.11e-16
c6821 1641 2151 1.361e-15
c6822 1635 1694 5.5e-16
c6823 4726 0 1.6462e-14
c6824 1666 0 8e-16
c6825 3393 707 3.15e-16
c6826 2434 1913 1.96e-16
c6827 2429 1919 1.96e-16
c6828 3822 3809 1.96e-16
c6829 3355 3344 1.58e-16
c6830 3033 0 1.5577e-14
c6831 657 3393 4.03e-16
c6832 4810 5051 1.96e-16
c6833 3898 4536 3.92e-16
c6834 3034 0 3.24424e-13
c6835 2882 2900 4.06e-16
c6836 2559 2803 3.92e-16
c6837 932 1 4.05e-16
c6838 752 26 7.12e-16
c6839 3989 0 1.5176e-14
c6840 1648 1646 1.6e-16
c6841 1643 1642 2.03e-16
c6842 3718 3707 1.58e-16
c6843 3886 1 4.57e-15
c6844 2860 858 5.03e-16
c6845 1 585 5.62e-16
c6846 4538 0 1.7575e-14
c6847 2013 1 6.15e-16
c6848 3858 3860 1.6e-16
c6849 3344 3854 1.96e-16
c6850 632 3095 1.84e-16
c6851 1845 2338 1.96e-16
c6852 234 1 1.456e-15
c6853 5326 5286 2.45e-16
c6854 2793 2407 5.66e-16
c6855 2620 2618 1.862e-15
c6856 1102 1103 7.46e-16
c6857 592 863 1.96e-16
c6858 1408 971 4.11e-16
c6859 3882 3503 1.58e-16
c6860 2557 2802 1.58e-16
c6861 2541 2790 1.58e-16
c6862 2196 647 3.15e-16
c6863 3228 747 1.58e-16
c6864 2557 2237 1.58e-16
c6865 3951 19 3.84e-16
c6866 3960 0 2.0707e-14
c6867 1331 1151 5.5e-16
c6868 747 754 1.6e-16
c6869 4351 1 1.716e-15
c6870 3116 2594 1.96e-16
c6871 3111 2600 1.96e-16
c6872 1026 0 3.7577e-14
c6873 4915 4917 9.29e-16
c6874 792 920 3.15e-16
c6875 3487 672 1.58e-16
c6876 4132 3404 1.96e-16
c6877 4915 31 3.84e-16
c6878 3645 3642 5.5e-16
c6879 2390 1 4.41e-15
c6880 2604 0 6.62e-16
c6881 812 802 6.38e-16
c6882 407 565 1.88e-16
c6883 642 3066 1.58e-16
c6884 4582 4813 1.58e-16
c6885 5481 410 5.5e-16
c6886 2527 2525 1.6e-16
c6887 881 1375 2.38e-15
c6888 3176 0 2.93e-15
c6889 2795 2792 3.01e-16
c6890 2791 2788 6.44e-16
c6891 3514 4336 1.58e-16
c6892 1794 662 3.15e-16
c6893 3560 1 2.054e-15
c6894 2559 762 3.58e-16
c6895 2015 2178 4.3e-16
c6896 674 0 7.709e-15
c6897 1708 1680 3.54e-16
c6898 3600 747 2.65e-16
c6899 4525 4526 1.6e-16
c6900 4521 3690 3.92e-16
c6901 2899 2897 1.186e-15
c6902 911 2175 1.58e-16
c6903 2764 807 1.58e-16
c6904 4799 4796 5.5e-16
c6905 2679 732 1.58e-16
c6906 1 554 4.92e-16
c6907 3409 3501 1.58e-16
c6908 2316 1800 1.136e-15
c6909 2223 1 5.808e-15
c6910 19 552 3.84e-16
c6911 3397 662 3.15e-16
c6912 4567 4605 3.92e-16
c6913 5409 468 5.5e-16
c6914 4725 497 1.88e-16
c6915 596 868 1.96e-16
c6916 617 2566 1.75e-16
c6917 920 737 3.69e-16
c6918 3310 837 1.58e-16
c6919 3321 858 1.58e-16
c6920 2559 2401 5.5e-16
c6921 2691 2299 2.38e-15
c6922 2015 2182 3.92e-16
c6923 2614 2612 1.6e-16
c6924 602 603 1.621e-15
c6925 3593 747 2.72e-16
c6926 1206 1207 8.58e-16
c6927 3882 4489 1.58e-16
c6928 3898 4501 1.58e-16
c6929 3690 4522 2.48e-16
c6930 1431 1786 1.58e-16
c6931 1718 1725 1.96e-16
c6932 1694 1335 1.58e-16
c6933 866 1 3.79e-16
c6934 3265 3272 6.73e-16
c6935 3175 2668 3.92e-16
c6936 1596 0 1.4092e-14
c6937 3174 3556 2.48e-16
c6938 3667 1 5.97e-15
c6939 2212 1 6.15e-16
c6940 2000 1999 1.6e-16
c6941 1992 1990 2.15e-16
c6942 480 477 2.142e-15
c6943 313 320 3.54e-16
c6944 308 303 1.482e-15
c6945 5148 5144 1.243e-15
c6946 497 495 6.01e-16
c6947 3473 3470 6.44e-16
c6948 3477 3474 3.01e-16
c6949 3174 722 1.75e-16
c6950 3364 852 2.8e-16
c6951 3048 858 3.15e-16
c6952 2308 1811 1.58e-16
c6953 894 732 8.34e-16
c6954 5323 5328 3.07e-16
c6955 5262 5200 6.96e-16
c6956 1431 702 1.58e-16
c6957 1011 1440 7.84e-16
c6958 3349 0 3.466e-15
c6959 397 407 1.88e-16
c6960 108 106 1.58e-16
c6961 3886 3463 5.5e-16
c6962 3707 858 3.69e-16
c6963 2787 822 5.73e-16
c6964 3152 2634 1.96e-16
c6965 1720 1315 4.11e-16
c6966 869 1 1.65e-16
c6967 627 980 1.85e-16
c6968 1426 1 2.054e-15
c6969 4497 3656 1.136e-15
c6970 1985 1986 9.1e-16
c6971 1708 1454 1.58e-16
c6972 1706 1448 5.5e-16
c6973 1694 1849 1.58e-16
c6974 1428 0 8e-16
c6975 362 364 1.58e-16
c6976 345 346 6.4e-16
c6977 2306 2317 1.96e-16
c6978 3034 3330 1.58e-16
c6979 2172 2456 1.58e-16
c6980 2194 2444 1.58e-16
c6981 393 9 4.88e-16
c6982 383 1 4.848e-15
c6983 384 0 1.4515e-14
c6984 4440 782 5.03e-16
c6985 5417 5478 6.38e-16
c6986 3304 1 5.97e-15
c6987 2680 2288 1.96e-16
c6988 4123 1 6.78e-16
c6989 1780 1 1.056e-15
c6990 4851 0 6.72e-16
c6991 2730 3254 4.36e-16
c6992 2102 2098 5.87e-16
c6993 3393 3022 5.5e-16
c6994 632 2631 4.81e-16
c6995 2196 1930 5.5e-16
c6996 3634 782 7.68e-16
c6997 909 858 3.15e-16
c6998 883 1216 1.88e-16
c6999 907 1209 1.58e-16
c7000 3882 662 3.15e-16
c7001 5450 5492 3.15e-16
c7002 2742 1 2.054e-15
c7003 1525 1537 2.32e-16
c7004 1331 952 1.58e-16
c7005 612 592 5.8e-16
c7006 2444 812 1.58e-16
c7007 1947 807 3.79e-16
c7008 1698 1701 2.109e-15
c7009 4070 26 4.48e-16
c7010 1691 1689 8.67e-16
c7011 642 1 4.1542e-14
c7012 2730 3247 4.11e-16
c7013 3173 702 2.4e-16
c7014 3034 3122 4.63e-16
c7015 3066 3061 1.642e-15
c7016 2066 2069 3.54e-16
c7017 3523 3535 2.32e-16
c7018 1694 1 4.57e-15
c7019 3627 782 5.03e-16
c7020 3542 707 5.03e-16
c7021 3347 858 1.58e-16
c7022 2149 0 1.7608e-14
c7023 2858 2469 2.386e-15
c7024 2841 2486 1.58e-16
c7025 2720 1 1.716e-15
c7026 894 1051 1.58e-16
c7027 907 1023 3.54e-16
c7028 5587 4531 3.38e-16
c7029 3303 1 8.43e-16
c7030 823 1 1.65e-16
c7031 3898 4264 3.92e-16
c7032 3250 3247 3.01e-16
c7033 3246 3243 6.44e-16
c7034 1595 1591 1.96e-16
c7035 792 796 2.19e-16
c7036 1396 1 8.43e-16
c7037 4687 4686 1.6e-16
c7038 2816 797 3.64e-16
c7039 3605 0 3.6368e-14
c7040 4946 4991 1.811e-15
c7041 4977 4978 5.88e-16
c7042 5277 354 3.54e-16
c7043 4936 4947 6.73e-16
c7044 617 2242 1.9e-16
c7045 3409 3202 5.5e-16
c7046 4824 1 1.013e-15
c7047 1059 707 1.58e-16
c7048 4708 1 1.8945e-14
c7049 5591 0 2.0051e-14
c7050 4804 497 1.88e-16
c7051 3722 3411 5.42e-16
c7052 3327 3387 1.58e-16
c7053 3882 4246 1.58e-16
c7054 1601 837 1.813e-15
c7055 1321 1076 5.5e-16
c7056 1331 1525 1.58e-16
c7057 3069 3067 1.6e-16
c7058 4260 1 1.868e-15
c7059 2724 722 1.9e-16
c7060 1864 1863 1.6e-16
c7061 1856 1854 2.15e-16
c7062 4250 0 2.93e-15
c7063 5011 5007 1.055e-15
c7064 792 1147 1.58e-16
c7065 4750 4747 3.01e-16
c7066 9 477 5.8e-16
c7067 245 250 1.482e-15
c7068 3219 3604 1.96e-16
c7069 3885 3401 5.8e-16
c7070 5160 5174 1.455e-15
c7071 1947 2464 2.38e-15
c7072 2463 822 2.72e-16
c7073 2172 2219 3.92e-16
c7074 1016 702 1.58e-16
c7075 1188 1202 1.96e-16
c7076 101 0 1.5696e-14
c7077 4205 4204 4.41e-16
c7078 1327 1324 1.123e-15
c7079 4044 1 4.64e-16
c7080 4482 4475 6.73e-16
c7081 4481 3639 1.96e-16
c7082 997 1 3.54e-16
c7083 3329 2821 2.48e-16
c7084 994 0 9.602e-15
c7085 3048 2566 1.58e-16
c7086 3046 2533 5.5e-16
c7087 3034 3087 1.58e-16
c7088 25 172 7.06e-16
c7089 0 169 6.224e-15
c7090 37 171 1.88e-16
c7091 465 570 1.88e-16
c7092 5197 1 1.23e-16
c7093 2082 0 3.0055e-14
c7094 107 508 1.88e-16
c7095 1117 767 6.38e-16
c7096 159 157 2.84e-16
c7097 2654 0 3.3717e-14
c7098 4107 4108 4.41e-16
c7099 4514 4864 2e-16
c7100 642 3463 3.79e-16
c7101 657 3446 1.58e-16
c7102 2545 2667 4.63e-16
c7103 778 1 1.65e-16
c7104 4015 37 1.88e-16
c7105 3394 3038 2.035e-15
c7106 1641 858 3.69e-16
c7107 1206 1343 1.58e-16
c7108 3906 0 3.22e-16
c7109 3387 762 3.15e-16
c7110 3135 2617 1.96e-16
c7111 3136 3129 6.73e-16
c7112 1708 1782 3.92e-16
c7113 1348 0 1.23e-16
c7114 3565 762 1.58e-16
c7115 911 3027 1.58e-16
c7116 5277 5387 1.58e-16
c7117 2485 1 8.43e-16
c7118 273 0 9.795e-15
c7119 3344 858 3.69e-16
c7120 2752 2367 1.96e-16
c7121 2536 2538 1.578e-15
c7122 2551 2544 7.06e-16
c7123 3061 1 2.054e-15
c7124 910 3034 5.03e-16
c7125 1086 1087 8.58e-16
c7126 3063 0 8e-16
c7127 1189 1190 7.51e-16
c7128 2541 2458 1.58e-16
c7129 596 0 2.62685e-13
c7130 4204 1 6.66e-16
c7131 3389 3388 6.67e-16
c7132 837 843 1.097e-15
c7133 3338 3333 1.642e-15
c7134 940 939 1.36e-16
c7135 1 248 1.65e-15
c7136 5073 91 3.54e-16
c7137 1190 837 1.85e-16
c7138 142 19 3.45e-16
c7139 3446 3452 1.418e-15
c7140 4283 4285 1.862e-15
c7141 4396 737 7.68e-16
c7142 5412 5407 7.46e-16
c7143 5410 5434 6.16e-16
c7144 1690 662 3.15e-16
c7145 919 980 3.92e-16
c7146 922 979 2.54e-16
c7147 543 552 1.58e-16
c7148 3383 1 2.346e-15
c7149 1493 1046 4.11e-16
c7150 3900 3882 4.312e-15
c7151 3876 3898 4.078e-15
c7152 3398 0 1.157e-14
c7153 3030 792 4.03e-16
c7154 2945 2944 1.6e-16
c7155 4834 4832 1.6e-16
c7156 2702 3211 7.84e-16
c7157 2015 852 3.15e-16
c7158 2016 2007 3.92e-16
c7159 1624 2010 5.66e-16
c7160 1690 1918 1.96e-16
c7161 479 204 1.88e-16
c7162 5159 5157 5.25e-16
c7163 2196 2359 1.58e-16
c7164 353 350 6.67e-16
c7165 303 345 9.5e-16
c7166 5388 5387 5.5e-16
c7167 221 222 2.84e-16
c7168 4821 1 2.7885e-14
c7169 4600 0 4.8442e-13
c7170 3898 3520 1.58e-16
c7171 1319 1744 4.36e-16
c7172 733 1 1.65e-16
c7173 4377 1 8.43e-16
c7174 4539 0 3.26e-15
c7175 1708 1718 1.58e-16
c7176 204 189 1.88e-16
c7177 1834 2345 5.66e-16
c7178 3491 662 5.03e-16
c7179 3030 737 3.15e-16
c7180 14 27 1.58e-16
c7181 4582 4830 1.58e-16
c7182 2705 2350 1.58e-16
c7183 2619 0 2.93e-15
c7184 2541 1 2.824e-15
c7185 64 410 1.88e-16
c7186 3616 797 1.58e-16
c7187 4702 5286 2.675e-15
c7188 632 995 5.74e-16
c7189 3514 4356 2.38e-15
c7190 1343 1606 3.92e-16
c7191 2705 2717 2.32e-16
c7192 4611 4231 1.96e-16
c7193 2545 2535 4.116e-15
c7194 1255 0 2.078e-15
c7195 3024 2849 5.5e-16
c7196 2194 807 3.15e-16
c7197 792 890 3.35e-16
c7198 747 592 5.8e-16
c7199 3117 672 1.813e-15
c7200 4880 4497 4.97e-16
c7201 4883 4879 1.96e-16
c7202 3282 3279 5.5e-16
c7203 3211 722 1.832e-15
c7204 2713 717 2.22e-16
c7205 3034 2662 5.5e-16
c7206 1 508 4.7546e-14
c7207 3642 3649 1.96e-16
c7208 1022 647 1.58e-16
c7209 3572 3191 3.92e-16
c7210 2243 1 2.054e-15
c7211 19 520 8.4e-16
c7212 3276 807 1.58e-16
c7213 4571 601 1.33e-16
c7214 4567 4622 3.92e-16
c7215 2406 1896 1.96e-16
c7216 2172 1800 1.58e-16
c7217 2178 1794 5.88e-16
c7218 1245 1248 7.1e-16
c7219 59 19 3.84e-16
c7220 55 37 1.88e-16
c7221 3373 2892 6.17e-16
c7222 3840 3842 3.92e-16
c7223 617 3101 3.64e-16
c7224 612 2594 2.22e-16
c7225 1345 1423 1.58e-16
c7226 4161 4158 1.76e-16
c7227 732 1 4.1542e-14
c7228 612 1375 1.58e-16
c7229 3898 4506 1.58e-16
c7230 3876 4518 1.58e-16
c7231 2464 827 1.84e-16
c7232 4134 19 7.04e-16
c7233 4149 0 1.5176e-14
c7234 1073 0 1.4198e-14
c7235 4796 4803 1.96e-16
c7236 2753 2764 1.58e-16
c7237 2104 2125 6.16e-16
c7238 2106 2105 1.624e-15
c7239 602 1721 1.58e-16
c7240 2559 722 3.15e-16
c7241 2221 1 1.716e-15
c7242 4580 3870 1.58e-16
c7243 4582 3873 1.58e-16
c7244 2182 1794 5.5e-16
c7245 3583 722 3.64e-16
c7246 5326 323 7.37e-16
c7247 5145 1 3.36e-16
c7248 2328 1811 2.38e-15
c7249 4838 5095 1.96e-16
c7250 2776 1 2.054e-15
c7251 2695 2299 1.96e-16
c7252 890 737 3.15e-16
c7253 907 1097 3.92e-16
c7254 812 807 2.77e-16
c7255 2778 0 8e-16
c7256 2597 1 1.056e-15
c7257 3321 3717 1.96e-16
c7258 5321 5333 8.45e-16
c7259 5284 5286 1.96e-16
c7260 2782 777 2.65e-16
c7261 2220 2602 2.48e-16
c7262 1837 692 1.832e-15
c7263 5577 5587 5.35e-16
c7264 4520 4582 1.58e-16
c7265 4514 4580 5.5e-16
c7266 4640 5450 5.37e-16
c7267 3170 1 9.28e-16
c7268 3588 4421 7.84e-16
c7269 2662 3176 4.97e-16
c7270 2294 677 1.84e-16
c7271 1637 1636 1.6e-16
c7272 1629 1627 2.15e-16
c7273 1684 1465 5.5e-16
c7274 1694 1854 1.58e-16
c7275 1909 1907 1.6e-16
c7276 1904 1903 2.03e-16
c7277 2866 2902 2.31e-16
c7278 632 1749 2.33e-16
c7279 3411 3638 3.92e-16
c7280 5239 178 9.42e-16
c7281 5096 0 1.65e-16
c7282 3034 707 3.15e-16
c7283 3748 3747 1.334e-15
c7284 3635 3634 1.6e-16
c7285 2494 1981 4.97e-16
c7286 2172 2461 1.58e-16
c7287 657 3034 7.99e-16
c7288 2535 2582 3.92e-16
c7289 1622 1623 9.1e-16
c7290 1343 1571 1.58e-16
c7291 1327 1559 1.58e-16
c7292 642 1321 3.15e-16
c7293 595 3877 9.02e-16
c7294 2765 752 3.64e-16
c7295 3359 2849 1.58e-16
c7296 2172 767 4.48e-16
c7297 1796 1 9.28e-16
c7298 4777 4395 1.443e-15
c7299 2545 858 3.15e-16
c7300 1 210 5.62e-16
c7301 4742 4361 5.2e-16
c7302 1862 1 5.97e-15
c7303 872 870 5.88e-16
c7304 3253 782 3.15e-16
c7305 5459 0 1.5617e-14
c7306 5141 5131 1.98e-16
c7307 2784 2782 1.6e-16
c7308 64 556 1.88e-16
c7309 4101 1 7.71e-16
c7310 3886 3622 1.58e-16
c7311 4506 4518 2.32e-16
c7312 2464 812 1.58e-16
c7313 822 1162 1.58e-16
c7314 627 592 5.8e-16
c7315 1047 0 6.29e-16
c7316 537 107 1.88e-16
c7317 1690 1624 1.58e-16
c7318 27 450 1.88e-16
c7319 479 175 1.88e-16
c7320 4580 4559 1.88e-16
c7321 5100 5101 3.54e-16
c7322 3503 702 5.73e-16
c7323 2746 1 8.43e-16
c7324 909 1038 3.54e-16
c7325 1176 827 2.33e-16
c7326 4028 4035 7.81e-16
c7327 3876 4281 3.92e-16
c7328 4763 4761 2.03e-16
c7329 602 1331 3.15e-16
c7330 3436 3055 3.92e-16
c7331 3440 3441 1.6e-16
c7332 1931 1 1.868e-15
c7333 175 189 1.88e-16
c7334 2296 2293 3.01e-16
c7335 2292 2289 6.44e-16
c7336 1921 0 2.93e-15
c7337 4759 236 5.8e-16
c7338 4022 4021 3.15e-16
c7339 3882 3486 1.58e-16
c7340 4519 842 7.38e-16
c7341 2851 2844 6.73e-16
c7342 687 692 2.77e-16
c7343 3882 4251 1.58e-16
c7344 3898 4263 1.58e-16
c7345 1971 827 1.339e-15
c7346 796 25 7.64e-16
c7347 1372 0 3.3846e-14
c7348 1178 1 4.59e-16
c7349 595 3876 1.511e-15
c7350 602 3898 4.46e-16
c7351 3429 1 5.97e-15
c7352 1175 0 1.0077e-14
c7353 3397 3407 3.92e-16
c7354 4563 4327 5.88e-16
c7355 4571 4333 1.58e-16
c7356 1208 858 1.58e-16
c7357 2840 2458 2.48e-16
c7358 1061 1517 4.36e-16
c7359 1515 1508 1.96e-16
c7360 3470 0 1.6491e-14
c7361 4063 1 6.66e-16
c7362 3650 3639 1.58e-16
c7363 2923 2880 2.15e-16
c7364 1783 1784 1.35e-16
c7365 3024 2577 5.5e-16
c7366 3034 3092 1.58e-16
c7367 1315 0 4.7664e-14
c7368 1548 1 6.15e-16
c7369 4599 1 8.43e-16
c7370 1694 1584 5.5e-16
c7371 193 187 5.8e-16
c7372 136 247 1.88e-16
c7373 3513 3506 1.96e-16
c7374 5452 439 7.37e-16
c7375 2375 1868 2.48e-16
c7376 1800 0 3.6368e-14
c7377 161 158 2.142e-15
c7378 281 273 1.58e-16
c7379 4324 662 1.09e-16
c7380 2670 2282 4.97e-16
c7381 921 647 3.15e-16
c7382 3898 3896 1.96e-16
c7383 3900 3890 5.5e-16
c7384 2674 0 1.4092e-14
c7385 1054 1055 7.51e-16
c7386 4514 4881 1.58e-16
c7387 2136 2117 1.58e-16
c7388 910 596 2.35e-16
c7389 4386 3548 4.97e-16
c7390 632 1414 1.58e-16
c7391 3888 0 5.86e-16
c7392 3411 777 3.58e-16
c7393 4661 4658 6.67e-16
c7394 1567 1539 2.64e-16
c7395 4537 4546 1.37e-16
c7396 5022 3839 3.54e-16
c7397 5009 4910 8.64e-16
c7398 911 3029 1.58e-16
c7399 421 426 1.88e-16
c7400 4753 4367 1.179e-15
c7401 4844 4850 5.87e-16
c7402 2542 2538 2.074e-15
c7403 2540 2536 1.988e-15
c7404 1042 1023 1.546e-15
c7405 3736 3729 8.3e-16
c7406 4103 4100 1.58e-16
c7407 1786 662 1.58e-16
c7408 5538 5535 5.88e-16
c7409 3243 0 1.6491e-14
c7410 1527 752 5.03e-16
c7411 1312 1306 8.89e-16
c7412 3079 0 6.72e-16
c7413 922 1160 3.92e-16
c7414 751 25 7.64e-16
c7415 537 1 3.4063e-14
c7416 4463 4458 1.642e-15
c7417 4265 4643 7.84e-16
c7418 3155 2645 1.58e-16
c7419 2718 707 1.58e-16
c7420 3046 2719 1.58e-16
c7421 1 150 4.92e-16
c7422 3219 3574 1.58e-16
c7423 3202 3591 2.386e-15
c7424 3600 3594 1.6e-16
c7425 2461 0 3.3692e-14
c7426 752 742 6.38e-16
c7427 3387 722 4.48e-16
c7428 4827 323 1.88e-16
c7429 2446 1930 4.11e-16
c7430 1291 1226 1.96e-16
c7431 5557 5556 1.08e-15
c7432 3829 3828 1.6e-16
c7433 3565 722 3.15e-16
c7434 5388 5356 1.58e-16
c7435 2559 822 3.58e-16
c7436 687 3393 4.03e-16
c7437 506 509 2.142e-15
c7438 140 129 2.45e-16
c7439 3612 0 6.72e-16
c7440 3431 1 9.28e-16
c7441 2196 868 3.58e-16
c7442 4006 1 7.08e-16
c7443 4462 4453 3.46e-16
c7444 767 0 2.8002e-13
c7445 1556 1557 1.35e-16
c7446 1684 1706 4.078e-15
c7447 1708 1690 4.312e-15
c7448 2713 3194 1.58e-16
c7449 617 1765 1.58e-16
c7450 3594 3593 1.6e-16
c7451 4566 1 2.56e-15
c7452 3124 662 1.339e-15
c7453 1706 1935 3.92e-16
c7454 44 49 1.88e-16
c7455 4572 0 5.86e-16
c7456 5036 5029 9.38e-16
c7457 2182 2180 5.93e-16
c7458 3803 3807 6.22e-16
c7459 632 2600 2.33e-16
c7460 285 1 2.87e-16
c7461 4298 647 7.38e-16
c7462 5324 5326 1.721e-15
c7463 4770 236 1.88e-16
c7464 2803 2435 1.96e-16
c7465 1854 732 1.58e-16
c7466 2136 2045 1.58e-16
c7467 2041 2044 1.887e-15
c7468 4205 3918 2.87e-16
c7469 4589 5535 6.5e-16
c7470 3402 0 6.35e-16
c7471 2933 2937 1.96e-16
c7472 2559 2807 1.58e-16
c7473 1598 797 1.09e-16
c7474 3882 3531 5.88e-16
c7475 3876 3537 1.58e-16
c7476 3616 4451 1.96e-16
c7477 2535 2248 5.5e-16
c7478 2545 2637 1.58e-16
c7479 934 0 1.1552e-14
c7480 2702 3209 3.92e-16
c7481 3214 3213 1.6e-16
c7482 3048 3041 3.54e-16
c7483 3030 3042 6.67e-16
c7484 2325 702 1.58e-16
c7485 1653 1644 3.92e-16
c7486 1191 1647 5.66e-16
c7487 1046 0 7.4292e-14
c7488 1281 1 4.17e-16
c7489 565 252 1.88e-16
c7490 3374 3048 1.96e-16
c7491 4923 1 4.69e-16
c7492 5157 0 3.6422e-14
c7493 3024 752 4.48e-16
c7494 216 1 2.946e-15
c7495 4827 5048 3.92e-16
c7496 230 37 5.71e-16
c7497 3397 852 7.99e-16
c7498 2282 0 6.9102e-14
c7499 2172 2196 4.383e-15
c7500 1321 732 3.15e-16
c7501 1398 966 1.96e-16
c7502 1399 1392 6.73e-16
c7503 4483 797 4.81e-16
c7504 1321 1623 3.92e-16
c7505 706 25 7.64e-16
c7506 4353 0 3.3724e-14
c7507 602 1706 4.46e-16
c7508 595 1684 1.511e-15
c7509 574 580 1.58e-16
c7510 4717 1 6.42e-16
c7511 4816 4813 5.5e-16
c7512 2161 1652 3.38e-16
c7513 15 291 5.8e-16
c7514 1 297 5.62e-16
c7515 2512 2196 3.25e-16
c7516 677 672 2.77e-16
c7517 895 898 5.05e-16
c7518 3918 3979 8.1e-16
c7519 4571 617 1.33e-16
c7520 4567 4639 3.92e-16
c7521 5546 526 1.58e-16
c7522 3003 1 6.636e-15
c7523 777 2418 2.22e-16
c7524 2194 1811 5.5e-16
c7525 5360 294 3.54e-16
c7526 2342 2354 2.32e-16
c7527 627 2594 3.79e-16
c7528 2708 2715 6.73e-16
c7529 4267 3435 2.48e-16
c7530 2469 852 1.58e-16
c7531 2486 827 1.58e-16
c7532 2299 677 3.15e-16
c7533 2908 2907 1.6e-16
c7534 3918 1 4.7861e-14
c7535 3288 2764 4.36e-16
c7536 3279 3286 1.96e-16
c7537 3046 3173 3.92e-16
c7538 762 752 3.28e-16
c7539 3649 3640 3.46e-16
c7540 3192 2679 1.532e-15
c7541 612 1735 1.58e-16
c7542 601 1721 1.84e-16
c7543 3185 3573 4.97e-16
c7544 4529 1 6.15e-16
c7545 2247 1 8.43e-16
c7546 19 549 8.4e-16
c7547 479 436 1.88e-16
c7548 310 508 1.88e-16
c7549 4567 4621 1.58e-16
c7550 4580 3874 5.5e-16
c7551 4582 4231 1.58e-16
c7552 883 752 6.45e-16
c7553 909 1112 4.35e-16
c7554 907 1111 1.88e-16
c7555 890 1104 1.58e-16
c7556 3397 3293 1.58e-16
c7557 2613 1 9.28e-16
c7558 1083 1084 1.21e-16
c7559 2785 2418 1.58e-16
c7560 1327 858 3.15e-16
c7561 1466 1460 1.6e-16
c7562 1031 1440 1.58e-16
c7563 657 596 1.96e-16
c7564 3369 0 8e-16
c7565 3183 1 6.15e-16
c7566 2895 2893 3.92e-16
c7567 3599 4433 1.58e-16
c7568 2401 752 1.58e-16
c7569 3919 37 1.88e-16
c7570 1708 1482 5.5e-16
c7571 1011 1 4.044e-15
c7572 1441 0 6.62e-16
c7573 602 595 5.95e-16
c7574 3089 3472 7.84e-16
c7575 2332 1811 1.96e-16
c7576 2327 1817 1.96e-16
c7577 3409 3654 1.58e-16
c7578 1732 2239 2.48e-16
c7579 1068 732 1.05e-15
c7580 4702 323 1.364e-15
c7581 113 71 9.5e-16
c7582 3882 852 4.03e-16
c7583 1345 692 3.15e-16
c7584 4338 3497 4.11e-16
c7585 5417 5511 7.46e-16
c7586 1321 1588 1.58e-16
c7587 1343 1576 1.58e-16
c7588 1211 1207 3.78e-16
c7589 1546 1544 1.6e-16
c7590 1541 1540 2.03e-16
c7591 3760 1 2.94e-16
c7592 3387 3089 1.58e-16
c7593 5103 62 5.5e-16
c7594 4037 4038 3.15e-16
c7595 1483 707 7.68e-16
c7596 1203 909 3.54e-16
c7597 392 49 1.88e-16
c7598 3900 702 3.58e-16
c7599 595 3896 2.13e-16
c7600 2954 2969 1.739e-15
c7601 2459 837 1.58e-16
c7602 602 1360 1.09e-16
c7603 4107 25 4.68e-16
c7604 3257 3258 9.1e-16
c7605 3046 3138 1.58e-16
c7606 3030 3126 1.58e-16
c7607 5220 5219 1.6e-16
c7608 792 1131 4e-16
c7609 552 545 3.54e-16
c7610 553 555 6.67e-16
c7611 479 349 1.88e-16
c7612 508 339 1.88e-16
c7613 3543 3540 5.5e-16
c7614 2175 1 8.766e-15
c7615 4827 265 1.88e-16
c7616 2391 1885 3.92e-16
c7617 2395 2396 1.6e-16
c7618 2196 2270 3.92e-16
c7619 5284 323 1.58e-16
c7620 3397 3409 4.369e-15
c7621 4362 702 2.65e-16
c7622 4133 4134 3.15e-16
c7623 4408 4407 5.65e-16
c7624 4402 3565 1.532e-15
c7625 4692 4316 3.92e-16
c7626 4704 4703 1.6e-16
c7627 601 1331 3.15e-16
c7628 1550 1 5.97e-15
c7629 2206 2218 2.32e-16
c7630 792 1920 1.58e-16
c7631 3411 3608 1.58e-16
c7632 3397 3621 4.63e-16
c7633 4708 410 1.88e-16
c7634 2553 1 1.002e-15
c7635 1073 707 3.57e-16
c7636 1053 1066 1.58e-16
c7637 596 790 2.45e-16
c7638 4657 439 1.88e-16
c7639 4056 4004 1.88e-16
c7640 3886 837 7.99e-16
c7641 4640 5461 1.96e-16
c7642 1091 767 1.58e-16
c7643 3898 4268 1.58e-16
c7644 3876 4280 1.58e-16
c7645 1988 868 1.58e-16
c7646 602 960 6.48e-16
c7647 612 954 2e-16
c7648 818 0 1.1363e-14
c7649 3387 822 3.15e-16
c7650 910 1315 1.58e-16
c7651 3073 2566 3.92e-16
c7652 3077 3078 1.6e-16
c7653 1392 0 1.4092e-14
c7654 601 3898 4.46e-16
c7655 4296 1 1.056e-15
c7656 1869 1880 1.96e-16
c7657 758 757 1.96e-16
c7658 3350 3351 5.65e-16
c7659 529 528 3.84e-16
c7660 2196 0 3.46872e-13
c7661 4563 4344 5.88e-16
c7662 4571 4350 1.58e-16
c7663 4810 33 1.88e-16
c7664 2487 1970 1.96e-16
c7665 2488 2481 6.73e-16
c7666 5584 5575 7.53e-16
c7667 3919 3921 1.06e-16
c7668 4872 91 1.88e-16
c7669 1031 1027 3.78e-16
c7670 920 1039 1.58e-16
c7671 618 0 7.86e-15
c7672 4219 4221 7.1e-16
c7673 4496 4489 1.96e-16
c7674 3650 4498 4.36e-16
c7675 3346 2832 4.97e-16
c7676 4616 1 8.43e-16
c7677 4361 4745 1.36e-15
c7678 4754 4748 1.6e-16
c7679 100 114 3.84e-16
c7680 602 26 7.12e-16
c7681 0 483 1.5723e-14
c7682 3910 3909 1.58e-16
c7683 91 0 1.2186e-13
c7684 146 368 1.88e-16
c7685 4347 677 4.81e-16
c7686 366 368 1.257e-15
c7687 2578 2169 1.96e-16
c7688 2579 2572 6.73e-16
c7689 3731 3728 3.54e-16
c7690 1629 837 2.72e-16
c7691 1420 1421 1.35e-16
c7692 1176 1179 1.58e-16
c7693 2541 2700 1.58e-16
c7694 4039 37 1.88e-16
c7695 4040 26 1.075e-15
c7696 3588 1 4.41e-15
c7697 3150 3143 1.96e-16
c7698 33 180 1.88e-16
c7699 4422 0 6.62e-16
c7700 3151 662 1.58e-16
c7701 4950 4923 1.37e-16
c7702 2269 1760 1.58e-16
c7703 165 247 1.88e-16
c7704 4861 4864 6.02e-16
c7705 2542 2540 8.67e-16
c7706 1062 692 4.98e-16
c7707 596 745 2.45e-16
c7708 79 71 2.218e-15
c7709 72 88 3.84e-16
c7710 2194 2389 3.92e-16
c7711 1091 1095 2.03e-16
c7712 3667 837 1.813e-15
c7713 4736 5262 1.96e-16
c7714 2831 2822 3.46e-16
c7715 1690 852 4.03e-16
c7716 2559 2475 1.58e-16
c7717 919 1174 1.58e-16
c7718 773 0 1.1445e-14
c7719 1708 1786 1.58e-16
c7720 4574 4566 1.6e-16
c7721 1488 0 3.6368e-14
c7722 1707 1 2.471e-15
c7723 276 49 1.88e-16
c7724 3393 3570 1.96e-16
c7725 2481 0 1.4092e-14
c7726 923 918 1.88e-16
c7727 3676 827 1.58e-16
c7728 2194 2191 1.58e-16
c7729 2172 2192 3.92e-16
c7730 5449 5451 9.16e-16
c7731 2923 2503 1.19e-16
c7732 919 807 3.15e-16
c7733 1708 702 3.58e-16
c7734 3444 1 6.15e-16
c7735 2646 2640 1.6e-16
c7736 2248 2637 2.386e-15
c7737 1504 1503 9.1e-16
c7738 537 310 1.88e-16
c7739 2316 717 1.813e-15
c7740 1211 1343 3.92e-16
c7741 1134 0 2.7186e-14
c7742 4201 37 3.84e-16
c7743 2407 782 2.33e-16
c7744 2178 702 4.03e-16
c7745 4851 4849 1.6e-16
c7746 641 640 6.67e-16
c7747 2040 2025 3.25e-16
c7748 2023 2026 6.71e-16
c7749 1 255 1.44e-16
c7750 3304 837 1.813e-15
c7751 4674 4675 9.93e-16
c7752 5410 439 1.58e-16
c7753 2271 0 3.6368e-14
c7754 2371 2359 2.32e-16
c7755 996 672 5.73e-16
c7756 1432 647 3.64e-16
c7757 1130 752 1.58e-16
c7758 4821 410 1.88e-16
c7759 2816 2424 1.96e-16
c7760 2254 2635 3.92e-16
c7761 2640 2639 1.6e-16
c7762 1874 732 1.58e-16
c7763 632 1389 1.58e-16
c7764 3401 0 8.1192e-14
c7765 3228 1 5.808e-15
c7766 2182 702 7.99e-16
c7767 1762 1761 1.6e-16
c7768 1196 1644 1.58e-16
c7769 931 0 3.7358e-14
c7770 1706 1934 1.58e-16
c7771 1690 1922 1.58e-16
c7772 303 346 1.88e-16
c7773 320 368 1.88e-16
c7774 3504 3117 1.532e-15
c7775 1845 2362 2.38e-15
c7776 2049 1 8.09e-16
c7777 1749 2255 3.92e-16
c7778 2260 2259 1.6e-16
c7779 890 977 1.96e-16
c7780 422 1 1.65e-15
c7781 227 216 2.45e-16
c7782 401 0 6.224e-15
c7783 407 19 3.84e-16
c7784 4719 33 1.88e-16
c7785 657 3470 1.58e-16
c7786 4070 4079 1.88e-16
c7787 2915 2917 6.87e-16
c7788 2940 2913 5.87e-16
c7789 1521 722 1.58e-16
c7790 4380 4373 6.73e-16
c7791 4379 3537 1.96e-16
c7792 4702 5324 3.54e-16
c7793 1694 837 7.99e-16
c7794 1345 1640 3.92e-16
c7795 2725 2722 5.5e-16
c7796 728 0 1.1593e-14
c7797 3600 1 1.868e-15
c7798 1331 1470 4.63e-16
c7799 1243 1 2.295e-15
c7800 4628 4248 1.96e-16
c7801 2773 782 1.58e-16
c7802 1694 1319 5.5e-16
c7803 4189 1 6.78e-16
c7804 4373 0 1.4092e-14
c7805 2688 692 1.832e-15
c7806 4889 4497 7.17e-16
c7807 4909 4897 1.74e-16
c7808 601 1706 4.46e-16
c7809 713 712 1.96e-16
c7810 367 366 2.84e-16
c7811 4734 1 6.42e-16
c7812 1824 0 6.72e-16
c7813 4 5 1.482e-15
c7814 3393 3506 1.58e-16
c7815 3659 3661 2.15e-16
c7816 3668 3669 1.6e-16
c7817 27 26 8.41e-16
c7818 3676 812 1.832e-15
c7819 3983 3974 1.88e-16
c7820 3027 1 8.766e-15
c7821 4567 4656 3.92e-16
c7822 5380 1 3.36e-16
c7823 4896 64 2.402e-15
c7824 2172 1828 5.5e-16
c7825 5514 5491 1.58e-16
c7826 1321 1011 1.58e-16
c7827 3376 1 1.052e-15
c7828 537 339 1.88e-16
c7829 4166 1 7.08e-16
c7830 3882 3690 1.58e-16
c7831 4150 37 1.88e-16
c7832 4159 25 4.68e-16
c7833 3997 1 6.78e-16
c7834 3024 3190 3.92e-16
c7835 4813 4820 1.96e-16
c7836 2104 2106 5.88e-16
c7837 2146 1249 1.33e-16
c7838 4715 4713 1.6e-16
c7839 627 1735 1.58e-16
c7840 307 308 6.67e-16
c7841 4567 4638 1.58e-16
c7842 4580 4242 5.5e-16
c7843 4582 4248 1.58e-16
c7844 2419 2413 1.6e-16
c7845 1896 2410 2.386e-15
c7846 1902 2418 1.136e-15
c7847 5363 0 2.078e-15
c7848 42 19 3.84e-16
c7849 392 194 1.88e-16
c7850 3373 3807 3.65e-16
c7851 2987 3847 1.389e-15
c7852 3866 3344 1.96e-16
c7853 4872 5106 1.984e-15
c7854 2707 2316 4.11e-16
c7855 2791 0 6.62e-16
c7856 5324 5284 5.69e-16
c7857 2231 2619 4.97e-16
c7858 3192 1 1.716e-15
c7859 3599 4438 2.386e-15
c7860 4447 4441 1.6e-16
c7861 3286 3277 3.46e-16
c7862 687 1823 1.58e-16
c7863 3937 19 3.84e-16
c7864 2844 842 1.84e-16
c7865 1466 1 1.868e-15
c7866 1456 0 2.93e-15
c7867 3100 3484 1.58e-16
c7868 601 595 2.77e-16
c7869 570 571 6.96e-16
c7870 5135 31 3.54e-16
c7871 5106 0 3.8894e-14
c7872 2787 797 2.33e-16
c7873 1988 0 1.6491e-14
c7874 3409 3659 1.58e-16
c7875 1096 1097 1.238e-15
c7876 5476 410 3.54e-16
c7877 5521 1 3.36e-16
c7878 687 3034 7.99e-16
c7879 1379 1370 3.46e-16
c7880 59 223 1.88e-16
c7881 676 1 4.03e-16
c7882 2594 3104 1.58e-16
c7883 4604 4592 2.62e-16
c7884 1914 1905 3.92e-16
c7885 1522 1908 5.66e-16
c7886 1690 1701 1.96e-16
c7887 4527 4525 1.6e-16
c7888 4864 4486 7.84e-16
c7889 5232 178 7.46e-16
c7890 3281 797 5.03e-16
c7891 3411 3106 1.58e-16
c7892 4794 4412 1.443e-15
c7893 2399 1 6.15e-16
c7894 2163 2078 4.06e-16
c7895 4776 4401 4.9e-16
c7896 4725 468 1.88e-16
c7897 2498 2495 5.5e-16
c7898 5308 1 7.49e-16
c7899 3950 3947 5.5e-16
c7900 3918 3934 6.32e-16
c7901 1046 707 3.15e-16
c7902 1493 717 2.72e-16
c7903 1056 1059 1.58e-16
c7904 1539 782 1.75e-16
c7905 687 1026 4e-16
c7906 3886 3650 5.5e-16
c7907 3024 3155 1.58e-16
c7908 3046 3143 1.58e-16
c7909 657 2282 2.22e-16
c7910 470 471 3.84e-16
c7911 4759 4767 1.81e-16
c7912 1995 1992 3.01e-16
c7913 1991 1988 6.44e-16
c7914 1597 0 6.72e-16
c7915 777 1136 4.21e-16
c7916 311 303 2.218e-15
c7917 316 320 1.58e-16
c7918 5139 5137 3.92e-16
c7919 2192 0 1.2366e-14
c7920 4244 4237 6.73e-16
c7921 4243 3384 1.96e-16
c7922 3531 702 3.79e-16
c7923 4353 707 1.58e-16
c7924 5136 149 1.96e-16
c7925 2589 2586 5.5e-16
c7926 1822 692 5.03e-16
c7927 1181 868 1.813e-15
c7928 1439 1440 2.48e-16
c7929 3882 4468 1.96e-16
c7930 101 99 2.84e-16
c7931 847 1 5.62e-16
c7932 692 19 1.676e-15
c7933 4108 25 1.88e-16
c7934 3915 1 4.64e-16
c7935 4104 19 7.35e-16
c7936 3886 3480 5.5e-16
c7937 2378 752 5.03e-16
c7938 4780 4778 2.03e-16
c7939 617 1331 3.15e-16
c7940 5103 5113 2.114e-15
c7941 910 2196 5.03e-16
c7942 3453 3066 1.532e-15
c7943 3459 3458 5.65e-16
c7944 2304 1794 1.96e-16
c7945 3693 868 1.58e-16
c7946 5160 5221 1.6e-16
c7947 602 3424 1.58e-16
c7948 1121 752 3.57e-16
c7949 3876 4285 1.58e-16
c7950 3900 4297 5.42e-16
c7951 4514 5575 1.477e-15
c7952 2865 2858 1.96e-16
c7953 2557 2554 1.58e-16
c7954 2535 2555 3.92e-16
c7955 1199 1 3.06e-16
c7956 617 3898 4.46e-16
c7957 3034 3309 4.63e-16
c7958 3046 662 4.46e-16
c7959 2112 178 9.36e-16
c7960 1919 1920 1.35e-16
c7961 1752 0 3.3874e-14
c7962 3397 3055 1.58e-16
c7963 3393 782 3.15e-16
c7964 4623 4248 4.9e-16
c7965 5204 5188 7.38e-16
c7966 3123 0 3.6368e-14
c7967 4424 767 1.84e-16
c7968 5479 5483 5.6e-16
c7969 5493 5452 3.18e-16
c7970 921 868 3.15e-16
c7971 920 827 3.69e-16
c7972 1907 767 5.03e-16
c7973 1535 1534 1.6e-16
c7974 1527 1525 2.15e-16
c7975 1345 1368 3.92e-16
c7976 2533 3074 4.97e-16
c7977 3030 2764 5.88e-16
c7978 4633 1 8.43e-16
c7979 4378 4745 1.58e-16
c7980 3393 3394 1.239e-15
c7981 2541 837 4.03e-16
c7982 276 194 1.88e-16
c7983 601 26 7.12e-16
c7984 3525 3523 2.15e-16
c7985 3533 3532 1.6e-16
c7986 5271 1 3.36e-16
c7987 1828 0 6.9481e-14
c7988 3883 3902 9.83e-16
c7989 5240 0 2.9101e-14
c7990 2557 2350 5.5e-16
c7991 3882 4433 1.58e-16
c7992 2770 0 3.5142e-14
c7993 2899 1 1.031e-15
c7994 4054 19 7.04e-16
c7995 2557 2717 1.58e-16
c7996 2541 2705 1.58e-16
c7997 1022 0 1.0003e-14
c7998 802 1 5.62e-16
c7999 1684 1986 3.92e-16
c8000 4447 1 1.868e-15
c8001 4595 0 1.4233e-14
c8002 4678 4675 6.67e-16
c8003 2559 672 3.58e-16
c8004 1694 1799 4.63e-16
c8005 25 346 7.06e-16
c8006 3518 3519 9.1e-16
c8007 2376 2388 2.32e-16
c8008 4437 0 2.93e-15
c8009 3526 692 1.84e-16
c8010 4905 4902 7.84e-16
c8011 2277 2283 1.6e-16
c8012 2274 1760 2.386e-15
c8013 907 662 4.8e-16
c8014 3397 3591 1.58e-16
c8015 4563 1 2.966e-15
c8016 4804 468 1.88e-16
c8017 2166 2571 4.11e-16
c8018 2136 2144 3.422e-15
c8019 4129 4126 1.76e-16
c8020 1623 837 2.4e-16
c8021 3264 0 3.466e-15
c8022 1330 1332 3.84e-16
c8023 1101 1108 7.95e-16
c8024 4390 4387 5.5e-16
c8025 4487 827 1.339e-15
c8026 5573 5569 1.243e-15
c8027 5536 5422 2.24e-16
c8028 2837 2836 9.1e-16
c8029 2559 2299 5.5e-16
c8030 4282 4660 7.84e-16
c8031 2790 807 1.58e-16
c8032 3628 777 1.58e-16
c8033 2705 732 1.58e-16
c8034 1859 1856 3.01e-16
c8035 1855 1852 6.44e-16
c8036 2821 827 2.33e-16
c8037 4989 0 1.63e-15
c8038 3024 2730 5.5e-16
c8039 3034 3245 1.58e-16
c8040 2173 2177 1.988e-15
c8041 1 454 9.8e-16
c8042 4580 4486 1.58e-16
c8043 5278 5280 5.62e-16
c8044 5302 5301 1.6e-16
c8045 601 2586 1.832e-15
c8046 245 251 5.8e-16
c8047 448 19 3.84e-16
c8048 4810 526 1.88e-16
c8049 2468 2459 3.46e-16
c8050 2194 1681 1.58e-16
c8051 3801 3805 5.87e-16
c8052 4402 752 1.339e-15
c8053 4725 64 1.88e-16
c8054 920 812 3.69e-16
c8055 598 1 7.18e-16
c8056 3453 1 1.716e-15
c8057 3624 0 2.93e-15
c8058 612 920 3.15e-16
c8059 4474 4470 1.96e-16
c8060 2172 717 3.15e-16
c8061 1769 1778 3.92e-16
c8062 1397 1764 1.58e-16
c8063 1683 1 2.259e-15
c8064 1 164 9.8e-16
c8065 117 37 1.88e-16
c8066 3674 827 1.339e-15
c8067 822 2435 1.813e-15
c8068 3611 752 1.58e-16
c8069 2292 0 6.62e-16
c8070 3811 3739 3.54e-16
c8071 3806 3775 1.58e-16
c8072 894 807 8.34e-16
c8073 2657 1 2.054e-15
c8074 3327 3710 7.84e-16
c8075 4188 4195 7.81e-16
c8076 632 1409 1.58e-16
c8077 4606 5422 6.17e-16
c8078 642 3480 2.22e-16
c8079 4282 4283 1.35e-16
c8080 3900 3548 5.5e-16
c8081 2798 3322 4.36e-16
c8082 2196 707 3.15e-16
c8083 4004 37 1.88e-16
c8084 4015 0 1.981e-14
c8085 2730 762 1.813e-15
c8086 1674 1664 7.29e-16
c8087 1659 1661 2.861e-15
c8088 967 0 1.8851e-14
c8089 4546 4540 9.61e-16
c8090 1684 1951 1.58e-16
c8091 1706 1939 1.58e-16
c8092 3128 3124 1.96e-16
c8093 657 2196 3.58e-16
c8094 1938 1556 2.48e-16
c8095 762 1525 1.58e-16
c8096 5031 5048 1.443e-15
c8097 3504 677 1.339e-15
c8098 602 1678 1.58e-16
c8099 612 1681 5.73e-16
c8100 2660 1 6.15e-16
c8101 883 992 3.92e-16
c8102 890 991 1.88e-16
c8103 880 878 3.54e-16
c8104 4302 647 1.832e-15
c8105 5384 5383 1.08e-15
c8106 4844 5032 2.69e-16
c8107 2807 2435 1.58e-16
c8108 287 19 3.45e-16
c8109 3293 3679 5.66e-16
c8110 3685 3676 3.92e-16
c8111 5538 1 3.39e-15
c8112 1413 1406 1.96e-16
c8113 2172 2371 1.58e-16
c8114 2334 707 7.68e-16
c8115 592 1 1.1755e-14
c8116 4200 1 6.03e-16
c8117 2508 858 7.38e-16
c8118 3134 692 1.58e-16
c8119 617 1706 4.46e-16
c8120 623 622 1.96e-16
c8121 4833 4830 5.5e-16
c8122 3237 737 3.64e-16
c8123 687 2654 1.58e-16
c8124 2444 1 5.808e-15
c8125 747 1499 1.813e-15
c8126 632 3117 1.58e-16
c8127 4567 4673 3.92e-16
c8128 2446 0 3.466e-15
c8129 902 891 2.933e-15
c8130 792 25 1.58e-16
c8131 3798 3785 3.92e-16
c8132 3996 4003 7.81e-16
c8133 3029 1 6.056e-15
c8134 792 1919 1.58e-16
c8135 1061 732 1.813e-15
c8136 3044 0 1.2366e-14
c8137 2545 2452 5.5e-16
c8138 2722 2729 1.96e-16
c8139 2662 2271 1.136e-15
c8140 1016 1015 3.94e-16
c8141 4284 3446 4.97e-16
c8142 1345 1026 1.58e-16
c8143 1331 1469 1.58e-16
c8144 3396 1 2.56e-15
c8145 3707 3898 1.58e-16
c8146 1987 868 1.58e-16
c8147 617 966 2.33e-16
c8148 617 4281 1.58e-16
c8149 3296 3298 2.15e-16
c8150 3048 3207 3.92e-16
c8151 3661 3657 1.96e-16
c8152 3230 737 1.9e-16
c8153 4711 0 3.485e-14
c8154 2009 1618 4.11e-16
c8155 627 1755 1.58e-16
c8156 1181 0 7.4292e-14
c8157 19 274 3.84e-16
c8158 3409 702 3.15e-16
c8159 4567 4655 1.58e-16
c8160 4580 4259 5.5e-16
c8161 4582 4265 1.58e-16
c8162 5152 5157 1.81e-15
c8163 3287 2770 1.136e-15
c8164 1178 837 1.58e-16
c8165 894 1126 1.58e-16
c8166 907 1098 3.54e-16
c8167 4268 4280 2.32e-16
c8168 5388 5365 1.58e-16
c8169 107 218 1.88e-16
c8170 4589 1 4.744e-15
c8171 687 596 1.96e-16
c8172 3976 1 5.1e-16
c8173 1879 767 1.58e-16
c8174 1708 1369 1.58e-16
c8175 3693 0 3.3874e-14
c8176 627 1733 1.58e-16
c8177 1031 1 5.821e-15
c8178 3100 3489 2.386e-15
c8179 3498 3492 1.6e-16
c8180 3876 762 3.15e-16
c8181 747 1506 1.58e-16
c8182 193 194 3.84e-16
c8183 5036 5035 5.87e-16
c8184 4915 4902 1.58e-16
c8185 2344 1828 4.11e-16
c8186 5120 122 5.93e-16
c8187 14 12 1.58e-16
c8188 5324 5340 1.23e-16
c8189 1104 737 8.3e-16
c8190 5253 5240 3.92e-16
c8191 4719 526 1.88e-16
c8192 617 3468 1.58e-16
c8193 2172 1987 1.58e-16
c8194 2178 1981 5.88e-16
c8195 4360 4351 3.46e-16
c8196 4804 64 1.88e-16
c8197 1327 1146 1.58e-16
c8198 4336 1 5.808e-15
c8199 4338 0 3.466e-15
c8200 921 0 3.20067e-13
c8201 3475 647 1.84e-16
c8202 4862 1 1.806e-15
c8203 3364 3372 2.15e-16
c8204 3301 797 1.09e-16
c8205 910 2192 1.58e-16
c8206 9 509 4.88e-16
c8207 5253 5254 1.6e-16
c8208 2182 1981 5.5e-16
c8209 88 89 7.03e-16
c8210 4006 857 1.88e-16
c8211 4895 64 8.9e-16
c8212 52 1 1.44e-16
c8213 3958 3951 2.45e-16
c8214 5514 5471 3.1e-16
c8215 5526 5522 1.243e-15
c8216 642 983 1.58e-16
c8217 2700 2701 9.1e-16
c8218 1948 782 3.64e-16
c8219 1551 1542 3.92e-16
c8220 1101 1545 5.66e-16
c8221 1106 1537 1.58e-16
c8222 3157 0 3.6368e-14
c8223 4590 4592 1.687e-15
c8224 4602 4595 6.73e-16
c8225 4601 3873 1.96e-16
c8226 4157 1 6.78e-16
c8227 1072 1 3.54e-16
c8228 4862 4873 1.96e-16
c8229 1069 0 9.602e-15
c8230 3409 3485 3.92e-16
c8231 3393 3134 5.88e-16
c8232 4776 4781 5.53e-16
c8233 3411 647 3.15e-16
c8234 3387 672 3.15e-16
c8235 4691 352 5.8e-16
c8236 5288 412 1.345e-15
c8237 910 2531 1.58e-16
c8238 3857 3855 1.96e-16
c8239 1162 797 1.58e-16
c8240 1143 1149 1.58e-16
c8241 78 508 1.88e-16
c8242 3385 3384 1.58e-16
c8243 4373 707 1.58e-16
c8244 5388 5299 1.58e-16
c8245 5303 5300 4.41e-16
c8246 601 594 1.74e-16
c8247 1842 692 1.09e-16
c8248 1647 858 1.84e-16
c8249 3898 4485 3.92e-16
c8250 4118 37 1.88e-16
c8251 4127 25 4.68e-16
c8252 4420 4421 2.48e-16
c8253 717 0 2.86312e-13
c8254 5588 4520 1.96e-16
c8255 2535 2769 3.92e-16
c8256 1632 1629 3.01e-16
c8257 1628 1625 6.44e-16
c8258 1962 1 6.15e-16
c8259 3409 3869 4.22e-16
c8260 3030 827 3.15e-16
c8261 2226 2223 5.5e-16
c8262 3387 3242 1.58e-16
c8263 612 3438 1.58e-16
c8264 601 3424 1.84e-16
c8265 4634 5459 7.87e-16
c8266 2557 2169 1.58e-16
c8267 1618 842 3.15e-16
c8268 2009 868 2.72e-16
c8269 1331 1106 5.5e-16
c8270 3090 2577 1.532e-15
c8271 3096 3095 5.65e-16
c8272 4300 1 1.716e-15
c8273 1895 1499 1.96e-16
c8274 1890 1505 1.96e-16
c8275 747 920 3.15e-16
c8276 4915 323 1.88e-16
c8277 3275 782 7.38e-16
c8278 1 218 2.1108e-14
c8279 15 193 6.58e-16
c8280 3381 3872 4.65e-16
c8281 4567 4745 1.58e-16
c8282 4571 4361 5.5e-16
c8283 1364 1358 1.6e-16
c8284 876 866 7.23e-16
c8285 5517 381 3.54e-16
c8286 3497 4302 1.58e-16
c8287 595 1322 9.02e-16
c8288 3728 1 1.23e-16
c8289 4508 4506 2.15e-16
c8290 4516 4515 1.6e-16
c8291 3046 2781 5.5e-16
c8292 1810 1414 1.96e-16
c8293 4097 0 9.4096e-14
c8294 1750 0 1.6491e-14
c8295 4650 1 8.43e-16
c8296 4395 4745 2e-16
c8297 4378 4762 1.36e-15
c8298 4771 4765 1.6e-16
c8299 3409 3421 1.58e-16
c8300 2668 702 1.58e-16
c8301 2082 2029 2.45e-16
c8302 1635 2007 1.58e-16
c8303 617 26 7.12e-16
c8304 26 433 1.03e-15
c8305 5151 236 7.38e-16
c8306 5112 5072 1.062e-15
c8307 866 867 6.67e-16
c8308 692 683 1.078e-15
c8309 890 827 3.15e-16
c8310 922 702 3.15e-16
c8311 957 954 1.791e-15
c8312 2535 2367 5.5e-16
c8313 2170 2166 1.58e-16
c8314 1816 677 7.38e-16
c8315 1625 842 1.339e-15
c8316 3882 4438 1.58e-16
c8317 3898 4450 1.58e-16
c8318 4501 4502 9.1e-16
c8319 2535 2734 1.58e-16
c8320 2557 2722 1.58e-16
c8321 2372 722 1.58e-16
c8322 1701 1693 1.606e-15
c8323 1708 2003 3.92e-16
c8324 4612 0 1.4233e-14
c8325 1954 1573 3.92e-16
c8326 1958 1959 1.6e-16
c8327 5096 5095 1.6e-16
c8328 4436 792 1.58e-16
c8329 3442 3440 1.6e-16
c8330 3437 3436 2.03e-16
c8331 5396 265 7.16e-16
c8332 3360 842 1.58e-16
c8333 3030 812 3.15e-16
c8334 762 1684 3.15e-16
c8335 777 1918 2.4e-16
c8336 2754 2373 3.92e-16
c8337 2707 0 3.466e-15
c8338 3321 3706 1.96e-16
c8339 1812 662 3.64e-16
c8340 3284 0 8e-16
c8341 2594 1 5.97e-15
c8342 612 3030 4.03e-16
c8343 595 3048 3.15e-16
c8344 602 3024 3.46e-16
c8345 1328 1347 9.83e-16
c8346 3886 3385 5.5e-16
c8347 4504 868 1.58e-16
c8348 2843 2839 1.96e-16
c8349 1851 732 1.58e-16
c8350 1249 1262 3.18e-16
c8351 794 0 7.709e-15
c8352 3155 3156 9.1e-16
c8353 1375 1 2.054e-15
c8354 2725 732 1.58e-16
c8355 1635 1176 1.136e-15
c8356 1377 0 8e-16
c8357 262 252 3.75e-16
c8358 2838 868 1.58e-16
c8359 2272 1760 1.532e-15
c8360 3048 2747 5.5e-16
c8361 1516 0 6.9481e-14
c8362 2179 2177 8.67e-16
c8363 4580 4503 1.58e-16
c8364 4878 4879 7.52e-16
c8365 617 2586 1.58e-16
c8366 1987 0 3.6368e-14
c8367 4838 352 1.88e-16
c8368 2474 2473 9.1e-16
c8369 2172 2405 1.58e-16
c8370 2194 2393 1.58e-16
c8371 2172 1715 1.58e-16
c8372 2178 1682 5.5e-16
c8373 4770 5205 5.91e-16
c8374 3006 2492 8.31e-16
c8375 3017 2503 1.58e-16
c8376 4306 4305 5.65e-16
c8377 4300 3463 1.532e-15
c8378 3479 1 8.43e-16
c8379 4215 3879 1.159e-15
c8380 1901 752 7.38e-16
c8381 1345 1348 1.6e-16
c8382 3623 792 1.58e-16
c8383 807 1 4.1542e-14
c8384 2703 732 1.58e-16
c8385 1148 0 1.4198e-14
c8386 627 920 3.15e-16
c8387 1769 1397 1.58e-16
c8388 1729 1 1.056e-15
c8389 2713 2719 1.418e-15
c8390 2559 797 3.15e-16
c8391 2730 2702 2.64e-16
c8392 2045 2056 3.92e-16
c8393 1 354 4.848e-15
c8394 3691 868 1.58e-16
c8395 3370 2855 1.958e-15
c8396 2196 1879 5.5e-16
c8397 2317 1 1.868e-15
c8398 2307 0 2.93e-15
c8399 0 369 1.0822e-14
c8400 2182 1682 5.5e-16
c8401 890 812 3.15e-16
c8402 907 1172 3.92e-16
c8403 842 868 3.28e-16
c8404 920 993 1.58e-16
c8405 3900 3903 1.6e-16
c8406 5358 5379 1.96e-16
c8407 612 890 3.35e-16
c8408 595 909 3.15e-16
c8409 602 883 3.03e-16
c8410 1767 1778 1.96e-16
c8411 2545 2288 1.58e-16
c8412 4361 4724 1.96e-16
c8413 3228 3227 2.48e-16
c8414 3165 677 1.09e-16
c8415 3034 3071 4.63e-16
c8416 1800 1801 1.35e-16
c8417 632 1769 1.832e-15
c8418 1523 0 1.6491e-14
c8419 5039 5026 1.96e-16
c8420 1862 1851 1.58e-16
c8421 3034 782 3.15e-16
c8422 612 2232 2.65e-16
c8423 601 1678 1.58e-16
c8424 910 3044 1.58e-16
c8425 2827 2435 2.38e-15
c8426 883 1006 1.88e-16
c8427 907 999 1.58e-16
c8428 596 933 2.397e-15
c8429 3733 3729 5.6e-16
c8430 3252 1 8.43e-16
c8431 2949 2959 8.28e-16
c8432 4028 3918 2.87e-16
c8433 1300 1218 5.88e-16
c8434 1828 707 3.15e-16
c8435 2344 717 2.72e-16
c8436 1661 1660 2.49e-16
c8437 749 0 7.709e-15
c8438 506 9 5.8e-16
c8439 3618 1 9.28e-16
c8440 1575 1131 2.48e-16
c8441 4645 4265 1.96e-16
c8442 687 1800 1.58e-16
c8443 3554 0 3.6368e-14
c8444 2172 842 4.48e-16
c8445 4546 3718 1.96e-16
c8446 3332 837 2.72e-16
c8447 1471 1 4.41e-15
c8448 1855 0 6.62e-16
c8449 3409 3151 5.5e-16
c8450 3685 3674 1.96e-16
c8451 2730 722 1.58e-16
c8452 687 2674 1.58e-16
c8453 2464 1 2.054e-15
c8454 1052 677 1.58e-16
c8455 1 130 1.073e-15
c8456 4567 4690 3.92e-16
c8457 5051 5049 4e-16
c8458 2466 0 8e-16
c8459 5530 5529 1.03e-16
c8460 4827 381 1.88e-16
c8461 1511 737 1.84e-16
c8462 1965 807 2.65e-16
c8463 1321 1031 5.5e-16
c8464 1331 1474 1.58e-16
c8465 529 526 4.6e-16
c8466 506 511 1.482e-15
c8467 146 143 3.54e-16
c8468 1981 852 1.58e-16
c8469 1998 827 1.58e-16
c8470 1818 1437 3.92e-16
c8471 1822 1823 1.6e-16
c8472 1122 0 6.29e-16
c8473 537 78 1.88e-16
c8474 4181 19 9.67e-16
c8475 4454 4456 2.03e-16
c8476 4830 4837 1.96e-16
c8477 4915 265 1.88e-16
c8478 1641 1706 1.58e-16
c8479 1879 1488 1.136e-15
c8480 4728 0 3.4813e-14
c8481 4732 4730 1.6e-16
c8482 0 43 1.5696e-14
c8483 28 34 1.059e-15
c8484 19 22 8.4e-16
c8485 27 49 1.88e-16
c8486 3589 3590 2.03e-16
c8487 4567 4672 1.58e-16
c8488 4580 4276 5.5e-16
c8489 4582 4282 1.58e-16
c8490 2818 1 1.056e-15
c8491 909 1113 3.54e-16
c8492 4390 732 1.58e-16
c8493 2729 2720 3.46e-16
c8494 4175 4167 9.33e-16
c8495 3751 3748 1.84e-16
c8496 3744 3747 1.887e-15
c8497 3380 0 2.0654e-14
c8498 910 921 1.58e-16
c8499 911 920 3.45e-16
c8500 4164 37 1.88e-16
c8501 3298 3294 1.96e-16
c8502 1913 752 1.58e-16
c8503 3989 19 9.67e-16
c8504 1646 1181 4.11e-16
c8505 4556 1 9.43e-16
c8506 4327 4714 2.196e-15
c8507 822 1151 1.813e-15
c8508 1502 1 1.056e-15
c8509 3900 777 3.58e-16
c8510 2007 1 5.808e-15
c8511 0 584 5.4938e-14
c8512 26 580 1.96e-16
c8513 5039 120 3.94e-16
c8514 2009 0 3.466e-15
c8515 226 1 1.44e-16
c8516 2265 1 5.97e-15
c8517 3708 3709 2.03e-16
c8518 4838 294 1.88e-16
c8519 2194 1998 5.5e-16
c8520 981 971 1.418e-15
c8521 1391 1387 1.96e-16
c8522 4736 5388 7.46e-16
c8523 3194 0 3.3874e-14
c8524 3960 19 7.35e-16
c8525 4366 4365 9.1e-16
c8526 1343 1161 1.58e-16
c8527 747 751 2.19e-16
c8528 704 0 7.709e-15
c8529 4356 1 2.054e-15
c8530 4358 0 8e-16
c8531 571 580 1.58e-16
c8532 4879 1 1.858e-15
c8533 4881 4503 1.527e-15
c8534 5010 33 1.88e-16
c8535 2987 2895 1.772e-15
c8536 2899 2896 1.84e-16
c8537 911 1681 1.88e-16
c8538 1008 1014 1.58e-16
c8539 1 302 4.59e-16
c8540 2714 2322 1.96e-16
c8541 2525 2512 3.92e-16
c8542 3876 722 4.48e-16
c8543 5514 381 6.06e-16
c8544 3010 1 1.106e-15
c8545 2789 2790 2.48e-16
c8546 1489 722 1.339e-15
c8547 2136 0 5.6075e-14
c8548 2557 2390 1.58e-16
c8549 1567 767 1.58e-16
c8550 4546 858 1.58e-16
c8551 687 1046 4.21e-16
c8552 1235 0 1.9454e-14
c8553 3690 4526 5.66e-16
c8554 4532 4523 3.92e-16
c8555 3030 2651 1.58e-16
c8556 1176 1 4.044e-15
c8557 3641 3643 2.03e-16
c8558 5036 180 1.345e-15
c8559 687 2282 1.813e-15
c8560 426 204 1.88e-16
c8561 1628 0 6.62e-16
c8562 5336 1 3.36e-16
c8563 722 716 1.74e-16
c8564 1715 0 3.5936e-14
c8565 2337 2338 9.1e-16
c8566 1162 1164 7.84e-16
c8567 59 305 1.88e-16
c8568 4258 4251 1.96e-16
c8569 3385 4260 4.36e-16
c8570 5388 5345 3.1e-16
c8571 4922 91 1.88e-16
c8572 1664 858 1.58e-16
c8573 3876 4502 3.92e-16
c8574 3938 1 4.738e-15
c8575 3886 4315 4.63e-16
c8576 3030 747 4.03e-16
c8577 4797 4795 2.03e-16
c8578 3919 0 2.0532e-14
c8579 3186 3177 3.92e-16
c8580 2668 3180 5.66e-16
c8581 2679 3172 1.58e-16
c8582 1607 1990 7.84e-16
c8583 1690 1867 1.96e-16
c8584 3471 3472 2.48e-16
c8585 4504 0 1.6491e-14
c8586 2208 0 3.466e-15
c8587 1971 1 1.716e-15
c8588 5072 1 1.021e-15
c8589 3046 852 3.15e-16
c8590 88 479 1.88e-16
c8591 5115 0 2.078e-15
c8592 3411 3259 1.58e-16
c8593 3781 852 1.58e-16
c8594 1085 732 1.85e-16
c8595 627 3438 1.58e-16
c8596 2838 0 3.5142e-14
c8597 396 395 2.84e-16
c8598 3898 3469 1.58e-16
c8599 4543 852 1.58e-16
c8600 4702 381 1.88e-16
c8601 1315 1318 1.576e-15
c8602 919 920 4.116e-15
c8603 3910 37 1.88e-16
c8604 3911 26 1.075e-15
c8605 3030 3342 1.58e-16
c8606 3168 2651 1.136e-15
c8607 2223 2230 1.96e-16
c8608 88 189 1.88e-16
c8609 596 817 3.134e-15
c8610 3397 3083 5.5e-16
c8611 2568 0 2.93e-15
c8612 2072 2095 1.96e-16
c8613 1 338 9.8e-16
c8614 9 303 5.8e-16
c8615 3387 797 4.48e-16
c8616 4166 857 1.88e-16
c8617 4567 4762 1.58e-16
c8618 4571 4378 5.5e-16
c8619 5098 62 3.54e-16
c8620 393 1 1.65e-15
c8621 386 0 2.87e-16
c8622 378 37 1.88e-16
c8623 3605 782 1.75e-16
c8624 1760 672 1.58e-16
c8625 2285 647 4.81e-16
c8626 3691 0 1.6491e-14
c8627 842 0 2.80434e-13
c8628 2977 2976 1.6e-16
c8629 2951 2954 3.54e-16
c8630 3708 1 1.716e-15
c8631 3024 2798 5.5e-16
c8632 2254 662 1.75e-16
c8633 747 890 3.35e-16
c8634 4667 1 8.43e-16
c8635 4395 4762 1.58e-16
c8636 2662 717 1.58e-16
c8637 3034 2611 5.5e-16
c8638 2098 2114 9.55e-16
c8639 5194 5197 3.54e-16
c8640 3538 3549 1.96e-16
c8641 552 546 1.58e-16
c8642 5104 5111 1.96e-16
c8643 5039 5098 3.54e-16
c8644 2397 2395 1.6e-16
c8645 2392 2391 2.03e-16
c8646 762 2376 1.58e-16
c8647 1457 702 1.58e-16
c8648 907 852 3.15e-16
c8649 5051 0 1.9278e-14
c8650 612 2529 1.58e-16
c8651 921 707 3.15e-16
c8652 1345 1372 1.58e-16
c8653 1464 1016 1.96e-16
c8654 657 921 3.15e-16
c8655 3834 1 1.88e-16
c8656 3839 3840 3.54e-16
c8657 4072 25 7.01e-16
c8658 2559 2751 5.42e-16
c8659 2535 2739 1.58e-16
c8660 3245 3243 1.862e-15
c8661 3048 2645 5.5e-16
c8662 3024 2628 5.5e-16
c8663 4465 1 9.28e-16
c8664 4629 0 1.4233e-14
c8665 4695 4692 6.67e-16
c8666 291 455 1.88e-16
c8667 5074 5073 5.01e-16
c8668 5072 5081 1.58e-16
c8669 3157 707 1.75e-16
c8670 5274 0 1.376e-15
c8671 3236 3231 1.642e-15
c8672 777 1708 3.58e-16
c8673 642 2557 3.15e-16
c8674 2727 0 8e-16
c8675 2216 2215 1.6e-16
c8676 1682 2168 1.58e-16
c8677 4563 4531 4.3e-16
c8678 1431 647 1.58e-16
c8679 1321 807 3.15e-16
c8680 4086 3918 2.48e-16
c8681 3300 0 6.72e-16
c8682 627 3030 4.03e-16
c8683 601 3024 4.48e-16
c8684 2178 777 4.03e-16
c8685 2764 792 1.813e-15
c8686 2781 777 2.22e-16
c8687 1591 1146 3.92e-16
c8688 1595 1596 1.6e-16
c8689 1321 1538 3.92e-16
c8690 1694 1803 1.58e-16
c8691 4196 4214 3.84e-16
c8692 3079 3077 1.6e-16
c8693 1867 1482 1.96e-16
c8694 1393 0 6.72e-16
c8695 5001 4980 1.96e-16
c8696 4972 4978 2.08e-16
c8697 2832 852 1.58e-16
c8698 1735 1 5.808e-15
c8699 3387 3604 3.92e-16
c8700 2186 2189 2.109e-15
c8701 3245 767 1.58e-16
c8702 596 772 3.134e-15
c8703 707 717 3.28e-16
c8704 3619 3617 1.6e-16
c8705 5434 1 7.49e-16
c8706 4776 0 3.19193e-13
c8707 5136 5133 7.46e-16
c8708 3370 3364 9.61e-16
c8709 617 2606 1.58e-16
c8710 2458 2486 2.64e-16
c8711 2480 2476 1.96e-16
c8712 2182 777 7.99e-16
c8713 3722 3409 1.58e-16
c8714 2879 1 1.55e-16
c8715 2194 1726 5.5e-16
c8716 1684 722 4.48e-16
c8717 1327 1537 1.58e-16
c8718 1471 1854 7.84e-16
c8719 2696 2305 1.136e-15
c8720 4747 4361 4.11e-16
c8721 4752 4743 3.46e-16
c8722 1 477 5.175e-15
c8723 130 131 1.88e-16
c8724 426 175 1.88e-16
c8725 1953 822 1.58e-16
c8726 1811 1 5.97e-15
c8727 2127 1 7.87e-16
c8728 3617 767 7.68e-16
c8729 909 1187 4.35e-16
c8730 907 1186 1.88e-16
c8731 890 1179 1.58e-16
c8732 104 1 4.22e-16
c8733 4708 5333 6.9e-16
c8734 5262 149 6.06e-16
c8735 595 2545 9.84e-16
c8736 367 368 3.84e-16
c8737 366 365 6.67e-16
c8738 4207 4204 5.5e-16
c8739 3455 0 3.3874e-14
c8740 2753 1 4.41e-15
c8741 627 890 3.35e-16
c8742 601 883 6.45e-16
c8743 4046 1 6.76e-16
c8744 657 4298 2.4e-16
c8745 3886 3571 1.58e-16
c8746 3340 3339 1.6e-16
c8747 4022 25 3.84e-16
c8748 2342 722 1.58e-16
c8749 2165 858 3.15e-16
c8750 4361 4741 1.96e-16
c8751 1690 1573 1.58e-16
c8752 3612 3610 1.6e-16
c8753 687 2196 3.58e-16
c8754 19 169 3.2e-16
c8755 30 181 6.83e-16
c8756 27 194 1.88e-16
c8757 3610 767 5.03e-16
c8758 3330 842 1.58e-16
c8759 2269 1777 1.58e-16
c8760 601 2234 4.81e-16
c8761 612 1726 3.79e-16
c8762 4922 5106 3.75e-16
c8763 2805 822 1.58e-16
c8764 890 993 3.54e-16
c8765 909 1014 1.58e-16
c8766 4107 4110 5.5e-16
c8767 1345 767 3.15e-16
c8768 2823 2825 2.03e-16
c8769 4024 37 5.71e-16
c8770 2154 852 1.58e-16
c8771 1331 1327 4.431e-15
c8772 1673 1677 1.96e-16
c8773 1482 1477 1.642e-15
c8774 777 784 1.6e-16
c8775 3876 822 3.15e-16
c8776 1939 1951 2.32e-16
c8777 1338 0 5.4701e-14
c8778 4219 1 5.1e-16
c8779 1880 1 1.868e-15
c8780 1870 0 2.93e-15
c8781 3387 3569 1.58e-16
c8782 2486 1 5.343e-15
c8783 842 833 1.078e-15
c8784 596 727 3.134e-15
c8785 5589 1 7.21e-16
c8786 2544 2546 3.84e-16
c8787 5417 468 3.94e-16
c8788 5356 1 9.493e-15
c8789 2482 0 6.72e-16
c8790 1947 792 2.22e-16
c8791 2282 1766 1.136e-15
c8792 911 3030 7.6e-16
c8793 2805 2807 1.862e-15
c8794 146 136 3.75e-16
c8795 5465 5444 5.87e-16
c8796 2739 2741 2.15e-16
c8797 1956 812 1.58e-16
c8798 1584 807 3.79e-16
c8799 1345 1046 5.5e-16
c8800 3139 2645 1.96e-16
c8801 627 986 4.21e-16
c8802 2707 707 1.9e-16
c8803 4201 0 2.0592e-14
c8804 777 1132 1.58e-16
c8805 2039 2023 9.43e-16
c8806 1 250 3.6e-16
c8807 13 247 1.88e-16
c8808 4567 4689 1.58e-16
c8809 4580 4293 5.5e-16
c8810 4810 207 1.88e-16
c8811 934 933 1.96e-16
c8812 3785 3796 3.92e-16
c8813 2834 1 9.28e-16
c8814 1016 647 3.57e-16
c8815 157 0 9.795e-15
c8816 4288 4285 5.5e-16
c8817 543 547 1.372e-15
c8818 537 535 1.88e-16
c8819 3038 3041 2.109e-15
c8820 1489 1491 1.862e-15
c8821 1046 1056 1.418e-15
c8822 642 1408 2.72e-16
c8823 3633 3605 2.64e-16
c8824 2882 2933 2.45e-16
c8825 1757 1754 3.01e-16
c8826 1753 1750 6.44e-16
c8827 954 1 3.56e-16
c8828 3046 3020 1.58e-16
c8829 3024 3023 1.58e-16
c8830 617 1754 1.9e-16
c8831 1694 1533 5.5e-16
c8832 5184 5174 3.92e-16
c8833 429 436 3.54e-16
c8834 2366 2357 3.46e-16
c8835 4531 4893 1.58e-16
c8836 4927 4900 1.79e-16
c8837 226 227 1.58e-16
c8838 2809 2418 4.11e-16
c8839 4081 4079 1.06e-16
c8840 4068 4070 4.33e-16
c8841 4188 3918 2.87e-16
c8842 4753 0 3.74587e-13
c8843 911 890 1.442e-15
c8844 3214 0 1.4092e-14
c8845 925 0 1.0812e-14
c8846 4372 4368 1.96e-16
c8847 1321 1176 1.58e-16
c8848 1327 1166 5.88e-16
c8849 687 2271 5.73e-16
c8850 1254 0 2.5968e-14
c8851 4374 0 6.72e-16
c8852 2987 2944 2.74e-16
c8853 3106 662 1.75e-16
c8854 5280 352 3.54e-16
c8855 5192 207 3.54e-16
c8856 822 1975 2.72e-16
c8857 1964 1959 1.642e-15
c8858 1027 1029 7.84e-16
c8859 15 27 5.8e-16
c8860 32 28 6.67e-16
c8861 3411 868 3.58e-16
c8862 4827 4833 5.87e-16
c8863 5229 5230 3.92e-16
c8864 5267 5257 1.98e-16
c8865 2333 2322 1.58e-16
c8866 3983 3985 1.06e-16
c8867 3996 3918 2.87e-16
c8868 3622 807 5.73e-16
c8869 1218 909 1.96e-16
c8870 920 1114 1.58e-16
c8871 2535 2407 1.58e-16
c8872 4607 4609 1.687e-15
c8873 4619 4612 6.73e-16
c8874 4618 4231 1.96e-16
c8875 3185 0 6.9481e-14
c8876 2535 3017 3.54e-16
c8877 2557 2541 4.274e-15
c8878 3701 4523 1.58e-16
c8879 4879 4890 1.96e-16
c8880 3046 2668 1.58e-16
c8881 3106 3107 1.35e-16
c8882 5232 5234 1.001e-15
c8883 5230 5227 3.54e-16
c8884 3191 3577 5.66e-16
c8885 3583 3574 3.92e-16
c8886 292 297 1.059e-15
c8887 302 310 1.58e-16
c8888 1248 1267 6.73e-16
c8889 3373 3847 5.5e-16
c8890 3370 2987 1.96e-16
c8891 3355 3393 4.3e-16
c8892 5348 0 1.65e-16
c8893 72 0 1.5696e-14
c8894 56 25 7.06e-16
c8895 4379 722 7.68e-16
c8896 3561 0 6.72e-16
c8897 3900 4519 3.92e-16
c8898 1803 1815 2.32e-16
c8899 3747 0 3.7361e-14
c8900 4149 19 9.67e-16
c8901 627 4249 1.58e-16
c8902 3278 3280 2.03e-16
c8903 2679 3177 1.58e-16
c8904 2837 827 7.38e-16
c8905 2557 732 3.15e-16
c8906 1618 1973 1.58e-16
c8907 1706 1884 3.92e-16
c8908 2866 2900 1.466e-15
c8909 2228 0 8e-16
c8910 1997 1 8.43e-16
c8911 3387 3270 5.5e-16
c8912 5131 0 1.1948e-14
c8913 5333 5331 3.92e-16
c8914 2603 2605 2.15e-16
c8915 890 879 3.84e-16
c8916 909 904 1.58e-16
c8917 907 882 1.58e-16
c8918 3327 3712 1.96e-16
c8919 627 3458 1.58e-16
c8920 1371 1373 2.03e-16
c8921 3599 4417 1.96e-16
c8922 4567 4571 4.116e-15
c8923 5577 4563 3.16e-16
c8924 2535 2773 1.58e-16
c8925 1319 1683 1.62e-16
c8926 2535 2170 5.5e-16
c8927 2545 2586 1.58e-16
c8928 673 1 1.65e-16
c8929 2291 662 1.832e-15
c8930 1176 1627 7.84e-16
c8931 1690 1866 1.58e-16
c8932 1907 1516 4.11e-16
c8933 822 1684 3.15e-16
c8934 3409 3638 3.92e-16
c8935 5151 178 3.54e-16
c8936 5047 120 9.42e-16
c8937 5010 526 1.88e-16
c8938 890 903 6.67e-16
c8939 894 893 1.167e-15
c8940 3242 3625 7.84e-16
c8941 4567 4779 1.58e-16
c8942 4571 4395 5.5e-16
c8943 5504 1 3.36e-16
c8944 2493 2504 1.96e-16
c8945 596 637 3.134e-15
c8946 2178 2286 1.58e-16
c8947 1321 1572 3.92e-16
c8948 3140 1 4.41e-15
c8949 1209 0 2.7376e-14
c8950 4302 0 3.3495e-14
c8951 3048 2815 5.5e-16
c8952 2230 2221 3.46e-16
c8953 4684 1 8.43e-16
c8954 4412 4762 2e-16
c8955 4395 4779 1.36e-15
c8956 4788 4782 1.6e-16
c8957 3194 707 1.832e-15
c8958 2696 702 2.22e-16
c8959 3017 858 3.15e-16
c8960 2072 2069 9.03e-16
c8961 426 436 3.75e-16
c8962 468 470 1.96e-16
c8963 2374 0 1.6491e-14
c8964 0 198 6.224e-15
c8965 3976 857 3.1e-16
c8966 3938 3934 1.76e-16
c8967 5025 5135 1.58e-16
c8968 2196 1766 1.58e-16
c8969 2182 2286 1.58e-16
c8970 1477 702 1.58e-16
c8971 592 837 5.8e-16
c8972 2671 2669 1.862e-15
c8973 4236 4232 1.96e-16
c8974 1327 966 1.58e-16
c8975 2584 2595 1.96e-16
c8976 1646 842 1.9e-16
c8977 3900 4455 1.58e-16
c8978 1023 0 4.6497e-14
c8979 849 1 5.57e-16
c8980 4478 1 6.15e-16
c8981 4582 3879 3.54e-16
c8982 4646 0 1.4233e-14
c8983 2837 812 1.58e-16
c8984 2535 692 4.48e-16
c8985 1971 1584 1.532e-15
c8986 1977 1976 5.65e-16
c8987 513 204 1.88e-16
c8988 5101 5103 1.387e-15
c8989 350 352 6.01e-16
c8990 3566 707 3.64e-16
c8991 4457 792 2.72e-16
c8992 110 117 3.54e-16
c8993 3696 3695 1.6e-16
c8994 3418 3419 1.35e-16
c8995 632 2559 3.15e-16
c8996 890 1067 1.96e-16
c8997 2743 0 6.72e-16
c8998 2584 2588 1.96e-16
c8999 1820 677 1.832e-15
c9000 1448 672 2.22e-16
c9001 2194 792 3.15e-16
c9002 3310 3397 1.58e-16
c9003 4031 4030 5.5e-16
c9004 4525 868 2.72e-16
c9005 3684 842 3.15e-16
c9006 3132 1 6.15e-16
c9007 617 3024 4.48e-16
c9008 3582 4399 1.58e-16
c9009 826 25 7.64e-16
c9010 3676 1 5.808e-15
c9011 595 1327 4.03e-16
c9012 3447 3438 3.92e-16
c9013 3055 3441 5.66e-16
c9014 3066 3433 1.58e-16
c9015 632 1732 1.75e-16
c9016 1755 1 2.054e-15
c9017 3265 767 1.58e-16
c9018 777 1922 1.58e-16
c9019 5589 4950 4.06e-16
c9020 4623 4627 1.81e-16
c9021 2178 1902 1.58e-16
c9022 1203 1204 1.21e-16
c9023 3665 1 6.15e-16
c9024 5499 5476 8.66e-16
c9025 1976 827 1.84e-16
c9026 3644 792 2.72e-16
c9027 1691 1324 1.939e-15
c9028 1695 1335 1.018e-15
c9029 1530 1527 3.01e-16
c9030 1526 1523 6.44e-16
c9031 2333 737 1.58e-16
c9032 1482 1866 1.58e-16
c9033 4266 0 1.6491e-14
c9034 2194 737 4.46e-16
c9035 1733 1 1.716e-15
c9036 3158 692 1.339e-15
c9037 426 349 1.88e-16
c9038 4567 4724 3.92e-16
c9039 2182 1902 1.58e-16
c9040 2353 1 1.056e-15
c9041 3528 3525 3.01e-16
c9042 338 339 3.84e-16
c9043 5200 1 1.021e-15
c9044 1879 2371 1.58e-16
c9045 5452 5410 3.41e-16
c9046 3879 3883 2.074e-15
c9047 1905 752 1.832e-15
c9048 657 1432 2.65e-16
c9049 1331 877 3.54e-16
c9050 3475 0 1.4092e-14
c9051 3288 1 1.868e-15
c9052 4680 4299 5.66e-16
c9053 2923 2929 1.572e-15
c9054 2435 797 3.15e-16
c9055 1793 1397 1.96e-16
c9056 1788 1403 1.96e-16
c9057 617 883 6.45e-16
c9058 4055 19 3.45e-16
c9059 3030 3104 1.58e-16
c9060 4378 4741 1.96e-16
c9061 2029 2033 1.96e-16
c9062 1706 1590 1.58e-16
c9063 1542 1 5.808e-15
c9064 1544 0 3.466e-15
c9065 4597 0 8e-16
c9066 777 1101 5.73e-16
c9067 687 3123 5.73e-16
c9068 5251 1 7.49e-16
c9069 2386 2385 1.6e-16
c9070 2378 2376 2.15e-16
c9071 4993 4992 3.92e-16
c9072 4944 4991 1.83e-15
c9073 2274 1777 1.58e-16
c9074 627 1726 1.813e-15
c9075 160 175 1.88e-16
c9076 4328 662 3.64e-16
c9077 2658 2656 1.6e-16
c9078 2653 2652 2.03e-16
c9079 883 1008 3.54e-16
c9080 894 1029 1.58e-16
c9081 4111 4118 2.45e-16
c9082 5580 1 1.871e-15
c9083 5558 5564 6.23e-16
c9084 2541 2684 1.96e-16
c9085 4385 4396 1.96e-16
c9086 2340 722 1.339e-15
c9087 3411 0 3.46872e-13
c9088 3409 777 3.15e-16
c9089 4662 4282 1.96e-16
c9090 687 1828 2.22e-16
c9091 4999 1 2.36e-16
c9092 4549 4980 1.805e-15
c9093 3328 842 1.339e-15
c9094 1499 1 5.97e-15
c9095 749 748 1.6e-16
c9096 427 431 1.372e-15
c9097 3387 3574 1.58e-16
c9098 3411 3586 5.42e-16
c9099 3393 3191 1.58e-16
c9100 1044 1051 2.27e-16
c9101 9 480 4.88e-16
c9102 4100 4101 7.45e-16
c9103 4108 4110 2.239e-15
c9104 5170 5183 9.34e-16
c9105 2542 2561 9.83e-16
c9106 2460 2462 2.03e-16
c9107 5558 5543 7.46e-16
c9108 1086 752 1.75e-16
c9109 1306 1236 1.586e-15
c9110 2533 0 6.9913e-14
c9111 1976 812 1.58e-16
c9112 1576 1588 2.32e-16
c9113 1414 1409 1.642e-15
c9114 599 1 1.65e-16
c9115 528 0 5.6917e-14
c9116 3621 777 2.4e-16
c9117 1835 1448 1.532e-15
c9118 1841 1840 5.65e-16
c9119 1695 1 3.009e-15
c9120 1696 0 5.86e-16
c9121 120 30 3.84e-16
c9122 4567 4706 1.58e-16
c9123 4580 4310 5.5e-16
c9124 4582 4316 1.58e-16
c9125 2442 2444 1.862e-15
c9126 1930 1936 1.418e-15
c9127 1947 1919 2.64e-16
c9128 3829 3773 9.34e-16
c9129 2847 1 6.15e-16
c9130 64 470 2.2e-16
c9131 2741 2737 1.96e-16
c9132 910 925 1.58e-16
c9133 151 152 3.84e-16
c9134 142 129 1.108e-15
c9135 146 165 1.88e-16
c9136 3321 3327 1.418e-15
c9137 4175 4184 3.84e-16
c9138 4189 4188 6.67e-16
c9139 1869 737 1.339e-15
c9140 4021 1 7.71e-16
c9141 4182 25 3.84e-16
c9142 3882 4383 1.96e-16
c9143 4466 4464 1.6e-16
c9144 975 1 3.06e-16
c9145 767 19 1.676e-15
c9146 4012 26 4.58e-16
c9147 4004 0 2.044e-14
c9148 1669 1659 7.53e-16
c9149 1663 1196 3.92e-16
c9150 1506 1 1.716e-15
c9151 4546 4548 3.2e-16
c9152 4344 4731 2.196e-15
c9153 3129 662 1.84e-16
c9154 513 175 1.88e-16
c9155 3604 752 7.38e-16
c9156 2356 2350 1.418e-15
c9157 3811 3807 3.54e-16
c9158 282 15 4.88e-16
c9159 245 9 5.8e-16
c9160 107 334 1.88e-16
c9161 4307 647 1.09e-16
c9162 5352 5291 6.38e-16
c9163 1125 752 6.48e-16
c9164 4092 4093 6.67e-16
c9165 4207 3918 6.32e-16
c9166 1602 797 3.64e-16
c9167 2541 2649 1.58e-16
c9168 939 26 2.65e-15
c9169 3990 25 3.84e-16
c9170 1533 1931 4.36e-16
c9171 1929 1922 1.96e-16
c9172 818 817 1.96e-16
c9173 3048 3024 4.383e-15
c9174 215 0 9.795e-15
c9175 3397 3535 1.58e-16
c9176 3393 858 3.15e-16
c9177 2635 0 1.6491e-14
c9178 632 3472 1.832e-15
c9179 2178 2355 1.96e-16
c9180 3734 3798 1.6e-16
c9181 3983 3992 3.84e-16
c9182 3997 3996 6.67e-16
c9183 4481 807 2.65e-16
c9184 1510 722 1.9e-16
c9185 2559 2424 1.58e-16
c9186 3121 2628 1.58e-16
c9187 4538 4540 2.861e-15
c9188 4553 4543 7.29e-16
c9189 580 581 7.03e-16
c9190 4714 1 2.378e-15
c9191 3024 2685 1.58e-16
c9192 3030 2679 5.88e-16
c9193 1690 1652 4.3e-16
c9194 1655 1 1.056e-15
c9195 1 308 3.6e-16
c9196 902 886 3.84e-16
c9197 4713 0 3.466e-15
c9198 2418 0 6.9484e-14
c9199 915 908 8.57e-16
c9200 0 304 1.5696e-14
c9201 3975 3976 6.4e-16
c9202 5412 468 7.46e-16
c9203 4878 439 1.88e-16
c9204 2182 2355 4.63e-16
c9205 3006 0 1.3715e-14
c9206 1177 1178 7.46e-16
c9207 986 985 3.94e-16
c9208 632 3387 4.48e-16
c9209 4270 4268 2.15e-16
c9210 4278 4277 1.6e-16
c9211 2786 792 2.4e-16
c9212 2629 2620 3.92e-16
c9213 2237 2623 5.66e-16
c9214 2541 3011 1.96e-16
c9215 1473 1041 2.48e-16
c9216 3048 762 3.58e-16
c9217 2879 2896 1.287e-15
c9218 1730 1319 1.58e-16
c9219 1097 0 1.0183e-14
c9220 4814 4812 2.03e-16
c9221 3117 2600 1.136e-15
c9222 2679 3197 2.38e-15
c9223 4523 1 5.808e-15
c9224 3107 647 1.339e-15
c9225 2854 868 2.4e-16
c9226 1684 1901 3.92e-16
c9227 888 893 6.01e-16
c9228 4525 0 3.466e-15
c9229 2244 0 6.72e-16
c9230 642 2583 5.73e-16
c9231 3411 3287 5.5e-16
c9232 6 4 2.84e-16
c9233 1837 717 1.58e-16
c9234 3177 1 5.808e-15
c9235 3886 4319 1.58e-16
c9236 893 1 2.56e-15
c9237 4569 64 1.88e-16
c9238 2559 2214 5.5e-16
c9239 3928 37 5.71e-16
c9240 4352 4354 2.03e-16
c9241 1181 1610 1.58e-16
c9242 1706 1883 1.58e-16
c9243 1690 1871 1.58e-16
c9244 1684 1703 1.58e-16
c9245 1708 1704 3.92e-16
c9246 920 1 3.33e-15
c9247 477 487 8.86e-16
c9248 3576 732 2.72e-16
c9249 3100 3468 1.96e-16
c9250 3048 3359 5.42e-16
c9251 3024 3347 1.58e-16
c9252 1973 0 3.3874e-14
c9253 777 922 3.15e-16
c9254 5074 0 4.4498e-14
c9255 2249 2250 1.6e-16
c9256 2240 2242 2.15e-16
c9257 2605 2601 1.96e-16
c9258 3253 3637 1.58e-16
c9259 4567 4796 1.58e-16
c9260 4571 4412 5.5e-16
c9261 5240 5237 3.92e-16
c9262 5200 5242 1.017e-15
c9263 4855 323 1.88e-16
c9264 91 93 3.84e-16
c9265 3776 3765 6.73e-16
c9266 3768 3769 2.67e-16
c9267 2798 822 1.813e-15
c9268 1343 702 3.15e-16
c9269 2978 1 7.87e-16
c9270 2194 2303 1.58e-16
c9271 2178 2291 1.58e-16
c9272 2231 1715 1.136e-15
c9273 3497 3503 1.418e-15
c9274 4334 4336 1.862e-15
c9275 3633 767 1.58e-16
c9276 4466 782 4.81e-16
c9277 5511 5515 1.202e-15
c9278 1345 1589 3.92e-16
c9279 3549 1 1.868e-15
c9280 1544 1091 4.11e-16
c9281 1331 1419 4.63e-16
c9282 4591 3870 4.97e-16
c9283 4594 4590 1.96e-16
c9284 2594 3088 1.96e-16
c9285 2957 3000 1.489e-15
c9286 2999 2995 1.243e-15
c9287 4144 1 3.79e-14
c9288 762 909 3.15e-16
c9289 4860 4480 1.96e-16
c9290 4701 1 8.43e-16
c9291 4412 4779 1.58e-16
c9292 2753 3262 7.84e-16
c9293 2103 2101 1.133e-15
c9294 2118 2119 3.92e-16
c9295 1 334 3.1683e-14
c9296 3393 3484 1.58e-16
c9297 2196 2490 5.42e-16
c9298 3559 3174 1.96e-16
c9299 3564 3168 1.96e-16
c9300 0 325 5.5081e-14
c9301 1681 1 4.044e-15
c9302 520 519 6.4e-16
c9303 4582 4586 1.6e-16
c9304 792 2384 1.58e-16
c9305 2390 2391 1.35e-16
c9306 2182 2291 1.58e-16
c9307 894 890 4.431e-15
c9308 909 883 4.291e-15
c9309 2015 2495 1.58e-16
c9310 687 685 3.327e-15
c9311 659 25 1.13e-15
c9312 1343 981 1.58e-16
c9313 1196 1200 2.03e-16
c9314 687 4338 2.72e-16
c9315 3882 3639 1.58e-16
c9316 2196 782 3.15e-16
c9317 595 877 1.655e-15
c9318 602 1364 3.64e-16
c9319 687 921 3.15e-16
c9320 1057 0 1.8851e-14
c9321 4119 37 1.88e-16
c9322 747 737 3.28e-16
c9323 3024 3139 3.92e-16
c9324 1845 1840 1.642e-15
c9325 4487 1 1.716e-15
c9326 4663 0 1.4233e-14
c9327 2198 1 2.86e-16
c9328 2402 2393 3.92e-16
c9329 1885 2396 5.66e-16
c9330 1896 2388 1.58e-16
c9331 3185 707 3.15e-16
c9332 2177 0 4.385e-14
c9333 4952 4949 3.92e-16
c9334 4940 4943 3.54e-16
c9335 2308 2306 1.862e-15
c9336 3865 3393 6.89e-16
c9337 3411 3863 1.96e-16
c9338 3397 3236 5.5e-16
c9339 2575 1 6.15e-16
c9340 5580 4950 7.85e-16
c9341 5283 5299 2.109e-15
c9342 2821 1 4.41e-15
c9343 3331 0 6.62e-16
c9344 3141 1 1.716e-15
c9345 1555 767 7.38e-16
c9346 3565 4407 2.38e-15
c9347 2384 737 1.58e-16
c9348 3739 0 5.6946e-14
c9349 1608 1151 1.532e-15
c9350 1614 1613 5.65e-16
c9351 4316 4694 7.84e-16
c9352 3539 3541 2.03e-16
c9353 4972 4988 9.55e-16
c9354 4979 4975 5.6e-16
c9355 3066 3438 1.58e-16
c9356 3367 858 1.58e-16
c9357 773 772 1.96e-16
c9358 3347 3359 2.32e-16
c9359 1937 0 1.6491e-14
c9360 3409 3608 1.58e-16
c9361 5286 5281 7.46e-16
c9362 5170 5158 1.75e-16
c9363 4915 381 1.88e-16
c9364 458 448 8.86e-16
c9365 4640 4642 4.93e-16
c9366 4651 439 1.88e-16
c9367 2194 1919 1.58e-16
c9368 3674 1 1.716e-15
c9369 2545 2546 1.027e-15
c9370 1345 1554 5.42e-16
c9371 1321 1542 1.58e-16
c9372 602 962 1.58e-16
c9373 641 1 5.57e-16
c9374 4564 3879 1.939e-15
c9375 3084 3075 3.92e-16
c9376 2566 3078 5.66e-16
c9377 2577 3070 1.58e-16
c9378 1331 1384 1.58e-16
c9379 2750 737 4.81e-16
c9380 642 2259 2.72e-16
c9381 1880 1874 1.6e-16
c9382 1482 1871 2.386e-15
c9383 1499 1854 1.58e-16
c9384 4507 4504 6.44e-16
c9385 4511 4508 3.01e-16
c9386 4840 1 8.85e-16
c9387 3350 2832 2.38e-15
c9388 1759 1 8.43e-16
c9389 4764 4378 4.11e-16
c9390 4769 4760 3.46e-16
c9391 2078 2086 1.96e-16
c9392 533 534 6.67e-16
c9393 1 439 3.36e-15
c9394 9 419 5.8e-16
c9395 4567 4741 3.92e-16
c9396 5462 1 3.36e-16
c9397 5165 5154 7.92e-16
c9398 3387 3018 3.54e-16
c9399 2369 1 9.28e-16
c9400 782 773 1.078e-15
c9401 2339 0 3.6368e-14
c9402 2911 1 1.88e-16
c9403 894 1201 1.58e-16
c9404 907 1173 3.54e-16
c9405 3900 647 3.15e-16
c9406 3876 672 3.15e-16
c9407 78 218 1.88e-16
c9408 3892 3885 7.06e-16
c9409 3877 3879 1.578e-15
c9410 614 25 1.13e-15
c9411 618 19 1.58e-16
c9412 542 117 1.88e-16
c9413 910 3411 5.03e-16
c9414 1436 1001 1.96e-16
c9415 3886 3599 5.5e-16
c9416 1029 1 2.972e-15
c9417 3345 3356 1.96e-16
c9418 1030 0 6.29e-16
c9419 1684 1607 1.58e-16
c9420 1690 1601 5.88e-16
c9421 4614 0 8e-16
c9422 1960 1958 1.6e-16
c9423 1955 1954 2.03e-16
c9424 762 1106 3.79e-16
c9425 612 25 1.58e-16
c9426 37 494 1.88e-16
c9427 513 436 1.88e-16
c9428 5073 5069 3.54e-16
c9429 2196 2253 3.92e-16
c9430 3908 3909 3.15e-16
c9431 2294 1777 2.38e-15
c9432 113 37 1.88e-16
c9433 59 450 1.88e-16
c9434 3497 662 3.15e-16
c9435 910 2533 3.45e-16
c9436 1134 782 1.58e-16
c9437 1176 837 4e-16
c9438 1430 986 1.96e-16
c9439 1425 996 1.96e-16
c9440 657 4302 1.58e-16
c9441 3882 4417 1.96e-16
c9442 2557 2701 3.92e-16
c9443 796 1 4.03e-16
c9444 1249 1252 1.062e-15
c9445 3428 3018 1.96e-16
c9446 3423 3021 1.96e-16
c9447 1916 1 1.056e-15
c9448 281 117 1.88e-16
c9449 2504 1 1.868e-15
c9450 1038 692 1.58e-16
c9451 79 88 1.58e-16
c9452 2494 0 2.93e-15
c9453 3582 3577 1.642e-15
c9454 2835 2833 1.6e-16
c9455 687 1036 1.35e-16
c9456 1971 837 1.58e-16
c9457 1331 1071 1.58e-16
c9458 779 26 2.65e-15
c9459 1147 1 3.54e-16
c9460 4240 1 6.15e-16
c9461 4378 3537 1.136e-15
c9462 4197 4566 5.8e-16
c9463 3401 3394 7.37e-16
c9464 1769 1414 1.58e-16
c9465 1144 0 9.602e-15
c9466 656 655 6.67e-16
c9467 3694 3691 6.44e-16
c9468 3698 3695 3.01e-16
c9469 1711 0 1.23e-16
c9470 954 955 2.643e-15
c9471 4855 265 1.88e-16
c9472 5177 0 1.9525e-14
c9473 2178 2179 1.239e-15
c9474 134 135 2.84e-16
c9475 3705 3397 1.58e-16
c9476 4328 3486 1.96e-16
c9477 2856 1 1.716e-15
c9478 1192 842 6.38e-16
c9479 284 285 1.58e-16
c9480 920 1010 3.92e-16
c9481 921 1009 2.54e-16
c9482 3886 3881 1.58e-16
c9483 3438 1 5.808e-15
c9484 3440 0 3.466e-15
c9485 4218 19 3.45e-16
c9486 1694 1420 1.58e-16
c9487 1765 1380 1.96e-16
c9488 989 1 3.06e-16
c9489 3506 3123 7.84e-16
c9490 1532 1 8.43e-16
c9491 2033 2025 3.54e-16
c9492 4674 4677 6.02e-16
c9493 513 349 1.88e-16
c9494 27 247 1.88e-16
c9495 2196 2199 1.6e-16
c9496 2084 1 3.36e-16
c9497 408 413 1.059e-15
c9498 404 390 3.84e-16
c9499 3733 3736 2.208e-15
c9500 1414 677 1.58e-16
c9501 1151 797 3.15e-16
c9502 2719 0 3.5142e-14
c9503 751 1 4.03e-16
c9504 1345 1181 5.5e-16
c9505 4396 1 1.868e-15
c9506 3509 3117 2.38e-15
c9507 4386 0 2.93e-15
c9508 728 727 1.96e-16
c9509 4902 4919 1.416e-15
c9510 1760 2252 1.58e-16
c9511 427 15 4.88e-16
c9512 215 217 2.84e-16
c9513 401 19 3.2e-16
c9514 404 37 5.71e-16
c9515 280 291 3.84e-16
c9516 3397 3540 1.58e-16
c9517 3287 3672 1.96e-16
c9518 5044 5273 1.33e-16
c9519 4872 33 1.88e-16
c9520 4085 4079 7.45e-16
c9521 1273 1272 6.09e-16
c9522 1280 1251 1.191e-15
c9523 1076 1080 2.03e-16
c9524 3650 807 3.79e-16
c9525 4472 812 1.58e-16
c9526 5540 5533 9.01e-16
c9527 5530 5535 1.493e-15
c9528 1106 1568 4.36e-16
c9529 1566 1559 1.96e-16
c9530 734 26 2.65e-15
c9531 4624 4626 1.687e-15
c9532 4636 4629 6.73e-16
c9533 4635 4248 1.96e-16
c9534 1706 1352 1.58e-16
c9535 1251 0 1.6532e-14
c9536 2497 858 5.03e-16
c9537 1824 1822 1.6e-16
c9538 1819 1818 2.03e-16
c9539 4731 1 2.378e-15
c9540 3048 2702 1.58e-16
c9541 3046 2696 5.5e-16
c9542 3034 3223 1.58e-16
c9543 2162 2154 7.29e-16
c9544 2149 2151 2.861e-15
c9545 1431 0 6.92e-14
c9546 1675 1 7.21e-16
c9547 1 18 2.87e-16
c9548 5265 5263 3.92e-16
c9549 4730 0 3.466e-15
c9550 595 2555 2.13e-16
c9551 926 930 9.66e-16
c9552 0 33 2.67922e-13
c9553 45 44 1.079e-15
c9554 3411 707 3.15e-16
c9555 5365 1 2.429e-15
c9556 2426 1919 2.48e-16
c9557 1243 1248 3.92e-16
c9558 4878 5136 5.5e-16
c9559 2721 2723 2.03e-16
c9560 657 3411 3.58e-16
c9561 1684 672 3.15e-16
c9562 1708 647 3.15e-16
c9563 3592 0 6.62e-16
c9564 3030 1 2.824e-15
c9565 4540 4539 2.49e-16
c9566 4843 812 1.23e-16
c9567 4172 26 4.58e-16
c9568 4164 0 2.061e-14
c9569 617 4270 1.9e-16
c9570 2545 2803 4.63e-16
c9571 2178 647 3.15e-16
c9572 1738 1744 1.6e-16
c9573 1735 1319 2.386e-15
c9574 1363 1718 1.58e-16
c9575 935 1 6.2e-16
c9576 2144 1257 9.94e-16
c9577 4710 4333 2.48e-16
c9578 15 580 3.92e-16
c9579 310 308 1.257e-15
c9580 2196 1834 1.58e-16
c9581 0 573 1.4803e-14
c9582 3202 732 3.79e-16
c9583 3866 3867 1.6e-16
c9584 3858 3857 9.13e-16
c9585 632 2577 1.58e-16
c9586 2620 1 5.808e-15
c9587 909 902 3.54e-16
c9588 596 875 5.28e-16
c9589 238 1 5.698e-15
c9590 2629 2618 1.96e-16
c9591 1857 717 1.58e-16
c9592 4219 857 3.1e-16
c9593 3011 3003 1.65e-16
c9594 4668 5515 2.137e-15
c9595 3197 1 2.054e-15
c9596 2882 2884 1.001e-15
c9597 1405 971 4.97e-16
c9598 3900 3497 5.5e-16
c9599 2182 647 3.15e-16
c9600 3942 37 1.88e-16
c9601 3237 747 2.65e-16
c9602 706 1 4.03e-16
c9603 2679 3201 1.96e-16
c9604 2685 3196 1.96e-16
c9605 2841 827 1.832e-15
c9606 1684 1900 1.58e-16
c9607 1706 1888 1.58e-16
c9608 1918 1917 9.1e-16
c9609 4491 822 2.72e-16
c9610 1993 0 1.4092e-14
c9611 792 919 3.15e-16
c9612 571 569 1.58e-16
c9613 5032 120 4.44e-16
c9614 3048 722 3.15e-16
c9615 890 888 3.15e-16
c9616 3270 3625 1.58e-16
c9617 3253 3642 2.386e-15
c9618 3651 3645 1.6e-16
c9619 4567 4813 1.58e-16
c9620 4571 4429 5.5e-16
c9621 5482 1 9.493e-15
c9622 2514 2515 9.13e-16
c9623 2511 2512 2.49e-16
c9624 1589 782 1.58e-16
c9625 1345 717 3.58e-16
c9626 1383 1381 1.6e-16
c9627 3966 3918 6.32e-16
c9628 2041 1 1.113e-15
c9629 2172 2320 1.58e-16
c9630 2194 2308 1.58e-16
c9631 1504 707 1.58e-16
c9632 3230 747 2.72e-16
c9633 2545 762 7.99e-16
c9634 668 0 1.1341e-14
c9635 3168 1 5.97e-15
c9636 890 1 2.665e-15
c9637 632 1760 3.15e-16
c9638 1694 1680 1.58e-16
c9639 4525 3684 4.11e-16
c9640 2671 677 1.832e-15
c9641 1223 0 1.8417e-14
c9642 4497 4860 1.96e-16
c9643 2242 2238 1.96e-16
c9644 4429 4779 2e-16
c9645 4412 4796 1.36e-15
c9646 4805 4799 1.6e-16
c9647 2685 722 1.75e-16
c9648 611 610 6.67e-16
c9649 15 541 6.58e-16
c9650 3393 3489 1.58e-16
c9651 3409 3106 1.58e-16
c9652 2393 1 5.808e-15
c9653 647 999 1.58e-16
c9654 2395 0 3.466e-15
c9655 2232 1 1.868e-15
c9656 747 25 1.58e-16
c9657 26 552 8.41e-16
c9658 3645 797 1.84e-16
c9659 3919 901 2.601e-15
c9660 4567 595 2.14e-16
c9661 4582 4604 1.58e-16
c9662 5492 0 2.9101e-14
c9663 5299 1 2.424e-15
c9664 4810 497 1.88e-16
c9665 777 1885 5.73e-16
c9666 1056 717 4e-16
c9667 2545 2401 5.5e-16
c9668 919 737 3.15e-16
c9669 920 1068 1.58e-16
c9670 3678 822 2.72e-16
c9671 2815 2810 1.642e-15
c9672 1666 858 6.67e-16
c9673 1206 1213 7.95e-16
c9674 3898 3656 1.58e-16
c9675 4521 4524 6.44e-16
c9676 2486 837 2.22e-16
c9677 601 1364 7.68e-16
c9678 3377 3367 7.29e-16
c9679 3925 1 7.71e-16
c9680 2753 3260 3.92e-16
c9681 3265 3264 1.6e-16
c9682 3048 3156 3.92e-16
c9683 1721 1722 5.65e-16
c9684 4513 1 8.43e-16
c9685 4680 0 1.4233e-14
c9686 1989 1990 2.48e-16
c9687 1136 0 7.4292e-14
c9688 310 334 1.88e-16
c9689 3555 3558 6.44e-16
c9690 3559 3562 3.01e-16
c9691 717 724 1.6e-16
c9692 497 500 4.6e-16
c9693 3034 858 3.15e-16
c9694 909 722 3.15e-16
c9695 883 1081 1.88e-16
c9696 907 1074 1.58e-16
c9697 966 969 1.58e-16
c9698 5286 5310 1.96e-16
c9699 3356 1 1.868e-15
c9700 1437 692 1.75e-16
c9701 1449 1011 1.96e-16
c9702 1450 1443 6.73e-16
c9703 4522 4524 2.03e-16
c9704 3346 0 2.93e-15
c9705 3141 2634 3.92e-16
c9706 3917 1 6.76e-16
c9707 1868 752 1.75e-16
c9708 1717 1315 4.97e-16
c9709 1694 1454 1.58e-16
c9710 986 1 5.821e-15
c9711 76 1 3.6e-16
c9712 4100 3027 2.573e-15
c9713 1016 0 7.4146e-14
c9714 3066 3458 2.38e-15
c9715 4847 4859 2.62e-16
c9716 2770 782 2.33e-16
c9717 4657 4664 1.81e-16
c9718 2172 1936 1.58e-16
c9719 2178 1930 5.88e-16
c9720 379 1 1.456e-15
c9721 3700 1 8.43e-16
c9722 5417 5476 3.54e-16
c9723 2541 2542 1.239e-15
c9724 1777 672 1.813e-15
c9725 601 962 1.58e-16
c9726 644 26 2.65e-15
c9727 2577 3075 1.58e-16
c9728 4107 1 6.66e-16
c9729 1197 0 6.29e-16
c9730 4857 1 8.85e-16
c9731 5010 207 1.88e-16
c9732 3264 782 5.03e-16
c9733 3411 3022 5.5e-16
c9734 4634 4629 1.536e-15
c9735 2182 1930 5.5e-16
c9736 5429 497 1.96e-16
c9737 5136 1 6.06e-15
c9738 909 1188 3.54e-16
c9739 5450 5481 1.58e-16
c9740 1522 767 1.75e-16
c9741 1086 1525 7.84e-16
c9742 4087 1 4.45e-16
c9743 2453 812 7.68e-16
c9744 3750 0 1.65e-16
c9745 2730 3244 4.97e-16
c9746 3048 3121 5.42e-16
c9747 3024 3109 1.58e-16
c9748 4764 4766 1.6e-16
c9749 2064 2069 7.25e-16
c9750 4631 0 8e-16
c9751 1584 1952 1.96e-16
c9752 627 25 1.58e-16
c9753 339 334 1.88e-16
c9754 3140 3523 7.84e-16
c9755 5072 5064 3.54e-16
c9756 5257 0 1.1948e-14
c9757 146 484 1.88e-16
c9758 2867 2469 4.36e-16
c9759 3898 4434 3.92e-16
c9760 2887 2949 3.54e-16
c9761 2535 2718 3.92e-16
c9762 2361 737 5.03e-16
c9763 2892 0 2.1139e-14
c9764 1597 1595 1.6e-16
c9765 1592 1591 2.03e-16
c9766 4438 777 1.58e-16
c9767 4954 4957 1.96e-16
c9768 4974 4910 2.249e-15
c9769 3349 858 5.03e-16
c9770 2298 1777 1.96e-16
c9771 165 163 1.257e-15
c9772 4793 1 2.3769e-14
c9773 1998 1 5.343e-15
c9774 1057 707 6.38e-16
c9775 2511 0 3.26e-15
c9776 4719 497 1.88e-16
c9777 1553 752 4.81e-16
c9778 3876 797 4.48e-16
c9779 4492 827 1.84e-16
c9780 3882 3384 1.58e-16
c9781 3628 0 1.4092e-14
c9782 3065 2529 1.96e-16
c9783 3060 2532 1.96e-16
c9784 4249 1 1.716e-15
c9785 1853 1854 2.48e-16
c9786 4546 5007 1.443e-15
c9787 3030 3257 1.58e-16
c9788 627 2599 2.4e-16
c9789 923 931 1.58e-16
c9790 15 485 4.88e-16
c9791 479 0 1.4669e-13
c9792 1 482 3.6e-16
c9793 268 263 1.059e-15
c9794 245 244 1.482e-15
c9795 118 123 1.059e-15
c9796 911 3392 1.58e-16
c9797 2472 2470 1.6e-16
c9798 2166 2167 1.76e-16
c9799 119 1 4.92e-16
c9800 3497 3486 1.58e-16
c9801 4407 752 1.84e-16
c9802 3093 0 6.62e-16
c9803 1129 1130 7.51e-16
c9804 3458 1 2.054e-15
c9805 1890 752 5.03e-16
c9806 1327 1339 6.67e-16
c9807 3460 0 8e-16
c9808 3900 4400 3.92e-16
c9809 4474 4475 1.6e-16
c9810 4470 3639 3.92e-16
c9811 3321 822 2.22e-16
c9812 3335 3332 3.01e-16
c9813 3331 3328 6.44e-16
c9814 3034 2566 1.58e-16
c9815 233 252 1.88e-16
c9816 0 189 5.9994e-14
c9817 19 171 3.45e-16
c9818 3361 3820 7.46e-16
c9819 2257 2269 2.32e-16
c9820 1117 1098 1.546e-15
c9821 3713 3710 5.5e-16
c9822 4191 4190 5.5e-16
c9823 161 167 1.372e-15
c9824 160 159 1.88e-16
c9825 156 157 6.67e-16
c9826 2742 2356 5.66e-16
c9827 3048 822 3.58e-16
c9828 3882 4387 1.58e-16
c9829 3898 4399 1.58e-16
c9830 4015 19 3.84e-16
c9831 4024 0 2.0707e-14
c9832 2559 2666 5.42e-16
c9833 2535 2654 1.58e-16
c9834 4578 0 1.1911e-14
c9835 3124 2617 3.92e-16
c9836 3128 3129 1.6e-16
c9837 1949 1948 1.6e-16
c9838 1941 1939 2.15e-16
c9839 1694 1782 4.63e-16
c9840 1508 0 3.3846e-14
c9841 320 484 1.88e-16
c9842 305 252 1.88e-16
c9843 3509 677 1.84e-16
c9844 2656 0 3.466e-15
c9845 944 902 7.05e-16
c9846 2529 1 5.329e-15
c9847 1270 1278 3.54e-16
c9848 1086 1093 7.95e-16
c9849 4492 812 1.58e-16
c9850 1211 1243 4.06e-16
c9851 2617 3125 2.48e-16
c9852 1327 1487 1.96e-16
c9853 762 760 3.327e-15
c9854 1690 1363 5.88e-16
c9855 4198 1 7.71e-16
c9856 2492 852 1.58e-16
c9857 2688 717 1.58e-16
c9858 1448 1816 1.96e-16
c9859 1295 0 3.5619e-14
c9860 592 700 6.34e-16
c9861 612 2569 1.58e-16
c9862 1936 0 3.6368e-14
c9863 1 251 9.8e-16
c9864 3676 837 1.58e-16
c9865 3781 3783 7.82e-16
c9866 3999 3998 5.5e-16
c9867 5543 0 3.3549e-14
c9868 5476 470 9.1e-16
c9869 2424 2435 1.58e-16
c9870 2178 2359 1.58e-16
c9871 4385 737 1.339e-15
c9872 5412 5427 1.96e-16
c9873 5410 5406 7.1e-16
c9874 921 782 3.15e-16
c9875 1016 1013 1.984e-15
c9876 4283 4294 1.96e-16
c9877 1490 1046 4.97e-16
c9878 4552 4556 1.96e-16
c9879 3886 3882 4.431e-15
c9880 3030 2634 1.58e-16
c9881 822 909 3.15e-16
c9882 4571 692 1.33e-16
c9883 2406 767 7.38e-16
c9884 2172 662 4.48e-16
c9885 4831 4829 2.03e-16
c9886 3220 2702 1.96e-16
c9887 3221 3214 6.73e-16
c9888 3128 647 1.9e-16
c9889 2005 2007 1.862e-15
c9890 1618 1624 1.418e-15
c9891 762 1327 4.03e-16
c9892 117 565 1.88e-16
c9893 2182 2359 1.58e-16
c9894 3594 737 1.58e-16
c9895 2358 2360 2.03e-16
c9896 3463 3458 1.642e-15
c9897 4736 1 2.6346e-14
c9898 2790 792 1.58e-16
c9899 1474 1486 2.32e-16
c9900 4640 0 3.55863e-13
c9901 3134 3123 1.58e-16
c9902 1733 1319 1.532e-15
c9903 3984 0 5.142e-14
c9904 908 0 1.5288e-14
c9905 2628 672 1.813e-15
c9906 2858 868 1.58e-16
c9907 1708 1917 5.42e-16
c9908 1684 1905 1.58e-16
c9909 1472 0 1.6491e-14
c9910 1221 1 2.87e-16
c9911 2186 1687 1.121e-15
c9912 2175 1698 7.84e-16
c9913 1694 1718 1.58e-16
c9914 5028 5026 5.62e-16
c9915 1828 1834 1.418e-15
c9916 1845 1817 2.64e-16
c9917 3397 3304 5.5e-16
c9918 2618 1 1.716e-15
c9919 12 15 6.58e-16
c9920 1 11 3.6e-16
c9921 4 0 9.795e-15
c9922 4567 4830 1.58e-16
c9923 4571 4446 5.5e-16
c9924 4872 526 1.88e-16
c9925 2333 2328 1.642e-15
c9926 632 3457 5.03e-16
c9927 3201 1 8.43e-16
c9928 2172 2325 1.58e-16
c9929 4364 4362 1.6e-16
c9930 1684 797 4.48e-16
c9931 3199 3196 3.01e-16
c9932 3585 1 1.056e-15
c9933 1555 1554 9.1e-16
c9934 1262 1 7.49e-16
c9935 4485 822 2.4e-16
c9936 4608 3874 4.97e-16
c9937 4611 4607 1.96e-16
c9938 4159 1 6.66e-16
c9939 3503 0 3.6368e-14
c9940 1431 1798 1.58e-16
c9941 1624 1625 1.35e-16
c9942 1250 0 2.078e-15
c9943 792 894 8.34e-16
c9944 542 378 1.88e-16
c9945 4877 4497 1.96e-16
c9946 3305 797 3.64e-16
c9947 3288 3282 1.6e-16
c9948 1804 0 6.62e-16
c9949 3645 3646 5.65e-16
c9950 3253 3640 1.532e-15
c9951 4429 4796 1.58e-16
c9952 3220 722 3.64e-16
c9953 1 509 1.65e-15
c9954 5151 5234 1.67e-16
c9955 0 526 1.271e-13
c9956 26 520 1.03e-15
c9957 1726 1 5.97e-15
c9958 3958 3960 3.54e-16
c9959 2984 1 1.81e-16
c9960 762 1896 3.79e-16
c9961 73 1 4.563e-15
c9962 397 117 1.88e-16
c9963 55 19 3.45e-16
c9964 59 26 8.41e-16
c9965 3373 3370 1.138e-15
c9966 1158 1159 1.21e-16
c9967 642 3397 7.99e-16
c9968 1321 986 5.5e-16
c9969 1331 1423 1.58e-16
c9970 4152 4150 3.54e-16
c9971 3882 3667 5.88e-16
c9972 3876 3673 1.58e-16
c9973 1947 827 1.58e-16
c9974 1813 1812 1.6e-16
c9975 1805 1803 2.15e-16
c9976 612 881 1.813e-15
c9977 4134 26 4.48e-16
c9978 2104 2100 6.22e-16
c9979 4697 0 1.4233e-14
c9980 2545 722 3.15e-16
c9981 3409 647 4.46e-16
c9982 4567 3873 1.58e-16
c9983 3338 3387 5.5e-16
c9984 1143 807 1.05e-15
c9985 894 737 3.15e-16
c9986 890 1068 3.54e-16
c9987 909 1089 1.58e-16
c9988 4838 5032 1.93e-15
c9989 1846 692 3.64e-16
c9990 1345 842 3.15e-16
c9991 601 593 5.58e-16
c9992 2887 2984 7.46e-16
c9993 5580 5577 5.5e-16
c9994 4520 4567 1.58e-16
c9995 717 19 1.41e-15
c9996 612 4234 1.58e-16
c9997 4431 4424 6.73e-16
c9998 4430 3588 1.96e-16
c9999 657 1431 2.22e-16
c10000 1626 1627 2.48e-16
c10001 2662 3173 1.96e-16
c10002 602 1723 1.09e-16
c10003 4489 0 3.3724e-14
c10004 1956 1 5.808e-15
c10005 5028 120 3.54e-16
c10006 5069 0 3.1318e-14
c10007 1958 0 3.466e-15
c10008 3393 3637 1.58e-16
c10009 3759 3748 3.92e-16
c10010 2491 1981 1.96e-16
c10011 2194 1947 5.5e-16
c10012 1559 767 1.832e-15
c10013 3900 868 3.58e-16
c10014 3143 0 3.3874e-14
c10015 1624 868 1.58e-16
c10016 1343 1116 1.58e-16
c10017 627 977 2.68e-16
c10018 392 146 1.88e-16
c10019 2577 3095 2.38e-15
c10020 372 378 1.58e-16
c10021 4305 1 2.054e-15
c10022 4307 0 8e-16
c10023 5231 178 3.54e-16
c10024 3030 3326 1.96e-16
c10025 3284 782 1.09e-16
c10026 2222 2224 2.03e-16
c10027 4786 4777 3.46e-16
c10028 2383 1 8.43e-16
c10029 978 992 1.96e-16
c10030 448 465 1.138e-15
c10031 466 471 1.059e-15
c10032 464 462 7.1e-16
c10033 426 425 3.84e-16
c10034 407 450 1.88e-16
c10035 4563 4757 1.58e-16
c10036 5221 5222 1.6e-16
c10037 3919 3926 2.45e-16
c10038 5522 381 7.16e-16
c10039 2860 2475 1.96e-16
c10040 2541 2356 1.58e-16
c10041 1091 1508 1.58e-16
c10042 642 3882 4.03e-16
c10043 4108 1 4.64e-16
c10044 3673 4506 7.84e-16
c10045 1947 812 3.15e-16
c10046 1043 1 4.59e-16
c10047 1040 0 1.0077e-14
c10048 1698 1707 1.846e-15
c10049 1131 1 4.044e-15
c10050 1708 1618 5.5e-16
c10051 4648 0 8e-16
c10052 1577 0 6.62e-16
c10053 0 442 1.4515e-14
c10054 33 441 3e-16
c10055 27 455 1.88e-16
c10056 3151 3535 1.58e-16
c10057 4563 4197 1.123e-15
c10058 5098 5101 1.18e-15
c10059 870 871 1.6e-16
c10060 88 426 1.88e-16
c10061 3893 3879 6.4e-16
c10062 1148 782 3.57e-16
c10063 1128 1141 1.58e-16
c10064 99 117 1.58e-16
c10065 1825 677 1.09e-16
c10066 1630 842 1.84e-16
c10067 1440 1001 2.386e-15
c10068 3876 4451 3.92e-16
c10069 662 0 2.8e-13
c10070 2559 2735 3.92e-16
c10071 824 0 7.709e-15
c10072 1965 1956 3.92e-16
c10073 1573 1959 5.66e-16
c10074 3440 3022 4.11e-16
c10075 1257 0 1.8887e-14
c10076 1920 1 1.716e-15
c10077 188 189 1.88e-16
c10078 158 169 2.45e-16
c10079 3540 702 1.58e-16
c10080 4936 4910 3.54e-16
c10081 281 479 1.88e-16
c10082 5283 5305 9.18e-16
c10083 4844 236 1.88e-16
c10084 2759 2373 5.66e-16
c10085 979 980 7.51e-16
c10086 4075 3918 8.1e-16
c10087 3898 3418 1.58e-16
c10088 2843 2844 1.6e-16
c10089 687 1023 1.05e-15
c10090 3107 0 1.6491e-14
c10091 920 1189 1.58e-16
c10092 4321 3480 4.11e-16
c10093 4275 1 8.43e-16
c10094 265 267 3.84e-16
c10095 4847 4846 2.48e-16
c10096 4850 4851 2.83e-16
c10097 3046 3274 1.58e-16
c10098 3030 3262 1.58e-16
c10099 2189 2181 1.606e-15
c10100 868 874 1.6e-16
c10101 3397 3383 1.58e-16
c10102 2322 1 4.41e-15
c10103 967 923 1.546e-15
c10104 4015 4023 3.45e-16
c10105 5136 5127 2.85e-16
c10106 2196 2406 3.92e-16
c10107 2325 0 3.3692e-14
c10108 392 320 1.88e-16
c10109 3108 0 2.93e-15
c10110 920 837 3.15e-16
c10111 3463 4305 2.38e-15
c10112 1910 752 1.09e-16
c10113 1506 1061 1.532e-15
c10114 1512 1511 5.65e-16
c10115 1345 1338 3.54e-16
c10116 657 1016 4.21e-16
c10117 3476 0 6.72e-16
c10118 2923 2920 9.03e-16
c10119 3231 3228 5.5e-16
c10120 2557 807 3.15e-16
c10121 4581 0 1.4914e-14
c10122 3510 3509 5.65e-16
c10123 2542 2175 1.939e-15
c10124 2546 2186 1.018e-15
c10125 2381 2378 3.01e-16
c10126 2377 2374 6.44e-16
c10127 4708 5335 1.96e-16
c10128 2858 0 3.3615e-14
c10129 1137 767 4.98e-16
c10130 922 647 5.14e-16
c10131 179 176 6.67e-16
c10132 3876 3875 1.58e-16
c10133 3898 3872 1.58e-16
c10134 2667 2282 1.96e-16
c10135 2166 2531 4.65e-16
c10136 4111 4119 3.45e-16
c10137 1778 1772 1.6e-16
c10138 4383 3548 1.96e-16
c10139 2559 2671 1.58e-16
c10140 3892 0 5.86e-16
c10141 1528 0 1.4092e-14
c10142 4414 1 9.28e-16
c10143 4991 4980 1.138e-15
c10144 421 422 7.08e-16
c10145 4563 4847 1.58e-16
c10146 4580 4859 1.58e-16
c10147 5170 5172 1.062e-15
c10148 1795 662 7.68e-16
c10149 3249 0 6.72e-16
c10150 3086 1 1.056e-15
c10151 1308 1306 1.095e-15
c10152 1294 1295 7.39e-16
c10153 146 276 1.88e-16
c10154 4487 837 1.58e-16
c10155 5536 5533 3.54e-16
c10156 1834 717 1.58e-16
c10157 1708 868 3.58e-16
c10158 536 9 6.48e-16
c10159 506 1 2.946e-15
c10160 1586 1585 1.6e-16
c10161 1578 1576 2.15e-16
c10162 4641 4643 1.687e-15
c10163 4653 4646 6.73e-16
c10164 4652 4265 1.96e-16
c10165 1708 1386 1.58e-16
c10166 1706 1380 5.5e-16
c10167 2708 717 1.58e-16
c10168 2178 868 4.03e-16
c10169 2194 827 4.46e-16
c10170 4910 4907 1.96e-16
c10171 2821 837 1.58e-16
c10172 3387 3553 3.92e-16
c10173 3304 3659 1.58e-16
c10174 3751 0 1.9795e-14
c10175 2165 1706 4.22e-16
c10176 15 100 5.8e-16
c10177 3598 3591 1.96e-16
c10178 3202 3600 4.36e-16
c10179 4749 0 6.72e-16
c10180 135 0 1.5723e-14
c10181 3397 732 7.99e-16
c10182 2443 1930 4.97e-16
c10183 1251 1226 2.537e-15
c10184 1292 1243 6.67e-16
c10185 4674 381 5.88e-16
c10186 3838 3834 9.07e-16
c10187 3355 3806 9.63e-16
c10188 3836 3725 1.58e-16
c10189 2541 2469 5.88e-16
c10190 2545 822 7.99e-16
c10191 687 3411 3.58e-16
c10192 1571 1572 9.1e-16
c10193 1327 1486 1.58e-16
c10194 1884 722 1.58e-16
c10195 146 139 3.54e-16
c10196 2686 717 1.58e-16
c10197 2182 868 7.99e-16
c10198 1829 1820 3.92e-16
c10199 1437 1823 5.66e-16
c10200 642 1690 4.03e-16
c10201 1098 0 4.6723e-14
c10202 3308 2798 1.58e-16
c10203 1694 1690 4.431e-15
c10204 4214 1 6.056e-15
c10205 4727 4350 2.48e-16
c10206 3145 672 2.72e-16
c10207 2535 767 4.48e-16
c10208 1661 0 3.8751e-14
c10209 777 1343 3.15e-16
c10210 33 34 3.84e-16
c10211 3202 3593 4.11e-16
c10212 3674 837 1.58e-16
c10213 595 2571 2.72e-16
c10214 2427 2439 2.32e-16
c10215 752 746 1.74e-16
c10216 5291 0 5.8577e-14
c10217 2733 2731 1.6e-16
c10218 890 1142 1.96e-16
c10219 921 923 3.15e-16
c10220 5357 5355 5.25e-16
c10221 3041 3033 1.606e-15
c10222 2172 2178 4.078e-15
c10223 2922 2913 1.873e-15
c10224 2545 2807 1.58e-16
c10225 1642 1644 1.862e-15
c10226 1181 1191 1.418e-15
c10227 2696 3213 4.11e-16
c10228 3596 3593 3.01e-16
c10229 3900 0 3.46872e-13
c10230 4930 1 2.73e-16
c10231 3364 3376 3.13e-16
c10232 1624 0 3.6368e-14
c10233 5326 5367 3.18e-16
c10234 2644 1 8.43e-16
c10235 909 962 4.78e-16
c10236 907 961 1.58e-16
c10237 890 955 1.58e-16
c10238 792 1 4.1542e-14
c10239 230 19 8.4e-16
c10240 5482 410 4.44e-16
c10241 2172 2182 4.116e-15
c10242 2178 2512 3.16e-16
c10243 632 3477 1.09e-16
c10244 1576 807 1.58e-16
c10245 1327 722 3.15e-16
c10246 1387 966 3.92e-16
c10247 1391 1392 1.6e-16
c10248 2535 2282 5.5e-16
c10249 2557 2265 5.5e-16
c10250 3109 3121 2.32e-16
c10251 4542 3701 3.92e-16
c10252 4548 4538 7.53e-16
c10253 2288 692 1.75e-16
c10254 2194 812 4.46e-16
c10255 3117 677 1.58e-16
c10256 2798 797 3.15e-16
c10257 4446 4796 2e-16
c10258 4429 4813 1.36e-15
c10259 4822 4816 1.6e-16
c10260 1008 672 1.05e-15
c10261 662 1013 1.58e-16
c10262 15 309 6.58e-16
c10263 1 311 1.607e-15
c10264 0 306 1.051e-14
c10265 3276 812 1.75e-16
c10266 5303 0 1.9525e-14
c10267 612 2194 3.15e-16
c10268 3981 3980 7.81e-16
c10269 3882 732 4.03e-16
c10270 2800 2793 6.73e-16
c10271 1494 722 1.84e-16
c10272 1226 1223 2.14e-15
c10273 632 992 1.58e-16
c10274 3008 0 8e-16
c10275 361 360 1.482e-15
c10276 5414 5411 2.05e-15
c10277 2708 2707 1.6e-16
c10278 4269 4266 6.44e-16
c10279 4273 4270 3.01e-16
c10280 737 1 3.1284e-14
c10281 1964 868 1.58e-16
c10282 2489 827 4.81e-16
c10283 627 881 1.58e-16
c10284 3282 3283 5.65e-16
c10285 26 549 1.03e-15
c10286 448 450 1.88e-16
c10287 465 449 3.84e-16
c10288 3185 3570 1.96e-16
c10289 4567 4231 1.58e-16
c10290 722 715 5.58e-16
c10291 971 647 1.58e-16
c10292 1171 1172 1.238e-15
c10293 883 1083 3.54e-16
c10294 894 1104 1.58e-16
c10295 612 614 5.59e-16
c10296 3378 1 7.21e-16
c10297 1465 692 3.15e-16
c10298 1464 1457 1.96e-16
c10299 612 4254 1.58e-16
c10300 3599 3588 1.58e-16
c10301 2404 752 4.81e-16
c10302 3919 19 3.84e-16
c10303 3928 0 2.0707e-14
c10304 2826 827 5.03e-16
c10305 1694 1482 5.5e-16
c10306 1446 1 6.15e-16
c10307 3482 3475 6.73e-16
c10308 3481 3089 1.96e-16
c10309 4509 0 1.4092e-14
c10310 1976 1 2.054e-15
c10311 561 562 6.67e-16
c10312 2324 1817 2.48e-16
c10313 4469 1 4.442e-15
c10314 4864 4876 2.62e-16
c10315 1978 0 8e-16
c10316 3393 3642 1.58e-16
c10317 3409 3259 1.58e-16
c10318 5286 5338 1.141e-15
c10319 5262 5259 7.46e-16
c10320 3777 3772 3.07e-16
c10321 4053 4054 3.15e-16
c10322 5200 5160 2.45e-16
c10323 2172 1964 5.5e-16
c10324 1331 692 3.15e-16
c10325 4855 381 1.88e-16
c10326 920 1238 3.54e-16
c10327 921 1237 3e-16
c10328 4335 3497 4.97e-16
c10329 1618 852 1.58e-16
c10330 1321 1131 1.58e-16
c10331 1327 1121 5.88e-16
c10332 85 25 7.06e-16
c10333 3046 3343 3.92e-16
c10334 1 303 5.175e-15
c10335 221 220 6.67e-16
c10336 4044 4038 1.96e-16
c10337 4563 4774 1.58e-16
c10338 5207 5198 1.58e-16
c10339 2178 2270 1.96e-16
c10340 384 30 6.83e-16
c10341 3886 702 7.99e-16
c10342 3898 692 4.46e-16
c10343 3031 2538 1.939e-15
c10344 3035 2549 1.018e-15
c10345 1472 707 1.339e-15
c10346 1223 1224 5.5e-16
c10347 4319 4331 2.32e-16
c10348 1933 767 4.81e-16
c10349 632 3876 4.48e-16
c10350 3874 4570 1.62e-16
c10351 2921 2968 1.836e-15
c10352 1065 1 3.06e-16
c10353 842 19 1.676e-15
c10354 4127 1 6.66e-16
c10355 3684 4489 1.58e-16
c10356 3046 2617 1.58e-16
c10357 632 2633 1.58e-16
c10358 4665 0 8e-16
c10359 3168 3523 1.58e-16
c10360 3151 3540 2.386e-15
c10361 3549 3543 1.6e-16
c10362 2395 1879 4.11e-16
c10363 2182 2270 4.63e-16
c10364 2190 1 1.002e-15
c10365 5323 323 5.5e-16
c10366 595 3058 1.58e-16
c10367 78 334 1.88e-16
c10368 5309 5308 1.6e-16
c10369 4140 4134 1.96e-16
c10370 911 881 1.88e-16
c10371 3839 3842 3.54e-16
c10372 3361 1 7.56e-16
c10373 4411 4402 3.46e-16
c10374 4640 5464 1.96e-16
c10375 2662 3143 1.58e-16
c10376 4696 4316 1.96e-16
c10377 2826 812 1.9e-16
c10378 1584 1956 1.58e-16
c10379 1684 1816 3.92e-16
c10380 5074 5095 1.96e-16
c10381 1708 0 3.46872e-13
c10382 1946 1 8.43e-16
c10383 4977 4972 1.291e-15
c10384 3369 858 6.67e-16
c10385 3360 852 2.4e-16
c10386 3030 837 4.03e-16
c10387 1681 2206 7.84e-16
c10388 3387 3219 5.5e-16
c10389 5284 5297 1.96e-16
c10390 4793 410 1.88e-16
c10391 160 88 1.88e-16
c10392 2178 0 3.63418e-13
c10393 2781 0 6.9481e-14
c10394 3882 3429 5.88e-16
c10395 3876 3435 1.58e-16
c10396 602 958 4.98e-16
c10397 3807 0 2.9272e-14
c10398 1602 1593 3.92e-16
c10399 1146 1596 5.66e-16
c10400 1690 1815 1.58e-16
c10401 3077 2533 4.11e-16
c10402 3022 3434 1.96e-16
c10403 3024 3291 1.58e-16
c10404 3046 3279 1.58e-16
c10405 3048 672 3.58e-16
c10406 2182 0 3.3139e-13
c10407 5425 1 2.424e-15
c10408 4922 33 1.88e-16
c10409 2476 1970 3.92e-16
c10410 2480 2481 1.6e-16
c10411 2015 2049 1.466e-15
c10412 1320 1340 2.07e-16
c10413 378 565 1.88e-16
c10414 1690 732 4.03e-16
c10415 919 1039 1.58e-16
c10416 3486 0 3.6368e-14
c10417 1172 0 1.0183e-14
c10418 4251 0 3.3724e-14
c10419 4493 4492 5.65e-16
c10420 4487 3650 1.532e-15
c10421 3343 2832 1.96e-16
c10422 2237 647 1.75e-16
c10423 1584 1131 1.136e-15
c10424 4752 4745 1.96e-16
c10425 4361 4754 1.914e-15
c10426 2662 662 1.58e-16
c10427 130 132 1.58e-16
c10428 3608 3615 1.96e-16
c10429 2323 0 1.6491e-14
c10430 1443 662 1.58e-16
c10431 890 837 3.35e-16
c10432 2277 2274 5.5e-16
c10433 1343 1340 1.58e-16
c10434 1321 1341 3.92e-16
c10435 2567 2169 3.92e-16
c10436 1176 1177 8.58e-16
c10437 3900 4404 1.58e-16
c10438 4037 0 1.5061e-14
c10439 4039 19 3.45e-16
c10440 2541 2305 1.58e-16
c10441 999 0 2.7376e-14
c10442 793 1 1.65e-16
c10443 3030 3088 1.96e-16
c10444 822 1327 4.03e-16
c10445 4427 1 6.15e-16
c10446 291 368 1.88e-16
c10447 5034 5048 1.455e-15
c10448 5158 0 3.0268e-14
c10449 1749 1760 1.58e-16
c10450 88 513 1.88e-16
c10451 909 672 3.15e-16
c10452 4563 4864 1.58e-16
c10453 4580 4876 1.58e-16
c10454 2333 747 1.58e-16
c10455 1055 692 5.74e-16
c10456 986 1418 1.58e-16
c10457 4012 4020 6.67e-16
c10458 4018 4008 7.1e-16
c10459 3102 1 9.28e-16
c10460 2194 747 3.15e-16
c10461 1327 1677 2e-16
c10462 2545 2475 1.58e-16
c10463 632 1772 1.58e-16
c10464 378 397 1.88e-16
c10465 1345 1504 3.92e-16
c10466 777 781 2.19e-16
c10467 1684 1397 5.5e-16
c10468 1694 1786 1.58e-16
c10469 2172 852 3.15e-16
c10470 3411 3570 3.92e-16
c10471 5010 497 1.88e-16
c10472 762 1888 1.58e-16
c10473 2765 2367 4.36e-16
c10474 3685 827 7.68e-16
c10475 4087 857 6.23e-16
c10476 5262 1 6.077e-15
c10477 5173 5175 3.92e-16
c10478 5039 91 3.54e-16
c10479 595 2170 2.22e-16
c10480 1964 0 6.9027e-14
c10481 2810 2807 5.5e-16
c10482 657 662 2.77e-16
c10483 2172 2168 3.54e-16
c10484 4406 737 1.9e-16
c10485 5442 5446 3.54e-16
c10486 2557 2486 5.5e-16
c10487 910 946 1.6e-16
c10488 1706 692 4.46e-16
c10489 1694 702 7.99e-16
c10490 1343 1503 1.58e-16
c10491 1327 1491 1.58e-16
c10492 2248 2646 4.36e-16
c10493 910 3900 5.03e-16
c10494 2512 852 2.8e-16
c10495 2196 858 3.15e-16
c10496 1448 1820 1.58e-16
c10497 632 1684 4.48e-16
c10498 1132 0 1.8851e-14
c10499 4201 19 3.84e-16
c10500 3316 3322 1.6e-16
c10501 3313 2798 2.386e-15
c10502 2815 3296 1.58e-16
c10503 4848 4846 2.03e-16
c10504 792 1321 3.15e-16
c10505 4674 4679 5.53e-16
c10506 2284 1 9.28e-16
c10507 2044 1 2.269e-15
c10508 0 246 1.5696e-14
c10509 5449 439 5.5e-16
c10510 657 3107 1.58e-16
c10511 827 1179 1.58e-16
c10512 5447 5458 9.85e-16
c10513 407 403 1.58e-16
c10514 4736 410 1.88e-16
c10515 2805 2424 3.92e-16
c10516 2535 2271 1.58e-16
c10517 2649 2265 1.58e-16
c10518 2637 2282 1.58e-16
c10519 2248 2639 4.11e-16
c10520 3392 1 6.056e-15
c10521 1482 732 1.813e-15
c10522 1494 1491 5.5e-16
c10523 642 981 4e-16
c10524 632 1398 7.68e-16
c10525 4092 4094 2.254e-15
c10526 3407 0 1.2366e-14
c10527 3237 1 1.868e-15
c10528 2410 767 1.832e-15
c10529 2325 707 1.58e-16
c10530 3390 3027 1.96e-16
c10531 3139 672 2.4e-16
c10532 3048 3047 1.866e-15
c10533 1706 1539 1.58e-16
c10534 2057 1 2.94e-16
c10535 449 450 1.88e-16
c10536 439 437 6.01e-16
c10537 441 442 3.84e-16
c10538 2370 2368 1.6e-16
c10539 4899 4902 3.54e-16
c10540 4929 4928 1.6e-16
c10541 413 1 5.62e-16
c10542 2642 2639 3.01e-16
c10543 2638 2635 6.44e-16
c10544 894 977 3.92e-16
c10545 909 976 1.88e-16
c10546 883 969 1.58e-16
c10547 407 26 8.41e-16
c10548 4634 33 1.88e-16
c10549 1321 737 4.48e-16
c10550 1271 1273 6.73e-16
c10551 3979 25 4.68e-16
c10552 4372 4373 1.6e-16
c10553 4368 3537 3.92e-16
c10554 1331 1640 4.63e-16
c10555 3589 1 1.716e-15
c10556 1276 1 3.15e-16
c10557 4625 4242 4.97e-16
c10558 4628 4624 1.96e-16
c10559 2782 782 7.68e-16
c10560 3531 0 6.9481e-14
c10561 5195 207 5.5e-16
c10562 822 1590 1.58e-16
c10563 1831 1 1.056e-15
c10564 3411 3506 1.58e-16
c10565 3397 3519 4.63e-16
c10566 3659 3658 2.48e-16
c10567 1 25 7.2697e-14
c10568 4446 4813 1.58e-16
c10569 4910 526 3.39e-16
c10570 1919 1 4.41e-15
c10571 2158 2149 7.53e-16
c10572 2153 1635 3.92e-16
c10573 747 1869 1.58e-16
c10574 1036 1037 1.238e-15
c10575 1035 662 6.48e-16
c10576 596 667 3.134e-15
c10577 7 5 1.88e-16
c10578 3409 868 3.15e-16
c10579 5239 5232 1.138e-15
c10580 5151 5261 1.58e-16
c10581 0 38 2.87e-16
c10582 3685 812 3.64e-16
c10583 2428 0 6.62e-16
c10584 627 2194 3.15e-16
c10585 397 479 1.88e-16
c10586 3042 1 1.002e-15
c10587 1939 797 1.58e-16
c10588 1363 1369 1.418e-15
c10589 1104 1 2.972e-15
c10590 3900 3684 5.5e-16
c10591 4542 4545 1.6e-16
c10592 1998 837 2.22e-16
c10593 4503 4884 6.24e-16
c10594 1105 0 6.29e-16
c10595 4150 19 7.04e-16
c10596 4712 4710 2.03e-16
c10597 2294 1783 5.66e-16
c10598 15 569 4.7e-16
c10599 1 568 3.6e-16
c10600 302 301 6.67e-16
c10601 310 311 6.96e-16
c10602 4567 4248 1.58e-16
c10603 1896 2419 4.36e-16
c10604 2417 2410 1.96e-16
c10605 732 730 3.327e-15
c10606 0 562 9.795e-15
c10607 2987 2899 1.761e-15
c10608 2796 1 6.15e-16
c10609 1179 812 8.3e-16
c10610 79 0 1.0822e-14
c10611 59 49 1.88e-16
c10612 2704 2316 4.97e-16
c10613 5324 5323 2.29e-16
c10614 2231 2616 1.96e-16
c10615 4184 4132 1.88e-16
c10616 3001 3006 2.029e-15
c10617 3882 4332 1.96e-16
c10618 4445 4438 1.96e-16
c10619 3599 4447 4.36e-16
c10620 687 1431 1.813e-15
c10621 2846 827 1.09e-16
c10622 1455 1 1.716e-15
c10623 3100 3089 1.58e-16
c10624 564 562 2.84e-16
c10625 5025 31 5.11e-16
c10626 1994 0 6.72e-16
c10627 792 1584 2.22e-16
c10628 1083 722 1.58e-16
c10629 909 914 1.6e-16
c10630 907 905 1.96e-16
c10631 1236 847 3.3e-16
c10632 3713 3712 1.6e-16
c10633 3752 3781 1.37e-16
c10634 4198 857 7.05e-16
c10635 2517 2514 1.6e-16
c10636 1369 1370 1.35e-16
c10637 4580 4563 4.274e-15
c10638 4571 5591 3.54e-16
c10639 2541 2598 1.58e-16
c10640 2594 2583 1.58e-16
c10641 1903 1905 1.862e-15
c10642 1516 1522 1.418e-15
c10643 1694 1693 1.357e-15
c10644 1230 1 3.64e-16
c10645 450 252 1.88e-16
c10646 632 1777 1.58e-16
c10647 1219 0 9.602e-15
c10648 4320 0 6.62e-16
c10649 4864 4862 1.687e-15
c10650 4867 4874 6.73e-16
c10651 5314 5316 1.77e-15
c10652 15 552 5.8e-16
c10653 4776 4777 9.93e-16
c10654 4563 4791 1.58e-16
c10655 5452 1 1.021e-15
c10656 5106 62 7.46e-16
c10657 4872 207 1.88e-16
c10658 4810 468 1.88e-16
c10659 2504 2498 1.6e-16
c10660 1981 2495 2.386e-15
c10661 1987 2503 1.136e-15
c10662 2194 2287 3.92e-16
c10663 3943 3951 9.33e-16
c10664 3944 3942 3.54e-16
c10665 3900 707 3.15e-16
c10666 1056 1057 8.58e-16
c10667 920 1085 3.92e-16
c10668 921 1084 2.54e-16
c10669 595 3393 4.03e-16
c10670 2559 2373 1.58e-16
c10671 657 3900 3.58e-16
c10672 852 0 2.94141e-13
c10673 2957 2969 1.697e-15
c10674 3372 3362 7.53e-16
c10675 3366 2849 3.92e-16
c10676 910 1708 5.03e-16
c10677 2036 2062 3.54e-16
c10678 1604 1 1.056e-15
c10679 418 419 1.482e-15
c10680 3393 3468 1.96e-16
c10681 4682 0 8e-16
c10682 479 478 1.88e-16
c10683 310 303 7.76e-16
c10684 0 207 1.21871e-13
c10685 19 198 3.2e-16
c10686 4844 178 1.88e-16
c10687 2379 0 1.4092e-14
c10688 910 2178 7.97e-16
c10689 911 2194 9.54e-16
c10690 3706 3393 1.96e-16
c10691 3873 3872 3.54e-16
c10692 4236 4237 1.6e-16
c10693 4232 3384 3.92e-16
c10694 4362 707 7.68e-16
c10695 4759 5173 8.41e-16
c10696 2595 2589 1.6e-16
c10697 2170 2586 2.386e-15
c10698 542 494 1.88e-16
c10699 1191 842 2.33e-16
c10700 1442 1438 1.96e-16
c10701 4103 37 1.88e-16
c10702 4104 26 1.075e-15
c10703 1522 1523 1.35e-16
c10704 692 26 7.12e-16
c10705 600 598 5.88e-16
c10706 595 1685 9.02e-16
c10707 1001 1 5.821e-15
c10708 3543 3544 5.65e-16
c10709 4472 1 5.808e-15
c10710 2541 702 4.03e-16
c10711 910 2182 5.03e-16
c10712 1584 1976 2.38e-15
c10713 1708 1833 3.92e-16
c10714 508 204 1.88e-16
c10715 4474 0 3.466e-15
c10716 5103 5130 9.6e-16
c10717 5128 5074 9.34e-16
c10718 5125 5114 3.92e-16
c10719 3462 3453 3.46e-16
c10720 3622 792 1.58e-16
c10721 103 100 2.142e-15
c10722 3871 3872 4.57e-16
c10723 1682 2218 1.58e-16
c10724 5259 149 5.5e-16
c10725 2769 2401 1.96e-16
c10726 2589 2588 1.6e-16
c10727 3749 3734 1.96e-16
c10728 602 3018 1.58e-16
c10729 612 3021 5.73e-16
c10730 3126 1 5.808e-15
c10731 394 1 4.22e-16
c10732 3886 4297 1.58e-16
c10733 3898 3446 5.5e-16
c10734 3900 3452 1.58e-16
c10735 3690 868 1.58e-16
c10736 2862 2861 5.65e-16
c10737 3128 0 3.466e-15
c10738 2559 2534 2.38e-16
c10739 2535 2531 3.54e-16
c10740 3163 3164 5.65e-16
c10741 2260 647 1.84e-16
c10742 1805 1420 1.96e-16
c10743 1151 1593 1.58e-16
c10744 3293 0 3.5724e-14
c10745 3048 3308 5.42e-16
c10746 3024 3296 1.58e-16
c10747 1922 0 3.3874e-14
c10748 1681 2204 3.92e-16
c10749 2209 2208 1.6e-16
c10750 76 78 1.257e-15
c10751 2095 2082 3.92e-16
c10752 2031 2078 2.851e-15
c10753 2080 2077 4.87e-16
c10754 3411 782 3.15e-16
c10755 4623 4624 9.93e-16
c10756 5429 468 1.58e-16
c10757 5558 497 5.5e-16
c10758 3582 767 1.58e-16
c10759 5501 5479 1.74e-16
c10760 5486 5478 3.54e-16
c10761 4878 149 1.88e-16
c10762 2931 1 1.3e-16
c10763 922 868 3.15e-16
c10764 919 827 3.15e-16
c10765 3661 0 3.466e-15
c10766 1524 1525 2.48e-16
c10767 1331 1368 4.63e-16
c10768 2533 3071 1.96e-16
c10769 687 1016 1.813e-15
c10770 4072 1 5.1e-16
c10771 4271 0 1.4092e-14
c10772 3163 692 1.84e-16
c10773 1740 0 8e-16
c10774 3411 3394 3.62e-16
c10775 642 2603 1.58e-16
c10776 2196 2410 1.58e-16
c10777 767 783 1.621e-15
c10778 335 333 1.58e-16
c10779 3769 3773 5.32e-16
c10780 5556 497 3.54e-16
c10781 762 2367 1.813e-15
c10782 747 2384 2.22e-16
c10783 5229 0 3.6193e-14
c10784 2841 2458 7.84e-16
c10785 2654 2661 1.96e-16
c10786 4566 3890 5.8e-16
c10787 1343 880 1.58e-16
c10788 2956 2959 1.931e-15
c10789 3882 3588 1.58e-16
c10790 2427 807 1.58e-16
c10791 4054 26 4.48e-16
c10792 3262 792 1.58e-16
c10793 3046 3105 3.92e-16
c10794 1101 0 3.7193e-14
c10795 4436 1 1.716e-15
c10796 3870 0 4.6935e-14
c10797 2545 672 7.99e-16
c10798 1708 1798 5.42e-16
c10799 1868 2376 7.84e-16
c10800 3048 797 3.15e-16
c10801 2274 2281 1.96e-16
c10802 151 180 3.75e-16
c10803 2689 0 6.62e-16
c10804 4120 4118 3.54e-16
c10805 4563 4881 1.58e-16
c10806 4580 4893 1.58e-16
c10807 4719 468 1.88e-16
c10808 2166 2568 4.97e-16
c10809 2136 2104 1.58e-16
c10810 4514 0 6.9906e-14
c10811 5562 5561 3.54e-16
c10812 3261 0 2.93e-15
c10813 2545 2299 5.5e-16
c10814 1326 1332 2.267e-15
c10815 3565 4370 1.58e-16
c10816 3548 4387 2.386e-15
c10817 4396 4390 1.6e-16
c10818 2345 722 1.84e-16
c10819 3409 0 3.5222e-13
c10820 4658 4660 1.687e-15
c10821 4670 4663 6.73e-16
c10822 4669 4282 1.96e-16
c10823 3253 762 2.22e-16
c10824 3236 777 1.813e-15
c10825 4549 4978 3.65e-16
c10826 5385 265 5.5e-16
c10827 4980 4546 1.589e-15
c10828 5009 5007 8.15e-16
c10829 1886 0 1.6491e-14
c10830 3409 3586 1.58e-16
c10831 3248 752 1.58e-16
c10832 762 1908 1.58e-16
c10833 1051 702 1.35e-16
c10834 1 480 1.65e-15
c10835 4861 4869 1.81e-16
c10836 5170 5174 2.95e-16
c10837 4922 526 1.88e-16
c10838 601 2595 3.64e-16
c10839 602 2214 1.58e-16
c10840 2308 1 5.808e-15
c10841 4038 3918 2.48e-16
c10842 910 3407 1.58e-16
c10843 1236 592 8.21e-16
c10844 1239 596 3.1e-16
c10845 919 812 3.15e-16
c10846 920 1143 1.58e-16
c10847 107 9 5.8e-16
c10848 3623 1 1.716e-15
c10849 4810 64 1.88e-16
c10850 1708 707 3.15e-16
c10851 532 0 2.87e-16
c10852 1448 1840 2.38e-15
c10853 657 1708 3.58e-16
c10854 612 919 3.15e-16
c10855 4022 1 7.08e-16
c10856 4471 4470 2.03e-16
c10857 4476 4474 1.6e-16
c10858 2178 707 3.15e-16
c10859 1769 1767 1.862e-15
c10860 792 1142 2.68e-16
c10861 1701 0 5.4794e-14
c10862 117 19 3.84e-16
c10863 3603 3604 9.1e-16
c10864 601 2588 1.9e-16
c10865 2447 2444 5.5e-16
c10866 2297 1 6.15e-16
c10867 657 2178 4.03e-16
c10868 3219 752 3.15e-16
c10869 3806 3773 1.58e-16
c10870 2841 1 5.808e-15
c10871 909 797 3.15e-16
c10872 883 1156 1.88e-16
c10873 907 1149 1.58e-16
c10874 2843 0 3.466e-15
c10875 3321 3713 2.38e-15
c10876 4183 4182 1.58e-16
c10877 1874 737 1.84e-16
c10878 3886 3548 5.5e-16
c10879 4600 5536 2.037e-15
c10880 2418 782 3.15e-16
c10881 2182 707 3.15e-16
c10882 3311 2798 1.532e-15
c10883 3887 1 3.009e-15
c10884 4004 19 3.84e-16
c10885 1676 1674 1.6e-16
c10886 2645 692 1.58e-16
c10887 1684 1556 1.58e-16
c10888 1690 1550 5.88e-16
c10889 1511 1 2.054e-15
c10890 657 2182 7.99e-16
c10891 1513 0 8e-16
c10892 1944 1941 3.01e-16
c10893 1940 1937 6.44e-16
c10894 833 832 1.96e-16
c10895 508 175 1.88e-16
c10896 3613 752 1.09e-16
c10897 632 2628 1.58e-16
c10898 3390 3396 5.8e-16
c10899 245 1 5.175e-15
c10900 64 180 2.52e-16
c10901 59 194 1.88e-16
c10902 4311 647 3.64e-16
c10903 3469 672 5.73e-16
c10904 1127 752 1.58e-16
c10905 894 991 1.58e-16
c10906 907 963 3.54e-16
c10907 3287 3293 1.418e-15
c10908 4086 4087 1.58e-16
c10909 1783 672 1.58e-16
c10910 1410 1409 5.65e-16
c10911 632 4268 1.58e-16
c10912 2557 2650 3.92e-16
c10913 2323 707 1.339e-15
c10914 1465 1026 1.136e-15
c10915 1299 1 7.308e-15
c10916 1270 0 4.4632e-14
c10917 3789 1 1.257e-15
c10918 4900 4907 8.3e-16
c10919 2299 1783 1.136e-15
c10920 1847 1 9.28e-16
c10921 4446 4830 1.36e-15
c10922 4839 4833 1.6e-16
c10923 2453 1 1.868e-15
c10924 224 0 1.0822e-14
c10925 5529 1 1.662e-15
c10926 2443 0 2.93e-15
c10927 149 1 3.36e-15
c10928 3991 3990 1.58e-16
c10929 4485 797 1.58e-16
c10930 1071 722 2.33e-16
c10931 657 999 1.58e-16
c10932 4281 3446 1.96e-16
c10933 2725 2726 5.65e-16
c10934 1331 1026 1.58e-16
c10935 4606 4600 1.605e-15
c10936 4623 4617 1.025e-15
c10937 4640 4634 1.997e-15
c10938 4657 4651 1.025e-15
c10939 4569 4589 9.14e-16
c10940 2503 842 1.58e-16
c10941 3296 3295 2.48e-16
c10942 3034 3207 4.63e-16
c10943 3658 3657 2.03e-16
c10944 3663 3661 1.6e-16
c10945 2006 1618 4.97e-16
c10946 0 296 5.7196e-14
c10947 4567 4265 1.58e-16
c10948 4725 439 1.88e-16
c10949 908 901 1.575e-15
c10950 891 898 1.682e-15
c10951 3984 3982 1.76e-16
c10952 986 983 1.984e-15
c10953 378 364 1.58e-16
c10954 392 368 1.88e-16
c10955 3435 4268 7.84e-16
c10956 5409 5425 2.109e-15
c10957 146 570 1.88e-16
c10958 4657 1 1.0869e-14
c10959 537 204 1.88e-16
c10960 642 1369 5.73e-16
c10961 1484 1483 1.6e-16
c10962 1476 1474 2.15e-16
c10963 3988 1 6.78e-16
c10964 3898 4349 3.92e-16
c10965 1694 1369 1.58e-16
c10966 4812 4811 2.03e-16
c10967 1481 1 8.43e-16
c10968 3718 4535 1.58e-16
c10969 3112 647 1.84e-16
c10970 2869 842 4.81e-16
c10971 822 1591 1.58e-16
c10972 3690 0 3.6368e-14
c10973 187 186 1.482e-15
c10974 3496 3489 1.96e-16
c10975 3100 3498 4.36e-16
c10976 3587 737 7.38e-16
c10977 4915 4929 9.34e-16
c10978 2341 1828 4.97e-16
c10979 4881 4893 2.62e-16
c10980 9 1 6.5814e-14
c10981 10 11 6.67e-16
c10982 3409 3287 5.5e-16
c10983 1102 737 1.58e-16
c10984 1083 1089 1.58e-16
c10985 4634 526 1.88e-16
c10986 2705 2322 7.84e-16
c10987 4242 4237 1.642e-15
c10988 3882 4331 1.58e-16
c10989 4719 64 1.88e-16
c10990 2668 0 3.5142e-14
c10991 2557 2615 1.58e-16
c10992 2541 2603 1.58e-16
c10993 617 978 1.58e-16
c10994 1345 1136 5.5e-16
c10995 4345 1 1.868e-15
c10996 1706 1691 1.632e-15
c10997 1690 1707 5.63e-16
c10998 3472 3117 1.58e-16
c10999 922 0 3.28459e-13
c11000 4335 0 2.93e-15
c11001 910 2168 1.58e-16
c11002 3083 647 1.58e-16
c11003 2072 2118 4.54e-16
c11004 1652 2117 8.82e-16
c11005 1 511 3.6e-16
c11006 4563 4808 1.58e-16
c11007 3768 3767 8.03e-16
c11008 93 89 6.38e-16
c11009 2172 2304 3.92e-16
c11010 59 15 5.8e-16
c11011 4339 4336 5.5e-16
c11012 2921 0 4.1103e-14
c11013 1540 1542 1.862e-15
c11014 1091 1101 1.418e-15
c11015 1345 1016 5.5e-16
c11016 1321 1001 5.5e-16
c11017 4594 4592 2.15e-16
c11018 4590 4601 1.96e-16
c11019 2041 2521 6.17e-16
c11020 2136 2518 1.96e-16
c11021 612 957 3.79e-16
c11022 1808 1805 3.01e-16
c11023 1804 1801 6.44e-16
c11024 2118 2125 3.92e-16
c11025 2072 2128 9.34e-16
c11026 1620 1 9.28e-16
c11027 3387 3117 5.5e-16
c11028 3411 3134 5.5e-16
c11029 5250 5227 2.12e-16
c11030 5234 5231 2.004e-15
c11031 4699 0 8e-16
c11032 523 513 1.88e-16
c11033 4776 352 1.88e-16
c11034 2406 2405 9.1e-16
c11035 3858 3855 5.5e-16
c11036 601 3075 1.832e-15
c11037 1160 807 1.85e-16
c11038 3719 868 2.65e-16
c11039 4372 717 2.72e-16
c11040 3531 707 3.15e-16
c11041 5388 5283 1.58e-16
c11042 78 73 1.88e-16
c11043 3522 0 2.93e-15
c11044 1181 858 1.58e-16
c11045 687 3503 1.58e-16
c11046 4118 19 7.04e-16
c11047 4423 4419 1.96e-16
c11048 4492 1 2.054e-15
c11049 2837 837 2.4e-16
c11050 2535 717 3.15e-16
c11051 4494 0 8e-16
c11052 5106 5113 1.138e-15
c11053 320 570 1.88e-16
c11054 4943 4936 8.94e-16
c11055 2874 352 1.163e-15
c11056 2569 1 5.808e-15
c11057 2232 2226 1.6e-16
c11058 1682 2223 2.386e-15
c11059 1726 2206 1.58e-16
c11060 3752 3748 6.35e-16
c11061 3605 3606 1.35e-16
c11062 612 3447 2.65e-16
c11063 601 3018 1.58e-16
c11064 3146 1 2.054e-15
c11065 1564 767 1.09e-16
c11066 3701 827 1.58e-16
c11067 3684 852 1.58e-16
c11068 3821 0 2.6642e-14
c11069 1151 1613 2.38e-15
c11070 1708 1832 5.42e-16
c11071 1684 1820 1.58e-16
c11072 3099 3090 3.46e-16
c11073 1887 1505 2.48e-16
c11074 3048 3313 1.58e-16
c11075 3157 3158 1.35e-16
c11076 1942 0 1.4092e-14
c11077 747 919 3.15e-16
c11078 466 468 6.01e-16
c11079 3236 3608 1.58e-16
c11080 2538 0 8.2814e-14
c11081 5410 1 1.0125e-14
c11082 4827 120 5.8e-16
c11083 4804 439 1.88e-16
c11084 3710 3338 1.58e-16
c11085 642 3046 3.15e-16
c11086 1327 672 4.03e-16
c11087 1343 647 4.46e-16
c11088 877 1364 4.36e-16
c11089 3919 3927 3.45e-16
c11090 921 858 3.15e-16
c11091 3616 752 1.58e-16
c11092 4449 767 4.81e-16
c11093 640 1 3.79e-16
c11094 3681 0 8e-16
c11095 4226 4217 1.96e-16
c11096 633 0 7.86e-15
c11097 4571 767 1.33e-16
c11098 2248 672 1.58e-16
c11099 2648 647 4.81e-16
c11100 4769 4762 1.96e-16
c11101 4378 4771 1.914e-15
c11102 2747 3240 1.58e-16
c11103 1756 0 6.72e-16
c11104 1 419 5.175e-15
c11105 4725 4731 5.87e-16
c11106 642 2623 1.58e-16
c11107 0 429 1.4803e-14
c11108 5039 5066 3.63e-16
c11109 687 3143 1.58e-16
c11110 894 827 3.15e-16
c11111 4725 5365 7.98e-16
c11112 910 3409 1.014e-15
c11113 3684 3293 1.136e-15
c11114 2739 762 1.58e-16
c11115 1181 1185 2.03e-16
c11116 537 175 1.88e-16
c11117 3898 3605 1.58e-16
c11118 3009 2929 3.01e-16
c11119 2957 2970 1.96e-16
c11120 2447 807 1.58e-16
c11121 3282 792 1.58e-16
c11122 1689 1701 3.225e-15
c11123 1685 1687 1.578e-15
c11124 1700 1693 7.06e-16
c11125 1028 0 1.4198e-14
c11126 826 1 4.03e-16
c11127 4757 4758 8.22e-16
c11128 1694 2003 4.63e-16
c11129 642 2601 1.58e-16
c11130 3521 3522 2.03e-16
c11131 3874 0 7.0527e-14
c11132 2559 677 3.15e-16
c11133 1249 1 1.113e-15
c11134 1958 1567 4.11e-16
c11135 508 436 1.88e-16
c11136 5094 5093 1.6e-16
c11137 158 171 1.58e-16
c11138 3551 692 4.81e-16
c11139 3350 868 1.58e-16
c11140 91 30 3.84e-16
c11141 93 33 1.88e-16
c11142 2714 1 1.868e-15
c11143 2704 0 2.93e-15
c11144 2764 1 5.97e-15
c11145 2756 2384 1.58e-16
c11146 642 907 3.15e-16
c11147 1338 1324 6.4e-16
c11148 3260 792 1.58e-16
c11149 3116 1 8.43e-16
c11150 595 3034 9.84e-16
c11151 2845 2843 1.6e-16
c11152 2840 2839 2.03e-16
c11153 687 1040 1.85e-16
c11154 2367 722 1.58e-16
c11155 788 0 1.1593e-14
c11156 881 1 5.68e-15
c11157 971 0 7.4292e-14
c11158 4950 4960 1.96e-16
c11159 2281 2272 3.46e-16
c11160 3034 2747 5.5e-16
c11161 4753 352 1.88e-16
c11162 4776 294 1.88e-16
c11163 3397 3396 1.357e-15
c11164 627 2220 1.58e-16
c11165 617 2595 7.68e-16
c11166 601 2214 3.15e-16
c11167 2172 1885 1.58e-16
c11168 2178 1879 5.88e-16
c11169 2328 1 2.054e-15
c11170 4008 4015 1.88e-16
c11171 911 3021 1.88e-16
c11172 4309 4300 3.46e-16
c11173 2518 2525 3.96e-16
c11174 1345 1508 1.58e-16
c11175 4234 1 5.808e-15
c11176 4236 0 3.466e-15
c11177 627 919 3.15e-16
c11178 660 659 1.6e-16
c11179 4196 1 4.608e-15
c11180 2545 797 3.15e-16
c11181 3370 3362 5.95e-16
c11182 3355 2838 1.136e-15
c11183 617 2588 5.03e-16
c11184 2182 1879 5.5e-16
c11185 2306 1 1.716e-15
c11186 657 3128 2.72e-16
c11187 2861 1 2.054e-15
c11188 1193 827 3.57e-16
c11189 894 812 3.15e-16
c11190 890 1143 3.54e-16
c11191 909 1164 1.58e-16
c11192 5412 5473 1.6e-16
c11193 280 282 1.58e-16
c11194 5356 5377 6.16e-16
c11195 5358 5357 5.68e-16
c11196 2863 0 8e-16
c11197 2649 2650 9.1e-16
c11198 919 993 1.58e-16
c11199 3055 0 3.5936e-14
c11200 612 894 8.34e-16
c11201 4858 4856 1.6e-16
c11202 987 0 6.29e-16
c11203 3855 1 6.636e-15
c11204 3048 3070 5.42e-16
c11205 3024 3058 1.58e-16
c11206 617 1397 1.58e-16
c11207 2033 2028 3.73e-16
c11208 1529 0 6.72e-16
c11209 0 256 6.224e-15
c11210 508 349 1.88e-16
c11211 565 494 1.88e-16
c11212 2196 2189 3.54e-16
c11213 410 413 4.6e-16
c11214 910 3020 1.58e-16
c11215 2652 2265 1.532e-15
c11216 909 978 3.54e-16
c11217 592 936 6.34e-16
c11218 3355 842 1.58e-16
c11219 632 4288 1.58e-16
c11220 3404 3038 5.8e-16
c11221 1635 827 1.58e-16
c11222 642 1771 2.72e-16
c11223 1343 1656 1.58e-16
c11224 1327 1644 1.58e-16
c11225 1581 1578 3.01e-16
c11226 1577 1574 6.44e-16
c11227 743 0 1.1593e-14
c11228 4642 4259 4.97e-16
c11229 4645 4641 1.96e-16
c11230 1337 0 5.86e-16
c11231 3398 3399 6.97e-16
c11232 3396 3400 1.71e-16
c11233 2022 207 1.707e-15
c11234 1860 1 6.15e-16
c11235 426 0 1.60597e-13
c11236 1947 1 5.97e-15
c11237 1023 1037 1.96e-16
c11238 1061 737 1.58e-16
c11239 1284 1231 1.96e-16
c11240 910 882 1.96e-16
c11241 911 879 4.84e-16
c11242 146 140 1.58e-16
c11243 3591 0 3.372e-14
c11244 1118 1 4.59e-16
c11245 4182 1 7.08e-16
c11246 1987 858 1.75e-16
c11247 1822 1431 4.11e-16
c11248 1811 1420 1.136e-15
c11249 1115 0 1.0077e-14
c11250 1671 1 2.48e-16
c11251 0 36 3.164e-15
c11252 4729 4727 2.03e-16
c11253 26 22 1.03e-15
c11254 41 49 1.58e-16
c11255 3409 707 4.46e-16
c11256 4567 4282 1.58e-16
c11257 5277 1 4.427e-15
c11258 2437 2436 1.6e-16
c11259 2429 2427 2.15e-16
c11260 3808 3809 1.624e-15
c11261 657 3409 3.15e-16
c11262 3446 4280 1.58e-16
c11263 3548 732 1.813e-15
c11264 921 965 1.96e-16
c11265 4174 4172 2.239e-15
c11266 4164 19 3.84e-16
c11267 3990 1 7.08e-16
c11268 617 3435 2.33e-16
c11269 3876 4366 3.92e-16
c11270 1550 1545 1.642e-15
c11271 911 919 3.45e-16
c11272 910 922 2.45e-16
c11273 3300 3298 1.6e-16
c11274 3295 3294 2.03e-16
c11275 927 0 1.4412e-14
c11276 3799 0 1.65e-16
c11277 1643 1181 4.97e-16
c11278 4722 4720 1.6e-16
c11279 889 893 5.5e-16
c11280 19 573 8.82e-16
c11281 3886 777 7.99e-16
c11282 5010 4992 1.58e-16
c11283 2016 1 1.868e-15
c11284 42 49 7.76e-16
c11285 2006 0 2.93e-15
c11286 5172 0 1.65e-16
c11287 1102 1104 7.84e-16
c11288 4172 4180 6.67e-16
c11289 4178 4168 7.1e-16
c11290 2237 0 3.6368e-14
c11291 4753 294 1.88e-16
c11292 1136 782 3.15e-16
c11293 1393 1391 1.6e-16
c11294 1388 1387 2.03e-16
c11295 3882 4336 1.58e-16
c11296 3898 4348 1.58e-16
c11297 4450 4451 9.1e-16
c11298 4668 5296 4.79e-16
c11299 2535 2632 1.58e-16
c11300 2557 2620 1.58e-16
c11301 3960 26 1.075e-15
c11302 3514 1 5.97e-15
c11303 3119 3118 1.6e-16
c11304 3111 3109 2.15e-16
c11305 2181 1687 1.176e-15
c11306 1457 0 3.3846e-14
c11307 3656 822 1.58e-16
c11308 4385 747 1.58e-16
c11309 2987 2879 1.58e-16
c11310 697 698 1.96e-16
c11311 3500 647 4.81e-16
c11312 3100 672 1.58e-16
c11313 4881 4879 1.23e-15
c11314 3046 732 3.15e-16
c11315 2252 1743 1.58e-16
c11316 1 307 4.22e-16
c11317 9 310 5.8e-16
c11318 4563 4825 1.58e-16
c11319 5452 410 1.58e-16
c11320 5388 1 6.077e-15
c11321 2703 2322 3.92e-16
c11322 2605 0 3.466e-15
c11323 1998 2515 5.69e-16
c11324 1025 672 1.85e-16
c11325 3622 3623 1.35e-16
c11326 3182 0 8e-16
c11327 777 2390 1.58e-16
c11328 1061 1065 2.03e-16
c11329 2792 2788 1.96e-16
c11330 2999 0 1.376e-15
c11331 674 26 2.65e-15
c11332 687 3900 3.58e-16
c11333 1690 1683 1.58e-16
c11334 3555 0 1.6491e-14
c11335 3594 747 1.58e-16
c11336 627 957 1.813e-15
c11337 1234 0 1.1947e-14
c11338 3684 3690 1.418e-15
c11339 4521 4523 1.862e-15
c11340 2892 2906 9.34e-16
c11341 2458 827 2.33e-16
c11342 2480 842 5.03e-16
c11343 1718 1730 2.32e-16
c11344 1633 1 6.15e-16
c11345 615 614 1.6e-16
c11346 1 540 3.6e-16
c11347 4793 4797 1.81e-16
c11348 1885 0 3.6012e-14
c11349 895 886 3.54e-16
c11350 33 557 4.6e-16
c11351 3387 677 4.48e-16
c11352 5426 468 7.94e-16
c11353 2407 2401 1.418e-15
c11354 617 3075 1.58e-16
c11355 4255 4254 5.65e-16
c11356 4249 3385 1.532e-15
c11357 1676 858 7.12e-16
c11358 537 436 1.88e-16
c11359 4523 4522 2.48e-16
c11360 3350 0 1.4092e-14
c11361 3770 1 6.62e-16
c11362 2373 752 2.33e-16
c11363 1721 1315 2.38e-15
c11364 863 1 5.62e-16
c11365 2764 3257 1.58e-16
c11366 3175 3177 1.862e-15
c11367 2662 2668 1.418e-15
c11368 2679 2651 2.64e-16
c11369 3557 3556 2.48e-16
c11370 1999 1607 1.96e-16
c11371 2000 1993 6.73e-16
c11372 897 893 1.36e-16
c11373 717 721 2.19e-16
c11374 4510 0 6.72e-16
c11375 5144 4915 1.407e-15
c11376 565 562 1.099e-15
c11377 478 494 3.84e-16
c11378 3474 3470 1.96e-16
c11379 3557 722 1.58e-16
c11380 3650 792 2.22e-16
c11381 3380 858 3.15e-16
c11382 2205 0 2.93e-15
c11383 907 732 3.15e-16
c11384 5111 0 2.078e-15
c11385 3763 3725 9.37e-16
c11386 601 3449 4.81e-16
c11387 612 3066 3.79e-16
c11388 3296 822 1.58e-16
c11389 3146 2634 5.66e-16
c11390 1716 1727 1.96e-16
c11391 3910 19 3.45e-16
c11392 3908 0 1.5061e-14
c11393 1766 662 1.75e-16
c11394 2009 858 5.03e-16
c11395 4563 3890 3.15e-16
c11396 1708 1837 1.58e-16
c11397 4564 4588 1.003e-15
c11398 1421 0 1.6491e-14
c11399 370 364 1.372e-15
c11400 4936 4946 1.021e-15
c11401 1794 2317 4.36e-16
c11402 3024 692 4.48e-16
c11403 1682 2221 1.532e-15
c11404 2226 2227 5.65e-16
c11405 592 820 6.34e-16
c11406 2773 2401 1.58e-16
c11407 9 339 5.8e-16
c11408 3397 807 7.99e-16
c11409 2540 0 4.3733e-14
c11410 3729 3734 7.46e-16
c11411 632 3048 3.15e-16
c11412 1345 662 3.15e-16
c11413 881 1317 1.58e-16
c11414 1487 692 1.58e-16
c11415 378 19 3.84e-16
c11416 4321 4319 2.15e-16
c11417 4329 4328 1.6e-16
c11418 5429 5427 3.63e-16
c11419 4804 5136 1.96e-16
c11420 659 1 7.18e-16
c11421 2680 2671 3.92e-16
c11422 2288 2674 5.66e-16
c11423 3516 1 9.28e-16
c11424 3697 0 6.72e-16
c11425 827 1 3.1284e-14
c11426 3718 842 1.58e-16
c11427 632 1743 3.15e-16
c11428 1173 0 4.6472e-14
c11429 747 894 8.34e-16
c11430 2730 3248 2.38e-15
c11431 2668 707 1.75e-16
c11432 2535 842 4.48e-16
c11433 5192 5197 7.25e-16
c11434 3409 3022 5.5e-16
c11435 552 553 7.03e-16
c11436 3628 782 1.84e-16
c11437 5025 5119 5.82e-16
c11438 1235 858 3.15e-16
c11439 890 1217 1.96e-16
c11440 5505 5492 3.92e-16
c11441 602 3060 1.9e-16
c11442 922 707 5.14e-16
c11443 921 1038 1.58e-16
c11444 1321 881 5.5e-16
c11445 1331 1372 1.58e-16
c11446 537 349 1.88e-16
c11447 4504 4505 2.03e-16
c11448 5404 528 1.188e-15
c11449 657 922 3.15e-16
c11450 837 25 1.58e-16
c11451 595 596 1.96e-16
c11452 2545 2751 1.58e-16
c11453 4403 4405 2.03e-16
c11454 3254 3243 1.96e-16
c11455 3034 2645 5.5e-16
c11456 1691 1687 2.074e-15
c11457 4384 4761 2.48e-16
c11458 2069 2067 1.462e-15
c11459 1828 1437 1.136e-15
c11460 3151 3519 1.96e-16
c11461 4242 0 6.8854e-14
c11462 323 326 4.6e-16
c11463 479 262 1.88e-16
c11464 2291 2293 2.15e-16
c11465 777 1694 7.99e-16
c11466 2333 1 5.97e-15
c11467 883 692 6.45e-16
c11468 909 1052 4.35e-16
c11469 907 1051 1.88e-16
c11470 890 1044 1.58e-16
c11471 2194 1 4.77e-16
c11472 1053 1054 1.21e-16
c11473 3307 1 1.056e-15
c11474 2737 762 1.58e-16
c11475 1327 797 3.15e-16
c11476 4685 4674 4.67e-16
c11477 4702 4691 4.67e-16
c11478 4719 4708 4.67e-16
c11479 4736 4725 4.67e-16
c11480 4753 4742 4.67e-16
c11481 4770 4759 4.67e-16
c11482 4787 4776 4.67e-16
c11483 4804 4793 4.67e-16
c11484 4821 4810 4.67e-16
c11485 4838 4827 4.67e-16
c11486 4855 4844 4.67e-16
c11487 4872 4861 4.67e-16
c11488 2887 2959 3.54e-16
c11489 632 909 3.15e-16
c11490 4092 3918 2.87e-16
c11491 3247 3243 1.96e-16
c11492 1851 737 1.75e-16
c11493 3276 1 4.41e-15
c11494 3847 0 1.5926e-14
c11495 1595 1136 4.11e-16
c11496 4675 4677 1.687e-15
c11497 4687 4680 6.73e-16
c11498 2810 797 1.58e-16
c11499 1400 1 1.056e-15
c11500 4438 0 3.3724e-14
c11501 2725 737 1.84e-16
c11502 4975 4980 7.46e-16
c11503 2838 858 1.75e-16
c11504 3254 767 7.68e-16
c11505 2524 1 1.052e-15
c11506 2186 2195 1.846e-15
c11507 852 854 5.59e-16
c11508 592 775 6.34e-16
c11509 3747 3745 3.92e-16
c11510 4861 0 2.71188e-13
c11511 4872 497 1.88e-16
c11512 617 2214 3.15e-16
c11513 2482 2480 1.6e-16
c11514 2477 2476 2.03e-16
c11515 3327 3393 1.58e-16
c11516 4175 3893 2.697e-15
c11517 3882 807 4.03e-16
c11518 1327 1086 1.58e-16
c11519 614 1 7.18e-16
c11520 812 1 3.1284e-14
c11521 4254 1 2.054e-15
c11522 1863 1471 1.96e-16
c11523 1864 1857 6.73e-16
c11524 687 1708 3.58e-16
c11525 4256 0 8e-16
c11526 3247 767 5.03e-16
c11527 3046 3258 3.92e-16
c11528 612 1 4.1688e-14
c11529 2332 1 8.43e-16
c11530 687 2178 4.03e-16
c11531 462 25 7.06e-16
c11532 471 0 1.4515e-14
c11533 128 130 2.84e-16
c11534 122 123 3.84e-16
c11535 2469 2464 1.642e-15
c11536 0 497 1.21701e-13
c11537 3606 767 1.339e-15
c11538 5224 238 9.1e-16
c11539 5078 5062 7.38e-16
c11540 1207 868 1.58e-16
c11541 883 1158 3.54e-16
c11542 894 1179 1.58e-16
c11543 111 1 2.87e-16
c11544 102 13 1.88e-16
c11545 2760 2759 5.65e-16
c11546 108 0 1.0822e-14
c11547 2288 2282 1.418e-15
c11548 4200 4208 1.88e-16
c11549 4201 4199 3.54e-16
c11550 1505 752 1.75e-16
c11551 1076 1503 1.58e-16
c11552 4036 1 2.259e-15
c11553 3650 4467 1.58e-16
c11554 3639 4475 5.66e-16
c11555 4481 4472 3.92e-16
c11556 627 894 8.34e-16
c11557 4028 25 1.88e-16
c11558 3048 3075 1.58e-16
c11559 687 2182 7.99e-16
c11560 1708 1567 5.5e-16
c11561 5062 5063 2.67e-16
c11562 3775 3821 4.54e-16
c11563 1749 1777 2.64e-16
c11564 1119 1126 2.27e-16
c11565 894 993 3.54e-16
c11566 4111 4103 9.33e-16
c11567 687 3486 5.73e-16
c11568 1331 767 3.15e-16
c11569 1001 1418 1.58e-16
c11570 4024 19 7.35e-16
c11571 1661 1345 3.25e-16
c11572 3393 762 4.03e-16
c11573 3135 3126 3.92e-16
c11574 2617 3129 5.66e-16
c11575 1556 1939 7.84e-16
c11576 1684 1414 5.5e-16
c11577 1344 0 1.4914e-14
c11578 1869 1 1.716e-15
c11579 3506 662 1.832e-15
c11580 5010 468 1.88e-16
c11581 288 25 7.06e-16
c11582 223 117 1.88e-16
c11583 3387 3174 1.58e-16
c11584 2489 1 1.056e-15
c11585 592 730 6.34e-16
c11586 3565 3174 1.136e-15
c11587 4072 857 3.1e-16
c11588 5569 0 1.5099e-14
c11589 1536 737 4.81e-16
c11590 1270 1226 3.105e-15
c11591 1218 1291 5.45e-16
c11592 3898 767 4.46e-16
c11593 2805 2816 1.96e-16
c11594 3056 0 1.6491e-14
c11595 2739 2738 2.48e-16
c11596 1965 812 7.68e-16
c11597 1331 1046 5.5e-16
c11598 2855 2856 1.35e-16
c11599 1323 0 5.96e-16
c11600 1140 1 3.06e-16
c11601 2525 858 1.58e-16
c11602 1 244 4.59e-16
c11603 5032 91 1.58e-16
c11604 4922 207 1.88e-16
c11605 2260 0 1.4092e-14
c11606 160 0 4.616e-14
c11607 4390 737 1.84e-16
c11608 5410 5409 3.92e-16
c11609 3446 4285 2.386e-15
c11610 4294 4288 1.6e-16
c11611 920 979 1.58e-16
c11612 4657 410 5.8e-16
c11613 1873 722 1.9e-16
c11614 1489 1500 1.96e-16
c11615 657 971 1.58e-16
c11616 3882 4556 2e-16
c11617 2947 2882 6.67e-16
c11618 2918 2929 1.211e-15
c11619 2541 2820 1.96e-16
c11620 2415 767 1.09e-16
c11621 4829 4828 2.03e-16
c11622 2798 3292 1.96e-16
c11623 2617 647 2.33e-16
c11624 2010 2007 5.5e-16
c11625 5540 584 1.345e-15
c11626 5154 236 3.54e-16
c11627 407 15 5.8e-16
c11628 408 1 1.456e-15
c11629 230 233 3.54e-16
c11630 223 215 1.58e-16
c11631 59 247 1.88e-16
c11632 2806 2418 4.97e-16
c11633 4668 0 4.441e-13
c11634 3633 3628 1.642e-15
c11635 911 894 3.45e-16
c11636 3898 4353 1.58e-16
c11637 3876 4365 1.58e-16
c11638 2696 0 6.9481e-14
c11639 4369 4368 2.03e-16
c11640 4374 4372 1.6e-16
c11641 4381 1 1.056e-15
c11642 1690 1730 1.58e-16
c11643 1477 0 1.4092e-14
c11644 1282 1 3.36e-16
c11645 3501 3502 9.1e-16
c11646 5031 5026 1.81e-15
c11647 5152 296 1.188e-15
c11648 890 889 5.85e-16
c11649 4872 4486 1.179e-15
c11650 5277 5314 5.48e-16
c11651 4827 4446 5.2e-16
c11652 4563 4842 1.58e-16
c11653 5258 5257 1.08e-15
c11654 2625 0 8e-16
c11655 632 3072 1.75e-16
c11656 4022 857 1.88e-16
c11657 3937 902 2.538e-15
c11658 3198 0 6.72e-16
c11659 1253 1264 1.96e-16
c11660 1221 1248 4.53e-16
c11661 1690 807 4.03e-16
c11662 3013 0 1.1956e-14
c11663 2541 777 4.03e-16
c11664 919 1114 1.58e-16
c11665 1321 1436 3.92e-16
c11666 4611 4609 2.15e-16
c11667 4607 4618 1.96e-16
c11668 1708 1318 1.58e-16
c11669 1706 1315 1.58e-16
c11670 601 1385 1.58e-16
c11671 3839 3731 1.58e-16
c11672 3030 2855 1.58e-16
c11673 4486 0 3.6274e-14
c11674 2131 2135 9.07e-16
c11675 2118 2106 1.697e-15
c11676 1 524 1.456e-15
c11677 4810 4812 4.93e-16
c11678 5230 5248 1.37e-16
c11679 3185 3191 1.418e-15
c11680 3572 3574 1.862e-15
c11681 0 513 1.96446e-13
c11682 3659 807 1.58e-16
c11683 48 1 9.8e-16
c11684 42 15 5.8e-16
c11685 5321 0 3.1318e-14
c11686 3373 2899 1.96e-16
c11687 3355 3411 3.92e-16
c11688 4368 722 1.339e-15
c11689 617 3095 1.58e-16
c11690 1327 1435 1.58e-16
c11691 1363 880 1.136e-15
c11692 3718 3747 1.048e-15
c11693 687 3531 2.22e-16
c11694 3886 4519 4.63e-16
c11695 2541 2785 1.58e-16
c11696 1074 0 2.7196e-14
c11697 4136 25 7.01e-16
c11698 3262 2764 1.58e-16
c11699 513 514 6.96e-16
c11700 4582 4592 1.58e-16
c11701 3577 722 1.58e-16
c11702 5133 1 1.81e-16
c11703 2698 2697 1.6e-16
c11704 592 702 5.8e-16
c11705 3397 3671 1.58e-16
c11706 2771 0 1.6491e-14
c11707 1100 722 1.58e-16
c11708 894 879 1.88e-16
c11709 5348 5347 1.6e-16
c11710 2776 777 1.58e-16
c11711 2603 2602 2.48e-16
c11712 1343 868 3.15e-16
c11713 1321 827 4.48e-16
c11714 627 3066 1.813e-15
c11715 3316 822 1.58e-16
c11716 2651 1 4.41e-15
c11717 1355 881 1.58e-16
c11718 3839 3820 1.58e-16
c11719 1636 1176 1.96e-16
c11720 1637 1630 6.73e-16
c11721 2841 837 1.58e-16
c11722 1690 1471 1.58e-16
c11723 595 1315 1.655e-15
c11724 602 1727 3.64e-16
c11725 632 2257 1.832e-15
c11726 1904 1516 4.97e-16
c11727 1573 0 3.6368e-14
c11728 5079 0 1.4815e-14
c11729 5031 120 5.5e-16
c11730 2593 1 8.43e-16
c11731 1082 732 2.68e-16
c11732 5291 5278 1.96e-16
c11733 3635 3628 6.73e-16
c11734 3634 3242 1.96e-16
c11735 747 1 4.1542e-14
c11736 5010 64 1.88e-16
c11737 3294 822 1.58e-16
c11738 3943 3937 1.58e-16
c11739 2178 1766 1.58e-16
c11740 921 1203 1.58e-16
c11741 1706 767 4.46e-16
c11742 3529 1 6.15e-16
c11743 4894 858 1.23e-16
c11744 687 1453 2.4e-16
c11745 2759 752 1.58e-16
c11746 1888 1900 2.32e-16
c11747 2955 2921 1.75e-16
c11748 1207 0 1.8851e-14
c11749 3034 2815 5.5e-16
c11750 1403 1 4.41e-15
c11751 1787 0 6.62e-16
c11752 3242 3627 1.96e-16
c11753 3236 3632 1.96e-16
c11754 4786 4779 1.96e-16
c11755 4395 4788 1.914e-15
c11756 3387 3467 1.58e-16
c11757 3203 707 3.64e-16
c11758 2384 1 5.97e-15
c11759 657 2237 5.73e-16
c11760 456 454 1.58e-16
c11761 422 436 1.58e-16
c11762 4580 4758 3.92e-16
c11763 0 209 5.5401e-14
c11764 2380 0 6.72e-16
c11765 294 325 1.88e-16
c11766 3928 3926 3.54e-16
c11767 3918 3909 2.48e-16
c11768 2182 1766 1.58e-16
c11769 1031 702 1.813e-15
c11770 601 3060 5.03e-16
c11771 2680 2669 1.96e-16
c11772 4233 4232 2.03e-16
c11773 4238 4236 1.6e-16
c11774 4110 1 6.76e-16
c11775 3886 4455 1.58e-16
c11776 3876 3616 5.5e-16
c11777 4086 25 3.84e-16
c11778 606 593 7.23e-16
c11779 597 598 1.6e-16
c11780 4774 4775 8.22e-16
c11781 632 2622 1.9e-16
c11782 2070 2062 3.54e-16
c11783 1706 2019 1.58e-16
c11784 1690 2007 1.58e-16
c11785 4259 0 6.9337e-14
c11786 1980 1971 3.46e-16
c11787 5115 5113 3.92e-16
c11788 3454 3456 2.03e-16
c11789 4940 4944 5.32e-16
c11790 632 2545 3.15e-16
c11791 105 100 1.482e-15
c11792 4336 702 1.58e-16
c11793 5296 5298 1.062e-15
c11794 2750 1 1.056e-15
c11795 894 1067 3.92e-16
c11796 909 1066 1.88e-16
c11797 883 1059 1.58e-16
c11798 5262 5160 1.58e-16
c11799 3323 1 9.28e-16
c11800 2584 2585 2.03e-16
c11801 1829 677 3.64e-16
c11802 1627 827 1.832e-15
c11803 1321 812 4.48e-16
c11804 4028 4022 1.96e-16
c11805 662 19 1.676e-15
c11806 3582 3554 2.64e-16
c11807 3685 1 1.868e-15
c11808 1416 1 9.28e-16
c11809 612 1321 3.15e-16
c11810 3436 3438 1.862e-15
c11811 3022 3055 1.418e-15
c11812 3066 3021 2.64e-16
c11813 1925 1 2.054e-15
c11814 181 178 4.6e-16
c11815 175 164 3.84e-16
c11816 186 194 1.58e-16
c11817 2293 2289 1.96e-16
c11818 2747 767 3.15e-16
c11819 1927 0 8e-16
c11820 777 1931 2.65e-16
c11821 2780 2384 1.96e-16
c11822 2850 2841 3.92e-16
c11823 3112 0 1.4092e-14
c11824 1584 827 1.58e-16
c11825 1179 1 2.972e-15
c11826 1482 1471 1.58e-16
c11827 4272 0 6.72e-16
c11828 1180 0 6.29e-16
c11829 792 1143 1.58e-16
c11830 3024 3275 3.92e-16
c11831 1913 1908 1.642e-15
c11832 627 1 4.1542e-14
c11833 969 976 2.27e-16
c11834 4023 4024 6.4e-16
c11835 4600 3873 1.179e-15
c11836 4708 4715 1.81e-16
c11837 4571 4711 1.58e-16
c11838 4582 4723 1.58e-16
c11839 5417 439 3.54e-16
c11840 5493 5494 1.6e-16
c11841 5452 5449 7.46e-16
c11842 1209 858 1.58e-16
c11843 399 393 1.372e-15
c11844 2557 2322 1.58e-16
c11845 1914 752 3.64e-16
c11846 1061 1511 2.38e-15
c11847 3083 0 6.9481e-14
c11848 3650 4472 1.58e-16
c11849 4293 4299 9.42e-16
c11850 2923 2882 2.45e-16
c11851 1785 1403 2.48e-16
c11852 911 1335 1.829e-15
c11853 993 1 1.56e-15
c11854 3030 2583 1.58e-16
c11855 1551 1 1.868e-15
c11856 4603 1 1.013e-15
c11857 1541 0 2.93e-15
c11858 33 352 1.88e-16
c11859 218 204 1.88e-16
c11860 27 368 1.88e-16
c11861 2375 2376 2.48e-16
c11862 1113 767 1.58e-16
c11863 157 158 1.482e-15
c11864 129 171 9.5e-16
c11865 288 245 1.88e-16
c11866 3898 3895 1.58e-16
c11867 4119 4120 6.4e-16
c11868 3258 777 2.4e-16
c11869 4659 4276 4.97e-16
c11870 4662 4658 1.96e-16
c11871 1567 1922 1.58e-16
c11872 2987 2978 8.15e-16
c11873 2093 0 2.28e-15
c11874 1895 1 8.43e-16
c11875 5362 354 8.44e-16
c11876 3326 827 7.38e-16
c11877 15 448 5.8e-16
c11878 3411 3191 1.58e-16
c11879 2552 2538 6.4e-16
c11880 4571 4860 3.92e-16
c11881 1043 1044 1.213e-15
c11882 3786 3785 1.96e-16
c11883 3756 3729 1.79e-16
c11884 4103 4102 1.58e-16
c11885 1306 1307 1.361e-15
c11886 3900 782 3.15e-16
c11887 920 1160 3.92e-16
c11888 921 1159 2.54e-16
c11889 536 1 1.073e-15
c11890 1584 812 3.15e-16
c11891 1131 1576 7.84e-16
c11892 1844 1835 3.46e-16
c11893 3241 752 7.38e-16
c11894 3024 3240 1.58e-16
c11895 3046 3228 1.58e-16
c11896 1688 0 6.78e-16
c11897 1 185 4.22e-16
c11898 3393 722 3.15e-16
c11899 4567 4316 1.58e-16
c11900 5051 5047 1.881e-15
c11901 4759 323 1.88e-16
c11902 2442 2453 1.96e-16
c11903 2743 2741 1.6e-16
c11904 2738 2737 2.03e-16
c11905 911 888 1.58e-16
c11906 687 3409 3.15e-16
c11907 3021 1 4.044e-15
c11908 3038 3047 1.846e-15
c11909 3422 0 6.62e-16
c11910 2557 2837 3.92e-16
c11911 767 26 7.12e-16
c11912 4188 25 1.88e-16
c11913 627 3463 2.22e-16
c11914 4457 3622 1.96e-16
c11915 4462 3616 1.96e-16
c11916 1343 0 3.5222e-13
c11917 911 1 2.9239e-14
c11918 4739 4737 1.6e-16
c11919 2611 662 1.58e-16
c11920 4575 0 5.86e-16
c11921 5053 5031 9.18e-16
c11922 5029 5033 5.6e-16
c11923 3828 3807 6.16e-16
c11924 632 3109 1.832e-15
c11925 5379 5326 3.18e-16
c11926 5377 5365 1.96e-16
c11927 4838 236 1.88e-16
c11928 4589 5546 6.02e-16
c11929 2541 2819 1.58e-16
c11930 1146 1148 7.72e-16
c11931 642 4287 2.72e-16
c11932 3876 4370 1.58e-16
c11933 3900 4382 5.42e-16
c11934 3996 25 1.88e-16
c11935 2541 2254 1.58e-16
c11936 2338 692 1.58e-16
c11937 1652 868 2.22e-16
c11938 1647 1644 5.5e-16
c11939 1211 1221 5.7e-16
c11940 3211 3209 1.862e-15
c11941 4562 0 6.78e-16
c11942 1920 1533 1.532e-15
c11943 1926 1925 5.65e-16
c11944 1706 1747 1.58e-16
c11945 1690 1735 1.58e-16
c11946 1681 1680 3.54e-16
c11947 30 584 3.84e-16
c11948 5010 5013 3.54e-16
c11949 4406 747 2.72e-16
c11950 3034 3024 4.116e-15
c11951 3364 3030 3.16e-16
c11952 3202 3197 1.642e-15
c11953 5174 0 2.8602e-14
c11954 4915 120 1.88e-16
c11955 3326 812 1.58e-16
c11956 3397 3140 1.58e-16
c11957 3659 3671 2.32e-16
c11958 3411 858 3.15e-16
c11959 2641 0 6.72e-16
c11960 2136 2028 1.58e-16
c11961 632 3481 3.64e-16
c11962 1398 1389 3.92e-16
c11963 966 1392 5.66e-16
c11964 792 2423 2.4e-16
c11965 1236 920 8.58e-16
c11966 2545 2424 1.58e-16
c11967 2557 792 3.15e-16
c11968 374 37 1.88e-16
c11969 2600 2628 2.64e-16
c11970 1345 1453 3.92e-16
c11971 3208 762 5.73e-16
c11972 4555 4553 1.6e-16
c11973 2491 868 2.4e-16
c11974 617 1385 7.38e-16
c11975 577 580 3.54e-16
c11976 568 563 1.482e-15
c11977 3134 662 3.15e-16
c11978 2255 1743 1.532e-15
c11979 1738 1735 5.5e-16
c11980 4327 1 6.275e-15
c11981 4503 0 3.6405e-14
c11982 1670 1667 1.138e-15
c11983 15 274 5.8e-16
c11984 426 565 1.88e-16
c11985 4827 4834 1.81e-16
c11986 912 891 1.132e-15
c11987 737 731 1.74e-16
c11988 0 314 6.224e-15
c11989 33 294 3.08e-16
c11990 3702 3703 1.6e-16
c11991 2196 2354 5.42e-16
c11992 5357 294 3.54e-16
c11993 361 362 5.8e-16
c11994 3310 868 5.73e-16
c11995 5435 5434 1.6e-16
c11996 5406 5409 3.54e-16
c11997 5427 5426 3.92e-16
c11998 2535 2418 5.5e-16
c11999 2705 2714 3.92e-16
c12000 2333 2700 1.58e-16
c12001 4267 4268 2.48e-16
c12002 2231 2237 1.418e-15
c12003 1867 707 1.58e-16
c12004 1479 1476 3.01e-16
c12005 1475 1472 6.44e-16
c12006 617 611 1.74e-16
c12007 3034 762 7.99e-16
c12008 879 1 2.061e-15
c12009 3282 2764 2.38e-15
c12010 3213 732 2.72e-16
c12011 4532 1 1.868e-15
c12012 3205 3203 1.6e-16
c12013 2557 737 4.46e-16
c12014 747 1321 3.15e-16
c12015 462 419 1.88e-16
c12016 470 439 1.88e-16
c12017 898 886 4.268e-15
c12018 4582 4609 1.58e-16
c12019 2251 1 1.056e-15
c12020 595 2196 3.15e-16
c12021 218 175 1.88e-16
c12022 4855 5103 9.43e-16
c12023 3397 3676 1.58e-16
c12024 2220 1 4.41e-15
c12025 8 16 1.372e-15
c12026 7 6 1.88e-16
c12027 1345 852 3.58e-16
c12028 2172 2491 3.92e-16
c12029 3186 1 1.868e-15
c12030 2905 2906 1.6e-16
c12031 2879 2876 3.54e-16
c12032 2896 2897 3.92e-16
c12033 903 1 6.93e-16
c12034 3928 19 7.35e-16
c12035 2545 2214 5.5e-16
c12036 617 995 1.58e-16
c12037 885 0 5.96e-16
c12038 1706 1488 1.58e-16
c12039 601 1727 7.68e-16
c12040 1440 1 5.808e-15
c12041 1442 0 3.466e-15
c12042 919 1 5.545e-15
c12043 1694 1704 3.92e-16
c12044 2335 2334 1.6e-16
c12045 3034 3359 1.58e-16
c12046 2240 2239 2.48e-16
c12047 2607 2605 1.6e-16
c12048 2602 2601 2.03e-16
c12049 3253 3242 1.58e-16
c12050 4182 857 1.88e-16
c12051 4770 323 1.88e-16
c12052 2178 2490 1.58e-16
c12053 2876 2877 5.67e-16
c12054 78 9 5.8e-16
c12055 392 136 1.88e-16
c12056 4334 4345 1.96e-16
c12057 5513 5511 1.167e-15
c12058 1708 782 3.15e-16
c12059 1331 1589 4.63e-16
c12060 632 1327 3.15e-16
c12061 3538 1 1.716e-15
c12062 1541 1091 4.97e-16
c12063 3731 1 1.55e-16
c12064 2178 782 3.15e-16
c12065 612 1355 1.58e-16
c12066 2781 782 3.15e-16
c12067 3271 2753 1.96e-16
c12068 3387 3472 1.58e-16
c12069 3411 3484 5.42e-16
c12070 3393 3089 1.58e-16
c12071 2696 707 3.15e-16
c12072 632 2248 3.15e-16
c12073 4759 4765 5.87e-16
c12074 4580 4775 3.92e-16
c12075 5074 62 1.58e-16
c12076 2196 1970 1.58e-16
c12077 2182 2490 1.58e-16
c12078 517 523 1.58e-16
c12079 3990 857 1.88e-16
c12080 5484 5492 1.725e-15
c12081 4742 5177 1.96e-16
c12082 1477 707 1.84e-16
c12083 1224 1234 2.74e-16
c12084 1232 909 1.96e-16
c12085 601 3080 1.09e-16
c12086 2756 1 5.808e-15
c12087 64 65 3.84e-16
c12088 3716 1 6.15e-16
c12089 3900 3633 5.5e-16
c12090 2923 2969 4.54e-16
c12091 1947 837 1.58e-16
c12092 2182 782 3.15e-16
c12093 822 1158 1.05e-15
c12094 687 922 3.15e-16
c12095 4119 19 3.45e-16
c12096 4401 4778 2.48e-16
c12097 3006 858 1.58e-16
c12098 4276 0 6.9337e-14
c12099 792 1576 1.58e-16
c12100 5106 5101 7.46e-16
c12101 5104 5072 1.75e-16
c12102 4759 265 1.88e-16
c12103 2391 2393 1.862e-15
c12104 1879 1885 1.418e-15
c12105 1896 1868 2.64e-16
c12106 3411 3865 6.7e-16
c12107 5298 0 1.65e-16
c12108 5286 323 1.58e-16
c12109 5084 1 3.36e-16
c12110 4945 4943 9.16e-16
c12111 2766 1 9.28e-16
c12112 4356 702 1.58e-16
c12113 5308 5300 3.92e-16
c12114 2214 2582 1.96e-16
c12115 3336 1 6.15e-16
c12116 1448 677 3.15e-16
c12117 4525 858 5.03e-16
c12118 3820 1 2.223e-15
c12119 4415 4413 1.6e-16
c12120 2387 737 4.81e-16
c12121 1617 1608 3.46e-16
c12122 4692 4694 1.687e-15
c12123 4704 4697 6.73e-16
c12124 4703 4316 1.96e-16
c12125 627 1321 3.15e-16
c12126 4944 4989 3.18e-16
c12127 3379 858 7.12e-16
c12128 1943 0 6.72e-16
c12129 792 1533 1.58e-16
c12130 777 1550 3.79e-16
c12131 5286 5301 1.96e-16
c12132 5284 5280 7.1e-16
c12133 1074 707 8.3e-16
c12134 596 787 3.134e-15
c12135 2475 2476 1.35e-16
c12136 595 931 8.22e-16
c12137 612 955 1.58e-16
c12138 1601 868 1.58e-16
c12139 2001 827 4.81e-16
c12140 1345 1101 1.58e-16
c12141 1343 1091 5.5e-16
c12142 1331 1554 1.58e-16
c12143 3393 822 4.03e-16
c12144 3073 3075 1.862e-15
c12145 2533 2566 1.418e-15
c12146 2577 2532 2.64e-16
c12147 1482 1880 4.36e-16
c12148 1878 1871 1.96e-16
c12149 3048 3292 3.92e-16
c12150 3397 3433 1.58e-16
c12151 2031 2086 1.141e-15
c12152 4606 4612 5.87e-16
c12153 4725 4733 1.81e-16
c12154 4571 4728 1.58e-16
c12155 4582 4740 1.58e-16
c12156 4742 33 1.88e-16
c12157 2487 2478 3.92e-16
c12158 1970 2481 5.66e-16
c12159 2178 2253 1.96e-16
c12160 3886 647 3.15e-16
c12161 2934 1 1.257e-15
c12162 1203 842 1.58e-16
c12163 2895 0 3.7361e-14
c12164 4219 4208 3.84e-16
c12165 4223 4224 6.67e-16
c12166 2535 2339 1.58e-16
c12167 1533 737 1.58e-16
c12168 1027 1 3.54e-16
c12169 3650 4492 2.38e-15
c12170 4310 4299 1.58e-16
c12171 1024 0 9.602e-15
c12172 4620 1 1.013e-15
c12173 3393 3404 1.96e-16
c12174 117 114 3.54e-16
c12175 19 494 3.84e-16
c12176 5068 5071 3.54e-16
c12177 5086 5034 1.141e-15
c12178 2182 2253 4.63e-16
c12179 2036 1 4.083e-15
c12180 3915 3909 1.96e-16
c12181 1652 0 5.7033e-14
c12182 1132 782 6.38e-16
c12183 113 19 3.45e-16
c12184 59 455 1.88e-16
c12185 102 27 1.88e-16
c12186 2578 2569 3.92e-16
c12187 2169 2572 5.66e-16
c12188 1422 996 2.48e-16
c12189 911 1317 1.88e-16
c12190 657 4311 2.65e-16
c12191 4037 19 9.67e-16
c12192 2355 732 2.4e-16
c12193 957 1 5.821e-15
c12194 4421 1 5.808e-15
c12195 4423 0 3.466e-15
c12196 3588 777 5.73e-16
c12197 3420 3021 2.48e-16
c12198 2987 2041 4.35e-16
c12199 601 2236 1.58e-16
c12200 246 262 3.84e-16
c12201 249 250 6.67e-16
c12202 3343 868 2.4e-16
c12203 2273 2275 2.03e-16
c12204 88 508 1.88e-16
c12205 276 136 1.88e-16
c12206 223 479 1.88e-16
c12207 2552 2540 3.225e-15
c12208 4770 4765 1.536e-15
c12209 4571 4877 3.92e-16
c12210 2493 1 1.716e-15
c12211 596 742 3.134e-15
c12212 4004 4008 3.84e-16
c12213 4012 4011 4.41e-16
c12214 4804 5262 7.46e-16
c12215 687 1028 1.58e-16
c12216 1204 1205 7.51e-16
c12217 4301 4303 2.03e-16
c12218 1136 1559 1.58e-16
c12219 910 1343 1.014e-15
c12220 911 1321 1.88e-16
c12221 4214 4197 1.083e-15
c12222 1850 1849 9.1e-16
c12223 3310 0 3.6368e-14
c12224 1871 0 3.3874e-14
c12225 3409 3570 3.92e-16
c12226 953 954 7.46e-16
c12227 5173 5182 1.96e-16
c12228 4770 265 1.88e-16
c12229 143 145 7.1e-16
c12230 4317 3486 3.92e-16
c12231 3571 737 2.33e-16
c12232 5469 5447 6.67e-16
c12233 1192 1173 1.546e-15
c12234 910 941 2.19e-16
c12235 919 1010 3.92e-16
c12236 922 1009 2.54e-16
c12237 3886 3885 1.357e-15
c12238 3447 1 1.868e-15
c12239 3437 0 2.93e-15
c12240 2535 2854 3.92e-16
c12241 3515 3123 1.96e-16
c12242 4846 4845 2.03e-16
c12243 3154 662 4.81e-16
c12244 117 305 1.88e-16
c12245 2196 2388 5.42e-16
c12246 5412 439 1.58e-16
c12247 1862 2355 1.96e-16
c12248 1426 647 1.58e-16
c12249 1423 672 1.58e-16
c12250 827 837 3.28e-16
c12251 408 410 6.01e-16
c12252 2810 2424 5.66e-16
c12253 2637 2635 1.862e-15
c12254 632 625 5.58e-16
c12255 2048 2031 1.541e-15
c12256 2557 2836 1.58e-16
c12257 2541 2824 1.58e-16
c12258 1151 1128 6.54e-16
c12259 1331 1181 5.5e-16
c12260 4385 1 1.716e-15
c12261 687 2304 2.4e-16
c12262 1684 1764 1.58e-16
c12263 1706 1752 1.58e-16
c12264 1682 1683 3.36e-16
c12265 336 337 6.67e-16
c12266 2367 2362 1.642e-15
c12267 3839 1 4.161e-15
c12268 2257 2255 1.862e-15
c12269 1749 1743 1.418e-15
c12270 595 2192 2.13e-16
c12271 1760 1732 2.64e-16
c12272 418 1 4.59e-16
c12273 215 233 1.58e-16
c12274 404 19 8.4e-16
c12275 412 0 5.7592e-14
c12276 4787 33 1.88e-16
c12277 596 697 3.134e-15
c12278 632 3100 3.15e-16
c12279 657 3083 1.58e-16
c12280 3229 0 6.62e-16
c12281 3537 4373 5.66e-16
c12282 4379 4370 3.92e-16
c12283 4481 812 7.68e-16
c12284 1811 702 1.813e-15
c12285 750 1 1.65e-16
c12286 3594 1 2.054e-15
c12287 1557 1106 1.532e-15
c12288 1563 1562 5.65e-16
c12289 4628 4626 2.15e-16
c12290 4624 4635 1.96e-16
c12291 4183 1 4.45e-16
c12292 2194 837 3.15e-16
c12293 762 596 1.96e-16
c12294 4571 842 1.33e-16
c12295 4913 4897 9.43e-16
c12296 3296 3308 2.32e-16
c12297 3034 2702 1.58e-16
c12298 3409 3506 1.58e-16
c12299 3662 3669 6.73e-16
c12300 4344 1 6.275e-15
c12301 2713 732 3.79e-16
c12302 2164 2162 1.6e-16
c12303 1037 662 1.58e-16
c12304 1 61 4.92e-16
c12305 4844 4852 1.81e-16
c12306 4582 4463 5.5e-16
c12307 0 50 1.0822e-14
c12308 45 51 1.372e-15
c12309 4036 857 1.88e-16
c12310 2432 2429 3.01e-16
c12311 2428 2425 6.44e-16
c12312 2178 1834 1.58e-16
c12313 642 647 2.77e-16
c12314 4389 722 1.9e-16
c12315 2559 2435 5.5e-16
c12316 2705 2333 1.58e-16
c12317 1001 1005 2.03e-16
c12318 1694 647 3.15e-16
c12319 1345 1452 5.42e-16
c12320 1321 1440 1.58e-16
c12321 3882 4523 1.58e-16
c12322 3898 4535 1.58e-16
c12323 2880 2905 7.65e-16
c12324 1103 0 1.4198e-14
c12325 926 1 1.503e-15
c12326 3991 1 4.45e-16
c12327 1735 1742 1.96e-16
c12328 2106 2148 1.57e-15
c12329 2137 1667 2.241e-15
c12330 3701 1 5.343e-15
c12331 4710 4709 2.03e-16
c12332 2559 752 3.15e-16
c12333 9 563 3.92e-16
c12334 304 305 1.88e-16
c12335 4582 4626 1.58e-16
c12336 2182 1834 1.58e-16
c12337 2267 1 9.28e-16
c12338 3338 3344 1.545e-15
c12339 2790 1 5.808e-15
c12340 2342 2351 3.92e-16
c12341 1845 2337 1.58e-16
c12342 62 33 1.88e-16
c12343 5410 5421 1.37e-16
c12344 2703 2714 1.96e-16
c12345 2792 0 3.466e-15
c12346 2629 1 1.868e-15
c12347 1465 717 1.813e-15
c12348 2679 1 5.97e-15
c12349 1402 971 1.96e-16
c12350 3886 3497 5.5e-16
c12351 3286 2764 1.96e-16
c12352 3942 19 7.04e-16
c12353 3957 0 1.5176e-14
c12354 2685 3193 2.48e-16
c12355 2850 827 3.64e-16
c12356 1684 1505 1.58e-16
c12357 1690 1499 5.88e-16
c12358 612 1319 1.813e-15
c12359 1460 1 2.054e-15
c12360 3114 3111 3.01e-16
c12361 1462 0 8e-16
c12362 3490 3488 2.03e-16
c12363 3576 737 5.03e-16
c12364 5139 31 3.54e-16
c12365 3296 797 1.832e-15
c12366 3034 722 3.15e-16
c12367 1601 0 6.9087e-14
c12368 894 888 1.58e-16
c12369 909 898 5.5e-16
c12370 3253 3651 4.36e-16
c12371 1343 707 4.46e-16
c12372 1331 717 7.99e-16
c12373 1379 881 1.96e-16
c12374 1374 952 1.96e-16
c12375 3969 3966 3.43e-16
c12376 2557 2599 3.92e-16
c12377 657 1343 3.15e-16
c12378 3564 1 8.43e-16
c12379 894 1 3.679e-15
c12380 2765 767 7.68e-16
c12381 1908 1905 5.5e-16
c12382 1706 1705 1.009e-15
c12383 1690 1695 8.56e-16
c12384 2680 677 3.64e-16
c12385 2892 2894 1.062e-15
c12386 2244 2242 1.6e-16
c12387 2239 2238 2.03e-16
c12388 3411 3489 1.58e-16
c12389 3397 3502 4.63e-16
c12390 4412 4805 1.914e-15
c12391 2402 1 1.868e-15
c12392 1641 2078 1.958e-15
c12393 647 997 6.38e-16
c12394 9 535 5.8e-16
c12395 4776 4779 6.02e-16
c12396 4580 4792 3.92e-16
c12397 0 560 2.87e-16
c12398 448 447 1.482e-15
c12399 3253 797 1.58e-16
c12400 4567 4604 1.58e-16
c12401 5481 0 3.6193e-14
c12402 4922 497 1.88e-16
c12403 2392 0 2.93e-15
c12404 3531 3526 1.642e-15
c12405 3898 717 3.15e-16
c12406 627 3094 2.72e-16
c12407 919 1068 1.58e-16
c12408 2305 2690 1.96e-16
c12409 1922 782 1.58e-16
c12410 392 165 1.88e-16
c12411 687 1457 1.58e-16
c12412 3587 747 2.4e-16
c12413 2955 2994 1.738e-15
c12414 2452 842 1.58e-16
c12415 601 1353 1.339e-15
c12416 852 19 1.41e-15
c12417 3379 3377 1.6e-16
c12418 2747 3264 4.11e-16
c12419 3034 3156 4.63e-16
c12420 747 1102 1.58e-16
c12421 4791 4792 8.22e-16
c12422 2196 1687 3.54e-16
c12423 4293 0 6.8896e-14
c12424 1992 1988 1.96e-16
c12425 309 320 3.84e-16
c12426 324 321 6.67e-16
c12427 513 565 1.88e-16
c12428 885 884 4.16e-16
c12429 3783 3775 3.54e-16
c12430 566 570 1.58e-16
c12431 909 1053 3.54e-16
c12432 966 967 8.58e-16
c12433 3384 4237 5.66e-16
c12434 4243 4234 3.92e-16
c12435 2858 2503 1.58e-16
c12436 3345 1 1.716e-15
c12437 1438 1011 3.92e-16
c12438 1442 1443 1.6e-16
c12439 406 404 7.1e-16
c12440 361 407 1.88e-16
c12441 3907 1 2.625e-15
c12442 3898 4298 3.92e-16
c12443 537 88 1.88e-16
c12444 3818 0 2.078e-15
c12445 3160 3172 2.32e-16
c12446 1430 1 8.43e-16
c12447 5074 5113 1.858e-15
c12448 3466 3464 1.6e-16
c12449 3639 0 3.6368e-14
c12450 360 368 1.58e-16
c12451 4945 4946 6.26e-16
c12452 4469 4847 7.84e-16
c12453 3736 3734 1.001e-15
c12454 5207 5205 3.92e-16
c12455 5580 5575 2.029e-15
c12456 5403 5497 5.82e-16
c12457 2617 0 3.5252e-14
c12458 2559 2549 5.5e-16
c12459 843 0 7.86e-15
c12460 660 1 1.65e-16
c12461 4320 4317 6.44e-16
c12462 4324 4321 3.01e-16
c12463 1667 1196 9.7e-16
c12464 1193 1 4.59e-16
c12465 1190 0 1.0077e-14
c12466 3397 3438 1.58e-16
c12467 3409 782 4.46e-16
c12468 4623 4626 6.02e-16
c12469 3876 677 4.48e-16
c12470 5486 5481 5.63e-16
c12471 5450 5504 9.34e-16
c12472 1223 858 2.03e-16
c12473 1203 1209 1.58e-16
c12474 2944 0 2.28e-15
c12475 921 1055 1.96e-16
c12476 1534 1086 1.96e-16
c12477 1535 1528 6.73e-16
c12478 1345 971 5.5e-16
c12479 1321 957 5.5e-16
c12480 4091 1 6.78e-16
c12481 2442 812 1.339e-15
c12482 4080 0 1.01356e-13
c12483 4637 1 1.013e-15
c12484 2730 3241 1.96e-16
c12485 3048 2600 1.58e-16
c12486 3046 2594 5.5e-16
c12487 3034 3121 1.58e-16
c12488 2060 2062 6.91e-16
c12489 1569 1 9.28e-16
c12490 3409 3394 1.632e-15
c12491 3533 3526 6.73e-16
c12492 3532 3140 1.96e-16
c12493 5259 1 1.81e-16
c12494 2350 0 6.9484e-14
c12495 1635 1 5.343e-15
c12496 3772 3775 9.03e-16
c12497 5492 5489 3.92e-16
c12498 5452 5494 1.017e-15
c12499 2150 0 3.26e-15
c12500 595 3044 2.13e-16
c12501 2856 2469 1.532e-15
c12502 2923 2970 3.18e-16
c12503 1612 827 5.03e-16
c12504 3279 0 3.3874e-14
c12505 3858 1 1.871e-15
c12506 3370 0 5.549e-14
c12507 4441 1 2.054e-15
c12508 4676 4293 4.97e-16
c12509 4679 4675 1.96e-16
c12510 2541 647 3.15e-16
c12511 291 484 1.88e-16
c12512 4443 0 8e-16
c12513 3140 702 5.73e-16
c12514 4447 777 2.65e-16
c12515 4940 4942 3.25e-16
c12516 5291 352 3.94e-16
c12517 3046 807 3.15e-16
c12518 617 2236 7.38e-16
c12519 3381 3382 1.76e-16
c12520 4571 4894 3.92e-16
c12521 4878 1 3.4618e-14
c12522 4872 468 1.88e-16
c12523 2866 3048 3.92e-16
c12524 2519 1 5.01e-16
c12525 1057 1038 1.546e-15
c12526 5587 0 1.2414e-14
c12527 4634 497 1.88e-16
c12528 3900 3381 1.58e-16
c12529 3650 827 1.58e-16
c12530 5561 5422 4.35e-16
c12531 2541 2492 1.58e-16
c12532 615 1 1.65e-16
c12533 3236 0 6.9194e-14
c12534 3057 2532 2.48e-16
c12535 2718 722 7.38e-16
c12536 1856 1852 1.96e-16
c12537 5013 3744 1.98e-16
c12538 4546 4978 2.206e-15
c12539 2987 2984 7.46e-16
c12540 3030 2736 1.58e-16
c12541 1891 0 1.4092e-14
c12542 2173 2175 1.578e-15
c12543 2188 2181 7.06e-16
c12544 468 0 1.24974e-13
c12545 4861 4480 5.2e-16
c12546 1 498 4.92e-16
c12547 3219 3603 1.58e-16
c12548 3387 752 4.48e-16
c12549 4742 526 1.88e-16
c12550 4838 178 1.88e-16
c12551 2468 1947 1.96e-16
c12552 2463 1953 1.96e-16
c12553 2457 822 2.4e-16
c12554 165 276 1.88e-16
c12555 2172 2218 1.58e-16
c12556 2194 2206 1.58e-16
c12557 107 1 8.25e-15
c12558 3801 3817 9.55e-16
c12559 3565 752 1.58e-16
c12560 1212 842 4.98e-16
c12561 1706 717 3.15e-16
c12562 3630 0 8e-16
c12563 3066 1 5.97e-15
c12564 528 30 3.84e-16
c12565 632 1419 1.58e-16
c12566 2559 2871 3.92e-16
c12567 595 921 1.089e-15
c12568 3886 4400 4.63e-16
c12569 4474 3633 4.11e-16
c12570 1769 1772 5.5e-16
c12571 4761 0 2.93e-15
c12572 1690 1952 1.96e-16
c12573 4563 4707 1.96e-16
c12574 4691 4316 4.9e-16
c12575 2293 0 3.466e-15
c12576 3828 3821 3.92e-16
c12577 5303 352 1.58e-16
c12578 5212 1 1.257e-15
c12579 5032 5043 1.37e-16
c12580 2196 1678 1.58e-16
c12581 907 807 3.15e-16
c12582 1749 2257 7.84e-16
c12583 1328 898 2.035e-15
c12584 3972 1338 1.96e-16
c12585 4188 4182 1.96e-16
c12586 4225 3918 6.32e-16
c12587 4600 5514 1.96e-16
c12588 3034 822 7.99e-16
c12589 2535 2853 1.58e-16
c12590 2557 2841 1.58e-16
c12591 1612 812 1.9e-16
c12592 3898 3554 1.58e-16
c12593 4006 37 1.88e-16
c12594 2545 2666 1.58e-16
c12595 1674 1661 3.92e-16
c12596 1335 1 8.822e-15
c12597 3128 2611 4.11e-16
c12598 3504 3507 6.44e-16
c12599 1938 1939 2.48e-16
c12600 1708 1781 5.42e-16
c12601 1684 1769 1.58e-16
c12602 3511 662 1.09e-16
c12603 3024 767 4.48e-16
c12604 612 2206 1.58e-16
c12605 4844 5034 2.45e-16
c12606 3397 3168 5.5e-16
c12607 3679 3676 5.5e-16
c12608 2866 3347 1.58e-16
c12609 2458 1 4.41e-15
c12610 2653 0 2.93e-15
c12611 279 0 9.795e-15
c12612 2751 2367 1.58e-16
c12613 3065 1 8.43e-16
c12614 1270 1272 5.5e-16
c12615 3650 812 3.15e-16
c12616 4804 149 7.84e-16
c12617 3124 3127 6.44e-16
c12618 4205 1 4.64e-16
c12619 5403 528 3.54e-16
c12620 777 592 5.8e-16
c12621 3231 737 1.58e-16
c12622 216 37 1.88e-16
c12623 602 2580 4.81e-16
c12624 792 2427 1.58e-16
c12625 2194 1851 1.58e-16
c12626 162 1 4.22e-16
c12627 3996 3990 1.96e-16
c12628 922 782 5.14e-16
c12629 921 1113 1.58e-16
c12630 151 0 5.5422e-14
c12631 2725 2333 2.38e-15
c12632 1684 677 4.48e-16
c12633 1345 1457 1.58e-16
c12634 719 25 1.13e-15
c12635 3125 3127 2.03e-16
c12636 534 552 1.58e-16
c12637 1487 1046 1.96e-16
c12638 4540 3900 3.25e-16
c12639 2299 692 3.15e-16
c12640 2690 702 2.72e-16
c12641 2495 868 1.58e-16
c12642 617 1389 1.832e-15
c12643 2920 2918 1.462e-15
c12644 2787 3305 1.96e-16
c12645 3299 3306 6.73e-16
c12646 762 767 2.77e-16
c12647 2005 2016 1.96e-16
c12648 4582 4643 1.58e-16
c12649 5154 5155 3.54e-16
c12650 447 449 2.84e-16
c12651 338 349 3.84e-16
c12652 3202 737 3.15e-16
c12653 5291 294 4.02e-16
c12654 2342 1845 1.58e-16
c12655 1179 837 1.58e-16
c12656 883 767 6.45e-16
c12657 909 1127 4.35e-16
c12658 907 1126 1.88e-16
c12659 890 1119 1.58e-16
c12660 4651 1 1.1647e-14
c12661 2799 792 2.65e-16
c12662 1041 1474 7.84e-16
c12663 4171 3918 8.1e-16
c12664 3222 1 1.056e-15
c12665 888 1 4.226e-15
c12666 3979 1 6.66e-16
c12667 2401 767 3.15e-16
c12668 1742 1733 3.46e-16
c12669 905 0 1.0868e-14
c12670 2867 868 2.65e-16
c12671 1708 1522 1.58e-16
c12672 1706 1516 5.5e-16
c12673 1694 1917 1.58e-16
c12674 627 1319 1.58e-16
c12675 1478 0 6.72e-16
c12676 747 1061 1.58e-16
c12677 3596 737 1.09e-16
c12678 2340 2351 1.96e-16
c12679 3387 3689 3.92e-16
c12680 7 0 8.958e-15
c12681 4787 526 1.88e-16
c12682 2172 2495 1.58e-16
c12683 1401 971 1.58e-16
c12684 4872 64 1.88e-16
c12685 2535 2616 3.92e-16
c12686 701 1 5.57e-16
c12687 4355 3520 1.96e-16
c12688 4360 3514 1.96e-16
c12689 1343 1605 1.58e-16
c12690 1327 1593 1.58e-16
c12691 4605 3874 1.96e-16
c12692 4873 1 1.749e-15
c12693 1743 2236 1.96e-16
c12694 1809 1 6.15e-16
c12695 4865 0 7.67e-16
c12696 4580 4809 3.92e-16
c12697 5240 5198 3.15e-16
c12698 0 517 6.224e-15
c12699 3670 797 4.81e-16
c12700 4468 782 1.58e-16
c12701 2887 1 4.083e-15
c12702 1246 1245 6.34e-16
c12703 642 984 1.58e-16
c12704 64 0 2.67409e-13
c12705 59 45 1.58e-16
c12706 4383 707 1.58e-16
c12707 1942 782 1.58e-16
c12708 1545 1542 5.5e-16
c12709 3873 4595 5.66e-16
c12710 4601 4592 3.92e-16
c12711 3540 0 3.3874e-14
c12712 4151 1 4.45e-16
c12713 2667 662 1.58e-16
c12714 1802 1803 2.48e-16
c12715 3752 0 1.7153e-14
c12716 4480 4486 9.42e-16
c12717 4418 4795 2.48e-16
c12718 3100 3095 1.642e-15
c12719 3409 3134 5.5e-16
c12720 4310 0 6.8946e-14
c12721 5252 5251 1.6e-16
c12722 523 508 1.88e-16
c12723 30 325 3.84e-16
c12724 3393 672 4.03e-16
c12725 3557 3569 2.32e-16
c12726 5324 323 5.5e-16
c12727 627 3088 2.4e-16
c12728 2780 1 8.43e-16
c12729 894 1068 3.54e-16
c12730 3385 4234 1.58e-16
c12731 3537 717 1.58e-16
c12732 5407 5404 1.075e-15
c12733 2693 2690 3.01e-16
c12734 2689 2686 6.44e-16
c12735 5325 5321 3.54e-16
c12736 1331 842 3.15e-16
c12737 1191 852 5.73e-16
c12738 1355 957 1.58e-16
c12739 602 4245 4.81e-16
c12740 4423 4424 1.6e-16
c12741 4419 3588 3.92e-16
c12742 1708 1324 3.54e-16
c12743 717 26 1.58e-16
c12744 1629 1625 1.96e-16
c12745 535 540 1.482e-15
c12746 1965 1 1.868e-15
c12747 1955 0 2.93e-15
c12748 107 363 1.88e-16
c12749 3387 3625 1.58e-16
c12750 3411 3637 5.42e-16
c12751 3393 3242 1.58e-16
c12752 1073 722 1.58e-16
c12753 2169 0 4.4783e-14
c12754 1568 767 3.64e-16
c12755 3886 868 7.99e-16
c12756 3898 842 4.46e-16
c12757 2535 2581 1.58e-16
c12758 2557 2569 1.58e-16
c12759 601 968 3.57e-16
c12760 1777 677 1.58e-16
c12761 911 1319 1.88e-16
c12762 3463 1 5.97e-15
c12763 3103 3101 1.6e-16
c12764 1898 1897 1.6e-16
c12765 1890 1888 2.15e-16
c12766 1215 1 3.06e-16
c12767 407 455 1.88e-16
c12768 4563 4367 1.58e-16
c12769 4742 4749 1.81e-16
c12770 392 291 1.88e-16
c12771 3927 3928 6.4e-16
c12772 1476 692 1.9e-16
c12773 2857 2475 2.48e-16
c12774 1327 1385 1.96e-16
c12775 629 25 1.13e-15
c12776 633 19 1.58e-16
c12777 4516 4509 6.73e-16
c12778 4515 3673 1.96e-16
c12779 4654 1 1.013e-15
c12780 3177 702 1.58e-16
c12781 1694 1618 5.5e-16
c12782 1363 0 6.9108e-14
c12783 1582 1 6.15e-16
c12784 3151 3140 1.58e-16
c12785 1972 1974 2.03e-16
c12786 0 451 1.051e-14
c12787 19 429 8.82e-16
c12788 4563 4576 6.67e-16
c12789 4582 4215 3.54e-16
c12790 920 702 3.15e-16
c12791 957 955 1.988e-15
c12792 107 131 1.88e-16
c12793 2722 0 3.3717e-14
c12794 3505 0 2.93e-15
c12795 3006 2929 8.32e-16
c12796 1166 842 1.58e-16
c12797 1632 827 1.09e-16
c12798 1449 1001 4.36e-16
c12799 3299 0 1.4092e-14
c12800 2545 2735 4.63e-16
c12801 1693 1695 3.84e-16
c12802 2535 662 4.48e-16
c12803 1954 1956 1.862e-15
c12804 1567 1573 1.418e-15
c12805 334 204 1.88e-16
c12806 175 172 3.54e-16
c12807 3549 702 2.65e-16
c12808 3599 792 1.58e-16
c12809 3437 3022 4.97e-16
c12810 2147 0 1.65e-16
c12811 868 866 3.327e-15
c12812 1806 662 1.58e-16
c12813 1423 1435 2.32e-16
c12814 3277 0 1.6491e-14
c12815 2178 2406 1.96e-16
c12816 4517 827 4.81e-16
c12817 3667 868 1.58e-16
c12818 2541 2316 5.88e-16
c12819 2359 732 1.58e-16
c12820 1249 1248 1.58e-16
c12821 3113 0 6.72e-16
c12822 919 1189 1.58e-16
c12823 794 26 2.65e-15
c12824 4318 3480 4.97e-16
c12825 1370 0 1.6491e-14
c12826 262 256 1.58e-16
c12827 247 252 1.88e-16
c12828 3421 3433 2.32e-16
c12829 2285 2283 1.6e-16
c12830 3046 2753 1.58e-16
c12831 2189 2177 3.225e-15
c12832 2179 2175 2.074e-15
c12833 233 479 1.88e-16
c12834 4589 4591 4.93e-16
c12835 2495 0 3.3605e-14
c12836 2182 2406 4.63e-16
c12837 2196 762 3.58e-16
c12838 2172 2223 1.58e-16
c12839 919 837 3.15e-16
c12840 4313 4311 1.6e-16
c12841 3599 737 1.58e-16
c12842 4432 752 4.81e-16
c12843 3003 2492 1.361e-15
c12844 3483 1 1.056e-15
c12845 1515 1506 3.46e-16
c12846 1345 1344 1.866e-15
c12847 2316 732 1.58e-16
c12848 822 596 1.96e-16
c12849 2921 2880 5.71e-16
c12850 1149 0 2.7376e-14
c12851 3384 0 4.4783e-14
c12852 2407 797 1.75e-16
c12853 1573 1574 1.35e-16
c12854 4778 0 2.93e-15
c12855 3237 3231 1.6e-16
c12856 2713 3228 2.386e-15
c12857 2730 3211 1.58e-16
c12858 2045 2049 6.35e-16
c12859 1706 1969 3.92e-16
c12860 1 363 2.3e-14
c12861 426 262 1.88e-16
c12862 3704 827 4.81e-16
c12863 3304 868 1.58e-16
c12864 3513 3504 3.46e-16
c12865 2313 0 8e-16
c12866 5424 0 1.65e-16
c12867 5450 439 5.5e-16
c12868 657 2617 1.58e-16
c12869 747 1851 5.73e-16
c12870 5221 0 2.285e-15
c12871 281 279 1.257e-15
c12872 1130 767 5.74e-16
c12873 1166 1170 2.03e-16
c12874 2559 2870 5.42e-16
c12875 2535 2858 1.58e-16
c12876 4293 3452 1.136e-15
c12877 3633 4468 1.96e-16
c12878 1380 1778 4.36e-16
c12879 2545 2671 1.58e-16
c12880 963 0 4.4793e-14
c12881 2719 3226 3.92e-16
c12882 3231 3230 1.6e-16
c12883 1076 0 7.4292e-14
c12884 19 256 3.2e-16
c12885 1862 2359 1.58e-16
c12886 3534 677 4.81e-16
c12887 4950 1 4.159e-15
c12888 612 2226 1.58e-16
c12889 890 1007 1.96e-16
c12890 4580 4469 1.58e-16
c12891 4855 120 1.88e-16
c12892 1784 662 1.339e-15
c12893 1606 812 7.38e-16
c12894 4031 3918 8.1e-16
c12895 4673 662 1.23e-16
c12896 5536 5551 1.37e-16
c12897 1293 1295 9.5e-16
c12898 2350 707 1.58e-16
c12899 1706 842 4.46e-16
c12900 1694 868 7.99e-16
c12901 642 1386 1.58e-16
c12902 632 1761 7.68e-16
c12903 1321 1657 3.92e-16
c12904 3225 1 4.41e-15
c12905 2739 2751 2.32e-16
c12906 1575 1576 2.48e-16
c12907 749 26 2.65e-15
c12908 1317 1 2.346e-15
c12909 3522 3134 4.97e-16
c12910 4645 4643 2.15e-16
c12911 4641 4652 1.96e-16
c12912 1694 1386 1.58e-16
c12913 4387 0 3.3724e-14
c12914 1836 1838 2.03e-16
c12915 1332 0 1.157e-14
c12916 595 2208 2.72e-16
c12917 612 2204 1.58e-16
c12918 1854 1 5.808e-15
c12919 3316 3313 5.5e-16
c12920 1856 0 3.466e-15
c12921 3676 3683 1.96e-16
c12922 4755 1 8.85e-16
c12923 827 821 1.74e-16
c12924 276 291 1.88e-16
c12925 1 131 8.25e-15
c12926 9 132 4.88e-16
c12927 122 0 5.8334e-14
c12928 136 27 1.88e-16
c12929 3589 3202 1.532e-15
c12930 2459 0 1.6491e-14
c12931 2440 1930 1.96e-16
c12932 5540 5543 1.96e-16
c12933 4759 381 1.88e-16
c12934 1327 898 3.15e-16
c12935 1251 1289 1.6e-16
c12936 1959 807 1.58e-16
c12937 1327 1041 1.58e-16
c12938 910 905 1.58e-16
c12939 146 142 1.58e-16
c12940 537 523 1.88e-16
c12941 2503 852 3.15e-16
c12942 1818 1820 1.862e-15
c12943 1431 1437 1.418e-15
c12944 1752 1754 2.15e-16
c12945 777 1126 1.35e-16
c12946 2787 2798 1.58e-16
c12947 3030 3224 1.96e-16
c12948 1321 1 3.564e-15
c12949 2151 1708 3.25e-16
c12950 76 71 1.482e-15
c12951 4727 4726 2.03e-16
c12952 33 30 7.67e-16
c12953 3202 3590 4.97e-16
c12954 4582 4660 1.58e-16
c12955 1919 2427 7.84e-16
c12956 642 2172 3.15e-16
c12957 632 3114 1.09e-16
c12958 894 1142 3.92e-16
c12959 909 1141 1.88e-16
c12960 883 1134 1.58e-16
c12961 2729 2333 1.96e-16
c12962 922 923 3.15e-16
c12963 4171 4166 1.96e-16
c12964 3405 1 1.002e-15
c12965 3025 3027 1.578e-15
c12966 3040 3033 7.06e-16
c12967 1852 732 1.58e-16
c12968 1046 1486 1.58e-16
c12969 4166 37 1.88e-16
c12970 3616 4450 1.58e-16
c12971 3298 2781 4.11e-16
c12972 2696 3210 4.97e-16
c12973 1642 1653 1.96e-16
c12974 3718 3900 3.92e-16
c12975 2628 677 1.58e-16
c12976 2858 858 1.58e-16
c12977 3886 0 3.3139e-13
c12978 0 585 1.4515e-14
c12979 334 175 1.88e-16
c12980 227 1 2.87e-16
c12981 3706 842 7.38e-16
c12982 2634 1 4.41e-15
c12983 1111 1112 1.238e-15
c12984 883 931 1.58e-16
c12985 894 955 1.58e-16
c12986 4164 4168 3.84e-16
c12987 230 26 1.03e-15
c12988 1406 971 2.386e-15
c12989 2559 2633 3.92e-16
c12990 1218 921 1.58e-16
c12991 1321 1622 1.58e-16
c12992 1343 1610 1.58e-16
c12993 687 1343 3.15e-16
c12994 1755 1369 5.66e-16
c12995 704 26 2.65e-15
c12996 4242 4605 1.96e-16
c12997 2600 3109 7.84e-16
c12998 4351 0 1.6491e-14
c12999 573 574 1.58e-16
c13000 4890 1 1.786e-15
c13001 4429 4822 1.914e-15
c13002 3654 3655 9.1e-16
c13003 4882 0 7.67e-16
c13004 2420 1 9.28e-16
c13005 1 310 1.9313e-14
c13006 4580 4826 3.92e-16
c13007 5540 526 3.54e-16
c13008 2390 0 3.6368e-14
c13009 3918 3980 2.87e-16
c13010 3015 1 7.21e-16
c13011 2792 2793 1.6e-16
c13012 1046 722 1.58e-16
c13013 5432 5414 6.67e-16
c13014 3560 0 1.4092e-14
c13015 601 1374 1.9e-16
c13016 1068 1 1.56e-15
c13017 4526 4523 5.5e-16
c13018 1970 842 1.75e-16
c13019 4497 4486 1.58e-16
c13020 4808 4809 8.22e-16
c13021 3046 3172 1.58e-16
c13022 3030 3160 1.58e-16
c13023 1627 1 5.808e-15
c13024 1629 0 3.466e-15
c13025 910 2169 3.75e-16
c13026 448 455 7.76e-16
c13027 5314 1 1.88e-16
c13028 2223 0 3.3692e-14
c13029 1158 797 1.58e-16
c13030 3385 4254 2.38e-15
c13031 2603 2615 2.32e-16
c13032 1661 858 9.97e-16
c13033 1674 852 3.64e-16
c13034 1461 1460 5.65e-16
c13035 3934 1 6.76e-16
c13036 612 3385 1.813e-15
c13037 3180 3177 5.5e-16
c13038 117 450 1.88e-16
c13039 3667 0 6.9037e-14
c13040 566 580 1.58e-16
c13041 490 494 1.58e-16
c13042 3474 3475 1.6e-16
c13043 3470 3089 3.92e-16
c13044 5127 1 7.87e-16
c13045 2330 2327 3.01e-16
c13046 2326 2323 6.44e-16
c13047 1584 1 5.97e-15
c13048 4776 5219 3.92e-16
c13049 3411 3642 1.58e-16
c13050 3397 3655 4.63e-16
c13051 1095 722 6.48e-16
c13052 5323 5318 7.25e-16
c13053 4183 857 6.23e-16
c13054 4139 3918 8.1e-16
c13055 1121 767 3.15e-16
c13056 396 407 3.84e-16
c13057 101 103 1.58e-16
c13058 3898 4302 1.58e-16
c13059 3876 4314 1.58e-16
c13060 3900 858 3.15e-16
c13061 4540 852 2.8e-16
c13062 4770 381 1.88e-16
c13063 1240 920 6.34e-16
c13064 919 1238 3.54e-16
c13065 617 968 1.58e-16
c13066 3908 19 9.67e-16
c13067 4332 3497 1.96e-16
c13068 1624 858 1.75e-16
c13069 4412 4407 1.642e-15
c13070 1426 0 1.4092e-14
c13071 668 667 1.96e-16
c13072 3030 702 4.03e-16
c13073 2072 2078 1.572e-15
c13074 1 339 2.3e-14
c13075 230 187 1.88e-16
c13076 3393 797 3.15e-16
c13077 4563 4384 1.58e-16
c13078 2574 0 8e-16
c13079 3991 857 6.23e-16
c13080 3147 0 6.72e-16
c13081 1046 1050 2.03e-16
c13082 383 0 5.6832e-14
c13083 4438 782 1.58e-16
c13084 5482 5450 1.75e-16
c13085 3304 0 6.9097e-14
c13086 1343 1402 3.92e-16
c13087 2583 3091 2.48e-16
c13088 2979 2978 1.6e-16
c13089 842 26 7.12e-16
c13090 3030 2804 1.58e-16
c13091 2637 662 1.58e-16
c13092 822 1175 1.85e-16
c13093 4671 1 1.013e-15
c13094 3008 858 6.67e-16
c13095 2541 868 4.03e-16
c13096 2557 827 4.46e-16
c13097 2518 852 1.58e-16
c13098 2116 2115 1.6e-16
c13099 5197 5195 1.373e-15
c13100 3387 3451 3.92e-16
c13101 3547 3540 1.96e-16
c13102 3151 3549 4.36e-16
c13103 692 708 1.621e-15
c13104 702 706 2.19e-16
c13105 2392 1879 4.97e-16
c13106 2196 2269 5.42e-16
c13107 595 3067 2.65e-16
c13108 602 2532 2.33e-16
c13109 971 923 6.54e-16
c13110 2742 0 1.4092e-14
c13111 4075 25 4.68e-16
c13112 2356 737 2.33e-16
c13113 1691 1710 9.83e-16
c13114 2029 2093 1.6e-16
c13115 1609 1611 2.03e-16
c13116 3622 1 4.41e-15
c13117 642 0 2.86786e-13
c13118 4693 4310 4.97e-16
c13119 4696 4692 1.96e-16
c13120 320 321 7.03e-16
c13121 4456 0 6.62e-16
c13122 5074 5032 3.41e-16
c13123 3168 702 3.79e-16
c13124 3540 707 1.58e-16
c13125 5059 1 3.36e-16
c13126 1694 0 3.3139e-13
c13127 890 702 3.35e-16
c13128 3397 3620 1.58e-16
c13129 2720 0 1.6491e-14
c13130 2215 1681 1.96e-16
c13131 2216 2209 6.73e-16
c13132 1682 2191 2.79e-16
c13133 4821 4435 1.179e-15
c13134 4878 410 1.88e-16
c13135 2194 2423 3.92e-16
c13136 2015 2044 1.048e-15
c13137 3701 837 2.22e-16
c13138 2557 2333 5.5e-16
c13139 910 3384 3.75e-16
c13140 3860 0 8e-16
c13141 1992 842 5.03e-16
c13142 1591 1593 1.862e-15
c13143 1136 1146 1.418e-15
c13144 4196 4197 3.01e-15
c13145 4564 4215 5.8e-16
c13146 4975 4978 5.5e-16
c13147 3024 2770 1.58e-16
c13148 3393 3604 1.96e-16
c13149 3034 672 7.99e-16
c13150 4606 4614 1.81e-16
c13151 4708 0 3.37468e-13
c13152 5136 5104 1.58e-16
c13153 2480 1964 4.11e-16
c13154 3710 3387 1.58e-16
c13155 5582 5579 1.6e-16
c13156 5427 0 2.156e-15
c13157 2896 1 2.386e-15
c13158 1470 677 1.58e-16
c13159 595 925 7.51e-16
c13160 624 1 5.57e-16
c13161 3499 1 9.28e-16
c13162 3643 0 6.62e-16
c13163 1701 1324 1.159e-15
c13164 3058 3070 2.32e-16
c13165 1521 1520 9.1e-16
c13166 4496 4487 3.46e-16
c13167 2172 732 3.15e-16
c13168 4795 0 2.93e-15
c13169 2557 812 4.46e-16
c13170 2031 2058 2.84e-16
c13171 1 487 1.44e-16
c13172 15 483 6.58e-16
c13173 3611 3612 5.65e-16
c13174 2461 822 1.58e-16
c13175 2329 0 6.72e-16
c13176 1658 1 7.56e-16
c13177 3611 767 1.84e-16
c13178 3907 857 1.88e-16
c13179 5039 5036 1.96e-16
c13180 894 837 8.34e-16
c13181 94 1 5.62e-16
c13182 64 441 1.88e-16
c13183 2898 0 1.65e-16
c13184 2837 2469 1.96e-16
c13185 612 2557 3.15e-16
c13186 602 2559 3.15e-16
c13187 600 25 7.64e-16
c13188 1345 1320 2.38e-16
c13189 1321 1317 3.54e-16
c13190 3262 1 5.808e-15
c13191 1176 1183 7.95e-16
c13192 3886 4404 1.58e-16
c13193 3876 3565 5.5e-16
c13194 2921 2939 1.23e-16
c13195 2196 722 3.15e-16
c13196 3339 2821 1.96e-16
c13197 2753 777 1.58e-16
c13198 997 0 1.8851e-14
c13199 1706 1968 1.58e-16
c13200 1690 1956 1.58e-16
c13201 3397 792 7.99e-16
c13202 3150 3141 3.46e-16
c13203 1355 1 5.808e-15
c13204 2070 1 1.021e-15
c13205 672 674 5.59e-16
c13206 310 363 1.88e-16
c13207 5064 5075 6.73e-16
c13208 5068 5067 2.67e-16
c13209 4903 1 9.49e-15
c13210 2681 1 9.28e-16
c13211 883 1022 3.92e-16
c13212 890 1021 1.88e-16
c13213 3355 852 3.15e-16
c13214 986 981 1.58e-16
c13215 73 71 1.88e-16
c13216 4736 5389 2.137e-15
c13217 2151 852 2.8e-16
c13218 1708 858 3.15e-16
c13219 632 1380 3.15e-16
c13220 1345 1343 4.506e-15
c13221 1331 1504 4.63e-16
c13222 1365 1 9.28e-16
c13223 4228 1 4.2638e-14
c13224 3390 3392 1.041e-15
c13225 2178 858 3.15e-16
c13226 1874 1 2.054e-15
c13227 3315 827 5.03e-16
c13228 1876 0 8e-16
c13229 3393 3569 1.58e-16
c13230 4772 1 8.85e-16
c13231 2754 2367 1.532e-15
c13232 3397 737 3.15e-16
c13233 5581 0 6.72e-16
c13234 5173 5171 3.92e-16
c13235 2172 1862 5.5e-16
c13236 4012 4013 7.81e-16
c13237 2816 2810 1.6e-16
c13238 3061 0 1.4092e-14
c13239 5444 5442 8.35e-16
c13240 2742 2749 6.73e-16
c13241 1343 1056 1.58e-16
c13242 3142 2628 4.97e-16
c13243 3788 1 3.36e-16
c13244 910 3886 5.03e-16
c13245 2182 858 3.15e-16
c13246 4200 37 1.88e-16
c13247 4201 26 1.075e-15
c13248 3313 3320 1.96e-16
c13249 3683 3674 3.46e-16
c13250 3145 677 5.03e-16
c13251 2032 2033 5.87e-16
c13252 1 266 4.92e-16
c13253 4582 4677 1.58e-16
c13254 1930 2439 1.58e-16
c13255 0 248 1.051e-14
c13256 827 1177 6.38e-16
c13257 165 27 1.88e-16
c13258 5412 5425 1.138e-15
c13259 4651 410 7.67e-16
c13260 2825 0 6.62e-16
c13261 2248 2636 4.97e-16
c13262 2254 2265 1.58e-16
c13263 536 535 5.8e-16
c13264 3031 3027 2.074e-15
c13265 3029 3025 1.988e-15
c13266 1488 722 2.33e-16
c13267 1500 1494 1.6e-16
c13268 1046 1491 2.386e-15
c13269 632 1387 1.339e-15
c13270 4092 4099 7.81e-16
c13271 3633 4438 1.58e-16
c13272 2928 2929 2.123e-15
c13273 2419 767 3.64e-16
c13274 1754 1750 1.96e-16
c13275 955 1 2.506e-15
c13276 951 0 1.23e-16
c13277 3046 3043 1.58e-16
c13278 3024 3044 3.92e-16
c13279 334 349 1.88e-16
c13280 449 455 3.84e-16
c13281 339 363 1.88e-16
c13282 513 262 1.88e-16
c13283 3882 792 4.03e-16
c13284 5157 236 5.5e-16
c13285 2366 1845 1.96e-16
c13286 2361 1851 1.96e-16
c13287 4531 1 9.42e-16
c13288 410 1 3.36e-15
c13289 223 224 6.96e-16
c13290 88 218 1.88e-16
c13291 415 0 2.87e-16
c13292 4191 3918 8.1e-16
c13293 4821 0 3.27376e-13
c13294 4606 33 1.88e-16
c13295 3976 37 5.71e-16
c13296 4372 3531 4.11e-16
c13297 2327 692 1.9e-16
c13298 1635 837 2.22e-16
c13299 1345 1639 5.42e-16
c13300 1321 1627 1.58e-16
c13301 1454 1455 1.35e-16
c13302 4622 4242 1.96e-16
c13303 2771 782 1.339e-15
c13304 1550 1917 1.58e-16
c13305 1706 1731 3.92e-16
c13306 3489 662 1.58e-16
c13307 4889 4885 2.24e-16
c13308 3315 812 1.9e-16
c13309 17 27 3.54e-16
c13310 13 44 1.88e-16
c13311 4580 4843 3.92e-16
c13312 2433 1 6.15e-16
c13313 592 670 6.34e-16
c13314 3999 3918 8.1e-16
c13315 3882 737 3.15e-16
c13316 4455 807 1.58e-16
c13317 1076 707 3.57e-16
c13318 1218 1235 1.58e-16
c13319 632 998 3.57e-16
c13320 2541 0 3.63418e-13
c13321 1948 797 7.68e-16
c13322 4231 4612 5.66e-16
c13323 4618 4609 3.92e-16
c13324 617 1374 5.03e-16
c13325 1102 1 3.54e-16
c13326 3886 3684 5.5e-16
c13327 4150 26 4.48e-16
c13328 4879 4884 1.106e-15
c13329 4497 4503 9.42e-16
c13330 1099 0 9.602e-15
c13331 4435 4812 2.48e-16
c13332 3291 3292 9.1e-16
c13333 3024 3189 1.58e-16
c13334 3046 3177 1.58e-16
c13335 2143 2104 1.738e-15
c13336 5230 5251 6.16e-16
c13337 5232 5231 5.68e-16
c13338 3577 3574 5.5e-16
c13339 0 508 1.40183e-13
c13340 306 305 7.08e-16
c13341 294 296 1.96e-16
c13342 30 526 3.84e-16
c13343 2408 1896 1.532e-15
c13344 2414 2413 5.65e-16
c13345 2196 2338 3.92e-16
c13346 5331 0 1.4815e-14
c13347 2243 0 1.4092e-14
c13348 42 45 2.142e-15
c13349 3851 3847 1.243e-15
c13350 3355 3409 3.92e-16
c13351 4373 722 1.84e-16
c13352 2701 2316 1.96e-16
c13353 1177 812 1.58e-16
c13354 1158 1164 1.58e-16
c13355 1856 707 1.9e-16
c13356 1384 1385 9.1e-16
c13357 3965 1 6.78e-16
c13358 627 3385 1.58e-16
c13359 4442 4441 5.65e-16
c13360 4436 3599 1.532e-15
c13361 732 0 2.86553e-13
c13362 2557 2786 3.92e-16
c13363 2221 0 1.6491e-14
c13364 2001 1 1.056e-15
c13365 4776 5198 5.37e-16
c13366 3393 3270 5.88e-16
c13367 2776 0 1.4092e-14
c13368 2240 2252 2.32e-16
c13369 2541 2203 1.58e-16
c13370 617 990 6.48e-16
c13371 4325 1 6.15e-16
c13372 1903 1914 1.96e-16
c13373 1694 1689 1.58e-16
c13374 762 921 3.15e-16
c13375 4864 4866 2.15e-16
c13376 3024 717 3.15e-16
c13377 1 556 5.848e-15
c13378 4563 4401 1.58e-16
c13379 4787 207 1.88e-16
c13380 4922 468 1.88e-16
c13381 2590 0 6.72e-16
c13382 1981 2504 4.36e-16
c13383 2502 2495 1.96e-16
c13384 3937 3941 7.45e-16
c13385 3948 3950 2.239e-15
c13386 1487 717 2.4e-16
c13387 1056 1063 7.95e-16
c13388 3497 4331 1.58e-16
c13389 3886 707 3.15e-16
c13390 2283 662 7.68e-16
c13391 2545 2373 1.58e-16
c13392 2557 747 3.15e-16
c13393 919 1085 3.92e-16
c13394 922 1084 2.54e-16
c13395 3523 1 5.808e-15
c13396 3718 852 3.15e-16
c13397 595 3411 3.15e-16
c13398 602 3387 3.46e-16
c13399 3525 0 3.466e-15
c13400 657 3886 7.99e-16
c13401 2957 2954 7.84e-16
c13402 3046 2821 1.58e-16
c13403 2458 837 1.58e-16
c13404 2654 672 1.58e-16
c13405 910 1694 5.03e-16
c13406 4688 1 1.013e-15
c13407 2535 852 3.15e-16
c13408 453 454 2.84e-16
c13409 421 419 1.88e-16
c13410 479 465 1.88e-16
c13411 3411 3468 3.92e-16
c13412 2196 822 3.58e-16
c13413 1862 0 6.9481e-14
c13414 0 210 1.4515e-14
c13415 448 491 1.88e-16
c13416 3706 3411 3.92e-16
c13417 2196 2274 1.58e-16
c13418 4351 707 1.339e-15
c13419 601 2532 1.75e-16
c13420 595 2533 2.22e-16
c13421 2557 2384 5.5e-16
c13422 2299 2654 1.58e-16
c13423 4236 3381 4.11e-16
c13424 1343 1401 1.58e-16
c13425 1327 1389 1.58e-16
c13426 2170 2595 4.36e-16
c13427 1444 1442 1.6e-16
c13428 1439 1438 2.03e-16
c13429 528 499 3.75e-16
c13430 3882 4467 1.58e-16
c13431 857 1 3.2438e-14
c13432 4101 0 1.5061e-14
c13433 4103 19 3.45e-16
c13434 1684 2020 3.92e-16
c13435 3170 3169 1.6e-16
c13436 4481 1 1.868e-15
c13437 1984 1982 1.6e-16
c13438 1694 1833 4.63e-16
c13439 30 442 6.83e-16
c13440 4471 0 2.93e-15
c13441 4580 4577 1.58e-16
c13442 4571 4578 3.92e-16
c13443 4563 4570 1.58e-16
c13444 349 345 1.58e-16
c13445 3560 707 1.58e-16
c13446 4903 4950 2.801e-15
c13447 4936 4944 3.54e-16
c13448 2303 1794 1.58e-16
c13449 792 1690 4.03e-16
c13450 102 100 1.88e-16
c13451 113 114 6.4e-16
c13452 3693 3695 2.15e-16
c13453 883 717 3.15e-16
c13454 596 672 1.96e-16
c13455 1682 1681 1.58e-16
c13456 2170 2588 4.11e-16
c13457 2172 2440 3.92e-16
c13458 409 1 4.92e-16
c13459 392 13 1.88e-16
c13460 3733 3734 4.61e-16
c13461 3135 1 1.868e-15
c13462 2865 2856 3.46e-16
c13463 911 3385 1.88e-16
c13464 3886 3452 1.58e-16
c13465 2545 2534 1.58e-16
c13466 1802 1420 2.48e-16
c13467 4480 3639 1.136e-15
c13468 3441 3438 5.5e-16
c13469 632 2240 1.58e-16
c13470 3048 2787 1.58e-16
c13471 3034 3308 1.58e-16
c13472 3048 677 3.15e-16
c13473 1678 2208 4.11e-16
c13474 2591 2588 3.01e-16
c13475 2096 2095 1.6e-16
c13476 4151 857 6.23e-16
c13477 4623 4628 5.53e-16
c13478 2194 2422 1.58e-16
c13479 2178 2410 1.58e-16
c13480 5476 5486 1.125e-15
c13481 4787 5229 9.43e-16
c13482 1690 737 3.15e-16
c13483 3658 0 2.93e-15
c13484 837 1 4.1542e-14
c13485 1527 1523 1.96e-16
c13486 1345 1367 5.42e-16
c13487 1321 1355 1.58e-16
c13488 4084 1 6.78e-16
c13489 3429 0 6.9058e-14
c13490 2457 797 1.58e-16
c13491 1178 0 1.4198e-14
c13492 1319 1 5.277e-15
c13493 4812 0 2.93e-15
c13494 3397 3392 1.58e-16
c13495 3411 3414 1.6e-16
c13496 2182 2410 1.58e-16
c13497 596 593 2.45e-16
c13498 3525 3521 1.96e-16
c13499 3765 3775 1.021e-15
c13500 858 852 3.28e-16
c13501 5452 5412 2.45e-16
c13502 3887 3881 2.267e-15
c13503 2850 2458 1.96e-16
c13504 2705 1 5.808e-15
c13505 2657 2658 5.65e-16
c13506 627 2557 3.15e-16
c13507 601 2559 3.15e-16
c13508 4214 3890 9.72e-16
c13509 657 1426 1.58e-16
c13510 3282 1 2.054e-15
c13511 3900 3582 5.5e-16
c13512 2921 2966 3.18e-16
c13513 1796 1795 1.6e-16
c13514 1788 1786 2.15e-16
c13515 2832 2821 1.58e-16
c13516 4060 26 4.58e-16
c13517 1684 1985 1.58e-16
c13518 1706 1973 1.58e-16
c13519 1694 1798 1.58e-16
c13520 777 1542 1.58e-16
c13521 200 204 1.58e-16
c13522 198 187 2.45e-16
c13523 2385 1868 1.96e-16
c13524 2386 2379 6.73e-16
c13525 4977 4991 2.09e-15
c13526 3034 797 3.15e-16
c13527 2277 2278 5.65e-16
c13528 288 290 7.1e-16
c13529 4322 662 1.58e-16
c13530 2836 2469 1.58e-16
c13531 2694 1 6.15e-16
c13532 909 677 3.15e-16
c13533 883 1036 1.88e-16
c13534 907 1029 1.58e-16
c13535 5577 1 6.744e-15
c13536 4634 468 1.88e-16
c13537 3260 1 1.716e-15
c13538 1343 782 4.46e-16
c13539 5560 5561 5.5e-16
c13540 1336 1330 1.6e-16
c13541 4394 4387 1.96e-16
c13542 3548 4396 4.36e-16
c13543 1828 722 1.58e-16
c13544 3636 1 1.056e-15
c13545 4662 4660 2.15e-16
c13546 4658 4669 1.96e-16
c13547 2788 807 1.58e-16
c13548 601 2225 1.9e-16
c13549 4549 5018 3.54e-16
c13550 2815 842 1.58e-16
c13551 3335 827 1.09e-16
c13552 4789 1 8.85e-16
c13553 2730 752 3.15e-16
c13554 762 1516 1.813e-15
c13555 1892 0 6.72e-16
c13556 747 1533 2.22e-16
c13557 3393 3574 1.58e-16
c13558 3409 3191 1.58e-16
c13559 5177 5185 9.34e-16
c13560 5262 5184 1.58e-16
c13561 692 1052 1.58e-16
c13562 1043 702 1.58e-16
c13563 4101 4102 3.15e-16
c13564 910 3383 1.58e-16
c13565 1525 752 1.58e-16
c13566 1091 732 4.21e-16
c13567 1295 1239 2.323e-15
c13568 1299 1236 1.028e-15
c13569 919 1143 1.58e-16
c13570 4922 64 1.88e-16
c13571 1694 707 3.15e-16
c13572 537 0 1.63838e-13
c13573 3401 3404 2.109e-15
c13574 1848 1846 1.6e-16
c13575 657 1694 7.99e-16
c13576 4028 1 4.64e-16
c13577 3250 752 1.09e-16
c13578 3048 3241 3.92e-16
c13579 1700 0 5.86e-16
c13580 1 191 4.22e-16
c13581 117 26 8.41e-16
c13582 4024 3972 1.88e-16
c13583 4691 4695 1.81e-16
c13584 4582 4694 1.58e-16
c13585 2453 2447 1.6e-16
c13586 1930 2444 2.386e-15
c13587 1936 2452 1.136e-15
c13588 1947 2427 1.58e-16
c13589 378 450 1.88e-16
c13590 2850 1 1.868e-15
c13591 909 1128 3.54e-16
c13592 2840 0 2.93e-15
c13593 149 152 4.6e-16
c13594 3031 3029 8.67e-16
c13595 1482 737 1.58e-16
c13596 3800 410 2.51e-16
c13597 4606 5564 1.628e-15
c13598 1913 767 3.15e-16
c13599 3320 3311 3.46e-16
c13600 1663 1664 9.13e-16
c13601 1061 1 5.821e-15
c13602 4546 4554 4.06e-16
c13603 4584 1 2.86e-16
c13604 5 18 2.45e-16
c13605 49 43 3.84e-16
c13606 4566 0 1.5582e-14
c13607 762 1523 1.58e-16
c13608 2033 236 1.098e-15
c13609 3773 3807 1.75e-16
c13610 910 2541 7.97e-16
c13611 911 2557 9.54e-16
c13612 1098 1112 1.96e-16
c13613 275 9 6.48e-16
c13614 276 13 1.88e-16
c13615 5366 5365 1.559e-15
c13616 285 0 6.224e-15
c13617 5570 1 1.65e-16
c13618 1596 797 1.58e-16
c13619 1413 1404 3.46e-16
c13620 632 4277 7.68e-16
c13621 642 3452 1.58e-16
c13622 941 19 1.96e-16
c13623 4259 4622 1.96e-16
c13624 1533 1925 2.38e-15
c13625 1684 1748 3.92e-16
c13626 1281 0 1.8523e-14
c13627 3571 747 1.58e-16
c13628 3024 3380 3.54e-16
c13629 3046 3030 4.274e-15
c13630 4563 4299 1.58e-16
c13631 4446 4839 1.914e-15
c13632 4923 0 1.7122e-14
c13633 216 0 4.6186e-14
c13634 281 508 1.88e-16
c13635 3409 858 1.58e-16
c13636 4719 4714 1.536e-15
c13637 2442 1 1.716e-15
c13638 5536 526 1.96e-16
c13639 3876 752 4.48e-16
c13640 4475 807 1.58e-16
c13641 657 997 1.58e-16
c13642 921 1130 1.96e-16
c13643 1121 1554 1.58e-16
c13644 4242 4621 1.58e-16
c13645 617 1394 1.09e-16
c13646 4553 4540 3.92e-16
c13647 2506 842 4.81e-16
c13648 581 584 6.38e-16
c13649 4825 4826 8.22e-16
c13650 3224 737 7.38e-16
c13651 3048 3206 5.42e-16
c13652 3024 3194 1.58e-16
c13653 737 730 5.58e-16
c13654 19 314 3.2e-16
c13655 0 297 1.4515e-14
c13656 4810 439 1.88e-16
c13657 5434 5426 3.92e-16
c13658 3003 0 3.9045e-14
c13659 1177 1179 7.84e-16
c13660 632 3393 3.15e-16
c13661 4278 4271 6.73e-16
c13662 4277 3435 1.96e-16
c13663 2623 2620 5.5e-16
c13664 1473 1474 2.48e-16
c13665 617 610 5.58e-16
c13666 3975 1 6.03e-16
c13667 1734 1736 2.03e-16
c13668 4571 662 1.33e-16
c13669 3918 0 2.99058e-13
c13670 3718 3690 2.64e-16
c13671 2594 647 1.58e-16
c13672 291 570 1.88e-16
c13673 3493 3492 5.65e-16
c13674 3487 3100 1.532e-15
c13675 2338 1828 1.96e-16
c13676 642 3092 1.58e-16
c13677 5110 122 8.44e-16
c13678 10 1 4.22e-16
c13679 4606 526 1.88e-16
c13680 4634 64 1.88e-16
c13681 2557 2220 1.58e-16
c13682 2321 677 1.58e-16
c13683 1331 1136 5.5e-16
c13684 1011 0 3.7037e-14
c13685 1238 1 8.48e-16
c13686 4334 1 1.716e-15
c13687 4524 0 6.62e-16
c13688 777 920 3.15e-16
c13689 2243 2250 6.73e-16
c13690 2127 2117 1.96e-16
c13691 2103 2072 1.58e-16
c13692 4563 4418 1.58e-16
c13693 5200 5241 3.18e-16
c13694 393 390 2.142e-15
c13695 2509 1 7.56e-16
c13696 78 1 4.563e-15
c13697 3514 4319 1.58e-16
c13698 3497 4336 2.386e-15
c13699 4345 4339 1.6e-16
c13700 3543 1 2.054e-15
c13701 601 3387 4.48e-16
c13702 1540 1551 1.96e-16
c13703 1331 1016 5.5e-16
c13704 3545 0 8e-16
c13705 4136 1 5.1e-16
c13706 2995 2041 1.666e-15
c13707 3024 2838 1.58e-16
c13708 3030 2832 5.88e-16
c13709 4705 1 1.013e-15
c13710 2036 2098 3.54e-16
c13711 216 219 2.142e-15
c13712 3409 3484 1.58e-16
c13713 5249 5234 6.67e-16
c13714 5224 5226 5.48e-16
c13715 596 650 5.28e-16
c13716 3559 3557 2.15e-16
c13717 3567 3566 1.6e-16
c13718 2206 1 5.808e-15
c13719 512 513 3.84e-16
c13720 0 329 2.87e-16
c13721 4580 4196 4.63e-16
c13722 4582 4564 3.62e-16
c13723 5278 412 1.188e-15
c13724 4861 352 1.88e-16
c13725 883 1235 3.54e-16
c13726 907 890 4.274e-15
c13727 3327 842 2.33e-16
c13728 5296 5308 3.18e-16
c13729 601 3084 3.64e-16
c13730 602 2577 1.58e-16
c13731 921 722 3.15e-16
c13732 1321 1418 1.58e-16
c13733 1343 1406 1.58e-16
c13734 64 60 6.38e-16
c13735 59 53 1.58e-16
c13736 3882 4472 1.58e-16
c13737 3898 4484 1.58e-16
c13738 602 1358 1.58e-16
c13739 2535 2768 1.58e-16
c13740 2557 2756 1.58e-16
c13741 3740 468 9.43e-16
c13742 3839 3838 5.5e-16
c13743 4118 26 4.48e-16
c13744 4420 4419 2.03e-16
c13745 4425 4423 1.6e-16
c13746 3196 717 2.72e-16
c13747 3650 1 5.97e-15
c13748 2541 707 3.15e-16
c13749 3552 3553 9.1e-16
c13750 2396 2393 5.5e-16
c13751 2175 0 8.275e-14
c13752 3024 842 4.48e-16
c13753 2311 2317 1.6e-16
c13754 2308 1794 2.386e-15
c13755 1811 2291 1.58e-16
c13756 657 2541 4.03e-16
c13757 2578 1 1.868e-15
c13758 1682 2232 4.36e-16
c13759 4134 4143 1.88e-16
c13760 5577 4950 9.61e-16
c13761 5300 5299 1.334e-15
c13762 1321 837 3.15e-16
c13763 3690 858 1.75e-16
c13764 3332 0 3.466e-15
c13765 2871 2870 9.1e-16
c13766 1621 1619 1.6e-16
c13767 1343 1555 3.92e-16
c13768 1708 1437 1.58e-16
c13769 1706 1431 5.5e-16
c13770 1694 1832 1.58e-16
c13771 3480 1 5.97e-15
c13772 3242 3243 1.35e-16
c13773 1893 1890 3.01e-16
c13774 1889 1886 6.44e-16
c13775 3377 852 3.64e-16
c13776 3034 3313 1.58e-16
c13777 1550 0 6.9168e-14
c13778 2560 1 2.86e-16
c13779 722 717 2.77e-16
c13780 5449 1 1.23e-16
c13781 5160 5212 1.141e-15
c13782 4719 439 1.88e-16
c13783 2491 2490 9.1e-16
c13784 2172 2439 1.58e-16
c13785 2194 2427 1.58e-16
c13786 4102 3918 2.48e-16
c13787 1353 877 1.532e-15
c13788 1359 1358 5.65e-16
c13789 922 858 1.58e-16
c13790 921 1188 1.58e-16
c13791 5509 381 3.54e-16
c13792 1684 752 4.48e-16
c13793 4223 4226 4.41e-16
c13794 3078 3075 5.5e-16
c13795 632 2238 1.339e-15
c13796 4086 1 7.08e-16
c13797 4508 4504 1.96e-16
c13798 3273 767 4.81e-16
c13799 1763 1 1.056e-15
c13800 2747 2719 2.64e-16
c13801 537 542 1.88e-16
c13802 4829 0 2.93e-15
c13803 3393 3018 1.58e-16
c13804 3188 692 4.81e-16
c13805 642 2231 1.813e-15
c13806 1851 1 4.41e-15
c13807 1 437 1.456e-15
c13808 4725 4344 5.2e-16
c13809 2196 1913 5.5e-16
c13810 3242 767 2.33e-16
c13811 2360 0 6.62e-16
c13812 3723 3397 4.63e-16
c13813 883 842 6.45e-16
c13814 909 1202 4.35e-16
c13815 907 1201 1.88e-16
c13816 890 1194 1.58e-16
c13817 5356 5170 2.24e-16
c13818 2725 1 2.054e-15
c13819 617 2559 3.15e-16
c13820 1128 1129 1.21e-16
c13821 4217 4218 1.58e-16
c13822 2282 672 3.79e-16
c13823 2265 647 3.15e-16
c13824 1930 807 1.813e-15
c13825 2832 3356 4.36e-16
c13826 1708 2002 5.42e-16
c13827 1684 1990 1.58e-16
c13828 1817 1818 1.35e-16
c13829 4469 4470 1.35e-16
c13830 2545 677 3.15e-16
c13831 1955 1567 4.97e-16
c13832 37 477 1.88e-16
c13833 33 499 3e-16
c13834 27 484 1.88e-16
c13835 617 1732 2.33e-16
c13836 2703 1 1.716e-15
c13837 2841 2469 1.58e-16
c13838 3286 1 8.43e-16
c13839 1627 837 1.58e-16
c13840 1433 1432 1.6e-16
c13841 1425 1423 2.15e-16
c13842 4004 1687 2.573e-15
c13843 4508 842 5.03e-16
c13844 1335 1330 4.17e-16
c13845 4038 25 3.84e-16
c13846 3898 4247 3.92e-16
c13847 2370 722 4.81e-16
c13848 1862 707 1.58e-16
c13849 1257 1258 2.24e-16
c13850 3652 1 9.28e-16
c13851 537 281 1.88e-16
c13852 1379 1 8.43e-16
c13853 3588 0 3.6012e-14
c13854 3431 3430 1.6e-16
c13855 3423 3421 2.15e-16
c13856 3022 3383 1.58e-16
c13857 617 2225 5.03e-16
c13858 262 263 7.03e-16
c13859 244 243 6.67e-16
c13860 3358 842 4.81e-16
c13861 2271 2272 1.35e-16
c13862 4806 1 8.85e-16
c13863 2498 1 2.054e-15
c13864 3355 3350 1.642e-15
c13865 617 2584 1.339e-15
c13866 2500 0 8e-16
c13867 4014 4011 5.5e-16
c13868 4861 294 1.88e-16
c13869 5417 5406 7.92e-16
c13870 3013 2503 3.38e-16
c13871 4299 4300 1.35e-16
c13872 1584 837 1.58e-16
c13873 1321 1061 5.5e-16
c13874 1331 1508 1.58e-16
c13875 781 19 1.96e-16
c13876 1507 1509 2.03e-16
c13877 4243 1 1.868e-15
c13878 2707 722 5.03e-16
c13879 4219 37 5.71e-16
c13880 4233 0 2.93e-15
c13881 3330 3332 2.15e-16
c13882 1896 1505 1.136e-15
c13883 3695 3691 1.96e-16
c13884 1707 0 1.4914e-14
c13885 2044 2046 3.92e-16
c13886 15 369 4.88e-16
c13887 3695 842 5.03e-16
c13888 4915 91 1.88e-16
c13889 0 357 2.87e-16
c13890 5160 1 3.986e-15
c13891 2178 2189 1.96e-16
c13892 129 135 5.8e-16
c13893 143 100 1.88e-16
c13894 4322 3486 5.66e-16
c13895 5447 5459 8.45e-16
c13896 5410 5412 1.96e-16
c13897 1194 1201 2.27e-16
c13898 894 1143 3.54e-16
c13899 1011 1013 7.72e-16
c13900 911 889 6.87e-16
c13901 3882 3887 8.56e-16
c13902 5356 5352 5.7e-16
c13903 1899 737 4.81e-16
c13904 1516 722 1.58e-16
c13905 983 1 4.59e-16
c13906 4854 4463 1.96e-16
c13907 980 0 1.0077e-14
c13908 3048 2532 1.58e-16
c13909 3046 2529 1.58e-16
c13910 3034 3070 1.58e-16
c13911 1536 1 1.056e-15
c13912 4361 4723 1.58e-16
c13913 822 1181 4.21e-16
c13914 0 255 1.4803e-14
c13915 2196 2195 1.866e-15
c13916 2060 1 1.88e-16
c13917 4537 4992 5.68e-16
c13918 59 368 1.88e-16
c13919 78 363 1.88e-16
c13920 2831 2435 1.96e-16
c13921 1783 677 1.75e-16
c13922 632 3446 3.15e-16
c13923 3228 0 3.372e-14
c13924 4383 4382 9.1e-16
c13925 2338 717 2.4e-16
c13926 1659 1662 6.71e-16
c13927 1343 1191 1.58e-16
c13928 4390 1 2.054e-15
c13929 4639 4259 1.96e-16
c13930 2792 782 1.9e-16
c13931 1708 1765 3.92e-16
c13932 1330 1 2.56e-15
c13933 419 432 1.108e-15
c13934 4392 0 8e-16
c13935 2049 0 1.7153e-14
c13936 4896 1 3.884e-15
c13937 4923 4918 7.46e-16
c13938 3326 837 2.4e-16
c13939 216 217 5.8e-16
c13940 233 224 1.58e-16
c13941 422 0 1.051e-14
c13942 280 274 5.8e-16
c13943 282 291 1.58e-16
c13944 5270 5274 1.243e-15
c13945 2735 2367 1.96e-16
c13946 2468 1 8.43e-16
c13947 5533 5537 5.6e-16
c13948 4719 5365 9.98e-16
c13949 2541 2441 1.58e-16
c13950 2734 2735 9.1e-16
c13951 736 19 1.96e-16
c13952 1106 1562 2.38e-15
c13953 4259 4621 1.58e-16
c13954 4248 4629 5.66e-16
c13955 4635 4626 3.92e-16
c13956 4188 1 4.64e-16
c13957 1819 1431 4.97e-16
c13958 1243 0 3.8691e-14
c13959 822 921 3.15e-16
c13960 4452 4829 2.48e-16
c13961 3048 3211 1.58e-16
c13962 2162 2151 3.92e-16
c13963 1206 1 4.58e-15
c13964 11 5 1.482e-15
c13965 4844 4463 5.2e-16
c13966 1665 0 6.72e-16
c13967 27 44 1.88e-16
c13968 2426 2427 2.48e-16
c13969 78 131 1.88e-16
c13970 3806 3809 7.84e-16
c13971 3027 0 8.1998e-14
c13972 3554 722 2.33e-16
c13973 4810 5136 1.96e-16
c13974 3446 3435 1.58e-16
c13975 922 965 3.92e-16
c13976 3593 0 3.466e-15
c13977 627 629 5.59e-16
c13978 3876 4536 3.92e-16
c13979 3376 0 1.1956e-14
c13980 3030 777 4.03e-16
c13981 3996 1 4.64e-16
c13982 4552 1 1.052e-15
c13983 4710 4711 2.48e-16
c13984 4715 4714 2.83e-16
c13985 4718 4327 1.96e-16
c13986 601 1748 1.58e-16
c13987 1 563 2.946e-15
c13988 1681 1679 3.54e-16
c13989 2005 1 1.716e-15
c13990 3853 3857 1.96e-16
c13991 919 889 1.58e-16
c13992 2620 2627 1.96e-16
c13993 4668 5484 2.039e-15
c13994 2882 2881 4.61e-16
c13995 2535 2802 1.58e-16
c13996 2557 2790 1.58e-16
c13997 1136 1113 6.54e-16
c13998 3898 3503 1.58e-16
c13999 3192 0 1.6491e-14
c14000 2196 672 3.58e-16
c14001 1363 1318 2.64e-16
c14002 3957 19 9.67e-16
c14003 3231 747 1.58e-16
c14004 2535 2237 1.58e-16
c14005 2541 2231 5.88e-16
c14006 371 1 1.44e-16
c14007 3194 3196 2.15e-16
c14008 2177 1687 7.67e-16
c14009 4360 1 8.43e-16
c14010 4881 4883 2.15e-16
c14011 5034 120 7.46e-16
c14012 5144 31 7.16e-16
c14013 1732 1743 1.58e-16
c14014 5368 5367 1.6e-16
c14015 1 292 1.456e-15
c14016 4563 4435 1.58e-16
c14017 2602 0 2.93e-15
c14018 2526 2525 1.6e-16
c14019 2527 1998 1.23e-16
c14020 2510 2004 3.92e-16
c14021 2514 2512 1.96e-16
c14022 2521 1 1.286e-15
c14023 2794 2792 1.6e-16
c14024 2789 2788 2.03e-16
c14025 690 1 1.65e-16
c14026 2015 2194 3.92e-16
c14027 617 3387 4.48e-16
c14028 687 3886 7.99e-16
c14029 3202 747 1.813e-15
c14030 4521 4532 1.96e-16
c14031 777 890 3.35e-16
c14032 2987 2897 1.58e-16
c14033 3409 3489 1.58e-16
c14034 3194 722 1.58e-16
c14035 1 535 5.851e-15
c14036 3259 807 5.73e-16
c14037 4742 497 1.88e-16
c14038 777 2393 1.58e-16
c14039 2226 1 2.054e-15
c14040 1491 717 1.58e-16
c14041 592 868 5.8e-16
c14042 3719 858 7.68e-16
c14043 627 2583 1.58e-16
c14044 617 3084 7.68e-16
c14045 601 2577 3.15e-16
c14046 2015 2524 3.38e-16
c14047 1175 797 1.58e-16
c14048 4258 4249 3.46e-16
c14049 1352 1353 1.35e-16
c14050 2613 2612 1.6e-16
c14051 3898 4489 1.58e-16
c14052 3876 4501 1.58e-16
c14053 601 1358 1.84e-16
c14054 3262 3260 1.862e-15
c14055 2764 2736 2.64e-16
c14056 4517 1 1.056e-15
c14057 3175 3186 1.96e-16
c14058 1988 1607 3.92e-16
c14059 1992 1993 1.6e-16
c14060 25 204 5.71e-16
c14061 30 207 3.84e-16
c14062 911 2536 2.09e-16
c14063 2204 1 1.716e-15
c14064 3471 3470 2.03e-16
c14065 3476 3474 1.6e-16
c14066 3253 3248 1.642e-15
c14067 498 495 6.67e-16
c14068 3566 722 7.68e-16
c14069 1157 807 2.68e-16
c14070 890 1082 1.96e-16
c14071 2598 2599 9.1e-16
c14072 1820 692 1.58e-16
c14073 1449 1440 3.92e-16
c14074 1011 1443 5.66e-16
c14075 107 106 3.84e-16
c14076 4553 858 1.58e-16
c14077 627 3436 1.58e-16
c14078 3352 0 8e-16
c14079 867 1 5.57e-16
c14080 702 25 1.58e-16
c14081 2376 752 1.58e-16
c14082 1879 732 2.22e-16
c14083 1684 1448 5.5e-16
c14084 1694 1837 1.58e-16
c14085 1427 0 6.72e-16
c14086 349 346 3.54e-16
c14087 362 368 3.84e-16
c14088 4949 4946 3.54e-16
c14089 2306 1794 1.532e-15
c14090 3279 782 1.832e-15
c14091 2564 0 2.96e-16
c14092 632 3034 3.15e-16
c14093 2492 2486 1.545e-15
c14094 2172 2444 1.58e-16
c14095 1327 677 3.15e-16
c14096 1331 662 3.15e-16
c14097 388 1 4.22e-16
c14098 378 26 8.41e-16
c14099 392 27 1.88e-16
c14100 3704 1 1.056e-15
c14101 4318 4319 2.48e-16
c14102 2271 672 1.58e-16
c14103 2541 2552 1.96e-16
c14104 839 25 1.13e-15
c14105 843 19 1.58e-16
c14106 646 19 1.96e-16
c14107 2748 752 7.68e-16
c14108 1779 1 9.28e-16
c14109 77 79 1.58e-16
c14110 3256 3254 1.6e-16
c14111 4846 0 2.93e-15
c14112 5188 5190 1.77e-15
c14113 2299 2271 2.64e-16
c14114 3236 782 1.58e-16
c14115 762 2374 1.58e-16
c14116 397 508 1.88e-16
c14117 3898 662 4.46e-16
c14118 5450 5452 1.721e-15
c14119 4804 5259 1.383e-15
c14120 1455 702 1.58e-16
c14121 1203 852 6.98e-16
c14122 894 1217 3.92e-16
c14123 909 1216 1.88e-16
c14124 883 1209 1.58e-16
c14125 922 1038 1.58e-16
c14126 1905 767 1.58e-16
c14127 5416 528 7.97e-16
c14128 2447 812 1.84e-16
c14129 4760 4761 2.03e-16
c14130 2062 2071 1.873e-15
c14131 2161 1 1.052e-15
c14132 3350 858 1.84e-16
c14133 2729 1 8.43e-16
c14134 2291 2290 2.48e-16
c14135 883 1023 3.54e-16
c14136 894 1044 1.58e-16
c14137 2861 2469 2.38e-15
c14138 5577 4531 1.58e-16
c14139 1161 827 1.75e-16
c14140 1328 1351 1.003e-15
c14141 3876 4264 3.92e-16
c14142 821 1 5.57e-16
c14143 3249 3247 1.6e-16
c14144 3244 3243 2.03e-16
c14145 2899 0 1.8423e-14
c14146 1592 1136 4.97e-16
c14147 4679 4677 2.15e-16
c14148 4675 4686 1.96e-16
c14149 2809 807 2.72e-16
c14150 911 1698 1.829e-15
c14151 617 2245 1.09e-16
c14152 1652 1191 1.136e-15
c14153 4946 4992 4.47e-16
c14154 4823 1 8.85e-16
c14155 3387 3603 1.58e-16
c14156 4725 1 1.7194e-14
c14157 2515 1 1.871e-15
c14158 1059 1066 2.27e-16
c14159 2514 0 3.792e-15
c14160 3327 3411 1.58e-16
c14161 3321 3387 5.5e-16
c14162 4563 0 3.62856e-13
c14163 4787 497 1.88e-16
c14164 3882 4234 1.58e-16
c14165 3898 4246 1.58e-16
c14166 2756 2758 2.15e-16
c14167 1345 1076 5.5e-16
c14168 3385 1 5.277e-15
c14169 3068 3067 1.6e-16
c14170 3060 3058 2.15e-16
c14171 2727 722 1.09e-16
c14172 1852 1471 3.92e-16
c14173 1856 1857 1.6e-16
c14174 1143 1 1.56e-15
c14175 687 1694 7.99e-16
c14176 4488 4490 2.03e-16
c14177 3744 5021 1.33e-16
c14178 2181 2183 3.84e-16
c14179 5280 5281 3.54e-16
c14180 3879 3401 7.84e-16
c14181 4749 4747 1.6e-16
c14182 923 961 1.58e-16
c14183 1 495 1.456e-15
c14184 454 0 1.5723e-14
c14185 135 137 1.58e-16
c14186 106 1 9.8e-16
c14187 71 9 5.8e-16
c14188 4861 62 5.8e-16
c14189 2763 2754 3.46e-16
c14190 1188 842 1.58e-16
c14191 3876 3877 1.487e-15
c14192 4205 4207 2.239e-15
c14193 598 0 7.709e-15
c14194 3453 0 1.6491e-14
c14195 1005 1 3.06e-16
c14196 3650 3622 2.64e-16
c14197 4051 1 6.78e-16
c14198 3633 3639 1.418e-15
c14199 4470 4472 1.862e-15
c14200 3332 3328 1.96e-16
c14201 4361 4740 1.58e-16
c14202 3024 2533 5.5e-16
c14203 3034 3075 1.58e-16
c14204 2929 852 1.58e-16
c14205 1694 1567 5.5e-16
c14206 216 259 1.88e-16
c14207 762 1544 2.72e-16
c14208 0 164 1.5723e-14
c14209 37 172 5.71e-16
c14210 25 175 5.71e-16
c14211 523 477 1.88e-16
c14212 5194 1 2.53e-16
c14213 5032 5036 1.96e-16
c14214 3773 3821 3.15e-16
c14215 1118 1119 1.213e-15
c14216 146 252 1.88e-16
c14217 161 165 1.58e-16
c14218 2657 0 1.4092e-14
c14219 59 102 1.88e-16
c14220 64 93 1.88e-16
c14221 1161 812 2.33e-16
c14222 3899 1 2.471e-15
c14223 4024 26 1.075e-15
c14224 2162 858 1.58e-16
c14225 1206 1321 1.58e-16
c14226 1196 1327 5.88e-16
c14227 776 1 5.57e-16
c14228 3411 762 3.58e-16
c14229 3905 0 2.96e-16
c14230 3124 3126 1.862e-15
c14231 2611 2617 1.418e-15
c14232 3506 3505 2.48e-16
c14233 4276 4639 1.96e-16
c14234 1948 1556 1.96e-16
c14235 1949 1942 6.73e-16
c14236 3599 747 2.22e-16
c14237 3515 662 3.64e-16
c14238 5165 207 3.54e-16
c14239 1981 1976 1.642e-15
c14240 88 334 1.88e-16
c14241 426 233 1.88e-16
c14242 5383 5387 8.88e-16
c14243 276 27 1.88e-16
c14244 3866 852 3.64e-16
c14245 2550 2544 1.6e-16
c14246 1281 1226 3.84e-16
c14247 1660 1662 1.6e-16
c14248 3062 0 6.72e-16
c14249 2557 2458 1.58e-16
c14250 3126 3125 2.48e-16
c14251 3138 2645 1.58e-16
c14252 1954 812 1.339e-15
c14253 4259 4638 1.58e-16
c14254 4207 1 6.76e-16
c14255 2701 707 7.38e-16
c14256 592 0 3.31034e-13
c14257 3675 3677 2.03e-16
c14258 4842 4843 8.22e-16
c14259 2444 0 3.3534e-14
c14260 926 889 1.081e-15
c14261 938 939 1.6e-16
c14262 5071 91 5.5e-16
c14263 3029 0 4.3406e-14
c14264 3548 737 1.58e-16
c14265 5440 5443 1.98e-16
c14266 1016 1014 1.931e-15
c14267 4292 4285 1.96e-16
c14268 3446 4294 4.36e-16
c14269 1706 662 4.46e-16
c14270 919 979 1.58e-16
c14271 3900 3898 4.506e-15
c14272 642 1402 2.4e-16
c14273 3396 0 1.5577e-14
c14274 3046 792 3.15e-16
c14275 2880 2944 1.6e-16
c14276 3134 2617 1.136e-15
c14277 3220 3211 3.92e-16
c14278 2702 3214 5.66e-16
c14279 2016 2010 1.6e-16
c14280 1618 2007 2.386e-15
c14281 1706 1918 3.92e-16
c14282 617 1748 7.38e-16
c14283 30 296 3.84e-16
c14284 5155 5157 1.441e-15
c14285 303 349 1.88e-16
c14286 5549 584 5.93e-16
c14287 4804 1 2.9721e-14
c14288 2803 2418 1.96e-16
c14289 4589 0 4.75679e-13
c14290 4071 4072 6.4e-16
c14291 2651 2652 1.35e-16
c14292 3882 3514 5.88e-16
c14293 3876 3520 1.58e-16
c14294 3616 4434 1.96e-16
c14295 1746 1744 1.6e-16
c14296 3976 0 2.0592e-14
c14297 2308 702 1.58e-16
c14298 917 0 3.8e-16
c14299 731 1 5.57e-16
c14300 3123 672 1.58e-16
c14301 1031 0 7.4292e-14
c14302 187 189 1.88e-16
c14303 2351 2345 1.6e-16
c14304 1834 2350 1.136e-15
c14305 5164 296 7.97e-16
c14306 3046 737 4.46e-16
c14307 822 1969 2.4e-16
c14308 2627 2618 3.46e-16
c14309 894 889 1.58e-16
c14310 13 27 3.75e-16
c14311 3397 827 3.15e-16
c14312 4563 4452 1.58e-16
c14313 2557 1 4.77e-16
c14314 1321 1606 3.92e-16
c14315 700 1 3.79e-16
c14316 693 0 7.86e-15
c14317 1694 1318 1.58e-16
c14318 4336 0 3.3724e-14
c14319 2545 2559 4.274e-15
c14320 2172 807 3.15e-16
c14321 792 907 3.15e-16
c14322 537 397 1.88e-16
c14323 3048 2849 5.5e-16
c14324 1803 1 5.808e-15
c14325 701 700 6.67e-16
c14326 1805 0 3.466e-15
c14327 4862 0 1.6462e-14
c14328 3214 722 1.58e-16
c14329 2141 2022 1.52e-16
c14330 2103 2106 7.84e-16
c14331 1022 672 2.68e-16
c14332 19 517 3.2e-16
c14333 306 312 1.372e-15
c14334 3572 3583 1.96e-16
c14335 3668 807 2.65e-16
c14336 2194 1794 5.5e-16
c14337 3918 3964 2.87e-16
c14338 1263 1262 1.6e-16
c14339 3373 3842 1.722e-15
c14340 617 2577 3.15e-16
c14341 52 0 1.4803e-14
c14342 4264 4263 9.1e-16
c14343 1327 996 1.58e-16
c14344 3876 4506 1.58e-16
c14345 3900 4518 5.42e-16
c14346 2469 827 3.15e-16
c14347 2196 797 3.15e-16
c14348 1813 1806 6.73e-16
c14349 1072 0 1.8851e-14
c14350 3952 1 4.738e-15
c14351 2106 2101 7.46e-16
c14352 612 1718 1.58e-16
c14353 518 514 1.372e-15
c14354 513 505 1.58e-16
c14355 4567 4592 1.58e-16
c14356 4571 3870 3.54e-16
c14357 2230 1 8.43e-16
c14358 3185 722 3.15e-16
c14359 3338 3393 5.88e-16
c14360 3344 3387 1.58e-16
c14361 5143 1 3.36e-16
c14362 687 2541 4.03e-16
c14363 907 737 4.8e-16
c14364 883 1097 3.92e-16
c14365 890 1096 1.88e-16
c14366 5388 5335 9.01e-16
c14367 4838 5034 2.665e-15
c14368 3397 3276 1.58e-16
c14369 5346 5345 1.6e-16
c14370 2777 0 6.72e-16
c14371 2596 1 9.28e-16
c14372 601 589 6.38e-16
c14373 83 79 1.372e-15
c14374 47 48 2.84e-16
c14375 53 42 2.45e-16
c14376 2997 2984 8.94e-16
c14377 1840 692 1.58e-16
c14378 3166 1 6.15e-16
c14379 4514 4571 5.5e-16
c14380 3599 4416 1.58e-16
c14381 3588 4424 5.66e-16
c14382 4430 4421 3.92e-16
c14383 1625 1176 3.92e-16
c14384 1629 1630 1.6e-16
c14385 2850 837 2.65e-16
c14386 1708 1465 5.5e-16
c14387 632 2266 3.64e-16
c14388 617 1760 1.58e-16
c14389 1901 1516 1.96e-16
c14390 5240 178 7.62e-16
c14391 5093 0 1.963e-15
c14392 2235 2236 9.1e-16
c14393 3409 3637 1.58e-16
c14394 3397 812 3.15e-16
c14395 2305 2306 1.35e-16
c14396 3882 827 3.15e-16
c14397 2559 2582 3.92e-16
c14398 922 1203 1.58e-16
c14399 2007 868 1.58e-16
c14400 1321 1571 1.58e-16
c14401 1343 1559 1.58e-16
c14402 642 1345 3.58e-16
c14403 602 3877 5.18e-16
c14404 612 3397 7.99e-16
c14405 1505 1888 7.84e-16
c14406 4300 0 1.6491e-14
c14407 3347 2849 1.58e-16
c14408 1792 1 6.15e-16
c14409 3387 3072 1.58e-16
c14410 3242 3624 2.48e-16
c14411 2387 1 1.056e-15
c14412 448 459 2.45e-16
c14413 9 204 5.8e-16
c14414 1 192 3.6e-16
c14415 0 218 6.1665e-14
c14416 3270 767 1.58e-16
c14417 3653 782 4.81e-16
c14418 3975 857 6.23e-16
c14419 5473 0 2.285e-15
c14420 3041 2538 1.159e-15
c14421 4451 767 1.58e-16
c14422 2783 2782 1.6e-16
c14423 2775 2773 2.15e-16
c14424 1041 692 2.33e-16
c14425 4366 692 1.58e-16
c14426 4196 3890 3.84e-16
c14427 1044 1 2.972e-15
c14428 4100 1 2.259e-15
c14429 2469 812 1.58e-16
c14430 2650 647 1.58e-16
c14431 4092 25 1.88e-16
c14432 1045 0 6.29e-16
c14433 1576 1 5.808e-15
c14434 1706 1624 1.58e-16
c14435 1578 0 3.466e-15
c14436 792 1116 5.73e-16
c14437 25 436 5.71e-16
c14438 4571 4559 3.84e-16
c14439 5111 5113 3.92e-16
c14440 5124 5101 2.12e-16
c14441 5108 5105 2.004e-15
c14442 3893 3883 5.8e-16
c14443 1149 782 8.3e-16
c14444 93 122 3.75e-16
c14445 687 3525 2.72e-16
c14446 1176 868 5.73e-16
c14447 1636 827 3.64e-16
c14448 3900 4281 3.92e-16
c14449 2857 2859 2.03e-16
c14450 662 26 7.12e-16
c14451 824 26 2.65e-15
c14452 1959 1956 5.5e-16
c14453 117 194 1.88e-16
c14454 3436 3447 1.96e-16
c14455 1533 1 5.97e-15
c14456 190 189 7.08e-16
c14457 3553 692 1.58e-16
c14458 5165 296 1.76e-16
c14459 2295 2293 1.6e-16
c14460 2290 2289 2.03e-16
c14461 5283 5288 3.73e-16
c14462 4776 236 1.88e-16
c14463 1053 692 1.58e-16
c14464 4136 857 3.1e-16
c14465 3898 3486 1.58e-16
c14466 3898 4251 1.58e-16
c14467 3876 4263 1.58e-16
c14468 3882 812 3.15e-16
c14469 2839 2841 1.862e-15
c14470 5403 5440 5.48e-16
c14471 2594 0 6.9481e-14
c14472 911 1680 1.88e-16
c14473 3638 792 2.4e-16
c14474 602 3876 3.46e-16
c14475 595 3900 3.15e-16
c14476 612 3882 4.03e-16
c14477 4279 1 1.056e-15
c14478 1375 0 1.4092e-14
c14479 1177 1 3.54e-16
c14480 1174 0 9.602e-15
c14481 4469 4845 3.92e-16
c14482 5010 439 1.88e-16
c14483 2179 2198 9.83e-16
c14484 412 352 3.45e-16
c14485 3397 3406 1.58e-16
c14486 968 969 1.213e-15
c14487 4567 4723 1.58e-16
c14488 4580 4327 5.5e-16
c14489 4582 4333 1.58e-16
c14490 747 2356 1.58e-16
c14491 5450 5410 5.69e-16
c14492 1459 677 1.9e-16
c14493 1207 858 6.38e-16
c14494 391 393 1.58e-16
c14495 911 3881 1.58e-16
c14496 1519 1517 1.6e-16
c14497 807 0 2.86609e-13
c14498 2921 2929 4.48e-16
c14499 1019 1 3.06e-16
c14500 1791 1788 3.01e-16
c14501 1787 1784 6.44e-16
c14502 4378 4740 1.58e-16
c14503 3048 2577 5.5e-16
c14504 1540 1 1.716e-15
c14505 3517 3515 1.6e-16
c14506 0 354 5.5097e-14
c14507 25 349 5.71e-16
c14508 218 219 1.079e-15
c14509 37 345 1.88e-16
c14510 2552 2175 1.159e-15
c14511 2373 2367 1.418e-15
c14512 2356 2384 2.64e-16
c14513 2378 2374 1.96e-16
c14514 921 672 3.15e-16
c14515 920 647 3.69e-16
c14516 160 158 1.88e-16
c14517 3876 3896 3.92e-16
c14518 2843 2452 4.11e-16
c14519 2136 2118 1.58e-16
c14520 910 592 5.8e-16
c14521 2541 2683 1.58e-16
c14522 2594 2203 1.136e-15
c14523 3571 1 4.41e-15
c14524 4656 4276 1.96e-16
c14525 4405 0 6.62e-16
c14526 421 418 1.099e-15
c14527 4861 5113 7.98e-16
c14528 1042 1043 7.46e-16
c14529 5177 5176 1.062e-15
c14530 2549 2544 4.17e-16
c14531 1789 662 1.84e-16
c14532 4086 857 1.88e-16
c14533 911 3390 1.58e-16
c14534 1218 1295 3.92e-16
c14535 1305 1306 3.92e-16
c14536 3886 782 3.15e-16
c14537 3650 837 1.58e-16
c14538 1690 827 3.15e-16
c14539 919 1160 3.92e-16
c14540 922 1159 2.54e-16
c14541 3143 2645 1.58e-16
c14542 1585 1131 1.96e-16
c14543 1586 1579 6.73e-16
c14544 4276 4638 1.58e-16
c14545 4265 4646 5.66e-16
c14546 4652 4643 3.92e-16
c14547 3024 2719 1.58e-16
c14548 3030 2713 5.88e-16
c14549 1471 0 3.583e-14
c14550 644 645 1.6e-16
c14551 3393 3553 1.96e-16
c14552 4986 526 9.36e-16
c14553 827 820 5.58e-16
c14554 1 132 1.65e-15
c14555 15 117 5.8e-16
c14556 9 175 5.8e-16
c14557 130 0 1.5696e-14
c14558 3411 722 3.15e-16
c14559 3202 3594 2.38e-15
c14560 5051 5031 1.58e-16
c14561 4844 323 1.88e-16
c14562 2464 0 1.4092e-14
c14563 1291 1231 3.92e-16
c14564 1243 1226 1.137e-15
c14565 3804 3803 3.54e-16
c14566 5388 5389 3.54e-16
c14567 4181 4175 7.45e-16
c14568 3427 1 6.15e-16
c14569 140 139 1.58e-16
c14570 143 142 6.4e-16
c14571 2299 717 1.58e-16
c14572 1823 1820 5.5e-16
c14573 1211 1657 1.96e-16
c14574 2662 2657 1.642e-15
c14575 4454 3622 2.48e-16
c14576 3312 3314 2.03e-16
c14577 2390 782 1.75e-16
c14578 1708 1706 4.506e-15
c14579 1666 1663 1.6e-16
c14580 76 88 1.58e-16
c14581 4197 1 4.709e-15
c14582 4727 4728 2.48e-16
c14583 4732 4731 2.83e-16
c14584 4735 4344 1.96e-16
c14585 1684 1935 3.92e-16
c14586 889 888 1.518e-15
c14587 2037 236 9.43e-16
c14588 5036 5028 3.54e-16
c14589 632 3118 3.64e-16
c14590 284 1 1.44e-16
c14591 4753 236 7.45e-16
c14592 3033 3035 3.84e-16
c14593 2041 2045 3.01e-16
c14594 1405 1407 2.03e-16
c14595 889 1 8.183e-15
c14596 4569 5535 9.43e-16
c14597 2918 2917 3.54e-16
c14598 4265 4266 1.35e-16
c14599 3886 4382 1.58e-16
c14600 3898 3531 5.5e-16
c14601 3900 3537 1.58e-16
c14602 2719 762 5.73e-16
c14603 2559 2248 5.5e-16
c14604 2328 702 1.58e-16
c14605 1653 1647 1.6e-16
c14606 1181 1644 2.386e-15
c14607 3220 3209 1.96e-16
c14608 2645 662 3.15e-16
c14609 3034 3035 1.027e-15
c14610 1794 1403 1.136e-15
c14611 3397 747 7.99e-16
c14612 4556 0 2.0654e-14
c14613 1929 1920 3.46e-16
c14614 1211 1 1.238e-15
c14615 647 641 1.74e-16
c14616 3048 752 3.15e-16
c14617 2007 0 3.3749e-14
c14618 235 1 4.92e-16
c14619 3276 3659 7.84e-16
c14620 2265 0 6.9068e-14
c14621 226 0 1.4803e-14
c14622 2041 2054 3.18e-16
c14623 1589 797 7.38e-16
c14624 1345 732 3.58e-16
c14625 1387 1389 1.862e-15
c14626 2178 2354 1.58e-16
c14627 2248 1732 1.136e-15
c14628 3989 3983 7.45e-16
c14629 3050 1 2.86e-16
c14630 1504 722 7.38e-16
c14631 719 1 7.18e-16
c14632 2306 702 1.58e-16
c14633 1690 812 3.15e-16
c14634 1345 1623 3.92e-16
c14635 374 19 3.45e-16
c14636 2611 3105 1.96e-16
c14637 1331 1453 4.63e-16
c14638 4356 0 1.4092e-14
c14639 4542 4543 9.13e-16
c14640 2475 842 2.33e-16
c14641 2671 692 1.58e-16
c14642 3502 647 1.58e-16
c14643 2987 2934 9.01e-16
c14644 2264 2255 3.46e-16
c14645 612 1690 4.03e-16
c14646 595 1708 3.15e-16
c14647 602 1684 3.46e-16
c14648 4718 1 8.43e-16
c14649 4879 0 1.6741e-14
c14650 2151 1652 1.66e-16
c14651 1670 2106 2.863e-15
c14652 662 1014 1.58e-16
c14653 1 301 4.22e-16
c14654 233 513 1.88e-16
c14655 2522 2196 1.96e-16
c14656 0 302 9.795e-15
c14657 3287 807 3.79e-16
c14658 3659 812 1.58e-16
c14659 2407 2408 1.35e-16
c14660 2182 2354 1.58e-16
c14661 2172 1811 5.5e-16
c14662 595 2178 4.03e-16
c14663 3918 3982 6.32e-16
c14664 3011 1 2.48e-16
c14665 2799 2790 3.92e-16
c14666 1056 732 5.73e-16
c14667 361 369 2.218e-15
c14668 4270 4266 1.96e-16
c14669 2705 2703 1.862e-15
c14670 2333 2305 2.64e-16
c14671 601 952 2.33e-16
c14672 2486 868 3.79e-16
c14673 3966 1 6.76e-16
c14674 601 4264 1.58e-16
c14675 3288 3290 1.6e-16
c14676 3024 3173 3.92e-16
c14677 762 1111 1.35e-16
c14678 1862 1857 1.642e-15
c14679 4521 1 1.716e-15
c14680 612 1738 1.58e-16
c14681 1176 0 3.7577e-14
c14682 4567 4609 1.58e-16
c14683 4571 3874 5.5e-16
c14684 1913 2405 1.58e-16
c14685 595 2182 9.84e-16
c14686 891 886 5.11e-16
c14687 722 712 6.38e-16
c14688 3452 3453 1.35e-16
c14689 909 752 3.15e-16
c14690 883 1111 1.88e-16
c14691 907 1104 1.58e-16
c14692 5262 5044 4.35e-16
c14693 2609 1 6.15e-16
c14694 2855 1 4.946e-15
c14695 1835 717 1.58e-16
c14696 1331 852 7.99e-16
c14697 1343 858 1.58e-16
c14698 657 592 5.8e-16
c14699 617 3457 1.9e-16
c14700 3368 0 6.72e-16
c14701 3175 1 1.716e-15
c14702 3599 4421 1.58e-16
c14703 2896 2893 3.92e-16
c14704 3938 0 2.6812e-14
c14705 3928 26 1.075e-15
c14706 601 1716 1.339e-15
c14707 1449 1 1.868e-15
c14708 1777 1772 1.642e-15
c14709 1439 0 2.93e-15
c14710 3089 3475 5.66e-16
c14711 3481 3472 3.92e-16
c14712 3882 747 4.03e-16
c14713 3100 3467 1.58e-16
c14714 485 484 6.96e-16
c14715 3570 732 2.4e-16
c14716 4847 1 4.832e-15
c14717 5072 0 4.0868e-14
c14718 2770 797 1.75e-16
c14719 1971 0 1.6491e-14
c14720 683 682 1.96e-16
c14721 3409 3642 1.58e-16
c14722 5262 5230 1.58e-16
c14723 1097 722 1.58e-16
c14724 601 3451 1.58e-16
c14725 2178 1970 1.58e-16
c14726 3898 852 3.15e-16
c14727 5403 5511 1.58e-16
c14728 2532 2530 3.54e-16
c14729 3909 25 3.84e-16
c14730 3176 3178 2.03e-16
c14731 1694 782 3.15e-16
c14732 1345 1588 5.42e-16
c14733 1321 1576 1.58e-16
c14734 1211 1215 2.03e-16
c14735 627 3397 7.99e-16
c14736 1538 1091 1.96e-16
c14737 2594 3087 1.58e-16
c14738 1516 1900 1.58e-16
c14739 4859 4480 1.58e-16
c14740 3411 3089 1.58e-16
c14741 217 218 1.88e-16
c14742 4036 4038 4.33e-16
c14743 4759 4378 5.2e-16
c14744 2182 1970 1.58e-16
c14745 0 338 1.5723e-14
c14746 762 2395 2.72e-16
c14747 393 0 1.051e-14
c14748 3321 3689 1.96e-16
c14749 5429 5425 1.866e-15
c14750 5484 5481 7.84e-16
c14751 4810 5262 5.5e-16
c14752 1031 707 1.58e-16
c14753 602 3896 1.58e-16
c14754 687 1011 5.73e-16
c14755 2978 2968 1.96e-16
c14756 2954 2923 1.58e-16
c14757 3744 3746 1.062e-15
c14758 687 4332 2.4e-16
c14759 3886 3633 5.5e-16
c14760 3708 0 1.6491e-14
c14761 4777 4778 2.03e-16
c14762 3024 3138 1.58e-16
c14763 3046 3126 1.58e-16
c14764 3083 2566 1.136e-15
c14765 3016 858 7.12e-16
c14766 5158 5219 1.6e-16
c14767 792 1585 2.65e-16
c14768 5404 468 3.54e-16
c14769 5104 5108 1.96e-16
c14770 4844 265 1.88e-16
c14771 2391 2402 1.96e-16
c14772 3514 702 1.813e-15
c14773 5311 5310 1.6e-16
c14774 4145 4143 1.06e-16
c14775 4132 4134 4.33e-16
c14776 4087 37 1.88e-16
c14777 4406 3571 1.96e-16
c14778 4411 3565 1.96e-16
c14779 2541 2752 1.96e-16
c14780 3834 0 1.2027e-14
c14781 4696 4694 2.15e-16
c14782 4692 4703 1.96e-16
c14783 642 19 1.41e-15
c14784 326 321 1.059e-15
c14785 4977 4975 1.133e-15
c14786 4944 5000 9.34e-16
c14787 1794 2287 1.96e-16
c14788 1950 1 1.056e-15
c14789 3875 3895 2.07e-16
c14790 3899 3904 9.6e-16
c14791 3393 3219 5.88e-16
c14792 4725 410 1.88e-16
c14793 2536 1 2.606e-15
c14794 1072 707 1.58e-16
c14795 1053 1059 1.58e-16
c14796 592 790 6.34e-16
c14797 687 3519 2.4e-16
c14798 3599 3594 1.642e-15
c14799 595 3407 2.13e-16
c14800 1106 752 3.15e-16
c14801 3876 4268 1.58e-16
c14802 3900 4280 5.42e-16
c14803 921 1205 1.96e-16
c14804 612 953 1.58e-16
c14805 629 1 7.18e-16
c14806 3411 822 3.58e-16
c14807 1607 842 1.75e-16
c14808 1596 1593 5.5e-16
c14809 1331 1101 1.58e-16
c14810 1698 1335 3.84e-16
c14811 601 3876 4.48e-16
c14812 627 3882 4.03e-16
c14813 4295 1 9.28e-16
c14814 3073 3084 1.96e-16
c14815 1869 1482 1.532e-15
c14816 1875 1874 5.65e-16
c14817 4989 4978 1.96e-16
c14818 642 2253 2.4e-16
c14819 3034 3292 4.63e-16
c14820 3151 3146 1.642e-15
c14821 3030 647 3.15e-16
c14822 1735 0 3.3874e-14
c14823 9 436 5.8e-16
c14824 3608 3620 2.32e-16
c14825 4606 3874 5.2e-16
c14826 4567 4740 1.58e-16
c14827 4580 4344 5.5e-16
c14828 4582 4350 1.58e-16
c14829 4827 33 1.88e-16
c14830 3397 3021 1.58e-16
c14831 2476 2478 1.862e-15
c14832 1964 1970 1.418e-15
c14833 1340 1341 1.736e-15
c14834 107 421 1.88e-16
c14835 4855 91 1.88e-16
c14836 1031 1035 2.03e-16
c14837 911 3397 3.45e-16
c14838 4500 4498 1.6e-16
c14839 2620 647 1.58e-16
c14840 2446 797 1.9e-16
c14841 4361 4748 2.196e-15
c14842 471 30 6.83e-16
c14843 131 132 7.08e-16
c14844 479 49 1.88e-16
c14845 3411 3404 3.54e-16
c14846 1811 0 6.9481e-14
c14847 0 477 4.6772e-14
c14848 26 494 8.41e-16
c14849 30 497 3.84e-16
c14850 5066 5071 7.25e-16
c14851 2196 2252 5.42e-16
c14852 1132 1113 1.546e-15
c14853 2567 2569 1.862e-15
c14854 2166 2169 1.576e-15
c14855 1428 1425 3.01e-16
c14856 1424 1421 6.44e-16
c14857 3882 4416 1.58e-16
c14858 2753 0 3.6007e-14
c14859 2339 722 2.33e-16
c14860 2557 2700 1.58e-16
c14861 2541 2688 1.58e-16
c14862 3154 3152 1.6e-16
c14863 4430 1 1.868e-15
c14864 4293 4656 1.96e-16
c14865 49 189 1.88e-16
c14866 4420 0 2.93e-15
c14867 248 262 1.58e-16
c14868 251 253 1.58e-16
c14869 3426 3423 3.01e-16
c14870 3422 3419 6.44e-16
c14871 2257 1760 1.58e-16
c14872 747 1690 4.03e-16
c14873 890 647 3.15e-16
c14874 592 745 6.34e-16
c14875 3722 3723 9.1e-16
c14876 4861 4867 5.87e-16
c14877 2542 2565 1.003e-15
c14878 73 88 1.88e-16
c14879 2172 2389 3.92e-16
c14880 4736 5170 4.79e-16
c14881 2583 1 4.41e-15
c14882 1706 852 3.15e-16
c14883 398 402 1.372e-15
c14884 392 389 1.099e-15
c14885 4276 4655 1.58e-16
c14886 1690 1403 1.58e-16
c14887 2804 827 1.75e-16
c14888 1698 1 8.822e-15
c14889 4219 0 2.0707e-14
c14890 2759 2367 2.38e-15
c14891 9 349 5.8e-16
c14892 3679 827 1.84e-16
c14893 2486 0 7.0011e-14
c14894 2178 2388 1.58e-16
c14895 5356 0 3.0503e-14
c14896 2172 2191 1.58e-16
c14897 921 797 3.15e-16
c14898 5442 5447 3.54e-16
c14899 1397 1392 1.642e-15
c14900 2248 2640 2.38e-15
c14901 3436 1 1.716e-15
c14902 911 3882 7.6e-16
c14903 2333 702 2.22e-16
c14904 1211 1321 3.92e-16
c14905 3504 3123 3.92e-16
c14906 2194 702 3.15e-16
c14907 1764 1380 1.58e-16
c14908 2541 782 3.15e-16
c14909 2023 2025 8.88e-16
c14910 2047 2046 1.6e-16
c14911 1 243 4.22e-16
c14912 822 2418 1.58e-16
c14913 2196 1868 1.58e-16
c14914 2182 2388 1.58e-16
c14915 2275 0 6.62e-16
c14916 0 250 9.795e-15
c14917 657 2594 1.58e-16
c14918 642 2611 3.79e-16
c14919 986 647 3.15e-16
c14920 5410 5461 1.191e-15
c14921 407 400 3.54e-16
c14922 404 403 6.4e-16
c14923 64 352 1.88e-16
c14924 4804 410 1.88e-16
c14925 2646 2635 1.96e-16
c14926 642 1406 1.58e-16
c14927 632 1392 1.84e-16
c14928 3789 3781 1.96e-16
c14929 4095 4094 5.5e-16
c14930 3231 1 2.054e-15
c14931 1151 1154 6.13e-16
c14932 954 0 1.8536e-14
c14933 3030 3031 1.239e-15
c14934 1652 858 3.15e-16
c14935 1684 1934 1.58e-16
c14936 1706 1922 1.58e-16
c14937 632 2196 3.15e-16
c14938 1316 1 1.96e-16
c14939 3513 3117 1.96e-16
c14940 1935 1934 9.1e-16
c14941 436 419 1.325e-15
c14942 508 262 1.88e-16
c14943 4931 4930 1.6e-16
c14944 2266 2255 1.96e-16
c14945 421 1 2.6688e-14
c14946 222 224 1.58e-16
c14947 2807 2418 2.386e-15
c14948 2639 2635 1.96e-16
c14949 907 977 3.92e-16
c14950 3287 3671 1.58e-16
c14951 404 26 1.03e-15
c14952 4702 33 1.88e-16
c14953 3234 1 6.15e-16
c14954 4470 812 1.339e-15
c14955 5550 5530 8.66e-16
c14956 3531 3537 1.418e-15
c14957 4368 4370 1.862e-15
c14958 1817 692 2.33e-16
c14959 3202 1 5.97e-15
c14960 1566 1557 3.46e-16
c14961 2776 782 1.84e-16
c14962 4187 1 6.78e-16
c14963 2691 692 1.58e-16
c14964 627 1690 4.03e-16
c14965 601 1684 4.48e-16
c14966 2804 812 2.33e-16
c14967 822 1973 1.58e-16
c14968 2787 3296 7.84e-16
c14969 3662 3661 1.6e-16
c14970 3276 3657 3.92e-16
c14971 4735 1 8.43e-16
c14972 2427 1 5.808e-15
c14973 2153 2154 9.13e-16
c14974 2150 2151 2.49e-16
c14975 747 1482 1.58e-16
c14976 1 40 4.22e-16
c14977 9 5 5.8e-16
c14978 4567 4463 5.5e-16
c14979 3679 812 1.58e-16
c14980 5377 1 7.49e-16
c14981 2429 0 3.466e-15
c14982 792 1902 5.73e-16
c14983 777 25 1.58e-16
c14984 3741 3739 6.16e-16
c14985 5514 5492 1.58e-16
c14986 1243 1246 1.001e-15
c14987 59 136 1.88e-16
c14988 2545 2435 5.5e-16
c14989 1345 1011 1.58e-16
c14990 1331 1452 1.58e-16
c14991 3364 1 6.636e-15
c14992 617 952 1.75e-16
c14993 4344 4339 1.642e-15
c14994 3898 3690 1.58e-16
c14995 4538 4541 6.71e-16
c14996 2669 692 1.339e-15
c14997 3995 1 6.78e-16
c14998 617 4264 7.38e-16
c14999 1738 1739 5.65e-16
c15000 3213 737 5.03e-16
c15001 3048 3190 3.92e-16
c15002 4547 1 5.01e-16
c15003 2545 752 3.15e-16
c15004 315 311 1.372e-15
c15005 3657 812 1.339e-15
c15006 4567 4626 1.58e-16
c15007 4571 4242 5.5e-16
c15008 1896 2413 2.38e-15
c15009 27 570 1.88e-16
c15010 3862 3338 1.96e-16
c15011 5364 0 1.65e-16
c15012 2799 1 1.868e-15
c15013 2342 2340 1.862e-15
c15014 56 5 1.88e-16
c15015 2789 0 2.93e-15
c15016 3014 3006 7.29e-16
c15017 3001 3003 2.861e-15
c15018 1471 707 2.33e-16
c15019 3599 4441 2.38e-15
c15020 732 19 1.41e-15
c15021 3942 26 4.48e-16
c15022 3192 3195 6.44e-16
c15023 3573 3575 2.03e-16
c15024 3100 3472 1.58e-16
c15025 4864 1 4.832e-15
c15026 909 891 4.02e-16
c15027 3710 3712 2.15e-16
c15028 5417 1 4.669e-15
c15029 617 3451 7.38e-16
c15030 2513 2510 6.71e-16
c15031 1371 952 2.48e-16
c15032 3224 747 2.4e-16
c15033 617 992 1.58e-16
c15034 2310 677 1.9e-16
c15035 4319 1 5.808e-15
c15036 2594 3092 1.58e-16
c15037 2754 767 1.339e-15
c15038 1914 1908 1.6e-16
c15039 1516 1905 2.386e-15
c15040 1233 1 1.23e-16
c15041 4321 0 3.466e-15
c15042 4497 4859 1.58e-16
c15043 4867 4486 5.66e-16
c15044 4864 4873 3.92e-16
c15045 5341 5316 5.87e-16
c15046 2178 1687 1.96e-16
c15047 2149 2078 5.95e-16
c15048 3387 3100 5.5e-16
c15049 5200 5195 7.37e-16
c15050 5151 5188 5.48e-16
c15051 4742 468 1.88e-16
c15052 2391 1 1.716e-15
c15053 993 1007 1.96e-16
c15054 5309 1 3.36e-16
c15055 3942 3947 1.96e-16
c15056 3918 3926 2.48e-16
c15057 1502 707 4.81e-16
c15058 64 294 1.88e-16
c15059 4250 4252 2.03e-16
c15060 595 3409 3.15e-16
c15061 2305 2687 2.48e-16
c15062 1931 782 7.68e-16
c15063 3672 822 2.4e-16
c15064 687 1466 2.65e-16
c15065 3140 0 3.6368e-14
c15066 852 26 1.58e-16
c15067 3366 3367 9.13e-16
c15068 911 1690 7.6e-16
c15069 2747 3261 4.97e-16
c15070 3048 3155 5.42e-16
c15071 3024 3143 1.58e-16
c15072 426 450 1.88e-16
c15073 4759 4766 1.81e-16
c15074 5198 5158 5.69e-16
c15075 3409 3468 3.92e-16
c15076 657 2265 3.79e-16
c15077 1994 1992 1.6e-16
c15078 1989 1988 2.03e-16
c15079 37 200 1.88e-16
c15080 30 209 3.84e-16
c15081 3706 3409 3.92e-16
c15082 3783 3773 1.58e-16
c15083 3772 3774 9.16e-16
c15084 4356 707 1.84e-16
c15085 1148 797 1.58e-16
c15086 966 973 7.95e-16
c15087 3381 3384 1.576e-15
c15088 4232 4234 1.862e-15
c15089 5044 149 1.96e-16
c15090 1644 842 1.832e-15
c15091 3898 4468 3.92e-16
c15092 3923 1 6.78e-16
c15093 4101 19 9.67e-16
c15094 2651 3160 7.84e-16
c15095 1420 1 4.41e-15
c15096 82 1 2.87e-16
c15097 479 194 1.88e-16
c15098 5103 5114 1.619e-15
c15099 4455 792 1.58e-16
c15100 5318 323 3.54e-16
c15101 4967 4950 1.96e-16
c15102 3462 3066 1.96e-16
c15103 3457 3072 1.96e-16
c15104 103 117 1.58e-16
c15105 2542 1 3.358e-15
c15106 5230 149 1.58e-16
c15107 5262 5241 2.85e-16
c15108 994 995 7.51e-16
c15109 398 1 1.607e-15
c15110 378 15 5.8e-16
c15111 4523 868 1.58e-16
c15112 5577 5576 2.49e-16
c15113 612 3421 1.58e-16
c15114 2869 2867 1.6e-16
c15115 3900 4285 1.58e-16
c15116 2713 2322 1.136e-15
c15117 2535 2554 1.58e-16
c15118 2559 2555 3.92e-16
c15119 3676 0 3.3874e-14
c15120 617 3876 4.48e-16
c15121 1667 1668 3.01e-16
c15122 189 194 1.88e-16
c15123 3024 662 4.48e-16
c15124 2206 2204 1.862e-15
c15125 2082 2078 1.583e-15
c15126 1755 0 1.4092e-14
c15127 982 963 1.546e-15
c15128 5536 497 1.58e-16
c15129 3127 0 6.62e-16
c15130 920 868 3.15e-16
c15131 5403 5475 4.25e-16
c15132 4810 149 5.88e-16
c15133 2654 2666 2.32e-16
c15134 922 1055 3.92e-16
c15135 1523 1086 3.92e-16
c15136 1527 1528 1.6e-16
c15137 1331 971 5.5e-16
c15138 4075 1 6.66e-16
c15139 3046 2764 5.5e-16
c15140 3746 0 1.65e-16
c15141 2651 702 5.73e-16
c15142 3034 2600 1.58e-16
c15143 2557 837 3.15e-16
c15144 1733 0 1.6491e-14
c15145 3393 3410 5.63e-16
c15146 3525 3526 1.6e-16
c15147 3521 3140 3.92e-16
c15148 2157 1 5.01e-16
c15149 344 340 1.372e-15
c15150 3772 3773 1.96e-16
c15151 5269 1 3.36e-16
c15152 5200 0 4.4446e-14
c15153 2535 2350 5.5e-16
c15154 2170 2534 1.62e-16
c15155 537 262 1.88e-16
c15156 3882 4421 1.58e-16
c15157 3898 4433 1.58e-16
c15158 2954 2973 7.95e-16
c15159 2618 647 1.339e-15
c15160 1403 1786 7.84e-16
c15161 2535 2717 1.58e-16
c15162 2557 2705 1.58e-16
c15163 2987 1 4.67e-15
c15164 4056 25 7.01e-16
c15165 1708 1986 3.92e-16
c15166 1542 0 3.3555e-14
c15167 3599 1 5.97e-15
c15168 4673 4293 1.96e-16
c15169 662 678 1.621e-15
c15170 37 346 5.71e-16
c15171 117 247 1.88e-16
c15172 4905 4932 2e-16
c15173 2277 1760 2.38e-15
c15174 149 180 1.88e-16
c15175 883 662 6.45e-16
c15176 2866 3034 3.92e-16
c15177 2690 0 3.466e-15
c15178 4580 1 3.69e-16
c15179 4787 468 1.88e-16
c15180 5580 0 1.3804e-14
c15181 4606 497 5.88e-16
c15182 3267 0 8e-16
c15183 1324 1332 3.84e-16
c15184 1316 1317 4.57e-16
c15185 3886 3381 3.54e-16
c15186 1834 732 5.73e-16
c15187 3884 0 4.64e-16
c15188 1327 1521 1.96e-16
c15189 4293 4655 1.58e-16
c15190 4282 4663 5.66e-16
c15191 4669 4660 3.92e-16
c15192 3063 3060 3.01e-16
c15193 3059 3056 6.44e-16
c15194 1858 1856 1.6e-16
c15195 1853 1852 2.03e-16
c15196 5018 4546 3.54e-16
c15197 5017 4978 1.537e-15
c15198 2821 868 5.73e-16
c15199 3339 827 3.64e-16
c15200 2987 2887 6.72e-16
c15201 3048 2730 5.5e-16
c15202 1499 0 6.9481e-14
c15203 1 470 5.698e-15
c15204 4563 4480 5.88e-16
c15205 4571 4486 1.58e-16
c15206 3219 3208 1.58e-16
c15207 4100 857 1.88e-16
c15208 5177 236 1.58e-16
c15209 5160 5162 1.001e-15
c15210 4827 526 1.88e-16
c15211 601 2589 1.58e-16
c15212 2460 1953 2.48e-16
c15213 3781 3855 9.61e-16
c15214 2015 1 1.492e-15
c15215 2172 1681 1.58e-16
c15216 2178 1678 1.58e-16
c15217 1205 842 5.74e-16
c15218 4742 64 1.88e-16
c15219 2755 2757 2.03e-16
c15220 600 1 4.03e-16
c15221 506 37 1.88e-16
c15222 3462 1 8.43e-16
c15223 4471 3633 4.97e-16
c15224 2545 2871 4.63e-16
c15225 2440 782 1.58e-16
c15226 1769 1380 2.386e-15
c15227 1397 1752 1.58e-16
c15228 595 922 3.15e-16
c15229 1680 1 2.346e-15
c15230 1695 0 1.157e-14
c15231 465 513 1.88e-16
c15232 4691 4692 9.93e-16
c15233 2300 1 1.868e-15
c15234 2290 0 2.93e-15
c15235 2080 1 1.3e-16
c15236 2182 1678 3.54e-16
c15237 890 1157 1.96e-16
c15238 2266 1749 1.96e-16
c15239 921 978 1.58e-16
c15240 3321 3710 2.386e-15
c15241 4455 4467 2.32e-16
c15242 4606 5569 5.5e-16
c15243 4600 5561 7.46e-16
c15244 4640 5514 1.596e-15
c15245 3324 3322 1.6e-16
c15246 4006 19 7.04e-16
c15247 4021 0 1.5176e-14
c15248 3881 1 6.056e-15
c15249 3018 3019 1.76e-16
c15250 632 1752 1.58e-16
c15251 1196 1664 5.69e-16
c15252 1708 1951 5.42e-16
c15253 1684 1939 1.58e-16
c15254 1941 1937 1.96e-16
c15255 1694 1781 1.58e-16
c15256 1506 0 1.6491e-14
c15257 3525 3134 4.11e-16
c15258 5058 5047 1.96e-16
c15259 1862 1834 2.64e-16
c15260 3846 3807 1.738e-15
c15261 602 2217 4.81e-16
c15262 275 1 1.073e-15
c15263 4302 672 1.58e-16
c15264 4305 647 1.58e-16
c15265 2652 1 1.716e-15
c15266 909 992 4.35e-16
c15267 907 991 1.88e-16
c15268 890 984 1.58e-16
c15269 3287 3676 2.386e-15
c15270 3685 3679 1.6e-16
c15271 285 19 3.2e-16
c15272 3370 858 1.58e-16
c15273 1788 647 1.9e-16
c15274 1327 752 3.15e-16
c15275 1417 1415 1.6e-16
c15276 1811 707 1.58e-16
c15277 1969 797 1.58e-16
c15278 1236 1 5.107e-15
c15279 1454 1 4.41e-15
c15280 617 1684 4.48e-16
c15281 5198 207 5.5e-16
c15282 2713 737 3.15e-16
c15283 1838 0 6.62e-16
c15284 216 19 3.84e-16
c15285 421 310 1.88e-16
c15286 236 33 3.08e-16
c15287 2447 1 2.054e-15
c15288 1023 672 1.58e-16
c15289 2741 2350 4.11e-16
c15290 612 2567 1.58e-16
c15291 2449 0 8e-16
c15292 792 2436 2.65e-16
c15293 902 908 3.54e-16
c15294 159 9 6.48e-16
c15295 152 1 5.62e-16
c15296 3734 3785 2.45e-16
c15297 1508 722 1.832e-15
c15298 922 1113 1.58e-16
c15299 1331 1457 1.58e-16
c15300 3390 1 8.766e-15
c15301 617 1398 3.64e-16
c15302 3701 3882 5.88e-16
c15303 3707 3876 1.58e-16
c15304 2504 868 2.65e-16
c15305 1981 827 3.15e-16
c15306 762 1098 1.05e-15
c15307 2787 3294 3.92e-16
c15308 3299 3298 1.6e-16
c15309 3233 737 1.09e-16
c15310 4714 0 1.4233e-14
c15311 0 308 9.795e-15
c15312 4567 4643 1.58e-16
c15313 4571 4259 5.5e-16
c15314 338 332 5.8e-16
c15315 383 352 1.88e-16
c15316 1186 1187 1.238e-15
c15317 1177 837 1.58e-16
c15318 883 1098 3.54e-16
c15319 894 1119 1.58e-16
c15320 986 984 1.931e-15
c15321 5426 5425 1.334e-15
c15322 5388 5366 1.58e-16
c15323 4569 1 4.325e-15
c15324 165 59 1.88e-16
c15325 1483 1041 1.96e-16
c15326 1484 1477 6.73e-16
c15327 687 592 5.8e-16
c15328 4539 4541 1.6e-16
c15329 3973 1 7.71e-16
c15330 1896 752 3.15e-16
c15331 601 1737 1.9e-16
c15332 1485 1 1.056e-15
c15333 1694 1522 1.58e-16
c15334 822 1136 1.58e-16
c15335 4523 0 3.3627e-14
c15336 192 191 6.67e-16
c15337 3100 3492 2.38e-15
c15338 3900 762 3.58e-16
c15339 5010 4930 1.58e-16
c15340 4881 1 4.623e-15
c15341 13 12 3.84e-16
c15342 2619 2621 2.03e-16
c15343 5253 5200 3.18e-16
c15344 4702 526 1.88e-16
c15345 2194 1981 5.5e-16
c15346 966 971 1.58e-16
c15347 4787 64 1.88e-16
c15348 3177 0 3.3874e-14
c15349 1218 1219 1.21e-16
c15350 893 0 1.5977e-14
c15351 4352 3520 2.48e-16
c15352 1343 1146 1.58e-16
c15353 4339 1 2.054e-15
c15354 476 484 1.58e-16
c15355 4341 0 8e-16
c15356 3030 3360 1.96e-16
c15357 4876 4497 1.58e-16
c15358 4870 1 6.42e-16
c15359 421 339 1.88e-16
c15360 4702 4697 1.536e-15
c15361 4793 4418 4.9e-16
c15362 5229 5198 1.58e-16
c15363 1017 647 4.98e-16
c15364 807 809 5.59e-16
c15365 3781 3770 1.211e-15
c15366 3958 3957 3.15e-16
c15367 1218 852 1.58e-16
c15368 47 1 3.6e-16
c15369 5482 5296 2.24e-16
c15370 642 982 1.58e-16
c15371 4197 857 2.573e-15
c15372 1550 782 3.15e-16
c15373 1551 1545 1.6e-16
c15374 1091 1542 2.386e-15
c15375 1106 1525 1.58e-16
c15376 4598 4592 7.25e-16
c15377 3870 3873 1.099e-15
c15378 687 1031 3.79e-16
c15379 1080 1 3.06e-16
c15380 3718 3752 1.466e-15
c15381 4155 1 6.78e-16
c15382 1981 812 1.58e-16
c15383 1805 1801 1.96e-16
c15384 4144 0 1.35812e-13
c15385 4862 4480 1.443e-15
c15386 4794 4795 2.03e-16
c15387 2036 2108 3.54e-16
c15388 1161 1 4.044e-15
c15389 3393 3117 5.88e-16
c15390 4776 4784 1.81e-16
c15391 1611 0 6.62e-16
c15392 3174 3557 7.84e-16
c15393 523 509 1.58e-16
c15394 0 334 9.2601e-14
c15395 37 303 1.88e-16
c15396 3411 672 3.58e-16
c15397 4708 352 1.88e-16
c15398 1681 0 4.4783e-14
c15399 3713 842 1.58e-16
c15400 3853 3855 2.861e-15
c15401 5388 5300 1.237e-15
c15402 5296 5299 1.817e-15
c15403 1170 797 6.48e-16
c15404 687 693 1.097e-15
c15405 3870 3871 1.76e-16
c15406 5320 5323 3.54e-16
c15407 601 591 1.74e-16
c15408 64 62 3.84e-16
c15409 687 4336 1.58e-16
c15410 3876 4485 3.92e-16
c15411 2992 2873 1.52e-16
c15412 4514 4520 1.52e-15
c15413 2559 2769 3.92e-16
c15414 612 4232 1.58e-16
c15415 595 4236 2.72e-16
c15416 4423 3582 4.11e-16
c15417 2662 3172 1.58e-16
c15418 1631 1629 1.6e-16
c15419 1626 1625 2.03e-16
c15420 1690 1850 1.96e-16
c15421 4487 0 1.6491e-14
c15422 4903 4967 1.6e-16
c15423 3030 868 4.03e-16
c15424 3046 827 4.46e-16
c15425 1954 1 1.716e-15
c15426 3411 3242 1.58e-16
c15427 4149 4143 7.45e-16
c15428 4634 5473 1.96e-16
c15429 612 3441 1.58e-16
c15430 2821 0 3.5142e-14
c15431 1116 1118 7.72e-16
c15432 3141 0 1.6491e-14
c15433 2535 2169 1.58e-16
c15434 2541 2166 1.58e-16
c15435 2018 842 4.81e-16
c15436 4309 1 8.43e-16
c15437 3099 2577 1.96e-16
c15438 3094 2583 1.96e-16
c15439 1887 1888 2.48e-16
c15440 3030 3325 1.58e-16
c15441 1 208 4.92e-16
c15442 3397 3066 5.5e-16
c15443 4640 4265 4.9e-16
c15444 4582 4361 5.5e-16
c15445 5412 1 3.986e-15
c15446 4872 439 1.88e-16
c15447 2356 1 4.41e-15
c15448 877 1358 2.38e-15
c15449 2778 2775 3.01e-16
c15450 2774 2771 6.44e-16
c15451 2003 827 1.58e-16
c15452 3674 0 1.6491e-14
c15453 3757 1 7.49e-16
c15454 4508 4509 1.6e-16
c15455 4504 3673 3.92e-16
c15456 602 1322 5.18e-16
c15457 3024 2781 5.5e-16
c15458 4378 4765 2.196e-15
c15459 3186 702 2.65e-16
c15460 2078 2067 1.211e-15
c15461 0 439 1.21385e-13
c15462 890 868 3.35e-16
c15463 907 827 4.8e-16
c15464 2291 2303 2.32e-16
c15465 3889 3885 1.71e-16
c15466 2559 2367 5.5e-16
c15467 919 702 3.15e-16
c15468 957 953 3.31e-16
c15469 1438 1001 1.532e-15
c15470 3898 4438 1.58e-16
c15471 3876 4450 1.58e-16
c15472 3016 2929 1.6e-16
c15473 2635 672 1.58e-16
c15474 632 921 3.15e-16
c15475 2559 2734 5.42e-16
c15476 2535 2722 1.58e-16
c15477 1029 0 2.7206e-14
c15478 1701 1687 6.4e-16
c15479 1689 1695 2.267e-15
c15480 4310 4673 1.96e-16
c15481 1954 1965 1.96e-16
c15482 5096 5034 6.67e-16
c15483 3046 812 4.46e-16
c15484 762 1708 3.58e-16
c15485 88 25 5.71e-16
c15486 2710 0 8e-16
c15487 1678 2168 4.65e-16
c15488 1070 692 1.58e-16
c15489 3747 3749 3.92e-16
c15490 996 1423 7.84e-16
c15491 2178 762 4.03e-16
c15492 4076 3918 2.87e-16
c15493 3673 842 1.75e-16
c15494 3283 0 6.72e-16
c15495 2764 777 3.79e-16
c15496 3120 1 1.056e-15
c15497 612 3046 3.15e-16
c15498 602 3048 3.15e-16
c15499 1328 1346 1.94e-16
c15500 810 1 1.65e-16
c15501 2368 732 2.65e-16
c15502 1249 1263 9.34e-16
c15503 4315 3480 1.96e-16
c15504 4293 4672 1.58e-16
c15505 1376 0 6.72e-16
c15506 3021 3421 7.84e-16
c15507 1482 1850 1.96e-16
c15508 262 255 3.54e-16
c15509 4905 4907 1.001e-15
c15510 3356 868 2.65e-16
c15511 2832 827 3.15e-16
c15512 2281 1760 1.96e-16
c15513 1718 1 5.808e-15
c15514 4563 4497 5.88e-16
c15515 4571 4503 1.58e-16
c15516 2045 2044 1.334e-15
c15517 4821 352 1.88e-16
c15518 2458 2469 1.58e-16
c15519 627 2603 1.58e-16
c15520 617 2589 1.84e-16
c15521 2182 762 7.99e-16
c15522 2172 2393 1.58e-16
c15523 2824 2836 2.32e-16
c15524 2194 1682 5.5e-16
c15525 4304 3469 1.96e-16
c15526 4309 3463 1.96e-16
c15527 4770 5207 7.87e-16
c15528 2541 2503 4.3e-16
c15529 1327 1520 1.58e-16
c15530 397 393 1.58e-16
c15531 4047 1 5.284e-15
c15532 2921 2920 1.96e-16
c15533 1147 0 1.8851e-14
c15534 3330 2821 7.84e-16
c15535 1728 1 9.28e-16
c15536 2713 3237 4.36e-16
c15537 3370 3377 3.96e-16
c15538 3171 677 4.81e-16
c15539 1794 1 5.97e-15
c15540 2044 2054 1.96e-16
c15541 1 342 1.44e-16
c15542 822 1936 5.73e-16
c15543 3818 3773 3.18e-16
c15544 1194 827 8.3e-16
c15545 1201 868 1.35e-16
c15546 907 812 4.8e-16
c15547 883 1172 3.92e-16
c15548 890 1171 1.88e-16
c15549 5459 5457 3.92e-16
c15550 5356 5355 3.92e-16
c15551 2856 0 1.6491e-14
c15552 2666 2282 1.58e-16
c15553 3898 3897 1.009e-15
c15554 3438 0 3.3874e-14
c15555 2736 1 4.41e-15
c15556 632 4298 1.58e-16
c15557 2545 2870 1.58e-16
c15558 1767 1380 1.532e-15
c15559 1773 1772 5.65e-16
c15560 612 907 3.15e-16
c15561 602 909 3.15e-16
c15562 3397 1 4.57e-15
c15563 2713 3230 4.11e-16
c15564 3156 662 1.58e-16
c15565 2030 2028 3.54e-16
c15566 19 255 8.82e-16
c15567 612 1682 1.813e-15
c15568 894 1007 3.92e-16
c15569 909 1006 1.88e-16
c15570 883 999 1.58e-16
c15571 592 933 1.96e-16
c15572 1270 1218 1.246e-15
c15573 765 1 1.65e-16
c15574 3394 3027 1.939e-15
c15575 3233 3230 3.01e-16
c15576 3229 3226 6.44e-16
c15577 2353 707 4.81e-16
c15578 1845 692 1.58e-16
c15579 632 1750 1.339e-15
c15580 3614 1 6.15e-16
c15581 1578 1574 1.96e-16
c15582 3145 2628 4.11e-16
c15583 3519 3134 1.96e-16
c15584 687 2317 2.65e-16
c15585 1863 1 1.868e-15
c15586 4910 4897 1.96e-16
c15587 2832 812 1.58e-16
c15588 1853 0 2.93e-15
c15589 1 128 4.59e-16
c15590 15 135 6.58e-16
c15591 412 30 3.84e-16
c15592 3387 3552 1.58e-16
c15593 3679 3680 5.65e-16
c15594 3287 3674 1.532e-15
c15595 2469 1 5.97e-15
c15596 3598 3589 3.46e-16
c15597 2465 0 6.72e-16
c15598 126 0 2.87e-16
c15599 5136 5049 4.2e-16
c15600 792 1930 3.79e-16
c15601 1278 1276 4.11e-16
c15602 5535 5546 1.33e-15
c15603 4844 381 1.88e-16
c15604 1567 807 1.813e-15
c15605 1345 1031 5.5e-16
c15606 506 523 1.138e-15
c15607 1119 1 2.972e-15
c15608 2690 707 5.03e-16
c15609 2495 858 1.58e-16
c15610 1998 868 3.79e-16
c15611 1818 1829 1.96e-16
c15612 4171 25 4.68e-16
c15613 1752 1751 2.48e-16
c15614 1120 0 6.29e-16
c15615 777 1118 1.58e-16
c15616 4839 4841 1.6e-16
c15617 1641 1684 1.58e-16
c15618 1635 1690 5.88e-16
c15619 85 71 3.84e-16
c15620 3202 3587 1.96e-16
c15621 4557 1 1.44e-16
c15622 4731 0 1.4233e-14
c15623 45 43 1.58e-16
c15624 27 21 1.58e-16
c15625 0 18 6.224e-15
c15626 4567 4660 1.58e-16
c15627 4571 4276 5.5e-16
c15628 2436 1919 1.96e-16
c15629 2437 2430 6.73e-16
c15630 5365 0 3.4847e-14
c15631 62 122 3.45e-16
c15632 2817 1 9.28e-16
c15633 996 998 7.72e-16
c15634 5352 5353 3.54e-16
c15635 1499 707 1.58e-16
c15636 1046 1041 1.58e-16
c15637 3030 0 3.5714e-13
c15638 4166 19 7.04e-16
c15639 617 4268 1.832e-15
c15640 3616 3605 1.58e-16
c15641 2918 2930 1.027e-15
c15642 910 920 1.58e-16
c15643 936 1 4.22e-16
c15644 3295 2781 4.97e-16
c15645 2696 3207 1.96e-16
c15646 617 1737 5.03e-16
c15647 1501 1 9.28e-16
c15648 3718 3886 3.92e-16
c15649 3882 1 2.824e-15
c15650 2867 858 7.68e-16
c15651 1921 1923 2.03e-16
c15652 5184 1 7.87e-16
c15653 2010 1 2.054e-15
c15654 2012 0 8e-16
c15655 5025 120 7.34e-16
c15656 5039 122 3.19e-16
c15657 5360 5350 1.125e-15
c15658 238 0 5.6676e-14
c15659 5417 410 4.02e-16
c15660 4821 294 1.88e-16
c15661 2620 0 3.358e-14
c15662 2172 1998 5.5e-16
c15663 2041 2042 3.18e-16
c15664 1574 807 1.58e-16
c15665 1415 971 4.36e-16
c15666 3197 0 1.4092e-14
c15667 1218 922 1.58e-16
c15668 2545 2633 4.63e-16
c15669 1321 1161 1.58e-16
c15670 1327 1151 5.88e-16
c15671 720 1 1.65e-16
c15672 3118 2600 1.96e-16
c15673 3119 3112 6.73e-16
c15674 2775 767 1.9e-16
c15675 4489 822 1.58e-16
c15676 4357 0 6.72e-16
c15677 3548 747 1.58e-16
c15678 2987 2896 1.58e-16
c15679 910 1681 3.75e-16
c15680 579 577 7.1e-16
c15681 570 580 1.88e-16
c15682 4887 1 6.42e-16
c15683 4881 4890 3.92e-16
c15684 4915 33 1.88e-16
c15685 2256 2258 2.03e-16
c15686 223 508 1.88e-16
c15687 281 334 1.88e-16
c15688 2316 2322 1.418e-15
c15689 1998 2512 1.885e-15
c15690 882 904 2.07e-16
c15691 5482 0 3.0503e-14
c15692 3900 722 3.15e-16
c15693 2041 0 2.1139e-14
c15694 2535 2390 1.58e-16
c15695 676 19 1.96e-16
c15696 3168 0 6.9481e-14
c15697 3874 3873 1.58e-16
c15698 3684 4523 2.386e-15
c15699 4532 4526 1.6e-16
c15700 627 1369 1.58e-16
c15701 890 0 3.53121e-13
c15702 1094 1 3.06e-16
c15703 3046 2651 1.58e-16
c15704 1636 1 1.868e-15
c15705 4793 4798 5.53e-16
c15706 687 2265 1.58e-16
c15707 1626 0 2.93e-15
c15708 3185 3569 1.58e-16
c15709 2393 0 3.3248e-14
c15710 722 714 1.74e-16
c15711 33 553 6.01e-16
c15712 3393 677 3.15e-16
c15713 3962 3960 7.1e-16
c15714 4563 4605 1.96e-16
c15715 5335 1 1.257e-15
c15716 5299 0 3.5057e-14
c15717 3327 852 5.73e-16
c15718 4262 4260 1.6e-16
c15719 3544 0 6.72e-16
c15720 2220 2603 7.84e-16
c15721 1464 1455 3.46e-16
c15722 612 619 1.6e-16
c15723 3900 4502 3.92e-16
c15724 3046 747 3.15e-16
c15725 1690 1335 3.15e-16
c15726 3925 0 1.5176e-14
c15727 3186 3180 1.6e-16
c15728 2662 3177 2.386e-15
c15729 2679 3160 1.58e-16
c15730 1999 1990 3.92e-16
c15731 1607 1993 5.66e-16
c15732 1706 1867 3.92e-16
c15733 117 455 1.88e-16
c15734 493 491 7.1e-16
c15735 478 477 5.8e-16
c15736 497 499 3.84e-16
c15737 3474 3083 4.11e-16
c15738 3024 852 3.15e-16
c15739 2211 0 8e-16
c15740 1980 1 8.43e-16
c15741 3387 3253 5.5e-16
c15742 101 102 1.88e-16
c15743 4058 4056 7.1e-16
c15744 3886 858 3.15e-16
c15745 4685 381 1.88e-16
c15746 1121 1098 6.54e-16
c15747 3882 3463 5.88e-16
c15748 3876 3469 1.58e-16
c15749 3582 4417 1.96e-16
c15750 1315 1727 4.36e-16
c15751 2274 662 1.58e-16
c15752 859 0 8.558e-15
c15753 822 824 5.59e-16
c15754 1690 1849 1.58e-16
c15755 986 0 7.4292e-14
c15756 76 0 9.795e-15
c15757 3046 3342 1.58e-16
c15758 3030 3330 1.58e-16
c15759 592 817 1.96e-16
c15760 1652 2095 7.46e-16
c15761 2072 2031 2.45e-16
c15762 3411 797 3.15e-16
c15763 4582 4378 5.5e-16
c15764 2196 2474 3.92e-16
c15765 3728 3732 6.9e-16
c15766 881 1340 2.79e-16
c15767 2178 2269 1.58e-16
c15768 4329 4322 6.73e-16
c15769 4447 782 7.68e-16
c15770 5482 5486 1.96e-16
c15771 4872 5136 7.46e-16
c15772 2674 2671 5.5e-16
c15773 3090 3093 6.44e-16
c15774 2921 2976 3.18e-16
c15775 2646 662 7.68e-16
c15776 1601 1146 1.136e-15
c15777 747 907 3.15e-16
c15778 3048 2798 5.5e-16
c15779 3177 707 1.58e-16
c15780 2679 702 3.79e-16
c15781 2080 2070 1.58e-16
c15782 5190 5199 2.177e-15
c15783 3538 3151 1.532e-15
c15784 5025 5098 2.02e-16
c15785 2389 1879 1.96e-16
c15786 2196 1749 1.58e-16
c15787 2182 2269 1.58e-16
c15788 883 852 3.15e-16
c15789 5136 0 5.8438e-14
c15790 4355 692 1.9e-16
c15791 920 707 3.69e-16
c15792 971 974 6.13e-16
c15793 1327 952 1.58e-16
c15794 3667 4505 4.97e-16
c15795 2639 662 5.03e-16
c15796 657 920 3.15e-16
c15797 2559 2739 1.58e-16
c15798 3839 3373 5.5e-16
c15799 4072 37 5.71e-16
c15800 3245 3252 1.96e-16
c15801 3048 2628 5.5e-16
c15802 3030 3122 1.96e-16
c15803 4762 4761 2.48e-16
c15804 4765 4766 2.83e-16
c15805 4461 1 6.15e-16
c15806 4690 4310 1.96e-16
c15807 2820 812 7.38e-16
c15808 323 321 6.01e-16
c15809 303 317 3.84e-16
c15810 5074 5071 7.46e-16
c15811 1690 1 2.824e-15
c15812 692 686 1.74e-16
c15813 3549 707 7.68e-16
c15814 642 2535 3.15e-16
c15815 2294 2301 6.73e-16
c15816 894 702 8.34e-16
c15817 3397 3225 1.58e-16
c15818 2726 0 6.72e-16
c15819 858 866 5.58e-16
c15820 4580 4531 3.92e-16
c15821 1431 672 3.79e-16
c15822 1345 807 3.58e-16
c15823 2194 777 3.15e-16
c15824 4095 3918 8.1e-16
c15825 627 3046 3.15e-16
c15826 601 3048 3.15e-16
c15827 820 1 3.79e-16
c15828 3565 4399 1.58e-16
c15829 2359 737 1.58e-16
c15830 3659 1 5.808e-15
c15831 3857 0 3.792e-15
c15832 1591 1602 1.96e-16
c15833 1345 1538 3.92e-16
c15834 813 0 7.86e-15
c15835 4310 4672 1.58e-16
c15836 4686 4677 3.92e-16
c15837 3259 792 1.58e-16
c15838 3022 3433 1.58e-16
c15839 601 1743 1.58e-16
c15840 761 760 6.67e-16
c15841 4974 4978 6.22e-16
c15842 410 470 3.45e-16
c15843 3248 767 1.84e-16
c15844 1738 1 2.054e-15
c15845 3411 3604 3.92e-16
c15846 1066 717 1.35e-16
c15847 592 772 1.96e-16
c15848 3618 3617 1.6e-16
c15849 1998 0 7.0008e-14
c15850 3327 3409 1.58e-16
c15851 5435 1 3.36e-16
c15852 4793 0 3.03219e-13
c15853 2477 1964 4.97e-16
c15854 2172 1726 5.5e-16
c15855 3648 1 6.15e-16
c15856 1708 722 3.15e-16
c15857 1343 1537 1.58e-16
c15858 1327 1525 1.58e-16
c15859 2532 3058 7.84e-16
c15860 2731 722 3.64e-16
c15861 1863 1854 3.92e-16
c15862 1471 1857 5.66e-16
c15863 1482 1849 1.58e-16
c15864 4249 0 1.6491e-14
c15865 2178 722 3.15e-16
c15866 3342 2832 1.58e-16
c15867 3606 3615 3.46e-16
c15868 2336 1 1.056e-15
c15869 15 494 5.8e-16
c15870 245 253 2.218e-15
c15871 128 131 1.099e-15
c15872 468 30 3.84e-16
c15873 2461 2473 2.32e-16
c15874 2470 822 2.65e-16
c15875 0 482 9.795e-15
c15876 3219 767 1.58e-16
c15877 2549 2186 3.84e-16
c15878 88 9 5.8e-16
c15879 71 1 5.175e-15
c15880 4708 5347 3.92e-16
c15881 4691 5286 5.87e-16
c15882 3003 2503 1.66e-16
c15883 2876 1 1.23e-16
c15884 2767 2765 1.6e-16
c15885 883 1186 1.88e-16
c15886 907 1179 1.58e-16
c15887 2305 1 4.41e-15
c15888 602 2545 3.15e-16
c15889 4199 4204 1.96e-16
c15890 2671 2282 2.386e-15
c15891 1888 752 1.58e-16
c15892 1331 1320 1.58e-16
c15893 3458 0 1.4092e-14
c15894 3271 1 1.868e-15
c15895 4038 1 7.08e-16
c15896 4475 4472 5.5e-16
c15897 2418 797 3.15e-16
c15898 2182 722 3.15e-16
c15899 911 1326 1.58e-16
c15900 627 907 3.15e-16
c15901 601 909 3.15e-16
c15902 3328 2821 3.92e-16
c15903 4022 37 1.88e-16
c15904 4031 25 4.68e-16
c15905 3030 3087 1.58e-16
c15906 1706 1573 1.58e-16
c15907 762 1101 4e-16
c15908 33 178 2.2e-16
c15909 5066 5067 8.03e-16
c15910 627 1682 1.58e-16
c15911 3333 842 1.84e-16
c15912 2257 1777 1.58e-16
c15913 767 1127 1.58e-16
c15914 894 1021 1.58e-16
c15915 907 993 3.54e-16
c15916 59 484 1.88e-16
c15917 4878 5104 3.65e-16
c15918 4107 4102 1.96e-16
c15919 2541 2667 1.96e-16
c15920 775 1 3.79e-16
c15921 3890 1 8.822e-15
c15922 1694 858 3.15e-16
c15923 1331 1343 4.369e-15
c15924 1673 1327 6.89e-16
c15925 768 0 7.86e-15
c15926 361 378 1.325e-15
c15927 537 223 1.88e-16
c15928 3409 762 3.15e-16
c15929 3129 3126 5.5e-16
c15930 3900 822 3.58e-16
c15931 687 1811 3.79e-16
c15932 3396 3394 3.67e-16
c15933 1482 1 5.97e-15
c15934 5398 5385 8.94e-16
c15935 762 1886 1.58e-16
c15936 245 37 1.88e-16
c15937 3387 3557 1.58e-16
c15938 3411 3569 5.42e-16
c15939 3393 3174 1.58e-16
c15940 3860 858 6.67e-16
c15941 5575 1 1.546e-15
c15942 2538 2546 3.84e-16
c15943 592 727 1.96e-16
c15944 4164 3879 2.573e-15
c15945 5403 468 7.38e-16
c15946 910 3030 7.97e-16
c15947 911 3046 9.54e-16
c15948 2814 2807 1.96e-16
c15949 4400 737 7.38e-16
c15950 5440 5444 1.088e-15
c15951 2529 0 4.79e-14
c15952 2742 2741 1.6e-16
c15953 3139 2628 1.96e-16
c15954 1959 812 1.84e-16
c15955 4208 1 4.997e-15
c15956 4361 3520 1.136e-15
c15957 2710 707 1.09e-16
c15958 1211 1206 1.58e-16
c15959 4198 0 1.5061e-14
c15960 4200 19 3.45e-16
c15961 3316 3317 5.65e-16
c15962 602 2582 1.58e-16
c15963 1 249 4.22e-16
c15964 4567 4677 1.58e-16
c15965 4571 4293 5.5e-16
c15966 5034 91 1.58e-16
c15967 4827 207 1.88e-16
c15968 1930 1919 1.58e-16
c15969 0 251 1.5723e-14
c15970 151 30 3.84e-16
c15971 5412 5409 7.84e-16
c15972 5446 5448 3.25e-16
c15973 2830 1 6.15e-16
c15974 1016 672 3.79e-16
c15975 1001 647 3.15e-16
c15976 1173 1187 1.96e-16
c15977 395 407 1.58e-16
c15978 2248 2633 1.96e-16
c15979 1046 1500 4.36e-16
c15980 1498 1491 1.96e-16
c15981 2944 2929 1.96e-16
c15982 953 1 3.54e-16
c15983 1756 1754 1.6e-16
c15984 1751 1750 2.03e-16
c15985 3048 3023 2.38e-16
c15986 3024 3020 3.54e-16
c15987 617 1757 1.09e-16
c15988 1662 0 6.78e-16
c15989 3126 647 1.832e-15
c15990 5157 5187 9.6e-16
c15991 425 419 5.8e-16
c15992 334 332 1.88e-16
c15993 441 439 3.84e-16
c15994 2358 1851 2.48e-16
c15995 4531 4881 2e-16
c15996 390 9 5.8e-16
c15997 223 216 7.76e-16
c15998 234 233 7.03e-16
c15999 4736 0 4.02382e-13
c16000 4080 4078 1.76e-16
c16001 2919 2917 3.25e-16
c16002 911 907 8.02e-16
c16003 910 890 5.75e-16
c16004 3980 25 1.88e-16
c16005 3976 19 7.35e-16
c16006 4369 3531 4.97e-16
c16007 1196 1640 1.96e-16
c16008 1345 1176 1.58e-16
c16009 1343 1166 5.5e-16
c16010 1331 1639 1.58e-16
c16011 930 0 3.36e-16
c16012 730 1 3.79e-16
c16013 723 0 7.86e-15
c16014 1558 1560 2.03e-16
c16015 1550 1522 2.64e-16
c16016 1221 0 1.8572e-14
c16017 2892 2882 1.58e-16
c16018 911 1682 1.88e-16
c16019 716 715 6.67e-16
c16020 3498 662 7.68e-16
c16021 2156 2153 1.6e-16
c16022 1 63 4.92e-16
c16023 12 27 3.84e-16
c16024 11 0 9.795e-15
c16025 3397 3518 1.58e-16
c16026 5010 149 1.88e-16
c16027 2618 0 1.6491e-14
c16028 632 3455 1.58e-16
c16029 2178 2338 1.96e-16
c16030 1218 1234 3.98e-16
c16031 78 421 1.88e-16
c16032 4353 4365 2.32e-16
c16033 2559 2407 1.58e-16
c16034 689 25 1.13e-15
c16035 693 19 1.58e-16
c16036 1937 797 1.339e-15
c16037 4242 3873 2.64e-16
c16038 4615 4609 7.25e-16
c16039 3874 4231 9.42e-16
c16040 2559 3017 3.54e-16
c16041 2535 2541 4.078e-15
c16042 4883 4884 2.4e-16
c16043 4879 4497 1.479e-15
c16044 4156 26 4.58e-16
c16045 3024 2668 1.58e-16
c16046 3030 2662 5.88e-16
c16047 2036 2133 7.46e-16
c16048 5230 5226 5.7e-16
c16049 3185 3574 2.386e-15
c16050 3583 3577 1.6e-16
c16051 0 509 1.051e-14
c16052 25 523 5.71e-16
c16053 294 297 4.6e-16
c16054 3672 797 1.58e-16
c16055 4563 4622 1.96e-16
c16056 2417 2408 3.46e-16
c16057 2182 2338 4.63e-16
c16058 79 15 4.88e-16
c16059 5345 0 1.963e-15
c16060 1726 0 6.9048e-14
c16061 73 0 2.5552e-14
c16062 59 44 1.88e-16
c16063 52 19 8.82e-16
c16064 56 37 5.71e-16
c16065 64 30 7.67e-16
c16066 3851 2899 9.75e-16
c16067 3531 722 1.58e-16
c16068 2231 2615 1.58e-16
c16069 1470 1469 9.1e-16
c16070 3010 3001 7.53e-16
c16071 4139 25 4.68e-16
c16072 601 4253 1.9e-16
c16073 4445 4436 3.46e-16
c16074 2535 732 3.15e-16
c16075 1777 1783 1.418e-15
c16076 1684 1884 3.92e-16
c16077 527 524 6.67e-16
c16078 505 508 1.099e-15
c16079 25 317 7.06e-16
c16080 2227 0 6.72e-16
c16081 788 787 1.96e-16
c16082 3191 732 1.58e-16
c16083 5104 1 9.493e-15
c16084 3411 3270 5.5e-16
c16085 1732 2240 7.84e-16
c16086 907 879 1.88e-16
c16087 883 882 1.58e-16
c16088 3321 3712 4.11e-16
c16089 2220 2601 3.92e-16
c16090 2606 2605 1.6e-16
c16091 4567 4582 4.274e-15
c16092 5585 4563 1.96e-16
c16093 3160 1 5.808e-15
c16094 2559 2773 1.58e-16
c16095 1578 782 1.9e-16
c16096 1319 1680 1.58e-16
c16097 2785 2786 9.1e-16
c16098 2559 2170 5.5e-16
c16099 2294 662 1.58e-16
c16100 1636 1627 3.92e-16
c16101 1176 1630 5.66e-16
c16102 671 1 5.57e-16
c16103 3180 3181 5.65e-16
c16104 1706 1866 1.58e-16
c16105 1690 1854 1.58e-16
c16106 3083 3468 1.96e-16
c16107 2769 752 1.58e-16
c16108 822 1708 3.58e-16
c16109 762 922 3.15e-16
c16110 5048 120 7.94e-16
c16111 4915 526 1.88e-16
c16112 3030 707 3.15e-16
c16113 1956 0 3.3633e-14
c16114 3242 3628 5.66e-16
c16115 3634 3625 3.92e-16
c16116 592 637 1.96e-16
c16117 4582 4395 5.5e-16
c16118 5450 1 1.021e-15
c16119 2493 1981 1.532e-15
c16120 2499 2498 5.65e-16
c16121 2178 822 4.03e-16
c16122 2781 822 1.58e-16
c16123 657 3030 4.03e-16
c16124 881 880 2.45e-16
c16125 3943 3942 1.58e-16
c16126 5493 0 2.078e-15
c16127 2194 2286 1.58e-16
c16128 2178 2274 1.58e-16
c16129 3616 767 3.15e-16
c16130 3038 2549 3.84e-16
c16131 2272 662 1.339e-15
c16132 1345 1572 3.92e-16
c16133 822 829 1.6e-16
c16134 3532 1 1.868e-15
c16135 4305 0 1.4092e-14
c16136 5414 528 1.345e-15
c16137 2663 672 2.65e-16
c16138 3369 3366 1.6e-16
c16139 1786 1 5.808e-15
c16140 1788 0 3.466e-15
c16141 3625 3627 2.15e-16
c16142 4395 4782 2.196e-15
c16143 3393 3467 1.58e-16
c16144 3197 707 1.58e-16
c16145 2541 858 3.15e-16
c16146 657 2620 1.58e-16
c16147 418 436 1.58e-16
c16148 1 204 4.22e-16
c16149 2182 822 7.99e-16
c16150 2196 2473 5.42e-16
c16151 5131 5135 8.88e-16
c16152 777 2384 1.813e-15
c16153 2182 2274 1.58e-16
c16154 3765 3774 1.873e-15
c16155 2311 2308 5.5e-16
c16156 2858 2475 7.84e-16
c16157 2671 2678 1.96e-16
c16158 4233 3381 4.97e-16
c16159 1343 966 1.58e-16
c16160 2584 2170 1.532e-15
c16161 1649 842 1.09e-16
c16162 702 1 4.1542e-14
c16163 3882 3622 1.58e-16
c16164 2656 672 2.72e-16
c16165 822 1172 2.68e-16
c16166 1043 0 1.4198e-14
c16167 3632 3623 3.46e-16
c16168 4470 1 1.716e-15
c16169 2559 692 3.15e-16
c16170 1980 1584 1.96e-16
c16171 1975 1590 1.96e-16
c16172 1131 0 3.7577e-14
c16173 37 419 1.88e-16
c16174 5100 5103 3.54e-16
c16175 5126 5125 1.6e-16
c16176 332 345 1.58e-16
c16177 3559 717 2.72e-16
c16178 3168 707 3.15e-16
c16179 3693 3692 2.48e-16
c16180 4952 4950 7.82e-16
c16181 890 707 3.15e-16
c16182 907 1067 3.92e-16
c16183 105 117 1.58e-16
c16184 5303 5302 1.062e-15
c16185 2768 2401 1.58e-16
c16186 2170 2585 4.97e-16
c16187 687 3140 1.58e-16
c16188 2804 1 4.41e-15
c16189 1823 677 1.58e-16
c16190 657 890 3.35e-16
c16191 4031 4022 1.96e-16
c16192 3314 0 6.62e-16
c16193 3124 1 1.716e-15
c16194 617 3048 3.15e-16
c16195 2172 792 3.15e-16
c16196 4534 842 4.81e-16
c16197 839 1 7.18e-16
c16198 3582 4387 1.58e-16
c16199 2367 752 3.15e-16
c16200 3679 1 2.054e-15
c16201 4310 4689 1.58e-16
c16202 981 1 4.044e-15
c16203 595 1343 3.15e-16
c16204 602 1327 3.15e-16
c16205 1407 0 6.62e-16
c16206 3447 3441 1.6e-16
c16207 3022 3438 2.386e-15
c16208 3066 3421 1.58e-16
c16209 632 2249 7.68e-16
c16210 617 1743 3.15e-16
c16211 1641 1642 1.35e-16
c16212 3034 2787 1.58e-16
c16213 3034 677 3.15e-16
c16214 1678 2205 4.97e-16
c16215 1920 0 1.6491e-14
c16216 777 1925 1.58e-16
c16217 5575 4950 5.95e-16
c16218 2194 1902 1.58e-16
c16219 4519 827 1.58e-16
c16220 2844 2841 5.5e-16
c16221 3657 1 1.716e-15
c16222 4319 3480 2.386e-15
c16223 392 59 1.88e-16
c16224 2533 3070 1.58e-16
c16225 1693 1335 5.8e-16
c16226 1707 1324 3.54e-16
c16227 1529 1527 1.6e-16
c16228 1524 1523 2.03e-16
c16229 1331 1367 1.58e-16
c16230 1482 1854 1.58e-16
c16231 4071 1 6.03e-16
c16232 2172 737 4.48e-16
c16233 4811 1 1.806e-15
c16234 1742 1 8.43e-16
c16235 3387 3386 1.58e-16
c16236 2352 1 9.28e-16
c16237 1964 822 3.79e-16
c16238 3527 3525 1.6e-16
c16239 3253 752 1.58e-16
c16240 2322 0 3.583e-14
c16241 3693 3338 1.58e-16
c16242 3765 3773 3.54e-16
c16243 4434 752 1.58e-16
c16244 1026 677 2.33e-16
c16245 3885 3887 3.84e-16
c16246 601 2545 3.15e-16
c16247 4349 677 1.58e-16
c16248 2839 2458 3.92e-16
c16249 1908 752 1.58e-16
c16250 4570 4577 2.07e-16
c16251 657 986 1.813e-15
c16252 2923 2933 7.84e-16
c16253 2952 2949 1.099e-15
c16254 617 909 3.15e-16
c16255 807 19 1.41e-15
c16256 3886 3582 5.5e-16
c16257 2425 807 1.58e-16
c16258 1785 1786 2.48e-16
c16259 1017 0 6.29e-16
c16260 3373 1 1.286e-15
c16261 3240 3241 9.1e-16
c16262 3046 3104 1.58e-16
c16263 3030 3092 1.58e-16
c16264 1545 1 2.054e-15
c16265 1684 1590 1.58e-16
c16266 1690 1584 5.88e-16
c16267 4596 0 6.72e-16
c16268 1547 0 8e-16
c16269 5158 236 4.44e-16
c16270 5252 1 3.36e-16
c16271 2374 1868 3.92e-16
c16272 2378 2379 1.6e-16
c16273 2196 2236 3.92e-16
c16274 743 742 1.96e-16
c16275 4944 4992 3.09e-16
c16276 910 2529 1.58e-16
c16277 909 1008 3.54e-16
c16278 2669 2282 1.532e-15
c16279 4117 4118 3.15e-16
c16280 1161 837 5.73e-16
c16281 3869 1 9.43e-16
c16282 4391 4390 5.65e-16
c16283 4385 3548 1.532e-15
c16284 2557 2684 3.92e-16
c16285 3889 0 6.35e-16
c16286 1899 1 1.056e-15
c16287 3536 677 1.58e-16
c16288 1 456 1.607e-15
c16289 3411 3574 1.58e-16
c16290 3397 3587 4.63e-16
c16291 2542 2560 1.94e-16
c16292 2540 2546 2.267e-15
c16293 4108 4102 1.96e-16
c16294 5136 5083 9.01e-16
c16295 1534 752 7.68e-16
c16296 5558 5529 1.58e-16
c16297 597 1 1.65e-16
c16298 506 0 4.6186e-14
c16299 1844 1448 1.96e-16
c16300 1839 1454 1.96e-16
c16301 1341 0 1.2366e-14
c16302 3034 3241 4.63e-16
c16303 1693 1 2.56e-15
c16304 601 2582 7.38e-16
c16305 1 175 4.22e-16
c16306 125 0 2.87e-16
c16307 122 30 3.84e-16
c16308 3409 722 4.46e-16
c16309 4567 4694 1.58e-16
c16310 4571 4310 5.5e-16
c16311 1930 2453 4.36e-16
c16312 2451 2444 1.96e-16
c16313 5556 5529 6.31e-16
c16314 378 455 1.88e-16
c16315 3804 3811 8.96e-16
c16316 3836 3739 7.46e-16
c16317 5388 5170 4.35e-16
c16318 3001 2486 1.477e-15
c16319 2839 1 1.716e-15
c16320 921 995 1.96e-16
c16321 3719 3327 1.96e-16
c16322 3421 1 5.808e-15
c16323 529 524 1.059e-15
c16324 506 514 2.218e-15
c16325 3423 0 3.466e-15
c16326 3839 3781 1.58e-16
c16327 4182 37 1.88e-16
c16328 4191 25 4.68e-16
c16329 4029 1 6.78e-16
c16330 3898 4383 3.92e-16
c16331 4457 4455 2.15e-16
c16332 4465 4464 1.6e-16
c16333 1380 1748 1.96e-16
c16334 3143 672 1.58e-16
c16335 1515 1 8.43e-16
c16336 4214 0 4.393e-14
c16337 5036 5031 3.73e-16
c16338 1328 886 1.939e-15
c16339 277 9 4.88e-16
c16340 268 1 5.62e-16
c16341 5355 5365 2.114e-15
c16342 4844 5086 1.96e-16
c16343 3749 3750 1.6e-16
c16344 4199 3918 2.48e-16
c16345 1136 797 3.15e-16
c16346 1595 807 2.72e-16
c16347 1146 1149 1.58e-16
c16348 632 4266 1.339e-15
c16349 3990 37 1.88e-16
c16350 3999 25 4.68e-16
c16351 2557 2649 1.58e-16
c16352 2541 2637 1.58e-16
c16353 1933 1931 1.6e-16
c16354 647 640 5.58e-16
c16355 30 585 6.83e-16
c16356 204 363 1.88e-16
c16357 4899 4914 3.25e-16
c16358 4900 4897 6.71e-16
c16359 224 15 4.88e-16
c16360 3397 3523 1.58e-16
c16361 3287 3655 1.96e-16
c16362 226 19 8.82e-16
c16363 5546 1 3.91e-16
c16364 632 3475 1.58e-16
c16365 792 0 2.85894e-13
c16366 1392 1389 5.5e-16
c16367 927 929 9.05e-16
c16368 3799 3798 1.6e-16
c16369 4047 857 1.88e-16
c16370 2194 2355 3.92e-16
c16371 1513 722 1.09e-16
c16372 59 276 1.88e-16
c16373 3633 807 1.813e-15
c16374 2803 2802 9.1e-16
c16375 1211 1248 4.41e-16
c16376 922 1130 3.92e-16
c16377 3109 2628 1.58e-16
c16378 4242 4231 1.58e-16
c16379 3591 762 1.58e-16
c16380 3701 4543 5.69e-16
c16381 3048 2685 1.58e-16
c16382 3046 2679 5.5e-16
c16383 3034 3206 1.58e-16
c16384 1654 1 9.28e-16
c16385 762 1115 1.85e-16
c16386 1706 1652 3.92e-16
c16387 662 672 3.28e-16
c16388 233 508 1.88e-16
c16389 4716 0 8e-16
c16390 0 311 1.0822e-14
c16391 3387 692 4.48e-16
c16392 4563 4639 1.96e-16
c16393 4922 439 1.88e-16
c16394 2423 2422 9.1e-16
c16395 3980 3988 6.67e-16
c16396 3986 3976 7.1e-16
c16397 5437 5436 1.6e-16
c16398 632 3411 3.15e-16
c16399 4270 4271 1.6e-16
c16400 4266 3435 3.92e-16
c16401 919 943 1.58e-16
c16402 3575 0 6.62e-16
c16403 2629 2623 1.6e-16
c16404 2231 2620 2.386e-15
c16405 1476 1472 1.96e-16
c16406 2299 662 1.58e-16
c16407 737 0 2.80402e-13
c16408 2907 2895 1.96e-16
c16409 617 4253 5.03e-16
c16410 2373 767 1.75e-16
c16411 1718 1319 1.58e-16
c16412 3969 0 5.617e-15
c16413 4526 1 2.054e-15
c16414 1708 1901 3.92e-16
c16415 465 451 1.58e-16
c16416 479 455 1.88e-16
c16417 3577 3578 5.65e-16
c16418 4563 4621 1.58e-16
c16419 2196 1817 1.58e-16
c16420 901 893 1.611e-15
c16421 3496 3487 3.46e-16
c16422 4528 0 8e-16
c16423 6 9 6.48e-16
c16424 8 13 1.58e-16
c16425 2603 1 5.808e-15
c16426 617 3072 2.33e-16
c16427 3180 1 2.054e-15
c16428 4606 64 1.88e-16
c16429 4327 4707 1.96e-16
c16430 2824 827 1.58e-16
c16431 1684 1883 1.58e-16
c16432 1706 1871 1.58e-16
c16433 1240 1 5.18e-16
c16434 1708 1703 1.58e-16
c16435 535 576 3.1e-16
c16436 2334 1817 1.96e-16
c16437 777 919 3.15e-16
c16438 3048 3347 1.58e-16
c16439 1732 2238 3.92e-16
c16440 2243 2242 1.6e-16
c16441 1976 0 1.4092e-14
c16442 3253 3625 1.58e-16
c16443 4469 0 3.563e-14
c16444 9 523 5.8e-16
c16445 3397 837 7.99e-16
c16446 4060 4062 2.254e-15
c16447 4582 4412 5.5e-16
c16448 4838 323 1.88e-16
c16449 1572 782 7.38e-16
c16450 1321 702 3.15e-16
c16451 2172 2303 1.58e-16
c16452 2194 2291 1.58e-16
c16453 5511 5517 6.23e-16
c16454 2979 1 3.36e-16
c16455 4343 4336 1.96e-16
c16456 3497 4345 4.36e-16
c16457 3151 1 5.97e-15
c16458 3293 822 1.58e-16
c16459 4148 1 6.78e-16
c16460 2955 2041 2.24e-16
c16461 2654 677 1.58e-16
c16462 4869 4866 3.01e-16
c16463 3271 3262 3.92e-16
c16464 2753 3265 5.66e-16
c16465 3393 3472 1.58e-16
c16466 3409 3089 1.58e-16
c16467 2103 2100 3.54e-16
c16468 2072 2119 3.18e-16
c16469 2196 2478 1.58e-16
c16470 523 511 1.58e-16
c16471 0 303 4.4191e-14
c16472 4582 4585 1.6e-16
c16473 5290 412 7.97e-16
c16474 762 1885 1.58e-16
c16475 2215 1 1.868e-15
c16476 707 723 1.621e-15
c16477 383 30 3.84e-16
c16478 1041 717 5.73e-16
c16479 894 907 4.452e-15
c16480 922 722 5.14e-16
c16481 921 1053 1.58e-16
c16482 4366 717 2.4e-16
c16483 1321 981 1.58e-16
c16484 661 25 7.64e-16
c16485 2756 777 1.58e-16
c16486 602 877 1.58e-16
c16487 612 880 5.73e-16
c16488 687 920 3.15e-16
c16489 868 25 1.58e-16
c16490 3898 3639 1.58e-16
c16491 2469 837 3.79e-16
c16492 4124 26 4.58e-16
c16493 3048 3139 3.92e-16
c16494 747 1096 1.35e-16
c16495 4779 4778 2.48e-16
c16496 4782 4783 2.83e-16
c16497 3003 858 9.97e-16
c16498 3014 852 3.64e-16
c16499 657 2618 1.58e-16
c16500 2100 2101 3.54e-16
c16501 4496 1 8.43e-16
c16502 1749 1750 1.35e-16
c16503 551 549 7.1e-16
c16504 310 204 1.88e-16
c16505 2402 2396 1.6e-16
c16506 1879 2393 2.386e-15
c16507 1885 2401 1.136e-15
c16508 1896 2376 1.58e-16
c16509 2197 1 2.86e-16
c16510 3387 3393 4.078e-15
c16511 5062 1 1.88e-16
c16512 2308 2315 1.96e-16
c16513 4821 5047 9.04e-16
c16514 2678 2669 3.46e-16
c16515 5283 5300 1.443e-15
c16516 2872 352 8.6e-16
c16517 2757 0 6.62e-16
c16518 2567 1 1.716e-15
c16519 3731 3748 1.287e-15
c16520 3339 1 1.868e-15
c16521 3329 0 2.93e-15
c16522 3150 1 8.43e-16
c16523 1355 1357 2.15e-16
c16524 3361 0 1.6878e-14
c16525 1617 1151 1.96e-16
c16526 1612 1161 1.96e-16
c16527 601 1327 3.15e-16
c16528 4316 4697 5.66e-16
c16529 4703 4694 3.92e-16
c16530 2824 812 1.832e-15
c16531 1694 1437 1.58e-16
c16532 3287 792 2.22e-16
c16533 2739 752 1.58e-16
c16534 363 175 1.88e-16
c16535 3553 717 2.4e-16
c16536 4972 4975 1.099e-15
c16537 2753 782 1.75e-16
c16538 2556 1 2.94e-16
c16539 1053 717 1.05e-15
c16540 2548 0 6.35e-16
c16541 461 448 1.58e-16
c16542 4640 4644 1.81e-16
c16543 4634 439 1.364e-15
c16544 2172 1919 1.58e-16
c16545 2178 1913 5.88e-16
c16546 1362 1353 3.46e-16
c16547 3882 837 4.03e-16
c16548 2545 2544 1.357e-15
c16549 922 1188 1.58e-16
c16550 639 1 5.57e-16
c16551 3683 1 8.43e-16
c16552 3409 822 3.15e-16
c16553 1345 1542 1.58e-16
c16554 4581 3879 3.54e-16
c16555 3084 3078 1.6e-16
c16556 2533 3075 2.386e-15
c16557 2577 3058 1.58e-16
c16558 1482 1874 2.38e-15
c16559 4092 1 4.64e-16
c16560 4510 4508 1.6e-16
c16561 4828 1 1.806e-15
c16562 3411 3018 1.58e-16
c16563 2365 1 6.15e-16
c16564 2082 2086 1.96e-16
c16565 1 436 4.22e-16
c16566 407 484 1.88e-16
c16567 4617 4612 1.536e-15
c16568 5461 1 1.257e-15
c16569 4674 33 1.88e-16
c16570 2481 2478 5.5e-16
c16571 2182 1913 5.5e-16
c16572 5425 0 3.5057e-14
c16573 3781 3858 8.32e-16
c16574 3900 672 3.58e-16
c16575 687 3141 1.58e-16
c16576 883 1173 3.54e-16
c16577 894 1194 1.58e-16
c16578 617 2545 3.15e-16
c16579 5356 5358 1.96e-16
c16580 616 25 7.64e-16
c16581 2955 2949 2.08e-16
c16582 3345 2832 1.532e-15
c16583 1936 797 2.33e-16
c16584 1635 2003 1.96e-16
c16585 1708 1607 1.58e-16
c16586 1706 1601 5.5e-16
c16587 1694 2002 1.58e-16
c16588 4613 0 6.72e-16
c16589 1952 1567 1.96e-16
c16590 19 477 3.84e-16
c16591 339 204 1.88e-16
c16592 5071 5069 1.373e-15
c16593 2133 1 1.81e-16
c16594 3907 3909 4.33e-16
c16595 2286 2287 9.1e-16
c16596 1134 1141 2.27e-16
c16597 2572 2569 5.5e-16
c16598 2873 2911 9.37e-16
c16599 1636 837 2.65e-16
c16600 1422 1423 2.48e-16
c16601 1016 1435 1.58e-16
c16602 910 1341 1.58e-16
c16603 1335 1326 5.71e-16
c16604 657 4305 1.58e-16
c16605 3898 4417 3.92e-16
c16606 4036 37 1.88e-16
c16607 2535 2701 3.92e-16
c16608 1499 1056 1.136e-15
c16609 657 1788 2.72e-16
c16610 1369 1 4.41e-15
c16611 250 262 1.58e-16
c16612 246 247 1.88e-16
c16613 4421 777 1.58e-16
c16614 3420 3421 2.48e-16
c16615 2987 2521 5.5e-16
c16616 1915 1 9.28e-16
c16617 1981 1 5.97e-15
c16618 1058 692 3.57e-16
c16619 1038 1051 1.58e-16
c16620 4007 4015 9.33e-16
c16621 4008 4006 3.54e-16
c16622 1091 737 3.15e-16
c16623 2834 2833 1.6e-16
c16624 2826 2824 2.15e-16
c16625 687 1029 1.58e-16
c16626 537 233 1.88e-16
c16627 4232 1 1.716e-15
c16628 1155 1 3.06e-16
c16629 3401 3410 1.846e-15
c16630 4219 19 7.35e-16
c16631 3330 3329 2.48e-16
c16632 3692 3691 2.03e-16
c16633 3697 3695 1.6e-16
c16634 2044 2042 3.92e-16
c16635 1 349 4.22e-16
c16636 5173 5157 2.109e-15
c16637 4838 265 1.88e-16
c16638 953 955 7.84e-16
c16639 5262 0 5.8479e-14
c16640 2194 2179 1.632e-15
c16641 2178 2195 5.63e-16
c16642 3582 732 2.22e-16
c16643 4404 737 1.832e-15
c16644 2865 1 8.43e-16
c16645 1436 647 1.58e-16
c16646 1193 1194 1.213e-15
c16647 3463 4297 1.58e-16
c16648 920 1009 1.58e-16
c16649 3983 1338 2.697e-15
c16650 3441 1 2.054e-15
c16651 3443 0 8e-16
c16652 2521 2015 1.96e-16
c16653 3509 3123 5.66e-16
c16654 2429 782 1.9e-16
c16655 651 640 7.23e-16
c16656 4361 4333 2.64e-16
c16657 3034 2532 1.58e-16
c16658 2023 2028 1.078e-15
c16659 4674 4680 5.87e-16
c16660 2083 1 1.257e-15
c16661 310 175 1.88e-16
c16662 160 49 1.88e-16
c16663 2044 0 3.7361e-14
c16664 401 400 1.58e-16
c16665 642 648 1.097e-15
c16666 632 622 6.38e-16
c16667 2136 2078 1.58e-16
c16668 3392 0 4.3741e-14
c16669 2322 707 2.33e-16
c16670 642 1765 2.4e-16
c16671 1326 1 6.056e-15
c16672 3548 1 5.97e-15
c16673 1694 1765 4.63e-16
c16674 451 450 1.079e-15
c16675 5005 1 1.88e-16
c16676 4930 4918 1.96e-16
c16677 4902 4889 4.53e-16
c16678 2257 1743 2.386e-15
c16679 1760 2240 1.58e-16
c16680 233 216 1.138e-15
c16681 1047 677 4.98e-16
c16682 413 0 1.4515e-14
c16683 287 291 1.58e-16
c16684 3639 3640 1.35e-16
c16685 3338 842 3.15e-16
c16686 4855 33 1.88e-16
c16687 902 927 3.53e-16
c16688 4475 812 1.84e-16
c16689 5540 5532 3.54e-16
c16690 5514 5511 7.46e-16
c16691 3230 0 3.466e-15
c16692 1221 1226 1.58e-16
c16693 4373 4370 5.5e-16
c16694 1690 837 4.03e-16
c16695 1958 797 1.9e-16
c16696 1570 1568 1.6e-16
c16697 1327 1470 1.96e-16
c16698 3589 0 1.6491e-14
c16699 4259 4231 2.64e-16
c16700 4632 4626 7.25e-16
c16701 4242 4248 9.42e-16
c16702 1684 1352 1.58e-16
c16703 1690 1319 5.5e-16
c16704 2475 852 5.73e-16
c16705 1816 1431 1.96e-16
c16706 822 922 3.15e-16
c16707 4906 4907 5.87e-16
c16708 3024 2696 5.5e-16
c16709 3034 3211 1.58e-16
c16710 1659 1 1.886e-15
c16711 236 296 3.45e-16
c16712 1635 2154 5.69e-16
c16713 1 5 5.175e-15
c16714 0 25 5.6444e-13
c16715 4733 0 8e-16
c16716 41 44 1.099e-15
c16717 28 31 6.01e-16
c16718 4038 857 1.88e-16
c16719 4563 4656 1.96e-16
c16720 5366 1 2.424e-15
c16721 2424 2418 1.418e-15
c16722 602 2555 1.58e-16
c16723 2407 2435 2.64e-16
c16724 1919 0 3.6368e-14
c16725 2429 2425 1.96e-16
c16726 927 928 8.05e-16
c16727 1327 886 1.96e-16
c16728 1243 1266 7.5e-16
c16729 1708 672 3.58e-16
c16730 3590 0 2.93e-15
c16731 3046 1 4.77e-16
c16732 3839 3748 1.58e-16
c16733 4543 4545 1.6e-16
c16734 2880 2879 3.92e-16
c16735 1104 0 2.7376e-14
c16736 3781 1 5.966e-15
c16737 617 4273 1.09e-16
c16738 2178 672 4.03e-16
c16739 2194 647 4.46e-16
c16740 1738 1319 2.38e-15
c16741 2106 1667 1.679e-15
c16742 2144 1249 1.573e-15
c16743 4543 1 1.871e-15
c16744 291 274 1.138e-15
c16745 4563 4638 1.58e-16
c16746 732 738 1.097e-15
c16747 4542 0 3.792e-15
c16748 2258 0 6.62e-16
c16749 0 568 9.795e-15
c16750 339 175 1.88e-16
c16751 3809 3807 5.88e-16
c16752 3858 3853 2.029e-15
c16753 2342 2345 5.5e-16
c16754 42 44 1.88e-16
c16755 2316 2714 4.36e-16
c16756 5326 5321 7.37e-16
c16757 5360 5359 5.87e-16
c16758 2623 1 2.054e-15
c16759 2231 2618 1.532e-15
c16760 2623 2624 5.65e-16
c16761 1136 1139 6.13e-16
c16762 4668 5517 5.5e-16
c16763 2880 2877 1.96e-16
c16764 2182 672 7.99e-16
c16765 2713 747 1.813e-15
c16766 3944 25 6.96e-16
c16767 4344 4707 1.96e-16
c16768 3194 3193 2.48e-16
c16769 2844 827 1.58e-16
c16770 2841 868 1.58e-16
c16771 1708 1900 5.42e-16
c16772 1684 1888 1.58e-16
c16773 3111 3107 1.96e-16
c16774 1455 0 1.6491e-14
c16775 4435 4436 1.35e-16
c16776 1828 1817 1.58e-16
c16777 570 569 3.84e-16
c16778 3486 672 1.58e-16
c16779 5106 31 1.58e-16
c16780 3191 3192 1.35e-16
c16781 2601 1 1.716e-15
c16782 890 901 1.96e-16
c16783 3253 3645 2.38e-15
c16784 3761 3734 2.84e-16
c16785 4208 857 1.88e-16
c16786 4582 4429 5.5e-16
c16787 5450 410 1.58e-16
c16788 687 3030 4.03e-16
c16789 2520 1998 1.96e-16
c16790 2517 2515 1.6e-16
c16791 1382 1381 1.6e-16
c16792 1374 1372 2.15e-16
c16793 2172 2308 1.58e-16
c16794 3958 3918 2.48e-16
c16795 2995 1 1.672e-15
c16796 1800 677 2.33e-16
c16797 3568 1 1.056e-15
c16798 3151 2634 1.136e-15
c16799 2759 767 1.84e-16
c16800 907 1 6e-16
c16801 2674 677 1.58e-16
c16802 777 894 8.34e-16
c16803 911 2173 2.09e-16
c16804 4412 4799 2.196e-15
c16805 3203 722 7.68e-16
c16806 2396 1 2.054e-15
c16807 596 655 2.45e-16
c16808 5452 0 4.4446e-14
c16809 5300 1 2.386e-15
c16810 4827 497 1.88e-16
c16811 2398 0 8e-16
c16812 1682 1 5.277e-15
c16813 1500 717 2.65e-16
c16814 617 3073 1.339e-15
c16815 2688 2690 2.15e-16
c16816 1456 1458 2.03e-16
c16817 601 877 1.58e-16
c16818 3751 3749 1.186e-15
c16819 3882 3650 5.88e-16
c16820 3876 3656 1.58e-16
c16821 4521 4522 2.03e-16
c16822 2849 3367 5.69e-16
c16823 3933 1 6.78e-16
c16824 3271 3260 1.96e-16
c16825 1992 1601 4.11e-16
c16826 304 320 3.84e-16
c16827 30 210 6.83e-16
c16828 468 499 1.88e-16
c16829 3555 3556 2.03e-16
c16830 3559 3561 1.6e-16
c16831 5106 5149 1.489e-15
c16832 2201 0 2.96e-16
c16833 552 570 1.88e-16
c16834 3555 722 1.339e-15
c16835 894 1082 3.92e-16
c16836 909 1081 1.88e-16
c16837 883 1074 1.58e-16
c16838 4237 4234 5.5e-16
c16839 5262 5253 2.85e-16
c16840 687 3168 2.22e-16
c16841 2832 1 5.97e-15
c16842 1829 692 7.68e-16
c16843 1438 1440 1.862e-15
c16844 687 890 3.35e-16
c16845 392 407 1.88e-16
c16846 361 404 1.88e-16
c16847 3909 1 7.44e-16
c16848 4102 25 3.84e-16
c16849 3882 3480 5.88e-16
c16850 2385 752 7.68e-16
c16851 1434 1 1.056e-15
c16852 617 1327 3.15e-16
c16853 90 1 4.92e-16
c16854 4472 0 3.3551e-14
c16855 4586 4581 9.6e-16
c16856 1001 0 7.4113e-14
c16857 369 368 6.96e-16
c16858 332 346 3.84e-16
c16859 352 354 1.96e-16
c16860 349 363 1.88e-16
c16861 2315 2306 3.46e-16
c16862 3288 782 3.64e-16
c16863 617 2248 1.58e-16
c16864 2563 0 1.23e-16
c16865 223 218 1.88e-16
c16866 4657 4659 4.93e-16
c16867 2194 1930 5.5e-16
c16868 391 9 6.48e-16
c16869 5577 5575 2.861e-15
c16870 5403 5476 1.03e-16
c16871 3126 0 3.3874e-14
c16872 2557 2542 1.632e-15
c16873 2541 2558 5.63e-16
c16874 4321 4317 1.96e-16
c16875 1803 1420 7.84e-16
c16876 2737 752 1.339e-15
c16877 1667 1664 8.32e-16
c16878 1194 1 2.972e-15
c16879 1195 0 6.29e-16
c16880 3030 3309 1.96e-16
c16881 4845 1 1.806e-15
c16882 4915 207 1.88e-16
c16883 984 991 2.27e-16
c16884 596 610 2.45e-16
c16885 5514 497 1.96e-16
c16886 5044 1 1.113e-15
c16887 3503 3504 1.35e-16
c16888 5483 5481 5.25e-16
c16889 1046 677 3.57e-16
c16890 1914 767 7.68e-16
c16891 1534 1525 3.92e-16
c16892 1086 1528 5.66e-16
c16893 2282 677 3.15e-16
c16894 1930 812 1.58e-16
c16895 4072 0 2.0592e-14
c16896 3048 3109 1.58e-16
c16897 2089 2062 5.87e-16
c16898 2064 2066 6.87e-16
c16899 1116 1 4.044e-15
c16900 1560 0 6.62e-16
c16901 3151 3518 1.58e-16
c16902 3140 3526 5.66e-16
c16903 3532 3523 3.92e-16
c16904 4630 0 6.72e-16
c16905 2154 1 1.871e-15
c16906 5230 1 9.493e-15
c16907 2153 0 3.792e-15
c16908 1128 767 1.58e-16
c16909 911 880 4.62e-16
c16910 3876 4434 3.92e-16
c16911 3853 1 1.886e-15
c16912 2559 2718 3.92e-16
c16913 792 790 3.327e-15
c16914 1690 1799 1.96e-16
c16915 4436 0 1.6491e-14
c16916 3523 702 1.58e-16
c16917 4441 777 1.58e-16
c16918 4943 4948 3.07e-16
c16919 5001 4991 1.96e-16
c16920 166 164 1.58e-16
c16921 3387 3208 1.58e-16
c16922 2866 3380 1.58e-16
c16923 2527 1 8e-16
c16924 1058 1059 1.213e-15
c16925 852 860 1.6e-16
c16926 4810 1 2.7943e-14
c16927 4702 497 1.88e-16
c16928 3898 3384 1.58e-16
c16929 3900 797 3.15e-16
c16930 5569 5514 1.383e-15
c16931 2756 2755 2.48e-16
c16932 595 905 3.03e-16
c16933 1331 1076 5.5e-16
c16934 4258 1 8.43e-16
c16935 3057 3058 2.48e-16
c16936 1856 1465 4.11e-16
c16937 1169 1 3.06e-16
c16938 4546 5011 3.92e-16
c16939 5013 5007 6.23e-16
c16940 3046 3257 1.58e-16
c16941 3030 3245 1.58e-16
c16942 2177 2183 2.267e-15
c16943 480 0 1.051e-14
c16944 1 500 5.62e-16
c16945 3393 752 3.15e-16
c16946 3899 3390 3.54e-16
c16947 5160 5184 1.96e-16
c16948 5051 5034 2.2e-16
c16949 4674 526 1.88e-16
c16950 2471 2470 1.6e-16
c16951 2463 2461 2.15e-16
c16952 3706 3705 9.1e-16
c16953 2308 0 3.3692e-14
c16954 3091 0 2.93e-15
c16955 108 15 4.88e-16
c16956 4770 5209 1.96e-16
c16957 590 0 1.1415e-14
c16958 367 369 1.58e-16
c16959 3623 0 1.6491e-14
c16960 4200 4199 1.58e-16
c16961 1331 1332 1.027e-15
c16962 3459 0 6.72e-16
c16963 4470 4481 1.96e-16
c16964 3334 3332 1.6e-16
c16965 3329 3328 2.03e-16
c16966 4361 4350 1.58e-16
c16967 1 180 5.798e-15
c16968 465 508 1.88e-16
c16969 4691 4694 6.02e-16
c16970 294 354 3.45e-16
c16971 647 663 1.621e-15
c16972 19 172 8.4e-16
c16973 64 499 1.88e-16
c16974 1338 898 5.8e-16
c16975 2841 0 3.3717e-14
c16976 1117 1118 7.46e-16
c16977 880 879 3.84e-16
c16978 4191 4182 1.96e-16
c16979 986 1402 1.96e-16
c16980 78 71 7.76e-16
c16981 3898 4387 1.58e-16
c16982 3876 4399 1.58e-16
c16983 4668 5514 7.46e-16
c16984 2887 2889 6.16e-16
c16985 2559 2654 1.58e-16
c16986 4021 19 9.67e-16
c16987 977 0 1.0003e-14
c16988 3887 0 1.157e-14
c16989 3124 3135 1.96e-16
c16990 1511 0 1.4092e-14
c16991 3140 3134 1.418e-15
c16992 1937 1556 3.92e-16
c16993 1941 1942 1.6e-16
c16994 910 25 1.58e-16
c16995 5383 5277 6.31e-16
c16996 911 3025 2.09e-16
c16997 2659 0 8e-16
c16998 245 0 4.1342e-14
c16999 5429 1 9.04e-16
c17000 1403 647 2.33e-16
c17001 4071 857 6.23e-16
c17002 4872 149 1.88e-16
c17003 3069 1 1.056e-15
c17004 1281 1289 6.19e-16
c17005 1817 717 5.73e-16
c17006 1343 1487 3.92e-16
c17007 4259 4248 1.58e-16
c17008 2617 2645 2.64e-16
c17009 1706 1363 5.5e-16
c17010 2514 858 1.58e-16
c17011 2804 837 5.73e-16
c17012 3208 3209 1.35e-16
c17013 1752 1764 2.32e-16
c17014 3387 3536 3.92e-16
c17015 2866 2838 2.64e-16
c17016 837 839 5.59e-16
c17017 596 710 5.28e-16
c17018 4563 4673 1.96e-16
c17019 5529 0 3.359e-14
c17020 595 2169 1.58e-16
c17021 2194 2359 1.58e-16
c17022 159 1 1.073e-15
c17023 3999 3990 1.96e-16
c17024 3053 0 2.96e-16
c17025 149 0 1.20749e-13
c17026 920 782 3.69e-16
c17027 1016 1012 3.78e-16
c17028 4289 4288 5.65e-16
c17029 4283 3446 1.532e-15
c17030 2541 2452 5.88e-16
c17031 1327 1469 1.58e-16
c17032 1380 952 1.136e-15
c17033 3413 1 2.86e-16
c17034 3046 2634 1.58e-16
c17035 1867 722 7.38e-16
c17036 4552 3882 6.89e-16
c17037 3886 3898 4.369e-15
c17038 943 1 3.444e-15
c17039 3296 3305 3.92e-16
c17040 2798 3291 1.58e-16
c17041 1660 1 4.03e-16
c17042 4531 4526 1.642e-15
c17043 2696 2702 1.418e-15
c17044 3131 647 1.09e-16
c17045 1618 2016 4.36e-16
c17046 2014 2007 1.96e-16
c17047 762 1343 3.15e-16
c17048 30 297 6.83e-16
c17049 4563 4655 1.58e-16
c17050 2196 1845 5.5e-16
c17051 339 349 1.88e-16
c17052 4719 1 1.7972e-14
c17053 2866 842 1.58e-16
c17054 2793 792 1.58e-16
c17055 4657 0 3.40595e-13
c17056 617 3100 1.58e-16
c17057 2196 677 3.15e-16
c17058 1742 1319 1.96e-16
c17059 1737 1352 1.96e-16
c17060 3117 3123 1.418e-15
c17061 601 1352 2.33e-16
c17062 595 1363 2.22e-16
c17063 2861 868 1.58e-16
c17064 1708 1905 1.58e-16
c17065 334 262 1.88e-16
c17066 1828 2351 4.36e-16
c17067 3393 3689 1.96e-16
c17068 2627 1 8.43e-16
c17069 777 1 4.1542e-14
c17070 9 0 2.10855e-13
c17071 8 27 1.58e-16
c17072 642 3474 2.72e-16
c17073 4582 4446 5.5e-16
c17074 5240 5239 1.559e-15
c17075 4855 526 1.88e-16
c17076 4702 5321 1.152e-15
c17077 1253 1255 3.92e-16
c17078 4355 4353 2.15e-16
c17079 4363 4362 1.6e-16
c17080 3198 3196 1.6e-16
c17081 1708 797 3.15e-16
c17082 3584 1 9.28e-16
c17083 1952 782 1.58e-16
c17084 1263 1 3.36e-16
c17085 1252 0 1.65e-16
c17086 3364 2855 1.361e-15
c17087 3034 2849 5.5e-16
c17088 2178 797 3.15e-16
c17089 1812 1 1.868e-15
c17090 4886 4883 3.01e-16
c17091 2781 797 3.15e-16
c17092 3298 807 2.72e-16
c17093 4866 0 3.466e-15
c17094 2696 722 3.15e-16
c17095 1802 0 2.93e-15
c17096 1 527 4.92e-16
c17097 3259 3644 1.96e-16
c17098 3253 3649 1.96e-16
c17099 993 647 1.58e-16
c17100 9 564 4.61e-16
c17101 0 511 9.795e-15
c17102 2409 2411 2.03e-16
c17103 1061 702 4.21e-16
c17104 1345 986 5.5e-16
c17105 4595 4592 5.5e-16
c17106 3748 1 2.386e-15
c17107 3886 4518 1.58e-16
c17108 3898 3667 5.5e-16
c17109 3900 3673 1.58e-16
c17110 3701 4519 1.96e-16
c17111 2182 797 3.15e-16
c17112 1805 1806 1.6e-16
c17113 822 1173 1.58e-16
c17114 4437 4439 2.03e-16
c17115 4796 4795 2.48e-16
c17116 4799 4800 2.83e-16
c17117 4412 4803 1.96e-16
c17118 2106 2119 1.96e-16
c17119 3185 3553 1.96e-16
c17120 523 524 7.03e-16
c17121 513 507 3.84e-16
c17122 3409 672 3.15e-16
c17123 2325 2327 2.15e-16
c17124 3338 3411 5.5e-16
c17125 2784 1 1.056e-15
c17126 1172 797 1.58e-16
c17127 894 1096 1.58e-16
c17128 907 1068 3.54e-16
c17129 4370 717 1.58e-16
c17130 2690 2686 1.96e-16
c17131 59 570 1.88e-16
c17132 4150 4143 2.45e-16
c17133 2873 2984 1.58e-16
c17134 1448 692 3.15e-16
c17135 1839 702 2.72e-16
c17136 1644 852 1.58e-16
c17137 3599 3571 2.64e-16
c17138 595 3384 1.58e-16
c17139 3582 3588 1.418e-15
c17140 4419 4421 1.862e-15
c17141 1879 737 3.15e-16
c17142 1629 1166 4.11e-16
c17143 1601 1986 1.96e-16
c17144 1694 1465 5.5e-16
c17145 657 25 1.58e-16
c17146 4492 0 1.4092e-14
c17147 1959 1 2.054e-15
c17148 1961 0 8e-16
c17149 3393 3625 1.58e-16
c17150 3409 3242 1.58e-16
c17151 5229 178 5.5e-16
c17152 5091 0 1.23e-16
c17153 1074 722 1.58e-16
c17154 2569 0 3.3553e-14
c17155 2172 1947 5.5e-16
c17156 1562 767 1.58e-16
c17157 3146 0 1.4092e-14
c17158 2545 2582 4.63e-16
c17159 601 969 8.3e-16
c17160 2271 677 1.75e-16
c17161 2287 647 1.58e-16
c17162 2016 868 2.65e-16
c17163 1618 827 3.15e-16
c17164 1321 1116 1.58e-16
c17165 1327 1106 5.88e-16
c17166 642 1331 7.99e-16
c17167 1897 1505 1.96e-16
c17168 1898 1891 6.73e-16
c17169 366 378 1.58e-16
c17170 4306 0 6.72e-16
c17171 3046 3326 3.92e-16
c17172 5227 178 9.15e-16
c17173 1930 1925 1.642e-15
c17174 9 219 4.88e-16
c17175 4563 4745 1.58e-16
c17176 4580 4757 1.58e-16
c17177 5160 5222 6.67e-16
c17178 3925 3926 3.15e-16
c17179 5410 0 3.0268e-14
c17180 2772 2773 2.48e-16
c17181 2557 2356 1.58e-16
c17182 537 465 1.88e-16
c17183 642 3898 3.15e-16
c17184 1042 1 3.54e-16
c17185 4115 1 6.78e-16
c17186 3673 4509 5.66e-16
c17187 4515 4506 3.92e-16
c17188 2472 812 4.81e-16
c17189 1964 797 1.58e-16
c17190 1039 0 9.602e-15
c17191 3190 692 1.58e-16
c17192 3072 3073 1.35e-16
c17193 1585 1 1.868e-15
c17194 3624 3626 2.03e-16
c17195 632 2616 7.38e-16
c17196 1575 0 2.93e-15
c17197 3151 3523 1.58e-16
c17198 4647 0 6.72e-16
c17199 870 869 1.6e-16
c17200 0 419 4.3431e-14
c17201 5123 5108 6.67e-16
c17202 5098 5100 5.48e-16
c17203 4334 702 1.58e-16
c17204 1147 782 1.58e-16
c17205 1128 1134 1.58e-16
c17206 1816 662 1.58e-16
c17207 1443 1001 2.38e-15
c17208 3003 2929 9.61e-16
c17209 3900 4451 3.92e-16
c17210 3886 4281 4.63e-16
c17211 840 1 1.65e-16
c17212 2809 812 5.03e-16
c17213 1965 1959 1.6e-16
c17214 1567 1956 2.386e-15
c17215 158 164 5.8e-16
c17216 3543 702 1.58e-16
c17217 1249 0 2.1171e-14
c17218 1929 1 8.43e-16
c17219 4759 5157 6.58e-16
c17220 5283 5304 1.6e-16
c17221 4861 236 1.88e-16
c17222 4922 4930 1.072e-15
c17223 4028 4029 6.67e-16
c17224 4078 3918 6.32e-16
c17225 2764 0 6.9021e-14
c17226 2839 2850 1.96e-16
c17227 3882 3385 5.5e-16
c17228 3876 3418 1.58e-16
c17229 1618 812 1.58e-16
c17230 595 932 1.11e-16
c17231 796 19 1.96e-16
c17232 595 3886 9.84e-16
c17233 4384 4385 1.35e-16
c17234 881 0 7.0343e-14
c17235 261 259 7.1e-16
c17236 3024 3274 1.58e-16
c17237 3046 3262 1.58e-16
c17238 2189 2175 6.4e-16
c17239 4469 4849 1.96e-16
c17240 4567 4333 1.58e-16
c17241 967 968 7.46e-16
c17242 4674 5303 1.96e-16
c17243 2328 0 1.4092e-14
c17244 1207 1188 1.546e-15
c17245 146 479 1.88e-16
c17246 5450 5449 2.29e-16
c17247 1515 1061 1.96e-16
c17248 1510 1071 1.96e-16
c17249 657 1001 3.79e-16
c17250 1327 1328 1.239e-15
c17251 4056 1 5.1e-16
c17252 4234 0 3.3555e-14
c17253 2832 3326 1.96e-16
c17254 661 659 5.88e-16
c17255 4378 4350 2.64e-16
c17256 3034 2577 5.5e-16
c17257 2535 807 3.15e-16
c17258 1 343 2.87e-16
c17259 5158 5155 3.54e-16
c17260 4196 0 3.9101e-14
c17261 2306 0 1.6491e-14
c17262 19 345 3.45e-16
c17263 657 3126 1.58e-16
c17264 2544 2186 5.8e-16
c17265 2558 2175 3.54e-16
c17266 2380 2378 1.6e-16
c17267 2375 2374 2.03e-16
c17268 747 2359 1.58e-16
c17269 146 189 1.88e-16
c17270 3721 842 4.81e-16
c17271 5358 5365 1.138e-15
c17272 2861 0 1.4092e-14
c17273 2840 2452 4.97e-16
c17274 922 672 3.15e-16
c17275 919 647 3.15e-16
c17276 3876 3872 3.54e-16
c17277 3882 3899 5.63e-16
c17278 3900 3875 2.38e-16
c17279 3667 3662 1.642e-15
c17280 2136 2103 1.58e-16
c17281 1380 1772 2.38e-15
c17282 2541 2288 1.58e-16
c17283 3228 3226 1.862e-15
c17284 3030 3071 1.96e-16
c17285 3855 0 3.931e-14
c17286 2028 2049 4.41e-16
c17287 4410 1 6.15e-16
c17288 1726 1318 1.136e-15
c17289 25 259 7.06e-16
c17290 33 267 2.68e-16
c17291 4423 762 2.72e-16
c17292 4992 4980 1.697e-15
c17293 3030 782 3.15e-16
c17294 3219 3214 1.642e-15
c17295 1 466 1.456e-15
c17296 4580 4847 1.58e-16
c17297 4571 4859 1.58e-16
c17298 1397 662 1.58e-16
c17299 986 1401 1.58e-16
c17300 2974 2959 6.67e-16
c17301 5538 5540 1.001e-15
c17302 5536 5532 5.7e-16
c17303 3085 1 9.28e-16
c17304 1297 1295 5.5e-16
c17305 2351 717 2.65e-16
c17306 3608 1 5.808e-15
c17307 1574 1131 3.92e-16
c17308 1578 1579 1.6e-16
c17309 751 19 1.96e-16
c17310 529 1 5.62e-16
c17311 542 9 5.8e-16
c17312 4276 4248 2.64e-16
c17313 4649 4643 7.25e-16
c17314 4259 4265 9.42e-16
c17315 1684 1380 5.5e-16
c17316 3225 777 5.73e-16
c17317 2194 868 3.15e-16
c17318 2172 827 4.48e-16
c17319 3339 837 2.65e-16
c17320 1679 1 1.96e-16
c17321 3411 3553 3.92e-16
c17322 4367 1 4.442e-15
c17323 2165 1684 3.54e-16
c17324 276 274 1.88e-16
c17325 273 291 1.58e-16
c17326 1 123 5.62e-16
c17327 9 188 6.48e-16
c17328 3602 3600 1.6e-16
c17329 4563 4690 1.96e-16
c17330 1947 0 6.9481e-14
c17331 4691 381 1.88e-16
c17332 1251 1231 2.45e-16
c17333 1276 1226 2.038e-15
c17334 5356 294 4.44e-16
c17335 2557 2469 5.5e-16
c17336 1343 1486 1.58e-16
c17337 1327 1474 1.58e-16
c17338 146 147 7.03e-16
c17339 1829 1823 1.6e-16
c17340 1431 1820 2.386e-15
c17341 642 1706 3.15e-16
c17342 4016 1 1.895e-14
c17343 4183 37 1.88e-16
c17344 4456 4453 6.44e-16
c17345 4460 4457 3.01e-16
c17346 1755 1762 6.73e-16
c17347 1118 0 1.4198e-14
c17348 4068 2538 2.573e-15
c17349 3296 2798 1.58e-16
c17350 1694 1706 4.369e-15
c17351 2161 1690 6.89e-16
c17352 85 88 3.54e-16
c17353 4576 1 1.002e-15
c17354 2559 767 3.15e-16
c17355 602 2571 1.9e-16
c17356 777 1321 3.15e-16
c17357 752 744 1.74e-16
c17358 50 49 6.96e-16
c17359 19 18 3.2e-16
c17360 479 320 1.88e-16
c17361 4563 4672 1.58e-16
c17362 3208 752 1.75e-16
c17363 3821 3809 1.697e-15
c17364 5277 0 5.7679e-14
c17365 890 782 3.15e-16
c17366 907 1142 3.92e-16
c17367 2732 2731 1.6e-16
c17368 281 9 5.8e-16
c17369 5353 5355 1.387e-15
c17370 2254 1 4.41e-15
c17371 920 923 3.15e-16
c17372 3041 3027 6.4e-16
c17373 1465 732 1.58e-16
c17374 642 966 5.73e-16
c17375 2172 2194 4.078e-15
c17376 642 4281 2.4e-16
c17377 3886 3537 1.58e-16
c17378 2920 2913 8.94e-16
c17379 2931 2932 2.12e-16
c17380 2918 2915 1.732e-15
c17381 3294 3305 1.96e-16
c17382 2545 2248 5.5e-16
c17383 3991 37 1.88e-16
c17384 617 1352 1.75e-16
c17385 1181 1653 4.36e-16
c17386 1651 1644 1.96e-16
c17387 3123 677 1.75e-16
c17388 3595 3593 1.6e-16
c17389 3718 4556 1.58e-16
c17390 4711 4723 2.62e-16
c17391 821 820 6.67e-16
c17392 4400 747 2.4e-16
c17393 5205 207 4.88e-16
c17394 3034 752 3.15e-16
c17395 883 961 1.58e-16
c17396 907 955 1.58e-16
c17397 217 9 6.48e-16
c17398 5277 5349 4.25e-16
c17399 3668 3276 1.96e-16
c17400 4168 4166 3.54e-16
c17401 3763 3767 1.845e-15
c17402 2178 2522 1.96e-16
c17403 1343 722 4.46e-16
c17404 1331 732 7.99e-16
c17405 1387 1398 1.96e-16
c17406 4474 797 1.9e-16
c17407 2559 2282 5.5e-16
c17408 2535 2265 5.5e-16
c17409 3964 25 1.88e-16
c17410 1828 677 1.58e-16
c17411 1331 1623 4.63e-16
c17412 1211 1259 2.31e-16
c17413 706 19 1.96e-16
c17414 3502 3134 1.96e-16
c17415 2747 2742 1.642e-15
c17416 3514 0 6.9481e-14
c17417 2680 692 7.68e-16
c17418 2172 812 4.48e-16
c17419 595 1694 9.84e-16
c17420 569 580 3.84e-16
c17421 4884 1 1.95e-15
c17422 822 1573 5.73e-16
c17423 4429 4816 2.196e-15
c17424 4883 0 3.466e-15
c17425 1670 2139 1.722e-15
c17426 2512 2524 3.13e-16
c17427 2004 2196 1.58e-16
c17428 1902 1 4.41e-15
c17429 662 1012 6.38e-16
c17430 642 3468 2.4e-16
c17431 2411 0 6.62e-16
c17432 612 2172 3.15e-16
c17433 904 905 6.57e-16
c17434 3668 812 7.68e-16
c17435 3310 3695 1.96e-16
c17436 5537 526 3.54e-16
c17437 5388 0 5.8479e-14
c17438 3898 732 3.15e-16
c17439 2788 2790 1.862e-15
c17440 3007 0 6.72e-16
c17441 4267 4266 2.03e-16
c17442 4272 4270 1.6e-16
c17443 5414 5407 9.38e-16
c17444 2478 842 1.58e-16
c17445 1981 837 3.79e-16
c17446 762 1103 1.58e-16
c17447 1092 0 6.29e-16
c17448 2770 3281 1.96e-16
c17449 3207 732 2.4e-16
c17450 616 614 5.88e-16
c17451 3643 3640 6.44e-16
c17452 3647 3644 3.01e-16
c17453 0 540 9.795e-15
c17454 3661 797 1.9e-16
c17455 1913 1885 2.64e-16
c17456 392 252 1.88e-16
c17457 909 1083 3.54e-16
c17458 981 983 7.72e-16
c17459 3362 1 1.886e-15
c17460 2231 2599 1.96e-16
c17461 1468 1466 1.6e-16
c17462 612 616 2.19e-16
c17463 3882 4315 1.96e-16
c17464 3925 19 9.67e-16
c17465 1438 1 1.716e-15
c17466 491 494 3.54e-16
c17467 490 477 1.108e-15
c17468 3083 3089 1.418e-15
c17469 3470 3472 1.862e-15
c17470 3100 3072 2.64e-16
c17471 2327 2323 1.96e-16
c17472 1977 0 6.72e-16
c17473 792 1567 3.79e-16
c17474 1068 1082 1.96e-16
c17475 5325 5316 2.177e-15
c17476 2792 2401 4.11e-16
c17477 2492 2493 1.35e-16
c17478 110 111 1.58e-16
c17479 107 88 1.88e-16
c17480 4556 858 3.15e-16
c17481 4838 381 1.88e-16
c17482 920 1237 2.86e-16
c17483 617 969 1.58e-16
c17484 854 25 1.13e-15
c17485 859 19 1.58e-16
c17486 3907 37 1.88e-16
c17487 2007 858 1.58e-16
c17488 1166 1623 1.96e-16
c17489 1345 1131 1.58e-16
c17490 1343 1121 5.5e-16
c17491 1331 1588 1.58e-16
c17492 2594 2566 2.64e-16
c17493 1516 1505 1.58e-16
c17494 85 37 5.71e-16
c17495 3024 3343 3.92e-16
c17496 4469 4480 1.58e-16
c17497 1 330 4.22e-16
c17498 233 218 1.88e-16
c17499 3409 797 4.46e-16
c17500 4668 4282 1.179e-15
c17501 4563 4762 1.58e-16
c17502 4580 4774 1.58e-16
c17503 5242 5241 1.6e-16
c17504 5072 62 1.58e-16
c17505 1998 2490 1.58e-16
c17506 2194 2270 3.92e-16
c17507 3876 692 4.48e-16
c17508 5417 5512 3.87e-16
c17509 5429 5409 1.58e-16
c17510 4742 5356 3.65e-16
c17511 3033 2549 5.8e-16
c17512 3047 2538 3.54e-16
c17513 921 1070 1.96e-16
c17514 659 0 7.709e-15
c17515 3092 3091 2.48e-16
c17516 632 3900 3.15e-16
c17517 827 0 2.8001e-13
c17518 3034 2549 1.58e-16
c17519 2921 2969 3.15e-16
c17520 4327 4299 2.64e-16
c17521 3024 2617 1.58e-16
c17522 3030 2611 5.88e-16
c17523 2098 2108 8.28e-16
c17524 3393 3451 1.96e-16
c17525 3151 3543 2.38e-15
c17526 4664 0 6.72e-16
c17527 2173 1 2.606e-15
c17528 552 541 3.84e-16
c17529 5320 323 6.67e-16
c17530 3855 3863 1.65e-16
c17531 3520 692 2.33e-16
c17532 595 3061 1.58e-16
c17533 602 3058 1.832e-15
c17534 2670 2672 2.03e-16
c17535 1069 1070 7.51e-16
c17536 2214 2581 1.58e-16
c17537 910 881 6.99e-16
c17538 4087 19 3.45e-16
c17539 4403 3571 2.48e-16
c17540 4455 1 5.808e-15
c17541 2829 812 1.09e-16
c17542 1708 1816 3.92e-16
c17543 642 26 1.58e-16
c17544 334 331 1.099e-15
c17545 117 368 1.88e-16
c17546 4457 0 3.466e-15
c17547 5074 5034 2.45e-16
c17548 4977 4974 3.54e-16
c17549 4976 4972 5.87e-16
c17550 3046 837 3.15e-16
c17551 776 775 6.67e-16
c17552 3899 3890 1.846e-15
c17553 3411 3219 5.5e-16
c17554 2333 0 6.9484e-14
c17555 2215 2206 3.92e-16
c17556 1681 2209 5.66e-16
c17557 1070 717 1.85e-16
c17558 4810 410 1.88e-16
c17559 2194 0 3.45254e-13
c17560 1354 1356 2.03e-16
c17561 1106 1083 6.54e-16
c17562 3886 4280 1.58e-16
c17563 3898 3429 5.5e-16
c17564 3900 3435 1.58e-16
c17565 922 1205 3.92e-16
c17566 1602 1596 1.6e-16
c17567 1136 1593 2.386e-15
c17568 809 25 1.13e-15
c17569 813 19 1.58e-16
c17570 1706 1815 1.58e-16
c17571 1690 1803 1.58e-16
c17572 1743 1352 1.136e-15
c17573 3276 0 3.6368e-14
c17574 1878 1869 3.46e-16
c17575 3048 3291 5.42e-16
c17576 3024 3279 1.58e-16
c17577 3409 3604 3.92e-16
c17578 1 425 9.8e-16
c17579 3225 3608 7.84e-16
c17580 3387 767 4.48e-16
c17581 4567 4350 1.58e-16
c17582 5426 1 2.386e-15
c17583 2524 0 1.1956e-14
c17584 2476 2487 1.96e-16
c17585 3710 3393 1.58e-16
c17586 5576 5575 1.6e-16
c17587 2178 2252 1.58e-16
c17588 1706 732 3.15e-16
c17589 614 0 7.709e-15
c17590 3106 1 4.41e-15
c17591 3644 0 3.466e-15
c17592 3490 0 6.62e-16
c17593 4254 0 1.4092e-14
c17594 4491 3656 1.96e-16
c17595 4496 3650 1.96e-16
c17596 812 0 2.80345e-13
c17597 2629 647 7.68e-16
c17598 4756 4754 1.6e-16
c17599 245 259 3.84e-16
c17600 276 252 1.88e-16
c17601 612 0 2.86378e-13
c17602 2117 1 2.223e-15
c17603 848 847 1.96e-16
c17604 3909 857 1.88e-16
c17605 5062 5064 1.783e-15
c17606 762 2350 1.58e-16
c17607 2196 1732 1.58e-16
c17608 2182 2252 1.58e-16
c17609 907 837 3.15e-16
c17610 88 1 4.22e-16
c17611 111 0 6.224e-15
c17612 3708 858 1.339e-15
c17613 4338 677 1.9e-16
c17614 2897 0 2.078e-15
c17615 595 2541 4.03e-16
c17616 921 677 3.15e-16
c17617 1321 1340 1.58e-16
c17618 1345 1341 3.92e-16
c17619 2567 2578 1.96e-16
c17620 2136 1670 5.5e-16
c17621 3882 3571 1.58e-16
c17622 2921 2917 5.32e-16
c17623 3262 777 1.58e-16
c17624 2557 2305 1.58e-16
c17625 791 1 5.57e-16
c17626 4044 26 4.58e-16
c17627 4036 0 2.061e-14
c17628 3046 3088 3.92e-16
c17629 1811 1806 1.642e-15
c17630 822 1343 3.15e-16
c17631 4419 1 1.716e-15
c17632 5071 5076 3.07e-16
c17633 251 262 3.84e-16
c17634 5218 0 1.23e-16
c17635 3330 827 1.832e-15
c17636 4878 5010 1.96e-16
c17637 894 647 3.15e-16
c17638 2672 0 6.62e-16
c17639 4580 4864 1.58e-16
c17640 4571 4876 1.58e-16
c17641 986 1406 1.58e-16
c17642 2172 747 3.15e-16
c17643 4007 4004 1.58e-16
c17644 4736 5358 2.039e-15
c17645 3098 1 6.15e-16
c17646 2829 2826 3.01e-16
c17647 2825 2822 6.44e-16
c17648 1845 717 3.79e-16
c17649 1343 1677 4.22e-16
c17650 764 25 1.13e-15
c17651 768 19 1.58e-16
c17652 378 375 3.54e-16
c17653 4276 4265 1.58e-16
c17654 1708 1397 5.5e-16
c17655 880 1 4.224e-15
c17656 3236 762 3.79e-16
c17657 1356 0 6.62e-16
c17658 4225 1 6.76e-16
c17659 4417 762 2.4e-16
c17660 2832 837 3.79e-16
c17661 4384 1 4.442e-15
c17662 4915 497 1.88e-16
c17663 1869 0 1.6491e-14
c17664 3409 3569 1.58e-16
c17665 612 2203 1.58e-16
c17666 602 2170 1.58e-16
c17667 2291 1 5.808e-15
c17668 9 332 5.8e-16
c17669 3287 827 1.58e-16
c17670 5417 470 3.19e-16
c17671 5170 1 1.113e-15
c17672 5025 91 3.54e-16
c17673 2178 1868 1.58e-16
c17674 3736 3739 1.96e-16
c17675 922 797 5.14e-16
c17676 921 1128 1.58e-16
c17677 146 135 3.84e-16
c17678 3480 4297 1.58e-16
c17679 4409 737 1.09e-16
c17680 2535 2486 5.5e-16
c17681 2739 2748 3.92e-16
c17682 1684 692 4.48e-16
c17683 1321 1503 1.58e-16
c17684 1343 1491 1.58e-16
c17685 2648 2646 1.6e-16
c17686 2714 707 3.64e-16
c17687 632 1708 3.15e-16
c17688 4198 19 9.67e-16
c17689 3316 2798 2.38e-15
c17690 601 2571 5.03e-16
c17691 2280 1 6.15e-16
c17692 632 2178 3.15e-16
c17693 792 1345 3.58e-16
c17694 1 253 1.607e-15
c17695 4674 4682 1.81e-16
c17696 4563 4689 1.58e-16
c17697 2182 1868 1.58e-16
c17698 0 244 9.795e-15
c17699 4514 3673 1.136e-15
c17700 5446 439 6.67e-16
c17701 1862 2354 1.58e-16
c17702 2045 1 2.386e-15
c17703 2824 1 5.808e-15
c17704 1421 672 1.58e-16
c17705 2826 0 3.466e-15
c17706 4719 410 1.88e-16
c17707 2559 2271 1.58e-16
c17708 2637 2265 1.58e-16
c17709 542 540 1.257e-15
c17710 3029 3041 3.225e-15
c17711 1871 722 1.832e-15
c17712 642 1415 2.65e-16
c17713 4092 4086 1.96e-16
c17714 2713 1 5.97e-15
c17715 1151 1150 3.94e-16
c17716 2413 767 1.58e-16
c17717 1754 1363 4.11e-16
c17718 3048 3038 5.5e-16
c17719 2328 707 1.84e-16
c17720 617 1761 3.64e-16
c17721 601 1380 1.58e-16
c17722 632 2182 3.15e-16
c17723 2019 2020 9.1e-16
c17724 1684 1539 1.58e-16
c17725 1690 1533 5.88e-16
c17726 457 451 1.372e-15
c17727 436 437 7.03e-16
c17728 5174 236 7.94e-16
c17729 2369 2368 1.6e-16
c17730 2361 2359 2.15e-16
c17731 2054 1 7.49e-16
c17732 2047 0 1.65e-16
c17733 731 730 6.67e-16
c17734 890 923 3.54e-16
c17735 909 969 1.58e-16
c17736 390 1 2.946e-15
c17737 226 233 3.54e-16
c17738 222 216 5.8e-16
c17739 2816 2418 4.36e-16
c17740 2641 2639 1.6e-16
c17741 2636 2635 2.03e-16
c17742 3287 3276 1.58e-16
c17743 4617 33 1.88e-16
c17744 3746 3745 1.6e-16
c17745 2938 2915 5.87e-16
c17746 1345 737 3.15e-16
c17747 4368 4379 1.96e-16
c17748 3598 1 8.43e-16
c17749 723 19 1.58e-16
c17750 1278 1 5.21e-16
c17751 4171 1 6.66e-16
c17752 1830 1 9.28e-16
c17753 720 719 1.6e-16
c17754 822 1982 2.65e-16
c17755 1 37 5.625e-14
c17756 15 50 4.88e-16
c17757 3270 3661 4.11e-16
c17758 5257 5261 8.88e-16
c17759 5240 5232 1.725e-15
c17760 2436 1 1.868e-15
c17761 592 667 1.96e-16
c17762 2426 0 2.93e-15
c17763 627 2172 3.15e-16
c17764 0 39 2.87e-16
c17765 407 570 1.88e-16
c17766 3548 3543 1.642e-15
c17767 3287 812 3.15e-16
c17768 3025 1 2.606e-15
c17769 4468 797 7.38e-16
c17770 5514 5481 1.58e-16
c17771 632 999 8.3e-16
c17772 4383 722 7.38e-16
c17773 3446 4264 1.96e-16
c17774 1942 797 1.84e-16
c17775 1331 1011 1.58e-16
c17776 4612 4609 5.5e-16
c17777 3744 3731 1.58e-16
c17778 4176 1 4.2638e-14
c17779 4542 4544 2.61e-16
c17780 2486 858 3.15e-16
c17781 4152 25 7.01e-16
c17782 4890 4884 3.47e-16
c17783 4813 4812 2.48e-16
c17784 4816 4817 2.83e-16
c17785 4429 4820 1.96e-16
c17786 3034 3190 4.63e-16
c17787 2139 2137 3.92e-16
c17788 302 305 1.099e-15
c17789 2421 2419 1.6e-16
c17790 803 802 1.96e-16
c17791 48 0 1.5723e-14
c17792 3856 3853 6.71e-16
c17793 3537 732 5.73e-16
c17794 4872 5133 1.383e-15
c17795 2788 1 1.716e-15
c17796 5324 5320 5.32e-16
c17797 3016 3014 1.6e-16
c17798 732 26 1.58e-16
c17799 4151 37 1.88e-16
c17800 3959 1 3.66e-16
c17801 595 3429 2.22e-16
c17802 601 3418 2.33e-16
c17803 3898 4332 3.92e-16
c17804 4449 4447 1.6e-16
c17805 3284 3281 3.01e-16
c17806 3280 3277 6.44e-16
c17807 1464 1 8.43e-16
c17808 687 25 1.58e-16
c17809 5010 1 3.7078e-14
c17810 3409 3270 5.5e-16
c17811 5131 31 3.54e-16
c17812 1088 737 1.58e-16
c17813 883 905 3.92e-16
c17814 64 581 6.01e-16
c17815 3713 3720 6.73e-16
c17816 2516 2514 2.61e-16
c17817 4571 4563 4.078e-15
c17818 4582 5591 3.54e-16
c17819 4634 5452 1.53e-15
c17820 1131 782 2.33e-16
c17821 1377 1374 3.01e-16
c17822 1373 1370 6.44e-16
c17823 2651 0 3.5142e-14
c17824 2557 2598 1.58e-16
c17825 2541 2586 1.58e-16
c17826 2532 2531 3.54e-16
c17827 670 1 3.79e-16
c17828 663 0 7.86e-15
c17829 4328 1 1.868e-15
c17830 1516 1914 4.36e-16
c17831 1912 1905 1.96e-16
c17832 1684 1685 1.487e-15
c17833 1694 1687 1.58e-16
c17834 5027 5026 5.87e-16
c17835 4318 0 2.93e-15
c17836 685 686 6.67e-16
c17837 4497 4469 2.64e-16
c17838 4864 4870 7.25e-16
c17839 88 363 1.88e-16
c17840 223 334 1.88e-16
c17841 3397 3501 1.58e-16
c17842 4563 4779 1.58e-16
c17843 4580 4791 1.58e-16
c17844 4855 207 1.88e-16
c17845 4827 468 1.88e-16
c17846 1981 2498 2.38e-15
c17847 797 788 1.078e-15
c17848 747 0 2.85991e-13
c17849 3918 3932 2.87e-16
c17850 3941 3942 3.15e-16
c17851 2172 2287 3.92e-16
c17852 920 1084 1.58e-16
c17853 602 3393 3.15e-16
c17854 1920 782 1.339e-15
c17855 2957 2923 1.58e-16
c17856 2747 3258 1.96e-16
c17857 3034 3155 1.58e-16
c17858 1403 0 3.5926e-14
c17859 1603 1 9.28e-16
c17860 465 454 3.84e-16
c17861 5198 5197 2.29e-16
c17862 4681 0 6.72e-16
c17863 2384 0 6.909e-14
c17864 910 2194 1.014e-15
c17865 911 2172 1.88e-16
c17866 2179 1 3.358e-15
c17867 480 478 1.58e-16
c17868 306 320 1.58e-16
c17869 0 213 2.87e-16
c17870 19 200 3.45e-16
c17871 3655 782 1.58e-16
c17872 5146 5133 8.94e-16
c17873 5143 5104 1.738e-15
c17874 4861 178 1.88e-16
c17875 3514 707 1.58e-16
c17876 601 3058 1.58e-16
c17877 4232 4243 1.96e-16
c17878 2170 2589 2.38e-15
c17879 2545 2186 1.58e-16
c17880 1653 842 3.64e-16
c17881 4809 782 1.23e-16
c17882 4475 1 2.054e-15
c17883 3169 2651 1.96e-16
c17884 3170 3163 6.73e-16
c17885 2557 702 3.15e-16
c17886 602 1685 5.18e-16
c17887 5072 5113 1.817e-15
c17888 702 700 3.327e-15
c17889 4464 792 2.65e-16
c17890 4477 0 8e-16
c17891 3454 3072 2.48e-16
c17892 360 362 2.84e-16
c17893 350 355 1.059e-15
c17894 3174 717 1.58e-16
c17895 4962 4944 1.23e-16
c17896 2307 2309 2.03e-16
c17897 102 117 1.88e-16
c17898 88 131 1.88e-16
c17899 1682 2206 1.58e-16
c17900 4838 4833 1.536e-15
c17901 397 9 5.8e-16
c17902 3684 827 3.15e-16
c17903 4532 868 2.65e-16
c17904 4514 5579 3.92e-16
c17905 602 3432 4.81e-16
c17906 3129 1 2.054e-15
c17907 2798 2407 1.136e-15
c17908 3886 4285 1.58e-16
c17909 3876 3446 5.5e-16
c17910 3131 0 8e-16
c17911 2545 2555 3.92e-16
c17912 2559 2531 3.54e-16
c17913 2651 3162 1.96e-16
c17914 2752 737 1.58e-16
c17915 1884 1883 9.1e-16
c17916 168 169 1.58e-16
c17917 3048 3296 1.58e-16
c17918 2215 2204 1.96e-16
c17919 1925 0 1.4092e-14
c17920 2031 2082 2.45e-16
c17921 5514 468 1.58e-16
c17922 2170 2171 3.36e-16
c17923 919 868 3.15e-16
c17924 5496 5481 7.95e-16
c17925 4922 149 1.88e-16
c17926 3664 0 8e-16
c17927 1527 1076 4.11e-16
c17928 687 1001 1.58e-16
c17929 4069 1 7.71e-16
c17930 1179 0 2.7216e-14
c17931 4480 4843 1.96e-16
c17932 2730 3240 1.58e-16
c17933 1739 0 6.72e-16
c17934 3411 3410 1.866e-15
c17935 596 589 3.134e-15
c17936 627 0 2.86543e-13
c17937 4563 4724 1.96e-16
c17938 338 340 1.58e-16
c17939 2373 2374 1.35e-16
c17940 3770 3775 7.46e-16
c17941 3883 3906 1.003e-15
c17942 2844 2458 5.66e-16
c17943 2663 2665 1.6e-16
c17944 1145 767 1.58e-16
c17945 4197 3890 7.84e-16
c17946 1321 880 1.58e-16
c17947 1327 877 1.58e-16
c17948 647 1 3.1284e-14
c17949 3898 3588 1.58e-16
c17950 2952 2959 8.96e-16
c17951 1795 1403 1.96e-16
c17952 1796 1789 6.73e-16
c17953 993 0 4.6723e-14
c17954 3024 3105 3.92e-16
c17955 1694 1986 4.63e-16
c17956 4445 1 8.43e-16
c17957 19 346 8.4e-16
c17958 192 204 1.58e-16
c17959 30 354 3.84e-16
c17960 2385 2376 3.92e-16
c17961 1868 2379 5.66e-16
c17962 4982 4910 3.54e-16
c17963 2697 1 1.868e-15
c17964 890 1037 1.96e-16
c17965 276 273 1.099e-15
c17966 88 310 1.88e-16
c17967 657 659 5.59e-16
c17968 3397 3202 5.5e-16
c17969 4580 4881 1.58e-16
c17970 4571 4893 1.58e-16
c17971 4702 468 1.88e-16
c17972 2492 1 4.946e-15
c17973 2687 0 2.93e-15
c17974 2136 2137 3.54e-16
c17975 3708 3717 3.46e-16
c17976 3684 812 1.58e-16
c17977 5564 5561 3.54e-16
c17978 1326 1330 5.8e-16
c17979 3548 4390 2.38e-15
c17980 2350 722 3.15e-16
c17981 4293 4265 2.64e-16
c17982 4666 4660 7.25e-16
c17983 4276 4282 9.42e-16
c17984 3145 3148 3.01e-16
c17985 3141 3144 6.44e-16
c17986 4549 4546 1.138e-15
c17987 5005 4896 7.59e-16
c17988 4401 1 4.442e-15
c17989 3330 3342 2.32e-16
c17990 3034 2730 5.5e-16
c17991 1 453 3.6e-16
c17992 3409 3574 1.58e-16
c17993 4861 4868 1.81e-16
c17994 1044 702 1.58e-16
c17995 3881 3390 7.67e-16
c17996 601 2170 3.15e-16
c17997 627 2203 5.73e-16
c17998 2311 1 2.054e-15
c17999 9 478 6.48e-16
c18000 473 0 2.87e-16
c18001 2466 2463 3.01e-16
c18002 2462 2459 6.44e-16
c18003 1239 592 3.6e-16
c18004 5561 5543 6.72e-16
c18005 4753 5173 9.04e-16
c18006 4827 64 1.88e-16
c18007 3632 1 8.43e-16
c18008 536 0 1.5696e-14
c18009 506 19 3.84e-16
c18010 3392 3388 1.988e-15
c18011 2333 707 3.15e-16
c18012 4031 1 6.66e-16
c18013 2194 707 4.46e-16
c18014 1769 1776 1.96e-16
c18015 792 782 3.28e-16
c18016 601 2591 1.09e-16
c18017 2289 1 1.716e-15
c18018 657 2194 3.15e-16
c18019 1 176 1.456e-15
c18020 4563 4706 1.58e-16
c18021 4691 4696 5.53e-16
c18022 3619 752 4.81e-16
c18023 2194 2193 1.009e-15
c18024 2178 2183 8.56e-16
c18025 2844 1 2.054e-15
c18026 2737 2748 1.96e-16
c18027 1425 662 5.03e-16
c18028 894 1157 3.92e-16
c18029 909 1156 1.88e-16
c18030 883 1149 1.58e-16
c18031 2846 0 8e-16
c18032 922 978 1.58e-16
c18033 3719 3713 1.6e-16
c18034 632 1417 4.81e-16
c18035 4600 5562 2.137e-15
c18036 4606 5538 1.344e-15
c18037 3021 0 4.4783e-14
c18038 3622 4455 7.84e-16
c18039 3320 2798 1.96e-16
c18040 3315 2804 1.96e-16
c18041 3885 1 2.56e-15
c18042 4006 26 4.48e-16
c18043 617 1380 3.15e-16
c18044 1675 1674 1.6e-16
c18045 1676 1196 1.23e-16
c18046 1659 1206 3.92e-16
c18047 1663 1661 1.96e-16
c18048 4546 3707 1.958e-15
c18049 4570 1 2.248e-15
c18050 4728 4740 2.62e-16
c18051 1708 1556 1.58e-16
c18052 1706 1550 5.5e-16
c18053 1694 1951 1.58e-16
c18054 911 0 3.0498e-13
c18055 1943 1941 1.6e-16
c18056 1938 1937 2.03e-16
c18057 762 1076 1.58e-16
c18058 747 1091 3.79e-16
c18059 1512 0 6.72e-16
c18060 5010 4950 1.58e-16
c18061 687 2308 1.58e-16
c18062 2182 2183 1.027e-15
c18063 662 656 1.74e-16
c18064 5299 352 9.42e-16
c18065 883 963 3.54e-16
c18066 894 984 1.58e-16
c18067 277 1 1.65e-15
c18068 88 339 1.88e-16
c18069 3463 647 3.15e-16
c18070 3287 3685 4.36e-16
c18071 5558 1 1.81e-16
c18072 3729 3726 6.71e-16
c18073 1146 807 4e-16
c18074 1408 981 1.96e-16
c18075 632 4271 1.84e-16
c18076 642 4285 1.58e-16
c18077 2535 2650 3.92e-16
c18078 1656 1657 9.1e-16
c18079 4404 747 1.58e-16
c18080 1843 1 6.15e-16
c18081 4899 4907 3.54e-16
c18082 822 1601 3.79e-16
c18083 4446 4833 2.196e-15
c18084 5556 1 1.88e-16
c18085 2738 2350 4.97e-16
c18086 1930 1 5.97e-15
c18087 792 19 1.41e-15
c18088 4056 857 3.1e-16
c18089 5535 0 3.7461e-14
c18090 3031 1 3.358e-15
c18091 1517 722 3.64e-16
c18092 134 1 3.6e-16
c18093 154 0 2.87e-16
c18094 538 552 1.58e-16
c18095 2684 702 2.4e-16
c18096 581 585 1.059e-15
c18097 1747 1748 9.1e-16
c18098 4327 0 6.9337e-14
c18099 908 898 2.303e-15
c18100 737 727 6.38e-16
c18101 3972 3976 3.84e-16
c18102 3980 3979 4.41e-16
c18103 4742 439 1.88e-16
c18104 5365 294 9.42e-16
c18105 378 368 3.75e-16
c18106 5409 5426 1.443e-15
c18107 5388 5355 1.58e-16
c18108 986 982 3.78e-16
c18109 632 3409 4.46e-16
c18110 3446 4263 1.58e-16
c18111 3435 4271 5.66e-16
c18112 4277 4268 3.92e-16
c18113 1472 1041 3.92e-16
c18114 1476 1477 1.6e-16
c18115 617 607 6.38e-16
c18116 737 19 1.676e-15
c18117 3980 1 4.64e-16
c18118 617 3418 1.75e-16
c18119 3876 4349 3.92e-16
c18120 4814 4811 6.67e-16
c18121 3718 4523 1.58e-16
c18122 3194 3206 2.32e-16
c18123 209 178 1.88e-16
c18124 3500 3498 1.6e-16
c18125 3886 762 7.99e-16
c18126 3387 3688 1.58e-16
c18127 1110 737 6.48e-16
c18128 921 924 3.54e-16
c18129 6 1 1.073e-15
c18130 4617 526 1.88e-16
c18131 2708 2322 5.66e-16
c18132 2220 0 3.6368e-14
c18133 3882 4319 1.58e-16
c18134 3898 4331 1.58e-16
c18135 3926 25 3.84e-16
c18136 4354 4351 6.44e-16
c18137 4358 4355 3.01e-16
c18138 4702 64 1.88e-16
c18139 2535 2615 1.58e-16
c18140 2557 2603 1.58e-16
c18141 2533 2534 3.36e-16
c18142 689 1 7.18e-16
c18143 1440 0 3.3846e-14
c18144 3387 3123 1.58e-16
c18145 3497 1 5.97e-15
c18146 3639 822 5.73e-16
c18147 4604 3874 1.58e-16
c18148 1690 1698 8.73e-16
c18149 483 484 3.84e-16
c18150 1743 2235 1.58e-16
c18151 1658 2117 7.46e-16
c18152 1 523 4.22e-16
c18153 4793 4794 9.93e-16
c18154 4563 4796 1.58e-16
c18155 4580 4808 1.58e-16
c18156 5229 5234 5.63e-16
c18157 1010 647 5.74e-16
c18158 3918 3947 8.1e-16
c18159 2968 1 2.223e-15
c18160 1256 1255 1.6e-16
c18161 65 1 5.62e-16
c18162 5482 5484 1.96e-16
c18163 601 3393 3.15e-16
c18164 1091 1551 4.36e-16
c18165 1549 1542 1.96e-16
c18166 1345 1001 5.5e-16
c18167 1327 1419 1.96e-16
c18168 3538 0 1.6491e-14
c18169 4594 4595 1.6e-16
c18170 4590 3870 1.443e-15
c18171 4139 1 6.66e-16
c18172 2041 2518 4.79e-16
c18173 2136 2048 1.761e-15
c18174 2995 2521 5.5e-16
c18175 2441 827 1.75e-16
c18176 1807 1805 1.6e-16
c18177 1802 1801 2.03e-16
c18178 602 1368 1.58e-16
c18179 4866 4480 4.11e-16
c18180 4871 4862 3.46e-16
c18181 1616 1 6.15e-16
c18182 3411 3117 5.5e-16
c18183 2117 2070 1.836e-15
c18184 4698 0 6.72e-16
c18185 5234 5227 9.81e-16
c18186 19 303 3.84e-16
c18187 3567 3560 6.73e-16
c18188 3566 3174 1.96e-16
c18189 4793 352 1.88e-16
c18190 2390 2401 1.58e-16
c18191 4381 707 4.81e-16
c18192 5414 5413 5.87e-16
c18193 5303 5310 3.18e-16
c18194 5296 5283 1.58e-16
c18195 4838 5086 1.96e-16
c18196 601 3078 1.58e-16
c18197 3874 3875 3.36e-16
c18198 2756 0 3.3437e-14
c18199 1196 842 3.15e-16
c18200 74 72 1.58e-16
c18201 687 4345 2.65e-16
c18202 2665 662 4.81e-16
c18203 2545 2769 4.63e-16
c18204 1067 0 1.0183e-14
c18205 3811 410 1.038e-15
c18206 4120 25 7.01e-16
c18207 4420 3582 4.97e-16
c18208 5041 180 5.93e-16
c18209 2662 2651 1.58e-16
c18210 2559 717 3.58e-16
c18211 479 368 1.88e-16
c18212 5106 5114 1.725e-15
c18213 2196 1760 5.5e-16
c18214 3633 792 3.79e-16
c18215 4493 0 6.72e-16
c18216 4903 4968 6.67e-16
c18217 4940 4941 3.54e-16
c18218 3429 3424 1.642e-15
c18219 1682 2226 2.38e-15
c18220 3321 3316 1.642e-15
c18221 2572 1 2.054e-15
c18222 3701 868 3.79e-16
c18223 4523 858 1.58e-16
c18224 4634 5410 1.925e-15
c18225 612 3022 1.813e-15
c18226 1355 880 7.84e-16
c18227 4404 4416 2.32e-16
c18228 3820 0 3.6242e-14
c18229 1708 1820 1.58e-16
c18230 367 378 3.84e-16
c18231 4299 1 4.442e-15
c18232 1890 1886 1.96e-16
c18233 4640 4641 9.93e-16
c18234 4567 4361 5.5e-16
c18235 4844 120 1.88e-16
c18236 4787 439 1.88e-16
c18237 642 3024 3.15e-16
c18238 1343 672 3.15e-16
c18239 1321 647 4.48e-16
c18240 1366 1364 1.6e-16
c18241 2557 2556 1.009e-15
c18242 2541 2546 8.56e-16
c18243 1470 692 7.38e-16
c18244 920 858 3.69e-16
c18245 3680 0 6.72e-16
c18246 4228 4225 1.76e-16
c18247 1327 1384 1.58e-16
c18248 4508 3667 4.11e-16
c18249 2441 812 2.33e-16
c18250 1590 1591 1.35e-16
c18251 2747 3228 1.58e-16
c18252 542 536 3.84e-16
c18253 4773 4771 1.6e-16
c18254 3409 3018 1.58e-16
c18255 2359 1 5.808e-15
c18256 4563 4741 1.96e-16
c18257 3625 767 1.832e-15
c18258 2361 0 3.466e-15
c18259 5422 5423 3.18e-16
c18260 4725 5366 3.92e-16
c18261 4708 5326 7.84e-16
c18262 894 868 8.34e-16
c18263 2949 294 1.108e-15
c18264 5400 5177 9.75e-16
c18265 2545 2367 5.5e-16
c18266 657 663 1.097e-15
c18267 3010 2929 3.2e-16
c18268 2955 2959 3.54e-16
c18269 632 922 5.14e-16
c18270 3882 3599 5.88e-16
c18271 3876 3605 1.58e-16
c18272 2452 807 2.22e-16
c18273 2196 752 3.15e-16
c18274 2545 2734 1.58e-16
c18275 1027 0 1.8851e-14
c18276 1699 1693 1.6e-16
c18277 4567 4565 5.93e-16
c18278 5032 5093 1.6e-16
c18279 2144 1 1.356e-15
c18280 617 2240 1.832e-15
c18281 2036 0 5.6946e-14
c18282 158 172 3.84e-16
c18283 4938 4910 4.39e-16
c18284 2316 1 5.97e-15
c18285 762 1694 7.99e-16
c18286 3290 1 1.056e-15
c18287 1432 996 1.96e-16
c18288 1433 1426 6.73e-16
c18289 642 883 3.15e-16
c18290 602 3034 3.15e-16
c18291 657 1403 1.58e-16
c18292 3259 1 4.41e-15
c18293 4293 4282 1.58e-16
c18294 911 1689 1.58e-16
c18295 1383 1 1.056e-15
c18296 957 0 7.4294e-14
c18297 4421 0 3.3268e-14
c18298 3430 3021 1.96e-16
c18299 3431 3424 6.73e-16
c18300 3022 3406 2.79e-16
c18301 2722 722 1.832e-15
c18302 4418 1 4.442e-15
c18303 2568 2570 2.03e-16
c18304 3397 3390 1.58e-16
c18305 627 2612 2.65e-16
c18306 617 2170 1.58e-16
c18307 612 2231 2.22e-16
c18308 2493 0 1.6491e-14
c18309 4793 294 1.88e-16
c18310 4736 352 1.88e-16
c18311 910 3021 3.75e-16
c18312 2194 1879 5.5e-16
c18313 2015 2010 1.642e-15
c18314 2518 1998 9.7e-16
c18315 384 381 4.6e-16
c18316 4301 3469 2.48e-16
c18317 1327 1071 1.58e-16
c18318 4237 1 2.054e-15
c18319 910 911 3.45e-16
c18320 3394 3392 8.67e-16
c18321 4239 0 8e-16
c18322 3333 3340 6.73e-16
c18323 666 655 7.23e-16
c18324 658 659 1.6e-16
c18325 3695 3304 4.11e-16
c18326 2315 1 8.43e-16
c18327 961 962 4.01e-16
c18328 9 364 4.88e-16
c18329 129 130 5.8e-16
c18330 3693 3387 1.58e-16
c18331 5474 5473 1.6e-16
c18332 1442 672 2.72e-16
c18333 1192 827 1.58e-16
c18334 842 1202 1.58e-16
c18335 1193 868 1.58e-16
c18336 894 1171 1.58e-16
c18337 907 1143 3.54e-16
c18338 1011 1014 1.58e-16
c18339 2862 0 6.72e-16
c18340 3882 3881 3.15e-16
c18341 5358 5353 7.46e-16
c18342 2826 2441 1.96e-16
c18343 1061 1503 1.58e-16
c18344 984 1 2.972e-15
c18345 3633 4467 1.58e-16
c18346 1919 782 2.33e-16
c18347 1690 1420 1.58e-16
c18348 1776 1767 3.46e-16
c18349 4857 4856 1.6e-16
c18350 985 0 6.29e-16
c18351 2713 3227 4.97e-16
c18352 3048 3058 1.58e-16
c18353 25 262 5.71e-16
c18354 27 252 1.88e-16
c18355 596 947 5.28e-16
c18356 5356 5374 1.37e-16
c18357 2661 2265 1.96e-16
c18358 1414 662 3.15e-16
c18359 1281 1218 1.58e-16
c18360 1635 868 3.79e-16
c18361 1206 1660 1.96e-16
c18362 1321 1656 1.58e-16
c18363 1343 1644 1.58e-16
c18364 1580 1578 1.6e-16
c18365 1575 1574 2.03e-16
c18366 4385 0 1.6491e-14
c18367 1336 0 6.35e-16
c18368 3744 1 6.04e-16
c18369 1852 1 1.716e-15
c18370 3839 0 5.5835e-14
c18371 418 0 9.795e-15
c18372 282 274 2.218e-15
c18373 1 133 4.22e-16
c18374 3387 3157 1.58e-16
c18375 2472 1 1.056e-15
c18376 1023 677 1.58e-16
c18377 3882 3390 1.96e-16
c18378 1076 722 3.15e-16
c18379 657 993 1.05e-15
c18380 910 879 3.84e-16
c18381 1573 797 2.33e-16
c18382 1331 1031 5.5e-16
c18383 3594 0 1.4092e-14
c18384 4629 4626 5.5e-16
c18385 506 512 5.8e-16
c18386 4191 1 6.66e-16
c18387 2504 858 7.68e-16
c18388 1117 1 3.54e-16
c18389 4921 4920 1.6e-16
c18390 1114 0 9.602e-15
c18391 3030 3223 1.58e-16
c18392 4830 4829 2.48e-16
c18393 4833 4834 2.83e-16
c18394 4446 4837 1.96e-16
c18395 82 71 2.45e-16
c18396 4344 0 6.9337e-14
c18397 27 22 3.54e-16
c18398 31 33 1.96e-16
c18399 3387 717 3.15e-16
c18400 5383 1 1.88e-16
c18401 2425 1919 3.92e-16
c18402 2429 2430 1.6e-16
c18403 3565 717 2.22e-16
c18404 4387 722 1.832e-15
c18405 2727 2724 3.01e-16
c18406 2723 2720 6.44e-16
c18407 3446 4268 1.58e-16
c18408 920 965 3.92e-16
c18409 921 964 1.88e-16
c18410 1856 722 5.03e-16
c18411 632 971 3.15e-16
c18412 2882 2895 1.138e-15
c18413 2541 2803 1.96e-16
c18414 910 919 1.58e-16
c18415 3999 1 6.66e-16
c18416 4166 26 4.48e-16
c18417 601 3446 1.58e-16
c18418 617 4277 3.64e-16
c18419 3900 4366 3.92e-16
c18420 3292 2781 1.96e-16
c18421 926 0 1.8747e-14
c18422 4709 4333 3.92e-16
c18423 4721 4720 1.6e-16
c18424 2856 858 1.339e-15
c18425 49 508 1.88e-16
c18426 3701 0 7.0003e-14
c18427 1618 1 5.97e-15
c18428 5010 410 1.88e-16
c18429 5326 5331 3.84e-16
c18430 5324 5363 3.18e-16
c18431 2790 0 3.3717e-14
c18432 920 942 2.041e-15
c18433 4167 4164 1.58e-16
c18434 4736 294 1.88e-16
c18435 4668 5522 5.5e-16
c18436 1404 971 1.532e-15
c18437 3898 4336 1.58e-16
c18438 3876 4348 1.58e-16
c18439 2679 0 6.9481e-14
c18440 2559 2632 5.42e-16
c18441 2535 2620 1.58e-16
c18442 3107 2600 3.92e-16
c18443 3111 3112 1.6e-16
c18444 1460 0 1.4092e-14
c18445 747 745 3.327e-15
c18446 3106 3488 2.48e-16
c18447 4364 1 1.056e-15
c18448 4498 822 2.65e-16
c18449 4242 4604 1.58e-16
c18450 207 267 1.58e-16
c18451 2175 1687 1.96e-16
c18452 4881 4887 7.25e-16
c18453 3024 732 3.15e-16
c18454 2899 2907 1.077e-15
c18455 2240 1743 1.58e-16
c18456 2608 0 8e-16
c18457 4563 4813 1.58e-16
c18458 4580 4825 1.58e-16
c18459 5296 1 1.113e-15
c18460 2525 2004 1.96e-16
c18461 952 1372 7.84e-16
c18462 64 236 1.88e-16
c18463 3181 0 6.72e-16
c18464 3886 722 3.15e-16
c18465 2541 762 4.03e-16
c18466 617 3393 3.15e-16
c18467 2600 3108 2.48e-16
c18468 1690 1680 3.54e-16
c18469 1706 1683 1.58e-16
c18470 4530 4523 1.96e-16
c18471 3684 4532 4.36e-16
c18472 2458 868 5.73e-16
c18473 601 1368 7.38e-16
c18474 894 0 3.14247e-13
c18475 1625 1 1.716e-15
c18476 621 610 7.23e-16
c18477 613 614 1.6e-16
c18478 1 561 4.22e-16
c18479 233 334 1.88e-16
c18480 421 204 1.88e-16
c18481 3411 677 3.15e-16
c18482 3185 3174 1.58e-16
c18483 3642 807 1.58e-16
c18484 4674 497 1.88e-16
c18485 5283 0 3.6422e-14
c18486 627 3092 1.58e-16
c18487 617 3078 1.84e-16
c18488 4253 3418 1.96e-16
c18489 4258 3385 1.96e-16
c18490 2929 2486 9.7e-16
c18491 2541 2401 5.88e-16
c18492 2612 2220 1.96e-16
c18493 2613 2606 6.73e-16
c18494 1663 852 2.42e-16
c18495 687 3514 3.79e-16
c18496 3886 4502 4.63e-16
c18497 2518 2984 1.383e-15
c18498 2764 3245 1.58e-16
c18499 2662 3186 4.36e-16
c18500 3184 3177 1.96e-16
c18501 1988 1990 1.862e-15
c18502 1601 1607 1.418e-15
c18503 3471 3083 4.97e-16
c18504 500 495 1.059e-15
c18505 3560 722 1.84e-16
c18506 3030 858 3.15e-16
c18507 883 732 3.15e-16
c18508 5112 0 1.65e-16
c18509 3397 3654 1.58e-16
c18510 595 598 5.59e-16
c18511 1443 1440 5.5e-16
c18512 4140 3918 2.87e-16
c18513 627 3022 1.58e-16
c18514 3345 0 1.6491e-14
c18515 2178 2474 1.96e-16
c18516 1121 1124 6.13e-16
c18517 389 407 1.58e-16
c18518 1716 1315 1.532e-15
c18519 3915 26 4.58e-16
c18520 3907 0 2.2246e-14
c18521 4497 4492 1.642e-15
c18522 2824 837 1.58e-16
c18523 1690 1454 1.58e-16
c18524 3455 3467 2.32e-16
c18525 2319 2317 1.6e-16
c18526 3048 692 3.15e-16
c18527 1682 2230 1.96e-16
c18528 1715 2225 1.96e-16
c18529 596 830 5.28e-16
c18530 2565 0 3.22e-16
c18531 4567 4378 5.5e-16
c18532 2182 2474 4.63e-16
c18533 391 1 1.073e-15
c18534 2178 1749 1.58e-16
c18535 4436 782 1.339e-15
c18536 5514 5427 4.2e-16
c18537 5484 5493 1.96e-16
c18538 4804 5044 4.79e-16
c18539 661 1 4.03e-16
c18540 4321 4322 1.6e-16
c18541 2276 647 1.9e-16
c18542 3512 1 6.15e-16
c18543 2680 2674 1.6e-16
c18544 1538 1537 9.1e-16
c18545 868 1 4.1542e-14
c18546 2952 2956 5.6e-16
c18547 632 2268 4.81e-16
c18548 4111 1 5.284e-15
c18549 1193 0 1.4198e-14
c18550 3034 2798 5.5e-16
c18551 1386 1 4.41e-15
c18552 1770 0 6.62e-16
c18553 3387 3450 1.58e-16
c18554 3186 707 7.68e-16
c18555 2559 842 3.15e-16
c18556 632 2237 2.33e-16
c18557 5215 5190 5.87e-16
c18558 5192 5194 6.87e-16
c18559 566 572 1.372e-15
c18560 3547 3538 3.46e-16
c18561 3959 857 6.23e-16
c18562 762 1862 1.58e-16
c18563 747 1879 3.79e-16
c18564 2182 1749 1.58e-16
c18565 5505 5452 3.18e-16
c18566 5503 5491 1.96e-16
c18567 5482 5489 1.96e-16
c18568 4804 5230 2.037e-15
c18569 890 858 3.15e-16
c18570 907 1217 3.92e-16
c18571 602 3063 1.09e-16
c18572 919 707 3.15e-16
c18573 920 1038 1.58e-16
c18574 971 970 3.94e-16
c18575 1345 881 5.5e-16
c18576 657 919 3.15e-16
c18577 595 592 5.8e-16
c18578 3667 4502 1.96e-16
c18579 3831 1 3.36e-16
c18580 4076 25 1.88e-16
c18581 4072 19 7.35e-16
c18582 2545 2739 1.58e-16
c18583 1698 1693 4.17e-16
c18584 2730 3243 1.532e-15
c18585 3248 3249 5.65e-16
c18586 3034 2628 5.5e-16
c18587 3179 692 1.9e-16
c18588 632 2605 5.03e-16
c18589 2066 2067 3.54e-16
c18590 325 326 3.84e-16
c18591 3623 782 1.339e-15
c18592 5072 5032 5.69e-16
c18593 1635 0 7.0008e-14
c18594 3538 707 1.339e-15
c18595 3881 3890 5.71e-16
c18596 4996 4977 5.87e-16
c18597 2733 1 1.056e-15
c18598 2294 2293 1.6e-16
c18599 909 692 3.15e-16
c18600 883 1051 1.88e-16
c18601 907 1044 1.58e-16
c18602 5177 5173 1.866e-15
c18603 5136 62 1.58e-16
c18604 2172 1 3.564e-15
c18605 4668 4674 1.605e-15
c18606 4685 4691 1.025e-15
c18607 4702 4708 1.997e-15
c18608 4719 4725 1.025e-15
c18609 4736 4742 1.605e-15
c18610 4753 4759 1.025e-15
c18611 4770 4776 1.997e-15
c18612 4787 4793 1.025e-15
c18613 4804 4810 1.605e-15
c18614 4821 4827 1.025e-15
c18615 4838 4844 1.997e-15
c18616 4855 4861 1.025e-15
c18617 4872 4878 1.605e-15
c18618 3306 1 9.28e-16
c18619 1610 827 1.58e-16
c18620 1343 797 4.46e-16
c18621 1331 807 7.99e-16
c18622 601 3034 3.15e-16
c18623 3868 1 8e-16
c18624 3565 3554 1.58e-16
c18625 2368 737 7.68e-16
c18626 3668 1 1.868e-15
c18627 3858 0 1.3715e-14
c18628 1331 1538 4.63e-16
c18629 1399 1 9.28e-16
c18630 4310 4282 2.64e-16
c18631 4683 4677 7.25e-16
c18632 4441 0 1.4092e-14
c18633 1870 1872 2.03e-16
c18634 3022 3021 1.58e-16
c18635 4941 4951 8.86e-16
c18636 3356 858 7.68e-16
c18637 4435 1 4.442e-15
c18638 2730 767 1.58e-16
c18639 3393 3603 1.58e-16
c18640 2512 1 6.636e-15
c18641 707 1067 1.58e-16
c18642 1058 717 1.58e-16
c18643 858 859 1.621e-15
c18644 852 856 2.19e-16
c18645 596 785 5.28e-16
c18646 617 2614 4.81e-16
c18647 627 2231 3.79e-16
c18648 3321 3393 5.88e-16
c18649 5136 5039 6.72e-16
c18650 4878 0 2.68308e-13
c18651 4855 497 1.88e-16
c18652 911 3022 1.88e-16
c18653 2474 1964 1.96e-16
c18654 3898 807 3.15e-16
c18655 616 1 4.03e-16
c18656 1694 722 3.15e-16
c18657 1343 1086 1.58e-16
c18658 3067 2532 1.96e-16
c18659 3068 3061 6.73e-16
c18660 1852 1854 1.862e-15
c18661 1465 1471 1.418e-15
c18662 1482 1454 2.64e-16
c18663 1167 0 6.29e-16
c18664 4255 0 6.72e-16
c18665 3024 3258 3.92e-16
c18666 2031 2033 1.001e-15
c18667 462 37 5.71e-16
c18668 245 262 1.325e-15
c18669 136 117 1.88e-16
c18670 421 175 1.88e-16
c18671 3883 3401 2.035e-15
c18672 3890 3390 1.121e-15
c18673 687 2194 3.15e-16
c18674 767 761 1.74e-16
c18675 1953 2461 7.84e-16
c18676 110 1 1.44e-16
c18677 4708 5284 2.69e-16
c18678 909 1158 3.54e-16
c18679 107 0 7.5596e-14
c18680 4198 4199 3.15e-16
c18681 2680 2282 4.36e-16
c18682 1897 752 7.68e-16
c18683 1076 1491 1.58e-16
c18684 598 26 2.65e-15
c18685 537 49 1.88e-16
c18686 3066 0 6.9118e-14
c18687 3650 4455 1.58e-16
c18688 3633 4472 2.386e-15
c18689 4481 4475 1.6e-16
c18690 3332 2815 4.11e-16
c18691 3709 0 2.93e-15
c18692 4022 19 7.04e-16
c18693 3030 2566 1.58e-16
c18694 672 679 1.6e-16
c18695 519 477 9.5e-16
c18696 3830 3821 3.92e-16
c18697 3775 3820 1.817e-15
c18698 5034 5036 1.001e-15
c18699 157 165 1.58e-16
c18700 78 88 3.75e-16
c18701 1610 812 1.832e-15
c18702 1166 807 4.21e-16
c18703 1001 1406 1.58e-16
c18704 1671 1345 1.96e-16
c18705 3135 3129 1.6e-16
c18706 2611 3126 2.386e-15
c18707 3886 822 7.99e-16
c18708 1948 1939 3.92e-16
c18709 1556 1942 5.66e-16
c18710 1708 1414 5.5e-16
c18711 1690 1782 1.96e-16
c18712 508 194 1.88e-16
c18713 296 267 3.75e-16
c18714 1335 0 8.1171e-14
c18715 3509 662 1.58e-16
c18716 4915 468 1.88e-16
c18717 602 2219 1.58e-16
c18718 1878 1 8.43e-16
c18719 5291 5385 7.46e-16
c18720 3411 3174 1.58e-16
c18721 3688 3689 9.1e-16
c18722 2488 1 9.28e-16
c18723 596 740 5.28e-16
c18724 288 37 5.71e-16
c18725 245 19 3.84e-16
c18726 3857 858 1.58e-16
c18727 3338 852 1.13e-15
c18728 2458 0 3.6368e-14
c18729 1270 1231 7.84e-16
c18730 1218 1243 1.2e-16
c18731 146 426 1.88e-16
c18732 3876 767 4.48e-16
c18733 2811 2810 5.65e-16
c18734 921 1145 1.96e-16
c18735 1567 812 1.58e-16
c18736 1998 858 3.15e-16
c18737 9 262 5.8e-16
c18738 2196 2372 3.92e-16
c18739 3780 3783 4.87e-16
c18740 3446 4288 2.38e-15
c18741 1876 722 1.09e-16
c18742 1489 1046 1.532e-15
c18743 1495 1494 5.65e-16
c18744 3898 4556 4.22e-16
c18745 2557 2820 3.92e-16
c18746 617 3446 3.15e-16
c18747 4831 4828 6.67e-16
c18748 3214 3211 5.5e-16
c18749 2617 672 5.73e-16
c18750 3135 647 3.64e-16
c18751 3034 3023 1.58e-16
c18752 338 337 2.84e-16
c18753 2364 2361 3.01e-16
c18754 2360 2357 6.44e-16
c18755 234 236 6.01e-16
c18756 230 229 6.4e-16
c18757 4872 1 4.3446e-14
c18758 4651 0 4.34722e-13
c18759 3876 4353 1.58e-16
c18760 3900 4365 5.42e-16
c18761 910 894 5.33e-16
c18762 1254 1253 1.334e-15
c18763 3975 37 1.88e-16
c18764 3976 26 1.075e-15
c18765 4366 3531 1.96e-16
c18766 2321 692 7.38e-16
c18767 2078 852 1.58e-16
c18768 1331 1176 1.58e-16
c18769 888 0 3.854e-14
c18770 1280 1 1.257e-15
c18771 4380 1 9.28e-16
c18772 3667 822 3.79e-16
c18773 4545 0 8e-16
c18774 1706 1730 1.58e-16
c18775 1690 1718 1.58e-16
c18776 3487 662 1.339e-15
c18777 3309 812 7.38e-16
c18778 1 0 8.44442e-13
c18779 2624 0 6.72e-16
c18780 642 3089 1.58e-16
c18781 3387 842 4.48e-16
c18782 4563 4830 1.58e-16
c18783 4580 4842 1.58e-16
c18784 632 3464 7.68e-16
c18785 4453 807 1.58e-16
c18786 4702 5331 5.91e-16
c18787 1254 1264 3.92e-16
c18788 3520 4353 7.84e-16
c18789 1706 807 3.15e-16
c18790 2545 2407 1.58e-16
c18791 2557 777 3.15e-16
c18792 1345 1436 3.92e-16
c18793 4611 4612 1.6e-16
c18794 4607 3874 1.443e-15
c18795 1684 1315 3.54e-16
c18796 2545 3017 6.18e-16
c18797 4883 4497 4.11e-16
c18798 4888 4879 3.46e-16
c18799 3046 2855 1.58e-16
c18800 2702 732 1.58e-16
c18801 2072 2106 1.58e-16
c18802 2022 2036 5.12e-16
c18803 1 514 1.607e-15
c18804 426 320 1.88e-16
c18805 4810 4814 1.81e-16
c18806 1 564 1.073e-15
c18807 3581 3574 1.96e-16
c18808 3185 3583 4.36e-16
c18809 3662 807 1.58e-16
c18810 2196 2337 5.42e-16
c18811 69 1 4.22e-16
c18812 1265 1264 1.6e-16
c18813 3373 2987 1.96e-16
c18814 3370 3809 1.794e-15
c18815 5343 0 1.23e-16
c18816 2887 0 5.6946e-14
c18817 921 752 3.15e-16
c18818 67 0 2.87e-16
c18819 56 19 8.4e-16
c18820 2700 2316 1.58e-16
c18821 1343 1435 1.58e-16
c18822 1327 1423 1.58e-16
c18823 3304 822 3.79e-16
c18824 2231 2220 1.58e-16
c18825 1850 707 7.38e-16
c18826 1812 1803 3.92e-16
c18827 3944 1 5.1e-16
c18828 4136 37 5.71e-16
c18829 2557 2785 1.58e-16
c18830 2541 722 3.15e-16
c18831 507 508 1.88e-16
c18832 3640 807 1.58e-16
c18833 4563 3873 1.58e-16
c18834 3338 3409 5.5e-16
c18835 3344 3393 1.58e-16
c18836 2325 1817 7.84e-16
c18837 5409 5430 1.6e-16
c18838 2249 1732 1.96e-16
c18839 3397 3659 1.58e-16
c18840 5348 5286 6.67e-16
c18841 2214 2605 4.11e-16
c18842 2203 1 4.41e-15
c18843 72 70 2.84e-16
c18844 2984 2988 1.202e-15
c18845 1454 702 1.58e-16
c18846 1321 868 3.15e-16
c18847 1345 827 3.15e-16
c18848 3169 1 1.868e-15
c18849 3839 3775 1.58e-16
c18850 4424 4421 5.5e-16
c18851 4520 4563 1.58e-16
c18852 2545 2773 1.58e-16
c18853 2545 2170 5.5e-16
c18854 602 1315 1.58e-16
c18855 612 1318 5.73e-16
c18856 1625 1627 1.862e-15
c18857 1166 1176 1.418e-15
c18858 2844 837 1.58e-16
c18859 1706 1471 1.58e-16
c18860 632 2260 1.58e-16
c18861 822 1694 7.99e-16
c18862 5081 0 1.5617e-14
c18863 722 732 3.28e-16
c18864 3236 3242 1.418e-15
c18865 4047 4038 1.88e-16
c18866 4567 4395 5.5e-16
c18867 4915 64 1.88e-16
c18868 2502 2493 3.46e-16
c18869 2178 2473 1.58e-16
c18870 2194 1766 1.58e-16
c18871 920 1203 1.58e-16
c18872 2293 672 2.72e-16
c18873 2020 842 1.58e-16
c18874 1684 767 4.48e-16
c18875 1331 1572 4.63e-16
c18876 3521 1 1.716e-15
c18877 1935 767 1.58e-16
c18878 3092 3104 2.32e-16
c18879 2955 2956 3.54e-16
c18880 3463 0 6.9481e-14
c18881 1795 1 1.868e-15
c18882 2764 782 3.15e-16
c18883 2228 2225 3.01e-16
c18884 2224 2221 6.44e-16
c18885 4790 4788 1.6e-16
c18886 1785 0 2.93e-15
c18887 3625 3624 2.48e-16
c18888 3393 3072 1.58e-16
c18889 3411 3467 5.42e-16
c18890 3387 3455 1.58e-16
c18891 2679 707 3.15e-16
c18892 421 436 1.88e-16
c18893 1 219 1.65e-15
c18894 4571 4758 3.92e-16
c18895 2196 1953 1.58e-16
c18896 2182 2473 1.58e-16
c18897 5131 5025 6.31e-16
c18898 687 2651 1.58e-16
c18899 2783 2776 6.73e-16
c18900 1474 692 1.832e-15
c18901 612 3077 2.72e-16
c18902 2867 2475 1.96e-16
c18903 2674 2675 5.65e-16
c18904 3330 1 5.808e-15
c18905 4102 1 7.08e-16
c18906 3900 3616 5.5e-16
c18907 2849 2838 1.58e-16
c18908 4086 37 1.88e-16
c18909 4095 25 4.68e-16
c18910 1691 1714 1.003e-15
c18911 1684 2019 1.58e-16
c18912 1706 2007 1.58e-16
c18913 632 2625 1.09e-16
c18914 2545 692 3.15e-16
c18915 1972 1590 2.48e-16
c18916 792 1559 1.58e-16
c18917 30 439 3.84e-16
c18918 19 419 3.84e-16
c18919 5098 5103 1.493e-15
c18920 5115 5114 3.92e-16
c18921 2749 1 9.28e-16
c18922 894 707 3.15e-16
c18923 890 1038 3.54e-16
c18924 909 1059 1.58e-16
c18925 5170 5160 1.58e-16
c18926 2170 2582 1.96e-16
c18927 537 194 1.88e-16
c18928 3319 1 6.15e-16
c18929 1431 677 3.15e-16
c18930 1630 827 1.58e-16
c18931 1627 868 1.58e-16
c18932 1345 812 3.15e-16
c18933 657 894 8.34e-16
c18934 4028 4031 4.41e-16
c18935 617 3034 3.15e-16
c18936 1862 722 3.15e-16
c18937 826 19 1.96e-16
c18938 3287 1 5.97e-15
c18939 1412 1 6.15e-16
c18940 612 1345 3.58e-16
c18941 3022 3447 4.36e-16
c18942 3445 3438 1.96e-16
c18943 2849 842 3.15e-16
c18944 1926 0 6.72e-16
c18945 4452 1 4.442e-15
c18946 777 1533 1.813e-15
c18947 762 1550 2.22e-16
c18948 868 873 1.097e-15
c18949 5283 5285 5.25e-16
c18950 4022 4023 1.58e-16
c18951 2850 2844 1.6e-16
c18952 602 934 1.078e-15
c18953 4328 3480 4.36e-16
c18954 1151 1589 1.96e-16
c18955 1689 1335 9.72e-16
c18956 2533 2532 1.58e-16
c18957 3048 3275 3.92e-16
c18958 4847 4845 1.687e-15
c18959 4850 4857 6.73e-16
c18960 4469 4856 1.96e-16
c18961 421 349 1.88e-16
c18962 4589 3873 4.9e-16
c18963 4708 4710 4.93e-16
c18964 4582 4711 1.58e-16
c18965 5136 5113 1.58e-16
c18966 3409 3408 1.009e-15
c18967 1964 2473 1.58e-16
c18968 5403 439 3.54e-16
c18969 5253 1 7.87e-16
c18970 2178 2236 1.96e-16
c18971 1209 1216 2.27e-16
c18972 4302 4314 2.32e-16
c18973 2535 2322 1.58e-16
c18974 1516 752 3.15e-16
c18975 1013 1 4.59e-16
c18976 807 26 1.58e-16
c18977 1947 782 1.58e-16
c18978 1788 1784 1.96e-16
c18979 1010 0 1.0077e-14
c18980 4602 1 8.85e-16
c18981 3173 677 1.58e-16
c18982 3046 2583 1.58e-16
c18983 1091 1 5.821e-15
c18984 777 1540 1.58e-16
c18985 677 668 1.078e-15
c18986 0 363 1.12079e-13
c18987 198 197 1.58e-16
c18988 200 201 6.4e-16
c18989 2378 1862 4.11e-16
c18990 2182 2236 4.63e-16
c18991 165 117 1.88e-16
c18992 5242 0 1.65e-16
c18993 279 278 6.67e-16
c18994 129 172 1.88e-16
c18995 1133 767 3.57e-16
c18996 1113 1126 1.58e-16
c18997 3882 3890 8.73e-16
c18998 3876 3895 1.58e-16
c18999 3711 3708 6.44e-16
c19000 1799 647 1.58e-16
c19001 3863 1 2.48e-16
c19002 4394 4385 3.46e-16
c19003 1488 1489 1.35e-16
c19004 4404 1 5.808e-15
c19005 2792 797 5.03e-16
c19006 4406 0 3.466e-15
c19007 3588 762 1.58e-16
c19008 601 2219 7.38e-16
c19009 2094 0 1.65e-16
c19010 420 426 3.84e-16
c19011 3387 3185 5.5e-16
c19012 4950 0 6.278e-14
c19013 1042 1044 7.84e-16
c19014 4753 4748 1.536e-15
c19015 4582 4860 3.92e-16
c19016 5177 5175 3.63e-16
c19017 1523 752 1.339e-15
c19018 1306 1309 5.78e-16
c19019 920 1159 1.58e-16
c19020 542 1 3.4063e-14
c19021 1984 812 4.81e-16
c19022 1601 797 1.58e-16
c19023 1585 1576 3.92e-16
c19024 1131 1579 5.66e-16
c19025 3225 0 3.6012e-14
c19026 4646 4643 5.5e-16
c19027 1836 1454 2.48e-16
c19028 1689 1 6.056e-15
c19029 3325 3326 9.1e-16
c19030 3048 3240 5.42e-16
c19031 3024 3228 1.58e-16
c19032 1854 0 3.3874e-14
c19033 3409 3553 3.92e-16
c19034 827 817 6.38e-16
c19035 1686 0 5.96e-16
c19036 1 188 1.073e-15
c19037 131 0 4.2857e-14
c19038 5136 5047 1.58e-16
c19039 5051 5048 4.69e-16
c19040 4776 323 1.88e-16
c19041 2442 1930 1.532e-15
c19042 2448 2447 5.65e-16
c19043 944 950 6.67e-16
c19044 943 889 3.92e-16
c19045 5559 5543 3.87e-16
c19046 3355 3361 9.59e-16
c19047 1016 677 3.15e-16
c19048 5388 5358 1.604e-15
c19049 2541 822 4.03e-16
c19050 922 995 3.92e-16
c19051 506 505 1.482e-15
c19052 146 160 1.88e-16
c19053 3430 1 1.868e-15
c19054 3420 0 2.93e-15
c19055 2535 2837 3.92e-16
c19056 4182 19 7.04e-16
c19057 4454 4455 2.48e-16
c19058 910 1 4.2163e-14
c19059 4726 4350 3.92e-16
c19060 4738 4737 1.6e-16
c19061 3152 672 2.65e-16
c19062 1321 0 3.17834e-13
c19063 44 43 1.88e-16
c19064 22 21 6.4e-16
c19065 4574 0 6.35e-16
c19066 2023 236 1.163e-15
c19067 836 835 6.67e-16
c19068 5052 5031 1.6e-16
c19069 632 3112 1.58e-16
c19070 281 1 1.9313e-14
c19071 64 178 1.88e-16
c19072 3480 647 3.15e-16
c19073 5355 5382 9.6e-16
c19074 5380 5326 9.34e-16
c19075 5377 5366 3.92e-16
c19076 4821 236 1.88e-16
c19077 2866 852 3.15e-16
c19078 1122 752 4.98e-16
c19079 3736 3726 9.99e-16
c19080 1146 1147 8.58e-16
c19081 3900 4370 1.58e-16
c19082 4569 5546 1.067e-15
c19083 2557 2819 1.58e-16
c19084 2541 2807 1.58e-16
c19085 3228 762 1.58e-16
c19086 2557 2254 1.58e-16
c19087 3990 19 7.04e-16
c19088 3211 3218 1.96e-16
c19089 3030 3041 1.96e-16
c19090 4560 0 5.96e-16
c19091 1929 1533 1.96e-16
c19092 1924 1539 1.96e-16
c19093 1684 1747 1.58e-16
c19094 1706 1735 1.58e-16
c19095 4918 1 3.66e-16
c19096 3034 3048 4.274e-15
c19097 3374 3030 1.96e-16
c19098 1970 1971 1.35e-16
c19099 217 1 1.073e-15
c19100 216 15 5.8e-16
c19101 2634 0 3.5142e-14
c19102 227 0 6.224e-15
c19103 238 30 3.84e-16
c19104 632 3083 3.15e-16
c19105 3782 3770 1.027e-15
c19106 2724 2339 1.96e-16
c19107 2528 2196 3.54e-16
c19108 2048 2056 1.077e-15
c19109 2041 2028 1.58e-16
c19110 1398 1392 1.6e-16
c19111 3639 797 2.33e-16
c19112 3212 0 6.62e-16
c19113 1236 1240 9.24e-16
c19114 372 1 2.87e-16
c19115 3531 4365 1.58e-16
c19116 1794 702 1.58e-16
c19117 2535 792 3.15e-16
c19118 4542 4540 1.96e-16
c19119 4538 3707 3.92e-16
c19120 4555 3701 1.23e-16
c19121 4554 4553 1.6e-16
c19122 3117 662 3.15e-16
c19123 2264 1743 1.96e-16
c19124 3034 2685 1.58e-16
c19125 4722 1 1.013e-15
c19126 1670 1257 1.96e-16
c19127 4827 4829 4.93e-16
c19128 0 310 1.28913e-13
c19129 3397 702 7.99e-16
c19130 2196 2342 1.58e-16
c19131 2178 1817 1.58e-16
c19132 737 729 1.74e-16
c19133 2793 2790 5.5e-16
c19134 1491 732 1.58e-16
c19135 5353 294 9.15e-16
c19136 146 513 1.88e-16
c19137 4270 3429 4.11e-16
c19138 2559 2418 5.5e-16
c19139 2708 2714 1.6e-16
c19140 2705 2316 2.386e-15
c19141 2333 2688 1.58e-16
c19142 2231 2629 4.36e-16
c19143 617 609 1.74e-16
c19144 1478 1476 1.6e-16
c19145 1473 1472 2.03e-16
c19146 601 1372 1.832e-15
c19147 4535 4536 9.1e-16
c19148 1068 0 4.6723e-14
c19149 906 1 3.14e-16
c19150 3204 3203 1.6e-16
c19151 1627 0 3.3846e-14
c19152 3684 1 5.97e-15
c19153 2535 737 4.48e-16
c19154 2250 1 9.28e-16
c19155 602 2196 3.15e-16
c19156 1694 1901 4.63e-16
c19157 747 1345 3.58e-16
c19158 888 884 2.235e-15
c19159 37 535 1.88e-16
c19160 4563 4231 1.58e-16
c19161 2182 1817 1.58e-16
c19162 3486 3487 1.35e-16
c19163 3191 737 1.75e-16
c19164 642 3090 1.58e-16
c19165 2337 1828 1.58e-16
c19166 890 1112 1.96e-16
c19167 3 4 6.67e-16
c19168 2612 1 1.868e-15
c19169 1448 717 1.58e-16
c19170 2662 1 5.97e-15
c19171 1385 971 1.96e-16
c19172 884 1 2.392e-15
c19173 873 0 7.86e-15
c19174 3189 3190 9.1e-16
c19175 601 1315 1.58e-16
c19176 1443 1 2.054e-15
c19177 2833 827 7.68e-16
c19178 1684 1488 1.58e-16
c19179 1690 1482 5.88e-16
c19180 1694 1703 1.58e-16
c19181 1445 0 8e-16
c19182 3475 3472 5.5e-16
c19183 3259 3260 1.35e-16
c19184 2323 1817 3.92e-16
c19185 3034 3347 1.58e-16
c19186 1584 0 6.9481e-14
c19187 3279 797 1.58e-16
c19188 1726 2242 4.11e-16
c19189 3771 3769 3.25e-16
c19190 4060 4067 7.81e-16
c19191 4567 4412 5.5e-16
c19192 4753 323 1.88e-16
c19193 2508 2507 9.1e-16
c19194 2194 2490 1.58e-16
c19195 2178 2478 1.58e-16
c19196 1327 692 3.15e-16
c19197 2904 2877 1.79e-16
c19198 2884 2881 2.208e-15
c19199 4457 782 1.9e-16
c19200 4340 4339 5.65e-16
c19201 4334 3497 1.532e-15
c19202 1431 996 1.136e-15
c19203 632 1343 4.46e-16
c19204 3547 1 8.43e-16
c19205 4597 4594 3.01e-16
c19206 4135 1 6.03e-16
c19207 2663 677 7.68e-16
c19208 2194 782 4.46e-16
c19209 2747 2753 1.418e-15
c19210 2103 2122 7.95e-16
c19211 1 353 4.92e-16
c19212 3411 3472 1.58e-16
c19213 3397 3485 4.63e-16
c19214 4571 4775 3.92e-16
c19215 2182 2478 1.58e-16
c19216 3559 3555 1.96e-16
c19217 512 511 2.84e-16
c19218 0 339 1.3976e-13
c19219 3882 702 4.03e-16
c19220 5484 5452 1.58e-16
c19221 4742 5262 1.96e-16
c19222 1203 890 3.54e-16
c19223 1232 1234 1.66e-16
c19224 922 1053 1.58e-16
c19225 687 1440 1.58e-16
c19226 707 1 3.1284e-14
c19227 2509 2968 7.46e-16
c19228 687 919 3.15e-16
c19229 827 19 1.676e-15
c19230 2656 677 5.03e-16
c19231 747 1088 1.58e-16
c19232 657 1 4.1542e-14
c19233 3190 717 2.4e-16
c19234 3034 3139 4.63e-16
c19235 2193 1 2.94e-16
c19236 792 1579 1.58e-16
c19237 707 701 1.74e-16
c19238 552 549 3.54e-16
c19239 548 535 4.67e-16
c19240 513 320 1.88e-16
c19241 3644 782 1.9e-16
c19242 4776 265 1.88e-16
c19243 1879 2402 4.36e-16
c19244 2400 2393 1.96e-16
c19245 2196 1777 5.5e-16
c19246 5083 1 1.257e-15
c19247 4938 4943 7.25e-16
c19248 2311 2312 5.65e-16
c19249 2185 0 6.35e-16
c19250 3411 3387 4.383e-15
c19251 3397 3869 6.18e-16
c19252 4821 5031 9.82e-16
c19253 612 3071 2.4e-16
c19254 2762 1 6.15e-16
c19255 3328 1 1.716e-15
c19256 1355 1354 2.48e-16
c19257 3775 1 1.021e-15
c19258 4406 4404 2.15e-16
c19259 4414 4413 1.6e-16
c19260 1609 1161 2.48e-16
c19261 627 1345 3.58e-16
c19262 4700 4694 7.25e-16
c19263 4310 4316 9.42e-16
c19264 2833 812 3.64e-16
c19265 3622 0 3.6368e-14
c19266 374 361 1.108e-15
c19267 4974 4972 3.54e-16
c19268 4944 4999 3.18e-16
c19269 3366 852 2.42e-16
c19270 780 779 1.6e-16
c19271 3896 3895 1.736e-15
c19272 3409 3219 5.5e-16
c19273 592 787 1.96e-16
c19274 5464 1 1.257e-15
c19275 2543 0 4.64e-16
c19276 1990 842 1.58e-16
c19277 1618 837 3.79e-16
c19278 1321 1091 5.5e-16
c19279 1331 1542 1.58e-16
c19280 911 1318 1.88e-16
c19281 3452 1 4.41e-15
c19282 2533 3084 4.36e-16
c19283 3082 3075 1.96e-16
c19284 2741 737 1.9e-16
c19285 1882 1880 1.6e-16
c19286 4286 0 6.62e-16
c19287 3347 3349 2.15e-16
c19288 1 441 4.848e-15
c19289 479 136 1.88e-16
c19290 281 363 1.88e-16
c19291 3236 3604 1.96e-16
c19292 4725 4732 1.81e-16
c19293 4582 4728 1.58e-16
c19294 4759 33 1.88e-16
c19295 3397 3421 1.58e-16
c19296 2487 2481 1.6e-16
c19297 1964 2478 2.386e-15
c19298 1970 2486 1.136e-15
c19299 963 976 1.58e-16
c19300 5409 0 3.6422e-14
c19301 5165 238 3.19e-16
c19302 2194 2253 3.92e-16
c19303 3886 672 7.99e-16
c19304 2896 0 2.703e-14
c19305 2559 2339 1.58e-16
c19306 1035 1 3.06e-16
c19307 812 19 1.676e-15
c19308 3354 3345 3.46e-16
c19309 4619 1 8.85e-16
c19310 1694 1607 1.58e-16
c19311 2022 1 4.493e-15
c19312 612 19 1.41e-15
c19313 0 487 1.4803e-14
c19314 136 189 1.88e-16
c19315 5064 5073 2.177e-15
c19316 1658 0 1.6392e-14
c19317 111 19 3.2e-16
c19318 94 0 1.4515e-14
c19319 3503 677 2.33e-16
c19320 1133 1134 1.213e-15
c19321 2578 2572 1.6e-16
c19322 2166 2569 2.386e-15
c19323 1425 1421 1.96e-16
c19324 657 3463 1.813e-15
c19325 910 1317 1.58e-16
c19326 77 76 2.84e-16
c19327 3262 0 3.3874e-14
c19328 790 1 3.79e-16
c19329 4036 19 3.84e-16
c19330 4424 1 2.054e-15
c19331 4426 0 8e-16
c19332 1355 0 3.3608e-14
c19333 257 253 1.372e-15
c19334 248 247 7.08e-16
c19335 244 262 1.58e-16
c19336 3423 3419 1.96e-16
c19337 2987 2995 3.422e-15
c19338 2070 0 4.1103e-14
c19339 2502 1 8.43e-16
c19340 592 742 1.96e-16
c19341 4582 4877 3.92e-16
c19342 2752 2384 1.96e-16
c19343 4111 857 1.88e-16
c19344 4004 4005 7.45e-16
c19345 4012 4014 2.239e-15
c19346 3092 1 5.808e-15
c19347 2823 2824 2.48e-16
c19348 1091 1068 6.54e-16
c19349 687 1027 1.58e-16
c19350 3094 0 3.466e-15
c19351 3904 0 1.23e-16
c19352 2541 2475 1.58e-16
c19353 1690 1786 1.58e-16
c19354 911 1345 3.45e-16
c19355 910 1321 5.22e-16
c19356 4228 0 1.63249e-13
c19357 4219 26 1.075e-15
c19358 1874 0 1.4092e-14
c19359 1 332 2.946e-15
c19360 4753 265 1.88e-16
c19361 911 3388 2.09e-16
c19362 2371 2372 9.1e-16
c19363 1192 1193 7.46e-16
c19364 3463 3452 1.58e-16
c19365 4413 737 3.64e-16
c19366 5451 5447 3.54e-16
c19367 1690 702 4.03e-16
c19368 919 1009 1.58e-16
c19369 3886 3879 1.58e-16
c19370 3022 1 5.277e-15
c19371 4199 25 3.84e-16
c19372 2559 2854 3.92e-16
c19373 1768 1770 2.03e-16
c19374 1142 0 1.0183e-14
c19375 4848 4845 6.67e-16
c19376 3143 677 1.58e-16
c19377 4674 4293 5.2e-16
c19378 2196 2376 1.58e-16
c19379 2276 0 3.466e-15
c19380 2196 2171 2.38e-16
c19381 107 565 1.88e-16
c19382 4872 410 1.88e-16
c19383 2637 2644 1.96e-16
c19384 3650 3259 1.136e-15
c19385 3416 0 2.96e-16
c19386 2136 2031 1.58e-16
c19387 1595 812 5.03e-16
c19388 1151 1148 1.984e-15
c19389 4276 3435 1.136e-15
c19390 2535 2836 1.58e-16
c19391 2557 2824 1.58e-16
c19392 1380 1352 2.64e-16
c19393 955 0 2.4253e-14
c19394 745 1 3.79e-16
c19395 4394 1 8.43e-16
c19396 2786 782 7.38e-16
c19397 1708 1764 5.42e-16
c19398 1684 1752 1.58e-16
c19399 436 432 1.58e-16
c19400 451 455 1.58e-16
c19401 1851 2359 7.84e-16
c19402 602 2192 1.58e-16
c19403 735 734 1.6e-16
c19404 4910 1 5.265e-15
c19405 2266 1743 4.36e-16
c19406 2257 2264 1.96e-16
c19407 228 224 1.372e-15
c19408 632 626 1.74e-16
c19409 3397 3151 5.5e-16
c19410 410 0 1.2388e-13
c19411 4531 0 5.8003e-14
c19412 2441 1 4.41e-15
c19413 1040 677 5.74e-16
c19414 592 697 1.96e-16
c19415 4770 33 1.88e-16
c19416 2734 2367 1.58e-16
c19417 2913 2917 3.82e-16
c19418 3633 812 1.58e-16
c19419 5547 5535 7.95e-16
c19420 5530 5540 1.125e-15
c19421 3227 0 2.93e-15
c19422 1277 1275 8.86e-16
c19423 657 1010 1.85e-16
c19424 748 1 1.65e-16
c19425 3531 4370 2.386e-15
c19426 4379 4373 1.6e-16
c19427 3218 3209 3.46e-16
c19428 1327 1640 1.96e-16
c19429 1566 1106 1.96e-16
c19430 1561 1116 1.96e-16
c19431 4628 4629 1.6e-16
c19432 4624 4242 1.443e-15
c19433 1226 1 4.915e-15
c19434 2305 702 1.58e-16
c19435 2172 837 3.15e-16
c19436 762 592 5.8e-16
c19437 2815 807 2.22e-16
c19438 4739 1 1.013e-15
c19439 2163 2162 1.6e-16
c19440 2164 1635 1.23e-16
c19441 2149 1641 3.92e-16
c19442 2153 2151 1.96e-16
c19443 1 34 5.62e-16
c19444 3659 3657 1.862e-15
c19445 4844 4851 1.81e-16
c19446 5272 5259 8.94e-16
c19447 5269 5230 1.738e-15
c19448 27 28 7.03e-16
c19449 2431 2429 1.6e-16
c19450 2426 2425 2.03e-16
c19451 792 2410 1.58e-16
c19452 2194 1834 1.58e-16
c19453 3836 3370 1.383e-15
c19454 3037 0 6.35e-16
c19455 4392 722 1.09e-16
c19456 1694 672 7.99e-16
c19457 1345 1440 1.58e-16
c19458 627 634 1.6e-16
c19459 1046 1470 1.96e-16
c19460 617 1372 1.58e-16
c19461 3898 4523 1.58e-16
c19462 3876 4535 1.58e-16
c19463 3707 4539 1.96e-16
c19464 1102 0 1.8851e-14
c19465 2139 1667 5.5e-16
c19466 2104 1249 2.24e-16
c19467 3586 3587 9.1e-16
c19468 4555 1 8e-16
c19469 4712 4709 6.67e-16
c19470 2871 842 1.58e-16
c19471 2263 1 6.15e-16
c19472 601 2196 3.15e-16
c19473 314 313 1.58e-16
c19474 4563 4248 1.58e-16
c19475 2418 2413 1.642e-15
c19476 2342 1828 2.386e-15
c19477 1845 2325 1.58e-16
c19478 2793 1 2.054e-15
c19479 2703 2316 1.532e-15
c19480 223 9 5.8e-16
c19481 2795 0 8e-16
c19482 2231 1 5.97e-15
c19483 601 618 1.621e-15
c19484 3014 3003 3.92e-16
c19485 1854 707 1.832e-15
c19486 1482 702 2.22e-16
c19487 3205 1 1.056e-15
c19488 1136 1135 3.94e-16
c19489 3964 1 4.64e-16
c19490 4657 5484 4.06e-16
c19491 2384 782 1.58e-16
c19492 2662 2634 2.64e-16
c19493 3192 3196 1.96e-16
c19494 1708 1505 1.58e-16
c19495 1706 1499 5.5e-16
c19496 1694 1900 1.58e-16
c19497 3113 3111 1.6e-16
c19498 1461 0 6.72e-16
c19499 3387 3672 3.92e-16
c19500 3310 3311 1.35e-16
c19501 3299 797 1.58e-16
c19502 3653 3651 1.6e-16
c19503 4567 4429 5.5e-16
c19504 5486 410 3.54e-16
c19505 2511 2004 1.96e-16
c19506 3731 3732 3.92e-16
c19507 4922 4878 3.41e-16
c19508 1321 707 4.48e-16
c19509 1371 1372 2.48e-16
c19510 2955 1 4.651e-15
c19511 2535 2599 3.92e-16
c19512 657 1321 3.15e-16
c19513 663 19 1.58e-16
c19514 1690 1693 1.96e-16
c19515 1224 1 4.895e-15
c19516 689 690 1.6e-16
c19517 3277 797 1.339e-15
c19518 4807 4805 1.6e-16
c19519 3192 722 1.339e-15
c19520 2162 2078 3.96e-16
c19521 1 565 5.2833e-14
c19522 3393 3100 5.88e-16
c19523 4776 4782 5.87e-16
c19524 4571 4792 3.92e-16
c19525 5200 5219 4.78e-16
c19526 4674 468 1.88e-16
c19527 1879 1 5.97e-15
c19528 0 556 5.6012e-14
c19529 747 19 1.41e-15
c19530 3723 3355 1.96e-16
c19531 5414 468 3.54e-16
c19532 687 2679 2.22e-16
c19533 777 2391 1.58e-16
c19534 3876 717 3.15e-16
c19535 2688 2687 2.48e-16
c19536 1925 782 1.84e-16
c19537 687 1460 1.58e-16
c19538 3523 0 3.3874e-14
c19539 3378 3377 1.6e-16
c19540 3379 2849 1.23e-16
c19541 3362 2855 3.92e-16
c19542 1851 1852 1.35e-16
c19543 426 424 1.257e-15
c19544 1989 1601 4.97e-16
c19545 305 303 1.88e-16
c19546 314 320 1.58e-16
c19547 25 201 7.06e-16
c19548 49 218 1.88e-16
c19549 489 485 1.372e-15
c19550 2200 0 1.23e-16
c19551 3520 717 5.73e-16
c19552 1149 797 1.58e-16
c19553 3381 4234 2.386e-15
c19554 4243 4237 1.6e-16
c19555 5284 5308 6.16e-16
c19556 3354 1 8.43e-16
c19557 1818 692 1.339e-15
c19558 1438 1449 1.96e-16
c19559 687 894 8.34e-16
c19560 99 107 1.58e-16
c19561 4542 858 1.58e-16
c19562 854 1 7.18e-16
c19563 4100 37 1.88e-16
c19564 3876 4298 3.92e-16
c19565 2374 752 1.339e-15
c19566 857 0 5.118e-14
c19567 1973 1985 2.32e-16
c19568 81 1 1.44e-16
c19569 117 484 1.88e-16
c19570 5074 5114 4.39e-16
c19571 349 342 3.54e-16
c19572 3457 3455 2.15e-16
c19573 3465 3464 1.6e-16
c19574 2552 1 7.228e-15
c19575 4469 4850 5.66e-16
c19576 1068 707 1.58e-16
c19577 397 1 2.6688e-14
c19578 4536 842 1.58e-16
c19579 5588 5590 1.6e-16
c19580 3882 4297 1.58e-16
c19581 4318 4317 2.03e-16
c19582 4323 4321 1.6e-16
c19583 1812 1420 1.96e-16
c19584 612 923 1.05e-15
c19585 658 1 1.65e-16
c19586 1192 1 3.54e-16
c19587 1667 1676 1.6e-16
c19588 3450 3451 9.1e-16
c19589 1189 0 9.602e-15
c19590 5026 120 3.54e-16
c19591 4623 4629 5.87e-16
c19592 983 984 1.213e-15
c19593 3944 857 3.1e-16
c19594 5561 497 6.06e-16
c19595 1459 692 5.03e-16
c19596 1230 858 9.11e-16
c19597 3900 677 3.15e-16
c19598 2945 0 1.65e-16
c19599 920 1055 3.92e-16
c19600 921 1054 2.54e-16
c19601 1903 767 1.339e-15
c19602 1523 1525 1.862e-15
c19603 1076 1086 1.418e-15
c19604 1345 957 5.5e-16
c19605 1327 1368 1.96e-16
c19606 837 0 2.86563e-13
c19607 3024 2594 5.5e-16
c19608 3034 3109 1.58e-16
c19609 1319 0 6.969e-14
c19610 1565 1 6.15e-16
c19611 4636 1 8.85e-16
c19612 3160 702 1.58e-16
c19613 2079 2067 1.027e-15
c19614 3893 3401 5.8e-16
c19615 3521 3523 1.862e-15
c19616 2164 1 8e-16
c19617 777 1561 2.72e-16
c19618 627 19 1.41e-15
c19619 325 323 3.84e-16
c19620 2389 2388 9.1e-16
c19621 165 479 1.88e-16
c19622 3883 3901 1.94e-16
c19623 602 3044 1.58e-16
c19624 2865 2469 1.96e-16
c19625 2705 0 3.3717e-14
c19626 3488 0 2.93e-15
c19627 3282 0 1.4092e-14
c19628 2545 2718 4.63e-16
c19629 1349 1344 9.6e-16
c19630 809 1 7.18e-16
c19631 3861 1 5.01e-16
c19632 3856 0 6.78e-16
c19633 2803 807 2.4e-16
c19634 2541 672 4.03e-16
c19635 2557 647 4.46e-16
c19636 3599 777 1.813e-15
c19637 4442 0 6.72e-16
c19638 4905 4923 4.06e-16
c19639 5277 352 7.38e-16
c19640 4940 4939 2.67e-16
c19641 3024 807 3.15e-16
c19642 165 189 1.88e-16
c19643 2520 1 1.106e-15
c19644 1057 1058 7.46e-16
c19645 4582 4894 3.92e-16
c19646 4922 1 3.3585e-14
c19647 4855 468 1.88e-16
c19648 2572 2573 5.65e-16
c19649 2136 1667 7.46e-16
c19650 5577 0 3.9123e-14
c19651 4617 497 1.88e-16
c19652 3722 3397 1.58e-16
c19653 3886 797 3.15e-16
c19654 5573 5429 9.7e-16
c19655 5561 5569 2.78e-15
c19656 3260 0 1.6491e-14
c19657 2541 2299 5.88e-16
c19658 1544 752 1.9e-16
c19659 2557 2492 1.58e-16
c19660 613 1 1.65e-16
c19661 4663 4660 5.5e-16
c19662 3143 3142 2.48e-16
c19663 3060 3056 1.96e-16
c19664 1853 1465 4.97e-16
c19665 3046 2736 1.58e-16
c19666 2187 2181 1.6e-16
c19667 1 475 4.22e-16
c19668 15 454 6.58e-16
c19669 1 478 1.073e-15
c19670 136 135 3.84e-16
c19671 3219 3591 1.58e-16
c19672 3411 752 3.15e-16
c19673 4102 857 1.88e-16
c19674 5160 5159 5.25e-16
c19675 4821 178 1.88e-16
c19676 4759 526 1.88e-16
c19677 2460 2461 2.48e-16
c19678 2172 2206 1.58e-16
c19679 99 1 4.59e-16
c19680 3582 737 3.15e-16
c19681 4674 64 1.88e-16
c19682 1684 717 3.15e-16
c19683 3629 0 6.72e-16
c19684 3466 1 1.056e-15
c19685 1837 1849 2.32e-16
c19686 595 920 3.47e-16
c19687 602 921 3.15e-16
c19688 4763 0 7.67e-16
c19689 1706 1952 3.92e-16
c19690 15 164 6.58e-16
c19691 114 25 7.06e-16
c19692 4580 4707 3.92e-16
c19693 762 1538 2.4e-16
c19694 26 172 1.03e-15
c19695 5388 352 1.58e-16
c19696 5211 1 3.36e-16
c19697 2296 0 8e-16
c19698 3822 3821 3.92e-16
c19699 3828 3820 1.96e-16
c19700 996 662 1.75e-16
c19701 883 807 3.15e-16
c19702 2266 2257 3.92e-16
c19703 1749 2260 5.66e-16
c19704 4315 647 1.58e-16
c19705 4188 4191 4.41e-16
c19706 4217 3918 2.48e-16
c19707 1615 812 1.09e-16
c19708 3882 3548 5.88e-16
c19709 3876 3554 1.58e-16
c19710 4600 5422 4.79e-16
c19711 2559 2853 5.42e-16
c19712 2535 2841 1.58e-16
c19713 2401 807 1.58e-16
c19714 2668 2669 1.35e-16
c19715 2545 2654 1.58e-16
c19716 764 1 7.18e-16
c19717 4008 25 7.01e-16
c19718 2342 717 1.58e-16
c19719 2153 858 1.58e-16
c19720 1196 1661 1.885e-15
c19721 1941 1550 4.11e-16
c19722 1708 1769 1.58e-16
c19723 1715 1716 1.35e-16
c19724 1061 0 7.4292e-14
c19725 911 19 1.676e-15
c19726 3504 3505 2.03e-16
c19727 662 655 5.58e-16
c19728 595 1681 1.58e-16
c19729 3330 837 1.58e-16
c19730 3048 767 3.15e-16
c19731 5386 5291 3.87e-16
c19732 2739 2367 1.58e-16
c19733 3667 797 1.58e-16
c19734 4500 812 4.81e-16
c19735 3404 3027 1.159e-15
c19736 3128 3130 1.6e-16
c19737 3124 3125 2.03e-16
c19738 4212 1 6.78e-16
c19739 1837 1 5.808e-15
c19740 4902 4907 3.73e-16
c19741 1839 0 3.466e-15
c19742 233 25 5.71e-16
c19743 612 2166 1.58e-16
c19744 2442 0 1.6491e-14
c19745 3287 837 1.58e-16
c19746 3996 3999 4.41e-16
c19747 792 2430 1.58e-16
c19748 1930 2423 1.96e-16
c19749 2172 1851 1.58e-16
c19750 2178 1845 5.88e-16
c19751 156 1 4.22e-16
c19752 627 2611 2.22e-16
c19753 3052 0 1.23e-16
c19754 919 782 3.15e-16
c19755 920 1113 1.58e-16
c19756 721 25 7.64e-16
c19757 4292 4283 3.46e-16
c19758 1708 677 3.15e-16
c19759 1327 1026 1.58e-16
c19760 617 1392 1.58e-16
c19761 4550 3900 1.96e-16
c19762 2699 692 4.81e-16
c19763 2498 868 1.58e-16
c19764 2178 677 3.15e-16
c19765 3296 3294 1.862e-15
c19766 2787 2781 1.418e-15
c19767 3030 3207 1.96e-16
c19768 2798 2770 2.64e-16
c19769 901 888 2.878e-15
c19770 617 2196 3.15e-16
c19771 2005 1618 1.532e-15
c19772 2011 2010 5.65e-16
c19773 3304 797 1.58e-16
c19774 3687 812 4.81e-16
c19775 3982 3979 5.5e-16
c19776 4563 4265 1.58e-16
c19777 5162 5159 2.05e-15
c19778 2182 1845 5.5e-16
c19779 339 332 7.76e-16
c19780 3602 737 4.81e-16
c19781 5277 294 3.54e-16
c19782 3287 3282 1.642e-15
c19783 642 3111 2.72e-16
c19784 1408 647 5.03e-16
c19785 909 767 3.15e-16
c19786 883 1126 1.88e-16
c19787 907 1119 1.58e-16
c19788 234 239 1.059e-15
c19789 4634 1 1.5399e-14
c19790 2632 2633 9.1e-16
c19791 1483 1474 3.92e-16
c19792 1041 1477 5.66e-16
c19793 1046 1469 1.58e-16
c19794 4174 3918 6.32e-16
c19795 3221 1 9.28e-16
c19796 901 1 9.155e-15
c19797 3982 1 6.76e-16
c19798 3616 4433 1.58e-16
c19799 2182 677 3.15e-16
c19800 1690 1369 1.58e-16
c19801 1734 1352 2.48e-16
c19802 3958 25 3.84e-16
c19803 1684 1516 5.5e-16
c19804 1694 1905 1.58e-16
c19805 439 499 1.58e-16
c19806 325 265 1.58e-16
c19807 218 194 1.88e-16
c19808 2340 1828 1.532e-15
c19809 2346 2345 5.65e-16
c19810 3411 3689 3.92e-16
c19811 3486 677 1.75e-16
c19812 1112 737 1.58e-16
c19813 32 1 4.92e-16
c19814 3723 858 7.38e-16
c19815 4567 4446 5.5e-16
c19816 5229 5239 2.114e-15
c19817 4770 526 1.88e-16
c19818 1389 971 1.58e-16
c19819 1253 1250 3.92e-16
c19820 4352 4353 2.48e-16
c19821 4855 64 1.88e-16
c19822 2559 2616 3.92e-16
c19823 1694 797 3.15e-16
c19824 1321 1605 1.58e-16
c19825 1343 1593 1.58e-16
c19826 699 1 5.57e-16
c19827 4614 4611 3.01e-16
c19828 657 2276 2.72e-16
c19829 1238 0 1.7331e-14
c19830 4152 1 5.1e-16
c19831 4334 0 1.6491e-14
c19832 3364 3362 2.861e-15
c19833 1801 1 1.716e-15
c19834 4480 1 6.275e-15
c19835 3259 3641 2.48e-16
c19836 4793 4796 6.02e-16
c19837 4571 4809 3.92e-16
c19838 5200 5198 1.721e-15
c19839 5388 294 1.58e-16
c19840 2873 1 4.493e-15
c19841 60 1 1.456e-15
c19842 392 117 1.88e-16
c19843 5429 5412 1.92e-16
c19844 5526 5303 9.75e-16
c19845 78 0 5.8699e-14
c19846 59 41 1.58e-16
c19847 3355 3855 1.66e-16
c19848 2509 0 1.6878e-14
c19849 2821 2822 1.35e-16
c19850 1331 986 5.5e-16
c19851 3543 0 1.4092e-14
c19852 3870 4592 1.36e-15
c19853 4601 4595 1.6e-16
c19854 3886 3673 1.58e-16
c19855 4480 4873 1.914e-15
c19856 4136 0 2.0592e-14
c19857 687 1 4.1542e-14
c19858 1610 1 5.808e-15
c19859 3409 3117 5.5e-16
c19860 5198 5251 3.18e-16
c19861 1612 0 3.466e-15
c19862 310 565 1.88e-16
c19863 33 323 1.88e-16
c19864 3951 3953 1.06e-16
c19865 2325 2324 2.48e-16
c19866 2206 0 3.3538e-14
c19867 3710 842 1.832e-15
c19868 3854 3855 2.49e-16
c19869 4379 717 2.65e-16
c19870 5406 5404 5.62e-16
c19871 5427 5428 1.6e-16
c19872 2692 2690 1.6e-16
c19873 2687 2686 2.03e-16
c19874 1143 1157 1.96e-16
c19875 3327 3708 3.92e-16
c19876 3719 3721 1.6e-16
c19877 4152 4151 6.4e-16
c19878 5323 5321 1.373e-15
c19879 59 42 1.138e-15
c19880 2873 2887 5.12e-16
c19881 4520 5580 8.67e-16
c19882 612 3381 1.58e-16
c19883 4419 4430 1.96e-16
c19884 1626 1166 4.97e-16
c19885 3650 0 6.9481e-14
c19886 4936 4941 3.54e-16
c19887 4968 4967 1.6e-16
c19888 1567 1 5.97e-15
c19889 3411 3625 1.58e-16
c19890 3397 3638 4.63e-16
c19891 1072 722 6.38e-16
c19892 2494 2496 2.03e-16
c19893 4047 4049 1.06e-16
c19894 3876 842 4.48e-16
c19895 1106 767 3.15e-16
c19896 1116 1119 1.58e-16
c19897 921 1220 1.96e-16
c19898 3497 4315 1.96e-16
c19899 2559 2581 5.42e-16
c19900 2535 2569 1.58e-16
c19901 1610 1622 2.32e-16
c19902 601 967 1.58e-16
c19903 910 1319 3.45e-16
c19904 3102 3101 1.6e-16
c19905 3094 3092 2.15e-16
c19906 4313 1 1.056e-15
c19907 1886 1505 3.92e-16
c19908 1890 1891 1.6e-16
c19909 3480 0 6.91e-14
c19910 5002 4946 9.34e-16
c19911 466 470 6.38e-16
c19912 410 441 1.88e-16
c19913 4640 4643 6.02e-16
c19914 4580 4367 1.58e-16
c19915 1479 692 1.09e-16
c19916 2775 2771 1.96e-16
c19917 1144 1145 7.51e-16
c19918 631 25 7.64e-16
c19919 3087 3088 9.1e-16
c19920 1343 1385 3.92e-16
c19921 3667 3673 1.418e-15
c19922 4504 4506 1.862e-15
c19923 1574 1 1.716e-15
c19924 4653 1 8.85e-16
c19925 3387 3434 3.92e-16
c19926 3180 702 1.58e-16
c19927 2078 2093 1.96e-16
c19928 565 339 1.88e-16
c19929 4567 4568 9.48e-16
c19930 1851 0 3.6368e-14
c19931 88 421 1.88e-16
c19932 101 100 5.8e-16
c19933 3531 677 1.58e-16
c19934 2959 294 1.038e-15
c19935 2725 0 1.4092e-14
c19936 3886 4451 4.63e-16
c19937 2611 2220 1.136e-15
c19938 1687 1695 3.84e-16
c19939 1679 1680 4.57e-16
c19940 1257 1253 3.03e-16
c19941 1690 2003 1.96e-16
c19942 2559 662 3.15e-16
c19943 1567 1965 4.36e-16
c19944 1963 1956 1.96e-16
c19945 508 455 1.88e-16
c19946 2196 1743 5.5e-16
c19947 3151 702 1.813e-15
c19948 5177 265 1.96e-16
c19949 4804 4418 1.179e-15
c19950 5283 5278 1.81e-15
c19951 2703 0 1.6491e-14
c19952 3748 3757 3.92e-16
c19953 4135 857 6.23e-16
c19954 2194 2406 3.92e-16
c19955 3684 837 3.79e-16
c19956 4506 842 1.58e-16
c19957 595 3030 4.03e-16
c19958 2557 2316 5.5e-16
c19959 2362 732 1.58e-16
c19960 1257 1264 1.077e-15
c19961 602 937 1.11e-16
c19962 3393 3038 3.15e-16
c19963 1635 1630 1.642e-15
c19964 263 267 6.38e-16
c19965 2284 2283 1.6e-16
c19966 3024 2753 1.58e-16
c19967 3030 2747 5.88e-16
c19968 2186 2181 4.17e-16
c19969 276 117 1.88e-16
c19970 596 760 2.45e-16
c19971 2498 0 1.4092e-14
c19972 4589 4593 1.81e-16
c19973 4742 5388 5.5e-16
c19974 1453 677 7.38e-16
c19975 4304 4302 2.15e-16
c19976 4312 4311 1.6e-16
c19977 5450 5466 1.23e-16
c19978 911 923 1.58e-16
c19979 3482 1 9.28e-16
c19980 4566 3879 1.151e-15
c19981 1507 1071 2.48e-16
c19982 1345 1335 5.5e-16
c19983 822 592 5.8e-16
c19984 601 921 3.15e-16
c19985 4571 737 1.33e-16
c19986 1318 1 4.044e-15
c19987 2713 3231 2.38e-15
c19988 1719 0 6.62e-16
c19989 4780 0 7.67e-16
c19990 2541 797 3.15e-16
c19991 2044 2028 2.062e-15
c19992 1684 1969 3.92e-16
c19993 1 364 1.65e-15
c19994 479 291 1.88e-16
c19995 822 2444 1.58e-16
c19996 1726 1721 1.642e-15
c19997 2312 0 6.72e-16
c19998 657 3135 2.65e-16
c19999 1011 672 4e-16
c20000 5160 0 3.8102e-14
c20001 280 279 2.84e-16
c20002 3886 3875 1.58e-16
c20003 2837 2452 1.96e-16
c20004 3245 1 5.808e-15
c20005 2559 2858 1.58e-16
c20006 1780 1778 1.6e-16
c20007 595 890 3.69e-16
c20008 2736 777 5.73e-16
c20009 983 0 1.4198e-14
c20010 4386 4388 2.03e-16
c20011 3237 3226 1.96e-16
c20012 3397 777 7.99e-16
c20013 33 265 1.88e-16
c20014 5010 4967 2.19e-16
c20015 2029 1 1.0179e-14
c20016 907 1007 3.92e-16
c20017 4571 4469 1.58e-16
c20018 4838 120 1.88e-16
c20019 2136 2119 8.15e-16
c20020 3255 1 9.28e-16
c20021 1684 842 4.48e-16
c20022 1345 1657 3.92e-16
c20023 3230 3226 1.96e-16
c20024 642 1778 2.65e-16
c20025 632 1363 1.58e-16
c20026 3617 1 1.868e-15
c20027 1578 1121 4.11e-16
c20028 4645 4646 1.6e-16
c20029 4641 4259 1.443e-15
c20030 2790 782 1.832e-15
c20031 1330 0 1.5577e-14
c20032 4390 0 1.4092e-14
c20033 3396 3404 1.606e-15
c20034 2705 707 1.832e-15
c20035 602 2208 1.9e-16
c20036 1857 1 2.054e-15
c20037 4743 1 1.806e-15
c20038 4896 0 5.5632e-14
c20039 4972 526 1.108e-15
c20040 2719 752 1.75e-16
c20041 1859 0 8e-16
c20042 413 30 6.83e-16
c20043 3393 3552 1.58e-16
c20044 3685 3687 1.6e-16
c20045 827 819 1.74e-16
c20046 596 715 2.45e-16
c20047 3598 3202 1.96e-16
c20048 1766 1 4.41e-15
c20049 9 158 5.8e-16
c20050 1251 1290 6.67e-16
c20051 5540 5529 1.67e-16
c20052 4776 381 1.88e-16
c20053 3849 3836 8.94e-16
c20054 1343 1041 1.58e-16
c20055 506 519 1.58e-16
c20056 3050 3031 9.83e-16
c20057 1431 1829 4.36e-16
c20058 1827 1820 1.96e-16
c20059 1211 1656 1.58e-16
c20060 4183 19 3.45e-16
c20061 1755 1754 1.6e-16
c20062 777 1119 1.58e-16
c20063 3046 3224 3.92e-16
c20064 2159 1708 1.96e-16
c20065 1879 1874 1.642e-15
c20066 1345 1 2.222e-15
c20067 82 88 1.58e-16
c20068 617 1752 1.832e-15
c20069 1206 0 3.7888e-14
c20070 4729 4726 6.67e-16
c20071 2545 767 3.15e-16
c20072 4563 4282 1.58e-16
c20073 2436 2427 3.92e-16
c20074 1919 2430 5.66e-16
c20075 1930 2422 1.58e-16
c20076 5050 5049 1.6e-16
c20077 378 484 1.88e-16
c20078 3469 3470 1.35e-16
c20079 894 782 3.15e-16
c20080 890 1113 3.54e-16
c20081 909 1134 1.58e-16
c20082 996 999 1.58e-16
c20083 2808 0 6.62e-16
c20084 919 923 3.15e-16
c20085 3388 1 2.606e-15
c20086 1471 722 1.75e-16
c20087 1046 1474 1.58e-16
c20088 3039 3033 1.6e-16
c20089 2880 2934 1.191e-15
c20090 933 1 6.14e-16
c20091 3732 1 1.0179e-14
c20092 4168 25 7.01e-16
c20093 3616 4438 1.58e-16
c20094 3991 19 3.45e-16
c20095 1642 1181 1.532e-15
c20096 1648 1647 5.65e-16
c20097 4333 4711 7.84e-16
c20098 2861 858 1.84e-16
c20099 1056 1 4.044e-15
c20100 4552 0 1.1956e-14
c20101 2179 1698 2.035e-15
c20102 1492 0 6.62e-16
c20103 0 563 4.1771e-14
c20104 37 576 1.88e-16
c20105 3882 777 4.03e-16
c20106 632 3105 7.38e-16
c20107 2005 0 1.6491e-14
c20108 909 931 1.58e-16
c20109 233 9 5.8e-16
c20110 4164 4165 7.45e-16
c20111 5355 5370 7.95e-16
c20112 3855 858 9.97e-16
c20113 2178 2004 1.58e-16
c20114 1121 807 1.58e-16
c20115 1409 971 2.38e-15
c20116 1218 920 1.58e-16
c20117 2545 2282 5.5e-16
c20118 2310 692 5.03e-16
c20119 1345 1622 5.42e-16
c20120 1321 1610 1.58e-16
c20121 687 1321 3.15e-16
c20122 371 0 1.4803e-14
c20123 3118 3109 3.92e-16
c20124 2600 3112 5.66e-16
c20125 2611 3104 1.58e-16
c20126 1533 1917 1.58e-16
c20127 564 563 5.8e-16
c20128 4881 4884 5.5e-16
c20129 4497 1 6.299e-15
c20130 3298 812 5.03e-16
c20131 4824 4822 1.6e-16
c20132 5373 5350 8.66e-16
c20133 4571 4826 3.92e-16
c20134 2515 2512 5.5e-16
c20135 2004 2182 1.58e-16
c20136 2416 1 6.15e-16
c20137 1008 1022 1.96e-16
c20138 3310 3692 2.48e-16
c20139 3696 3693 5.5e-16
c20140 3001 1 1.886e-15
c20141 777 2412 2.72e-16
c20142 1061 707 3.15e-16
c20143 2788 2799 1.96e-16
c20144 642 978 1.05e-15
c20145 2521 0 2.7161e-14
c20146 3874 4592 1.58e-16
c20147 2487 842 7.68e-16
c20148 2480 827 1.9e-16
c20149 601 1377 1.09e-16
c20150 1088 1 4.59e-16
c20151 1085 0 1.0077e-14
c20152 2770 3278 2.48e-16
c20153 3024 3172 1.58e-16
c20154 3046 3160 1.58e-16
c20155 1630 1 2.054e-15
c20156 687 2634 5.73e-16
c20157 1632 0 8e-16
c20158 0 535 4.226e-14
c20159 3387 662 4.48e-16
c20160 3409 677 4.46e-16
c20161 3951 3960 3.84e-16
c20162 3965 3964 6.67e-16
c20163 2196 2321 3.92e-16
c20164 2226 0 1.4092e-14
c20165 3548 702 2.22e-16
c20166 5303 5286 1.92e-16
c20167 4844 91 5.88e-16
c20168 2316 2684 1.96e-16
c20169 1163 812 1.58e-16
c20170 1839 707 5.03e-16
c20171 1196 852 1.13e-15
c20172 1459 1026 1.96e-16
c20173 537 455 1.88e-16
c20174 3926 1 7.44e-16
c20175 2395 752 1.9e-16
c20176 1993 1990 5.5e-16
c20177 479 484 1.88e-16
c20178 3470 3481 1.96e-16
c20179 2204 0 1.6491e-14
c20180 1984 1 1.056e-15
c20181 485 483 1.58e-16
c20182 488 494 1.58e-16
c20183 5128 1 3.36e-16
c20184 2329 2327 1.6e-16
c20185 2324 2323 2.03e-16
c20186 3393 3253 5.88e-16
c20187 5320 5318 6.87e-16
c20188 5262 5165 6.72e-16
c20189 2789 2401 4.97e-16
c20190 1009 1010 7.51e-16
c20191 398 390 2.218e-15
c20192 109 103 1.372e-15
c20193 4047 4056 3.84e-16
c20194 4061 4060 6.67e-16
c20195 4142 3918 6.32e-16
c20196 4753 381 1.88e-16
c20197 3310 3338 2.64e-16
c20198 2874 2884 9.99e-16
c20199 3876 4302 1.58e-16
c20200 3900 4314 5.42e-16
c20201 3907 19 3.84e-16
c20202 2016 858 7.68e-16
c20203 1331 1131 1.58e-16
c20204 627 982 1.58e-16
c20205 617 967 6.38e-16
c20206 364 363 7.08e-16
c20207 342 343 1.58e-16
c20208 85 19 8.4e-16
c20209 1798 1799 9.1e-16
c20210 3046 702 3.15e-16
c20211 3168 3163 1.642e-15
c20212 2573 0 6.72e-16
c20213 2072 2082 7.84e-16
c20214 997 978 1.546e-15
c20215 596 625 2.45e-16
c20216 15 338 6.58e-16
c20217 4039 4040 6.4e-16
c20218 4580 4384 1.58e-16
c20219 5108 62 3.54e-16
c20220 1998 1970 2.64e-16
c20221 762 2389 2.4e-16
c20222 3321 3688 1.58e-16
c20223 1223 1222 7.46e-16
c20224 4328 4319 3.92e-16
c20225 4441 782 1.84e-16
c20226 922 1070 3.92e-16
c20227 653 0 1.1353e-14
c20228 3506 1 5.808e-15
c20229 1924 767 1.9e-16
c20230 1321 1402 3.92e-16
c20231 3508 0 3.466e-15
c20232 632 3886 3.15e-16
c20233 4120 1 5.1e-16
c20234 2921 2954 1.58e-16
c20235 2441 837 5.73e-16
c20236 2640 662 1.84e-16
c20237 3046 2804 1.58e-16
c20238 3245 3257 2.32e-16
c20239 4670 1 8.85e-16
c20240 3411 3451 3.92e-16
c20241 2557 868 3.15e-16
c20242 2535 827 4.48e-16
c20243 5194 5195 3.54e-16
c20244 3551 3549 1.6e-16
c20245 5039 5108 3.54e-16
c20246 2196 2257 1.58e-16
c20247 2203 2204 1.35e-16
c20248 5492 5491 1.559e-15
c20249 3855 3865 3.13e-16
c20250 595 2529 1.655e-15
c20251 602 3067 3.64e-16
c20252 2971 0 1.65e-16
c20253 971 968 1.984e-15
c20254 1327 1372 1.58e-16
c20255 1318 1317 3.54e-16
c20256 4135 4136 6.4e-16
c20257 2214 2169 2.64e-16
c20258 2541 2751 1.58e-16
c20259 3828 1 7.49e-16
c20260 4405 4402 6.44e-16
c20261 4409 4406 3.01e-16
c20262 3030 2645 5.88e-16
c20263 1691 1709 1.94e-16
c20264 1703 1683 2.07e-16
c20265 2029 2094 6.67e-16
c20266 4464 1 1.868e-15
c20267 1694 1816 4.63e-16
c20268 4454 0 2.93e-15
c20269 2161 0 1.1956e-14
c20270 3543 707 1.84e-16
c20271 4982 4979 1.931e-15
c20272 5056 1 7.49e-16
c20273 2291 2300 3.92e-16
c20274 1794 2286 1.58e-16
c20275 777 1690 4.03e-16
c20276 907 702 3.15e-16
c20277 5050 0 1.65e-16
c20278 1678 1681 1.576e-15
c20279 3397 3608 1.58e-16
c20280 4922 410 1.88e-16
c20281 858 863 6.38e-16
c20282 2172 2423 3.92e-16
c20283 1106 1109 6.13e-16
c20284 3886 3435 1.58e-16
c20285 2535 2333 5.5e-16
c20286 817 1 5.62e-16
c20287 1136 1602 4.36e-16
c20288 1600 1593 1.96e-16
c20289 4680 4677 5.5e-16
c20290 2807 807 1.58e-16
c20291 3642 792 1.58e-16
c20292 4581 4215 1.988e-15
c20293 4936 4934 6.91e-16
c20294 3048 2770 1.58e-16
c20295 3034 3291 1.58e-16
c20296 2179 2202 1.003e-15
c20297 3618 3611 6.73e-16
c20298 3617 3225 1.96e-16
c20299 2515 0 1.3715e-14
c20300 3710 3411 1.58e-16
c20301 4606 4613 1.81e-16
c20302 5136 5137 3.54e-16
c20303 4725 0 3.22058e-13
c20304 5581 5579 2.61e-16
c20305 2178 1732 1.58e-16
c20306 1220 842 1.58e-16
c20307 602 925 1.58e-16
c20308 2259 647 5.03e-16
c20309 3495 1 6.15e-16
c20310 3641 0 2.93e-15
c20311 608 0 1.1404e-14
c20312 1857 1854 5.5e-16
c20313 3385 0 6.9668e-14
c20314 4488 3656 2.48e-16
c20315 2696 2691 1.642e-15
c20316 2440 797 7.38e-16
c20317 1143 0 4.6723e-14
c20318 617 921 3.15e-16
c20319 3346 3348 2.03e-16
c20320 3225 3610 1.96e-16
c20321 3219 3615 1.96e-16
c20322 4749 4748 2.83e-16
c20323 4752 4361 1.96e-16
c20324 4797 0 7.67e-16
c20325 2535 812 4.48e-16
c20326 2031 2056 1.96e-16
c20327 767 760 5.58e-16
c20328 15 477 5.8e-16
c20329 465 25 5.71e-16
c20330 2464 822 1.58e-16
c20331 2182 1732 1.58e-16
c20332 93 1 2.79e-15
c20333 4770 5158 1.925e-15
c20334 2906 1 3.36e-16
c20335 1451 662 4.81e-16
c20336 890 1187 1.96e-16
c20337 2893 0 2.078e-15
c20338 2688 1 5.808e-15
c20339 612 2535 3.15e-16
c20340 922 677 5.14e-16
c20341 921 1008 1.58e-16
c20342 106 0 1.5723e-14
c20343 1331 1341 3.92e-16
c20344 1345 1317 3.54e-16
c20345 3265 1 2.054e-15
c20346 911 1324 1.58e-16
c20347 657 3480 3.79e-16
c20348 3900 3565 5.5e-16
c20349 2815 2821 1.418e-15
c20350 2832 2804 2.64e-16
c20351 3271 777 2.65e-16
c20352 1684 1968 1.58e-16
c20353 1706 1956 1.58e-16
c20354 1952 1951 9.1e-16
c20355 762 1542 1.58e-16
c20356 5034 5058 1.96e-16
c20357 672 676 2.19e-16
c20358 601 1715 2.33e-16
c20359 595 1726 2.22e-16
c20360 4943 1 1.23e-16
c20361 2677 1 6.15e-16
c20362 909 1022 4.35e-16
c20363 907 1021 1.88e-16
c20364 890 1014 1.58e-16
c20365 2836 2452 1.58e-16
c20366 2563 2558 9.6e-16
c20367 1038 1039 1.21e-16
c20368 1327 767 3.15e-16
c20369 4736 5391 5.5e-16
c20370 1345 1321 4.383e-15
c20371 772 1 5.62e-16
c20372 632 1780 4.81e-16
c20373 642 1397 3.79e-16
c20374 378 392 1.88e-16
c20375 3899 0 1.4914e-14
c20376 1361 1 6.15e-16
c20377 777 775 3.327e-15
c20378 1694 1397 5.5e-16
c20379 2194 858 1.58e-16
c20380 601 2208 5.03e-16
c20381 4760 1 1.806e-15
c20382 762 1499 1.58e-16
c20383 1875 0 6.72e-16
c20384 3393 3557 1.58e-16
c20385 3409 3174 1.58e-16
c20386 2763 2367 1.96e-16
c20387 5576 0 3.26e-15
c20388 5358 1 3.914e-15
c20389 2441 2442 1.35e-16
c20390 2282 2277 1.642e-15
c20391 2739 2737 1.862e-15
c20392 922 1128 1.58e-16
c20393 3480 3452 2.64e-16
c20394 1121 1572 1.96e-16
c20395 1321 1056 1.58e-16
c20396 1327 1046 5.88e-16
c20397 632 642 3.28e-16
c20398 782 1 3.1284e-14
c20399 2004 852 1.58e-16
c20400 632 1694 3.15e-16
c20401 2196 1783 1.58e-16
c20402 792 1331 7.99e-16
c20403 1 262 4.22e-16
c20404 1930 2427 1.58e-16
c20405 5444 439 3.54e-16
c20406 149 30 3.84e-16
c20407 5412 5426 1.455e-15
c20408 2833 1 1.868e-15
c20409 1192 837 1.58e-16
c20410 2823 0 2.93e-15
c20411 3394 1 3.358e-15
c20412 2545 2271 1.58e-16
c20413 1880 722 3.64e-16
c20414 1046 1494 2.38e-15
c20415 542 535 7.76e-16
c20416 3038 3033 4.17e-16
c20417 2931 2929 7.82e-16
c20418 1896 767 3.15e-16
c20419 1751 1363 4.97e-16
c20420 3024 3043 1.58e-16
c20421 3048 3044 3.92e-16
c20422 3898 792 3.15e-16
c20423 2025 1 1.23e-16
c20424 441 437 6.38e-16
c20425 2358 2359 2.48e-16
c20426 4900 4904 5.6e-16
c20427 4537 1 4.69e-16
c20428 894 923 3.54e-16
c20429 64 267 1.88e-16
c20430 59 252 1.88e-16
c20431 2805 2418 1.532e-15
c20432 4804 0 3.64784e-13
c20433 4623 33 1.88e-16
c20434 3321 3693 1.58e-16
c20435 3726 3742 9.43e-16
c20436 1331 737 3.15e-16
c20437 642 3435 5.73e-16
c20438 2330 692 1.09e-16
c20439 1345 1627 1.58e-16
c20440 727 1 5.62e-16
c20441 3210 3212 2.03e-16
c20442 1272 1 1.23e-16
c20443 4631 4628 3.01e-16
c20444 1550 1905 1.58e-16
c20445 1684 1731 3.92e-16
c20446 3492 662 1.84e-16
c20447 4889 4880 2.58e-16
c20448 5190 207 3.15e-16
c20449 3318 812 1.09e-16
c20450 2899 2882 1.541e-15
c20451 371 372 1.58e-16
c20452 3270 3658 4.97e-16
c20453 1 19 5.625e-14
c20454 2425 1 1.716e-15
c20455 2152 2149 6.71e-16
c20456 1032 662 4.98e-16
c20457 1028 677 1.58e-16
c20458 596 680 5.28e-16
c20459 4 44 1.3e-16
c20460 4571 4843 3.92e-16
c20461 5257 5151 6.31e-16
c20462 5229 5232 7.84e-16
c20463 1218 890 1.96e-16
c20464 3898 737 4.46e-16
c20465 632 997 1.58e-16
c20466 2557 0 3.5222e-13
c20467 1550 797 1.58e-16
c20468 1106 1554 1.58e-16
c20469 4242 4592 2e-16
c20470 3874 4609 1.36e-15
c20471 4618 4612 1.6e-16
c20472 1816 1815 9.1e-16
c20473 627 1391 2.72e-16
c20474 1110 1 3.06e-16
c20475 4497 4890 1.872e-15
c20476 3048 3189 5.42e-16
c20477 3024 3177 1.58e-16
c20478 1803 0 3.3874e-14
c20479 4810 4811 9.93e-16
c20480 5232 5227 7.46e-16
c20481 1 583 4.92e-16
c20482 2417 1896 1.96e-16
c20483 2412 1902 1.96e-16
c20484 5333 0 1.5617e-14
c20485 1185 812 6.48e-16
c20486 42 41 1.482e-15
c20487 1859 707 1.09e-16
c20488 3882 4519 1.96e-16
c20489 3005 3006 9.13e-16
c20490 3002 3003 2.49e-16
c20491 2535 2786 3.92e-16
c20492 3963 1 6.78e-16
c20493 4151 19 3.45e-16
c20494 4440 3605 1.96e-16
c20495 4445 3599 1.96e-16
c20496 3952 0 1.632e-14
c20497 602 1731 1.58e-16
c20498 49 334 1.88e-16
c20499 2866 2895 1.048e-15
c20500 2000 1 9.28e-16
c20501 3574 732 1.58e-16
c20502 5291 323 3.54e-16
c20503 1828 2321 1.96e-16
c20504 2603 2601 1.862e-15
c20505 890 904 1.58e-16
c20506 2511 2513 1.6e-16
c20507 4567 5591 6.18e-16
c20508 2730 2339 1.136e-15
c20509 2557 2203 1.58e-16
c20510 2304 677 7.38e-16
c20511 1630 1627 5.5e-16
c20512 4317 1 1.716e-15
c20513 1903 1516 1.532e-15
c20514 1909 1908 5.65e-16
c20515 762 920 3.15e-16
c20516 4867 4866 1.6e-16
c20517 3048 717 3.58e-16
c20518 3397 3106 1.58e-16
c20519 3628 3625 5.5e-16
c20520 1 557 5.62e-16
c20521 4580 4401 1.58e-16
c20522 5505 1 7.87e-16
c20523 4770 207 1.364e-15
c20524 2506 2504 1.6e-16
c20525 3948 3942 1.96e-16
c20526 3161 0 6.62e-16
c20527 3497 4319 1.58e-16
c20528 1760 662 1.58e-16
c20529 1211 868 4.21e-16
c20530 919 1084 1.58e-16
c20531 3526 1 2.054e-15
c20532 602 3411 3.15e-16
c20533 2535 747 3.15e-16
c20534 3528 0 8e-16
c20535 3191 747 5.73e-16
c20536 2657 672 1.58e-16
c20537 1217 0 1.0183e-14
c20538 3365 3362 6.71e-16
c20539 3024 2821 1.58e-16
c20540 3030 2815 5.88e-16
c20541 4687 1 8.85e-16
c20542 3409 3467 1.58e-16
c20543 2685 717 1.58e-16
c20544 2559 852 3.58e-16
c20545 2072 2067 7.46e-16
c20546 2022 2060 9.37e-16
c20547 5198 5214 1.23e-16
c20548 0 192 9.795e-15
c20549 5494 0 1.65e-16
c20550 5039 5133 7.46e-16
c20551 3770 3774 3.54e-16
c20552 612 2566 1.58e-16
c20553 601 3067 7.68e-16
c20554 602 2533 1.58e-16
c20555 78 565 1.88e-16
c20556 2535 2384 5.5e-16
c20557 1321 1401 1.58e-16
c20558 1343 1389 1.58e-16
c20559 2597 2595 1.6e-16
c20560 595 1341 2.13e-16
c20561 1191 1193 7.72e-16
c20562 3882 4455 1.58e-16
c20563 3898 4467 1.58e-16
c20564 1044 0 2.7376e-14
c20565 855 1 1.65e-16
c20566 4108 26 4.58e-16
c20567 4100 0 2.3527e-14
c20568 2070 2029 5.71e-16
c20569 1708 2020 3.92e-16
c20570 3633 1 5.97e-15
c20571 4563 3879 1.96e-16
c20572 3158 2651 3.92e-16
c20573 1983 1982 1.6e-16
c20574 1975 1973 2.15e-16
c20575 1576 0 3.3846e-14
c20576 37 432 1.88e-16
c20577 3157 3539 2.48e-16
c20578 4580 4570 1.58e-16
c20579 4571 4577 1.58e-16
c20580 4582 4578 3.92e-16
c20581 5128 5127 1.6e-16
c20582 3460 3457 3.01e-16
c20583 3456 3453 6.44e-16
c20584 632 2541 3.15e-16
c20585 2291 1794 1.58e-16
c20586 792 1706 3.15e-16
c20587 909 717 3.15e-16
c20588 592 672 5.8e-16
c20589 5303 5301 3.63e-16
c20590 3696 842 1.84e-16
c20591 5165 149 7.46e-16
c20592 1085 707 1.58e-16
c20593 687 3523 1.58e-16
c20594 4152 857 3.1e-16
c20595 595 3423 2.72e-16
c20596 612 3419 1.58e-16
c20597 3315 0 3.466e-15
c20598 2611 1 5.97e-15
c20599 910 3385 3.45e-16
c20600 2545 2531 1.58e-16
c20601 612 965 1.58e-16
c20602 637 1 5.62e-16
c20603 2651 3159 2.48e-16
c20604 1406 1 5.808e-15
c20605 1408 0 3.466e-15
c20606 632 2243 1.84e-16
c20607 363 262 1.88e-16
c20608 2289 2300 1.96e-16
c20609 3034 3296 1.58e-16
c20610 1533 0 6.9184e-14
c20611 2590 2588 1.6e-16
c20612 2096 2031 6.67e-16
c20613 4623 4631 1.81e-16
c20614 2172 2422 1.58e-16
c20615 2194 2410 1.58e-16
c20616 2880 1 1.0179e-14
c20617 1706 737 4.46e-16
c20618 1918 752 1.58e-16
c20619 1524 1076 4.97e-16
c20620 1345 1355 1.58e-16
c20621 3076 3074 2.03e-16
c20622 1177 0 1.8851e-14
c20623 4076 1 4.64e-16
c20624 1746 1 1.056e-15
c20625 2730 2719 1.58e-16
c20626 4814 0 7.67e-16
c20627 3387 3407 3.92e-16
c20628 3393 3386 1.58e-16
c20629 642 2214 1.58e-16
c20630 1834 1 4.41e-15
c20631 592 593 6.34e-16
c20632 2196 1896 5.5e-16
c20633 2343 0 6.62e-16
c20634 3705 3338 1.58e-16
c20635 3770 3773 9.58e-16
c20636 1457 677 1.832e-15
c20637 1031 672 4.21e-16
c20638 1216 852 1.35e-16
c20639 3885 3881 5.8e-16
c20640 2708 1 2.054e-15
c20641 627 2535 3.15e-16
c20642 3134 1 5.97e-15
c20643 1508 1520 2.32e-16
c20644 2921 2967 1.062e-15
c20645 1913 807 1.58e-16
c20646 1784 1403 3.92e-16
c20647 1788 1789 1.6e-16
c20648 4047 37 1.88e-16
c20649 2747 792 1.58e-16
c20650 2029 2026 1.96e-16
c20651 1708 1985 5.42e-16
c20652 1684 1973 1.58e-16
c20653 1540 0 1.6491e-14
c20654 3506 3518 2.32e-16
c20655 26 346 1.03e-15
c20656 200 187 1.108e-15
c20657 2374 2376 1.862e-15
c20658 1862 1868 1.418e-15
c20659 1879 1851 2.64e-16
c20660 617 1715 1.75e-16
c20661 4903 4900 2.48e-16
c20662 4977 4992 1.734e-15
c20663 2686 1 1.716e-15
c20664 1766 2276 1.96e-16
c20665 894 1037 3.92e-16
c20666 909 1036 1.88e-16
c20667 883 1029 1.58e-16
c20668 277 275 1.58e-16
c20669 159 175 3.84e-16
c20670 3712 842 1.9e-16
c20671 2841 2452 2.386e-15
c20672 2824 2469 1.58e-16
c20673 5585 1 3.82e-16
c20674 4617 468 7.45e-16
c20675 2741 747 2.72e-16
c20676 2136 2135 5.5e-16
c20677 3269 1 8.43e-16
c20678 1805 672 2.72e-16
c20679 1610 837 1.58e-16
c20680 1321 782 4.48e-16
c20681 4398 4396 1.6e-16
c20682 5564 5562 3.92e-16
c20683 3635 1 9.28e-16
c20684 4662 4663 1.6e-16
c20685 4658 4276 1.443e-15
c20686 3571 0 3.6368e-14
c20687 5291 265 7.46e-16
c20688 4980 5023 1.489e-15
c20689 4910 4896 1.594e-15
c20690 5012 5007 1.078e-15
c20691 3018 3383 4.65e-16
c20692 2987 2968 1.58e-16
c20693 601 2228 1.09e-16
c20694 4777 1 1.806e-15
c20695 3256 752 4.81e-16
c20696 2747 737 1.58e-16
c20697 1051 1052 1.238e-15
c20698 1042 702 1.58e-16
c20699 9 465 5.8e-16
c20700 13 479 1.88e-16
c20701 3885 3390 1.176e-15
c20702 4100 4102 4.33e-16
c20703 474 0 2.87e-16
c20704 1528 752 1.84e-16
c20705 1295 1314 1.532e-15
c20706 1307 1236 3.92e-16
c20707 1299 1239 3.56e-16
c20708 543 1 1.607e-15
c20709 1847 1846 1.6e-16
c20710 1839 1837 2.15e-16
c20711 1699 0 6.35e-16
c20712 1 195 1.607e-15
c20713 132 0 1.051e-14
c20714 13 189 1.88e-16
c20715 4563 4316 1.58e-16
c20716 1930 2447 2.38e-15
c20717 3725 3739 5.12e-16
c20718 3803 3811 3.54e-16
c20719 3806 3808 3.73e-16
c20720 3355 3820 8.82e-16
c20721 3014 2486 4.69e-16
c20722 1499 722 3.15e-16
c20723 3031 3054 1.003e-15
c20724 923 1 2.207e-15
c20725 4023 1 4.45e-16
c20726 4465 4458 6.73e-16
c20727 4464 3622 1.96e-16
c20728 3312 2804 2.48e-16
c20729 1669 1196 1.96e-16
c20730 1666 1664 1.6e-16
c20731 4546 4538 5.95e-16
c20732 4583 1 2.86e-16
c20733 4350 4728 7.84e-16
c20734 3398 3038 1.018e-15
c20735 1694 1556 1.58e-16
c20736 1519 1 1.056e-15
c20737 4197 0 4.2433e-14
c20738 840 839 1.6e-16
c20739 117 570 1.88e-16
c20740 310 262 1.88e-16
c20741 5010 4993 7.01e-16
c20742 5033 5031 5.25e-16
c20743 5283 352 5.5e-16
c20744 1338 886 1.159e-15
c20745 4300 672 1.58e-16
c20746 5326 5365 1.858e-15
c20747 910 2557 1.014e-15
c20748 911 2535 1.88e-16
c20749 1098 752 1.58e-16
c20750 284 0 1.4803e-14
c20751 1782 647 7.38e-16
c20752 1405 981 2.48e-16
c20753 632 3429 1.58e-16
c20754 642 4294 2.65e-16
c20755 889 0 7.5183e-14
c20756 1708 1748 3.92e-16
c20757 334 194 1.88e-16
c20758 4413 747 2.65e-16
c20759 4580 4299 1.58e-16
c20760 3048 3380 3.54e-16
c20761 3024 3030 4.078e-15
c20762 1211 0 6.9115e-14
c20763 5291 5350 3.54e-16
c20764 2451 1 8.43e-16
c20765 227 19 3.2e-16
c20766 3387 852 3.15e-16
c20767 2735 2350 1.96e-16
c20768 792 26 1.58e-16
c20769 177 1 4.92e-16
c20770 129 9 5.8e-16
c20771 3900 752 3.15e-16
c20772 1071 1073 7.72e-16
c20773 920 1130 3.92e-16
c20774 921 1129 2.54e-16
c20775 2541 2424 1.58e-16
c20776 719 0 7.709e-15
c20777 4284 4286 2.03e-16
c20778 1584 782 1.58e-16
c20779 1121 1542 1.58e-16
c20780 4242 4609 1.58e-16
c20781 3701 4540 1.885e-15
c20782 3048 3194 1.58e-16
c20783 1191 1 4.044e-15
c20784 1645 0 6.62e-16
c20785 3393 692 3.15e-16
c20786 5152 5162 9.99e-16
c20787 4827 439 1.88e-16
c20788 908 891 3.54e-16
c20789 913 888 8.91e-16
c20790 902 893 1.012e-15
c20791 146 508 1.88e-16
c20792 3429 3435 1.418e-15
c20793 4266 4268 1.862e-15
c20794 3446 3418 2.64e-16
c20795 3576 0 3.466e-15
c20796 1476 1031 4.11e-16
c20797 3030 762 4.03e-16
c20798 2900 2895 7.46e-16
c20799 913 1 2.86e-16
c20800 737 26 7.12e-16
c20801 3736 468 1.098e-15
c20802 3117 3112 1.642e-15
c20803 2685 3194 7.84e-16
c20804 2860 842 1.9e-16
c20805 601 1731 7.38e-16
c20806 454 455 3.84e-16
c20807 465 419 1.88e-16
c20808 3491 3106 1.96e-16
c20809 3496 3100 1.96e-16
c20810 4521 0 1.6491e-14
c20811 805 806 6.67e-16
c20812 339 262 1.88e-16
c20813 4 13 1.58e-16
c20814 3387 3293 1.58e-16
c20815 922 924 3.54e-16
c20816 617 3455 1.832e-15
c20817 4623 526 1.88e-16
c20818 2855 0 3.6813e-14
c20819 1391 957 4.11e-16
c20820 1384 1372 2.32e-16
c20821 1319 1318 1.58e-16
c20822 4617 64 1.88e-16
c20823 3175 0 1.6491e-14
c20824 2535 2220 1.58e-16
c20825 2541 2214 5.88e-16
c20826 897 0 6.35e-16
c20827 870 25 1.13e-15
c20828 873 19 1.58e-16
c20829 3932 25 1.88e-16
c20830 1237 1 1.336e-15
c20831 4343 1 8.43e-16
c20832 4522 0 2.93e-15
c20833 1690 1704 3.92e-16
c20834 1708 1712 1.6e-16
c20835 565 563 1.88e-16
c20836 494 484 3.75e-16
c20837 3030 3359 1.58e-16
c20838 2240 2238 1.862e-15
c20839 1743 1715 2.64e-16
c20840 4847 0 3.4756e-14
c20841 2127 2118 3.92e-16
c20842 2103 1652 9.63e-16
c20843 807 814 1.6e-16
c20844 1 512 9.8e-16
c20845 4063 4062 5.5e-16
c20846 4580 4418 1.58e-16
c20847 5151 5223 4.25e-16
c20848 71 88 1.325e-15
c20849 93 94 3.84e-16
c20850 2231 2226 1.642e-15
c20851 2866 3370 1.96e-16
c20852 3622 782 2.33e-16
c20853 3497 4339 2.38e-15
c20854 2302 662 4.81e-16
c20855 1794 647 1.58e-16
c20856 2020 852 2.4e-16
c20857 1327 1589 1.96e-16
c20858 601 3411 3.15e-16
c20859 2688 2700 2.32e-16
c20860 1540 1091 1.532e-15
c20861 1546 1545 5.65e-16
c20862 1331 1001 5.5e-16
c20863 3676 822 1.58e-16
c20864 4594 3870 4.11e-16
c20865 4599 4590 3.46e-16
c20866 2999 2048 9.75e-16
c20867 2955 2521 3.65e-16
c20868 3718 3731 4.68e-16
c20869 4133 1 7.71e-16
c20870 3048 2838 1.58e-16
c20871 3046 2832 5.5e-16
c20872 762 890 3.35e-16
c20873 3265 3262 5.5e-16
c20874 3409 3472 1.58e-16
c20875 4704 1 8.85e-16
c20876 2127 2128 1.6e-16
c20877 1 331 4.59e-16
c20878 3397 647 3.15e-16
c20879 3559 3560 1.6e-16
c20880 3555 3174 3.92e-16
c20881 4582 4581 1.866e-15
c20882 5514 439 1.58e-16
c20883 4878 352 1.88e-16
c20884 762 2393 1.58e-16
c20885 2178 1760 5.88e-16
c20886 2209 1 2.054e-15
c20887 381 33 1.88e-16
c20888 1474 717 1.58e-16
c20889 909 1235 3.54e-16
c20890 883 890 4.078e-15
c20891 3866 3855 3.92e-16
c20892 601 2533 3.15e-16
c20893 627 2566 5.73e-16
c20894 920 722 3.69e-16
c20895 3321 842 3.15e-16
c20896 5296 5309 9.34e-16
c20897 1345 1418 5.42e-16
c20898 1321 1406 1.58e-16
c20899 1196 1173 6.54e-16
c20900 3898 4472 1.58e-16
c20901 3876 4484 1.58e-16
c20902 3715 0 8e-16
c20903 2559 2768 5.42e-16
c20904 2535 2756 1.58e-16
c20905 4500 1 1.056e-15
c20906 2557 707 4.46e-16
c20907 2545 717 7.99e-16
c20908 508 320 1.88e-16
c20909 5106 5103 7.84e-16
c20910 2182 1760 5.5e-16
c20911 707 700 5.58e-16
c20912 3387 3409 4.078e-15
c20913 4945 4941 3.54e-16
c20914 4963 4936 5.87e-16
c20915 3048 842 3.15e-16
c20916 657 2557 3.15e-16
c20917 2311 1794 2.38e-15
c20918 2234 2232 1.6e-16
c20919 2758 0 3.466e-15
c20920 2166 1 5.329e-15
c20921 1448 662 1.58e-16
c20922 1345 837 3.58e-16
c20923 3335 0 8e-16
c20924 3154 1 1.056e-15
c20925 3571 4404 7.84e-16
c20926 4532 858 7.68e-16
c20927 4640 5471 3.92e-16
c20928 1620 1619 1.6e-16
c20929 1612 1610 2.15e-16
c20930 1321 1555 3.92e-16
c20931 4697 4694 5.5e-16
c20932 1684 1431 5.5e-16
c20933 1694 1820 1.58e-16
c20934 3097 3094 3.01e-16
c20935 1892 1890 1.6e-16
c20936 1887 1886 2.03e-16
c20937 374 375 6.4e-16
c20938 4950 4946 1.572e-15
c20939 2849 852 1.13e-15
c20940 3262 782 1.58e-16
c20941 3387 3621 3.92e-16
c20942 5262 5219 3.1e-16
c20943 2536 0 1.4835e-14
c20944 4640 4645 5.53e-16
c20945 5446 1 2.53e-16
c20946 4702 439 1.88e-16
c20947 2475 2486 1.58e-16
c20948 2172 2427 1.58e-16
c20949 1362 877 1.96e-16
c20950 1357 880 1.96e-16
c20951 4440 767 1.9e-16
c20952 919 858 3.15e-16
c20953 920 1188 1.58e-16
c20954 3687 1 1.056e-15
c20955 1708 752 3.15e-16
c20956 1605 1606 9.1e-16
c20957 1327 1554 1.58e-16
c20958 4219 4217 3.54e-16
c20959 629 0 7.709e-15
c20960 4095 1 6.66e-16
c20961 3347 2838 7.84e-16
c20962 2178 752 3.15e-16
c20963 1762 1 9.28e-16
c20964 4769 4378 1.96e-16
c20965 4831 0 7.67e-16
c20966 2036 2038 6.16e-16
c20967 537 534 1.099e-15
c20968 2368 1 1.868e-15
c20969 2358 0 2.93e-15
c20970 3634 767 3.64e-16
c20971 3926 857 1.88e-16
c20972 5116 5115 1.6e-16
c20973 3781 3853 5.95e-16
c20974 3919 3911 1.88e-16
c20975 3882 647 3.15e-16
c20976 4725 5355 6.5e-16
c20977 909 842 3.15e-16
c20978 883 1201 1.88e-16
c20979 907 1194 1.58e-16
c20980 2961 294 9.02e-16
c20981 5358 5401 1.617e-15
c20982 687 3480 1.58e-16
c20983 4489 4501 2.32e-16
c20984 3358 3356 1.6e-16
c20985 2265 672 1.813e-15
c20986 2444 797 1.832e-15
c20987 2182 752 3.15e-16
c20988 1708 1990 1.58e-16
c20989 2104 1 4.651e-15
c20990 595 25 1.58e-16
c20991 19 487 8.82e-16
c20992 3627 767 1.9e-16
c20993 3542 692 1.9e-16
c20994 3347 842 1.832e-15
c20995 617 2249 3.64e-16
c20996 71 37 1.88e-16
c20997 2712 1 8.43e-16
c20998 782 1142 1.58e-16
c20999 1630 837 1.58e-16
c21000 1421 996 3.92e-16
c21001 1425 1426 1.6e-16
c21002 1335 1324 4.097e-15
c21003 4038 37 1.88e-16
c21004 3876 4247 3.92e-16
c21005 3143 3155 2.32e-16
c21006 4903 4916 1.96e-16
c21007 3419 3021 3.92e-16
c21008 3423 3424 1.6e-16
c21009 2279 2276 3.01e-16
c21010 2275 2272 6.44e-16
c21011 627 2242 2.72e-16
c21012 1522 1 4.41e-15
c21013 1906 0 6.62e-16
c21014 4794 1 1.806e-15
c21015 4967 0 1.666e-15
c21016 2503 1 1.387e-15
c21017 1059 692 8.3e-16
c21018 4120 857 3.1e-16
c21019 4878 294 1.88e-16
c21020 2499 0 6.72e-16
c21021 4006 4011 1.96e-16
c21022 4062 3918 6.32e-16
c21023 2834 2827 6.73e-16
c21024 2583 0 3.5142e-14
c21025 2518 2519 3.01e-16
c21026 4303 4300 6.44e-16
c21027 4307 4304 3.01e-16
c21028 1345 1061 5.5e-16
c21029 3381 1 5.329e-15
c21030 4378 4373 1.642e-15
c21031 2533 3023 1.62e-16
c21032 537 146 1.88e-16
c21033 3333 3332 1.6e-16
c21034 3692 3304 4.97e-16
c21035 1698 0 8.1192e-14
c21036 2045 2046 3.92e-16
c21037 1 352 3.36e-15
c21038 5173 5174 1.334e-15
c21039 2869 1 1.056e-15
c21040 1011 1012 8.58e-16
c21041 160 136 1.88e-16
c21042 5472 5471 1.6e-16
c21043 2823 2441 2.48e-16
c21044 3900 3883 3.62e-16
c21045 3882 3885 1.96e-16
c21046 1061 1056 1.58e-16
c21047 3436 0 1.6491e-14
c21048 982 1 3.54e-16
c21049 4208 37 1.88e-16
c21050 3633 3622 1.58e-16
c21051 979 0 9.602e-15
c21052 4361 4711 2e-16
c21053 2713 3224 1.96e-16
c21054 3024 2529 3.54e-16
c21055 3034 3058 1.58e-16
c21056 2025 2026 5.67e-16
c21057 1535 1 9.28e-16
c21058 2196 2186 5.5e-16
c21059 4537 4531 1.02e-15
c21060 4304 662 5.03e-16
c21061 1332 898 1.018e-15
c21062 5270 5136 1.389e-15
c21063 2531 2530 4.57e-16
c21064 1146 812 1.75e-16
c21065 632 4296 4.81e-16
c21066 3231 0 1.4092e-14
c21067 1659 1660 1.6e-16
c21068 1321 1191 1.58e-16
c21069 1327 1181 5.88e-16
c21070 1324 1 8.766e-15
c21071 762 768 1.097e-15
c21072 3518 3134 1.58e-16
c21073 4648 4645 3.01e-16
c21074 2795 782 1.09e-16
c21075 4391 0 6.72e-16
c21076 3582 747 3.79e-16
c21077 4923 4919 6.35e-16
c21078 421 0 1.29165e-13
c21079 287 274 1.58e-16
c21080 4079 4087 3.45e-16
c21081 5044 5230 2.24e-16
c21082 4011 3918 8.1e-16
c21083 5540 5535 5.63e-16
c21084 5514 5482 1.58e-16
c21085 1272 1269 7.59e-16
c21086 1076 1053 6.54e-16
c21087 2557 2441 1.58e-16
c21088 4036 2189 1.96e-16
c21089 4259 4609 2e-16
c21090 4242 4626 1.36e-15
c21091 4635 4629 1.6e-16
c21092 3202 0 6.9481e-14
c21093 1292 0 1.65e-16
c21094 2493 858 1.339e-15
c21095 822 920 3.15e-16
c21096 4571 827 1.33e-16
c21097 3030 2702 1.58e-16
c21098 1674 1 1.601e-15
c21099 1635 2151 1.885e-15
c21100 26 25 1.9927e-14
c21101 3202 3586 1.58e-16
c21102 2427 0 3.3692e-14
c21103 2429 1913 4.11e-16
c21104 4396 722 3.64e-16
c21105 4810 5044 6.17e-16
c21106 1690 647 3.15e-16
c21107 919 965 3.92e-16
c21108 922 964 1.88e-16
c21109 627 631 2.19e-16
c21110 537 320 1.88e-16
c21111 3596 0 8e-16
c21112 3900 4536 3.92e-16
c21113 3364 0 3.931e-14
c21114 3886 4366 4.63e-16
c21115 3046 777 3.15e-16
c21116 2882 2879 7.84e-16
c21117 940 1 1.65e-16
c21118 1257 1667 1.96e-16
c21119 2696 3206 1.58e-16
c21120 4540 1 6.636e-15
c21121 4713 4333 1.96e-16
c21122 2015 868 2.22e-16
c21123 2259 0 3.466e-15
c21124 2014 1 8.43e-16
c21125 2339 2340 1.35e-16
c21126 73 49 1.88e-16
c21127 4810 5230 3.65e-16
c21128 223 1 1.5625e-14
c21129 5326 5345 4.78e-16
c21130 890 902 1.96e-16
c21131 3763 3765 6.91e-16
c21132 1578 797 5.03e-16
c21133 1136 1133 1.984e-15
c21134 4248 4249 1.35e-16
c21135 3882 3497 5.88e-16
c21136 3876 3503 1.58e-16
c21137 2882 2877 7.46e-16
c21138 2559 2802 5.42e-16
c21139 2535 2790 1.58e-16
c21140 2559 2237 1.58e-16
c21141 2557 2231 5.5e-16
c21142 2545 2632 1.58e-16
c21143 3947 25 4.68e-16
c21144 3197 3196 1.6e-16
c21145 3111 2594 4.11e-16
c21146 2769 767 7.38e-16
c21147 3491 647 1.9e-16
c21148 3030 722 3.15e-16
c21149 704 705 1.6e-16
c21150 4864 0 3.4659e-14
c21151 812 803 1.078e-15
c21152 1 294 3.36e-15
c21153 3747 3734 1.138e-15
c21154 4580 4435 1.58e-16
c21155 5484 1 3.914e-15
c21156 2510 2525 1.96e-16
c21157 2508 2196 3.92e-16
c21158 1327 717 4.03e-16
c21159 1381 952 1.96e-16
c21160 1382 1375 6.73e-16
c21161 5417 0 5.8577e-14
c21162 2518 1 5.051e-15
c21163 642 995 1.85e-16
c21164 688 1 1.65e-16
c21165 1811 672 2.22e-16
c21166 617 3411 3.15e-16
c21167 2015 2172 3.92e-16
c21168 3107 3110 6.44e-16
c21169 4319 0 3.3724e-14
c21170 4527 4526 5.65e-16
c21171 4521 3684 1.532e-15
c21172 4571 812 1.33e-16
c21173 1618 1161 1.136e-15
c21174 777 907 3.15e-16
c21175 3197 722 1.84e-16
c21176 1 545 1.44e-16
c21177 647 1007 1.58e-16
c21178 596 652 3.134e-15
c21179 448 449 5.8e-16
c21180 4563 4604 1.58e-16
c21181 4759 497 1.88e-16
c21182 2391 0 1.6491e-14
c21183 1494 717 1.58e-16
c21184 627 3101 2.65e-16
c21185 617 2533 1.58e-16
c21186 2887 294 3.39e-16
c21187 2325 2337 2.32e-16
c21188 4250 3418 2.48e-16
c21189 2305 2697 1.96e-16
c21190 2691 2698 6.73e-16
c21191 2015 2512 1.66e-16
c21192 3108 3110 2.03e-16
c21193 3744 3757 3.18e-16
c21194 3876 4489 1.58e-16
c21195 3900 4501 5.42e-16
c21196 3684 4522 4.97e-16
c21197 2452 827 3.15e-16
c21198 3927 1 4.45e-16
c21199 602 4247 1.58e-16
c21200 1718 1720 2.15e-16
c21201 3262 3269 1.96e-16
c21202 3030 3156 1.96e-16
c21203 3175 2662 1.532e-15
c21204 3168 3556 4.97e-16
c21205 4516 1 9.28e-16
c21206 4327 4690 1.96e-16
c21207 910 2536 7.06e-16
c21208 2213 1 8.43e-16
c21209 1988 1999 1.96e-16
c21210 717 715 3.327e-15
c21211 37 204 1.88e-16
c21212 3168 722 1.58e-16
c21213 2202 0 3.22e-16
c21214 890 722 3.15e-16
c21215 907 1082 3.92e-16
c21216 797 807 3.28e-16
c21217 3397 3259 1.58e-16
c21218 2775 2390 1.96e-16
c21219 1823 692 1.84e-16
c21220 1449 1443 1.6e-16
c21221 601 3440 1.9e-16
c21222 3351 0 6.72e-16
c21223 1121 1120 3.94e-16
c21224 3582 4416 1.58e-16
c21225 3701 858 3.15e-16
c21226 2367 767 1.58e-16
c21227 2379 752 1.84e-16
c21228 1725 1716 3.46e-16
c21229 865 1 5.57e-16
c21230 857 19 3.563e-15
c21231 1708 1448 5.5e-16
c21232 4581 4564 3.54e-16
c21233 1516 1884 1.96e-16
c21234 1420 0 3.6368e-14
c21235 349 343 1.58e-16
c21236 82 0 6.224e-15
c21237 3072 3455 7.84e-16
c21238 4903 4946 2.15e-16
c21239 2315 1794 1.96e-16
c21240 2310 1800 1.96e-16
c21241 642 1749 1.58e-16
c21242 671 670 6.67e-16
c21243 3282 782 1.58e-16
c21244 3034 692 3.15e-16
c21245 1715 2222 2.48e-16
c21246 2542 0 4.1004e-14
c21247 4045 4044 7.81e-16
c21248 602 3434 1.58e-16
c21249 1343 677 4.46e-16
c21250 2858 2870 2.32e-16
c21251 398 0 1.0822e-14
c21252 5417 5486 3.54e-16
c21253 841 25 7.64e-16
c21254 3703 1 9.28e-16
c21255 1667 1661 9.61e-16
c21256 1775 1 6.15e-16
c21257 4856 1 1.749e-15
c21258 3260 782 1.339e-15
c21259 4848 0 7.67e-16
c21260 3175 707 1.339e-15
c21261 2545 842 3.15e-16
c21262 5206 5195 9.85e-16
c21263 3387 3055 1.58e-16
c21264 596 607 3.134e-15
c21265 557 556 3.84e-16
c21266 3253 767 3.15e-16
c21267 1026 692 1.75e-16
c21268 894 858 3.15e-16
c21269 1222 852 1.58e-16
c21270 890 1188 3.54e-16
c21271 909 1209 1.58e-16
c21272 3876 662 4.48e-16
c21273 4434 767 7.38e-16
c21274 378 570 1.88e-16
c21275 4349 692 7.38e-16
c21276 919 1038 1.58e-16
c21277 1908 767 1.84e-16
c21278 1528 1525 5.5e-16
c21279 1331 881 5.5e-16
c21280 837 19 1.41e-15
c21281 2452 812 3.15e-16
c21282 3355 1 1.387e-15
c21283 1698 1689 5.71e-16
c21284 4071 37 1.88e-16
c21285 4072 26 1.075e-15
c21286 4760 4763 6.67e-16
c21287 3030 3121 1.58e-16
c21288 2062 2069 8.94e-16
c21289 2064 2067 1.732e-15
c21290 1559 1 5.808e-15
c21291 1561 0 3.466e-15
c21292 3526 3523 5.5e-16
c21293 2151 1 6.636e-15
c21294 777 1116 4e-16
c21295 333 334 1.88e-16
c21296 339 331 1.58e-16
c21297 5072 5071 2.29e-16
c21298 3885 3890 4.17e-16
c21299 909 1023 3.54e-16
c21300 1619 827 7.68e-16
c21301 1328 1338 5.8e-16
c21302 3854 1 4.03e-16
c21303 3900 4264 3.92e-16
c21304 2357 737 1.339e-15
c21305 819 1 5.57e-16
c21306 2987 0 5.6075e-14
c21307 4679 4680 1.6e-16
c21308 4675 4293 1.443e-15
c21309 2818 797 4.81e-16
c21310 3599 0 6.9134e-14
c21311 3536 692 7.38e-16
c21312 4938 4961 5.87e-16
c21313 4954 4960 1.96e-16
c21314 4989 4991 3.92e-16
c21315 4946 4531 8.77e-16
c21316 3345 858 1.339e-15
c21317 3387 3591 1.58e-16
c21318 3411 3603 5.42e-16
c21319 3393 3208 1.58e-16
c21320 4742 1 2.1168e-14
c21321 4580 0 3.52217e-13
c21322 4770 497 1.88e-16
c21323 2517 0 8e-16
c21324 3321 3411 5.5e-16
c21325 1101 752 2.33e-16
c21326 3898 4234 1.58e-16
c21327 3876 4246 1.58e-16
c21328 4262 1 1.056e-15
c21329 3056 2532 3.92e-16
c21330 3060 3061 1.6e-16
c21331 1852 1863 1.96e-16
c21332 1163 1 4.59e-16
c21333 1160 0 1.0077e-14
c21334 2175 2183 3.84e-16
c21335 5288 5285 2.05e-15
c21336 462 19 8.4e-16
c21337 470 0 5.7133e-14
c21338 479 27 1.88e-16
c21339 223 363 1.88e-16
c21340 3409 752 4.46e-16
c21341 3397 3395 5.93e-16
c21342 2470 1953 1.96e-16
c21343 2471 2464 6.73e-16
c21344 923 955 1.58e-16
c21345 4164 3893 1.96e-16
c21346 1442 677 5.03e-16
c21347 1208 842 3.57e-16
c21348 1188 1201 1.58e-16
c21349 4878 62 1.88e-16
c21350 2015 0 6.102e-14
c21351 921 1025 1.96e-16
c21352 4205 4199 1.96e-16
c21353 1886 752 1.339e-15
c21354 3882 4400 1.96e-16
c21355 4479 4472 1.96e-16
c21356 3633 4481 4.36e-16
c21357 3329 2815 4.97e-16
c21358 4022 26 4.48e-16
c21359 4361 4728 1.58e-16
c21360 3048 2533 5.5e-16
c21361 37 175 1.88e-16
c21362 27 189 1.88e-16
c21363 3621 752 1.58e-16
c21364 3773 3820 1.836e-15
c21365 281 421 1.88e-16
c21366 4321 672 2.72e-16
c21367 1117 1119 7.84e-16
c21368 160 165 1.88e-16
c21369 3702 3696 1.6e-16
c21370 2534 2554 2.07e-16
c21371 1619 812 3.64e-16
c21372 3030 822 4.03e-16
c21373 2541 2666 1.58e-16
c21374 774 1 5.57e-16
c21375 3401 3038 3.84e-16
c21376 1635 858 3.15e-16
c21377 642 1414 2.22e-16
c21378 1661 1673 3.13e-16
c21379 1206 1345 1.58e-16
c21380 1196 1343 5.5e-16
c21381 3881 0 4.3835e-14
c21382 2611 3135 4.36e-16
c21383 3133 3126 1.96e-16
c21384 1937 1939 1.862e-15
c21385 1550 1556 1.418e-15
c21386 1694 1414 5.5e-16
c21387 296 265 1.88e-16
c21388 3523 3134 2.386e-15
c21389 5151 207 3.54e-16
c21390 2652 0 1.6491e-14
c21391 842 836 1.74e-16
c21392 288 19 8.4e-16
c21393 275 0 1.5696e-14
c21394 3858 858 1.58e-16
c21395 1786 647 1.832e-15
c21396 1406 1418 2.32e-16
c21397 2178 2372 1.96e-16
c21398 2814 2805 3.46e-16
c21399 1527 737 1.9e-16
c21400 1293 1296 5.87e-16
c21401 1281 1231 1.96e-16
c21402 922 1145 3.92e-16
c21403 2535 2458 1.58e-16
c21404 4259 4626 1.58e-16
c21405 3138 2628 1.58e-16
c21406 3126 2645 1.58e-16
c21407 1236 0 4.8679e-14
c21408 4199 1 7.08e-16
c21409 1454 0 3.6368e-14
c21410 426 291 1.88e-16
c21411 3393 3536 1.96e-16
c21412 15 251 6.58e-16
c21413 5486 470 1.345e-15
c21414 5068 91 6.67e-16
c21415 595 2569 1.58e-16
c21416 2447 0 1.4092e-14
c21417 2182 2372 4.63e-16
c21418 166 1 1.607e-15
c21419 3054 0 3.22e-16
c21420 152 0 1.4515e-14
c21421 4296 4294 1.6e-16
c21422 5440 5441 2.67e-16
c21423 1684 662 4.48e-16
c21424 2248 2632 1.58e-16
c21425 1498 1489 3.46e-16
c21426 3390 0 8.2949e-14
c21427 3900 3876 4.383e-15
c21428 2697 702 2.65e-16
c21429 822 890 3.35e-16
c21430 3024 792 3.15e-16
c21431 2880 2945 6.67e-16
c21432 3220 3214 1.6e-16
c21433 2696 3211 2.386e-15
c21434 2871 852 2.4e-16
c21435 1618 2010 2.38e-15
c21436 1684 1918 3.92e-16
c21437 5183 5182 1.6e-16
c21438 5154 5157 3.54e-16
c21439 5175 5174 3.92e-16
c21440 430 429 1.58e-16
c21441 425 436 3.84e-16
c21442 642 2600 1.58e-16
c21443 981 647 1.75e-16
c21444 238 236 1.96e-16
c21445 4787 1 2.4547e-14
c21446 4076 4084 6.67e-16
c21447 4082 4072 7.1e-16
c21448 4569 0 3.49037e-13
c21449 3886 4365 1.58e-16
c21450 3898 3514 5.5e-16
c21451 3900 3520 1.58e-16
c21452 2912 2911 2.67e-16
c21453 1745 1744 1.6e-16
c21454 729 1 5.57e-16
c21455 3973 0 1.5061e-14
c21456 3975 19 3.45e-16
c21457 1196 1639 1.58e-16
c21458 1690 1917 1.58e-16
c21459 4446 3605 1.136e-15
c21460 1828 2345 2.38e-15
c21461 3409 3689 3.92e-16
c21462 3718 1 1.492e-15
c21463 3024 737 4.48e-16
c21464 4881 0 3.5099e-14
c21465 5326 5316 1.021e-15
c21466 4 27 1.58e-16
c21467 3397 868 7.99e-16
c21468 4580 4452 1.58e-16
c21469 632 3453 1.339e-15
c21470 2178 2337 1.58e-16
c21471 3650 782 1.58e-16
c21472 5514 5493 2.85e-16
c21473 4702 5345 1.96e-16
c21474 2535 1 3.564e-15
c21475 4363 4356 6.73e-16
c21476 4362 3520 1.96e-16
c21477 1345 1606 3.92e-16
c21478 3191 1 4.41e-15
c21479 2708 2705 5.5e-16
c21480 1331 1436 4.63e-16
c21481 4611 3874 4.11e-16
c21482 4616 4607 3.46e-16
c21483 3013 2559 6.7e-16
c21484 4339 0 1.4092e-14
c21485 1806 1 2.054e-15
c21486 792 883 3.15e-16
c21487 3485 647 7.38e-16
c21488 2141 2131 1.98e-16
c21489 1808 0 8e-16
c21490 1 505 4.59e-16
c21491 3642 3644 2.15e-16
c21492 5165 5226 6.38e-16
c21493 2196 2507 5.42e-16
c21494 3572 3185 1.532e-15
c21495 3270 807 1.813e-15
c21496 4023 857 6.23e-16
c21497 3966 3964 2.254e-15
c21498 792 2401 1.813e-15
c21499 2182 2337 1.58e-16
c21500 2172 1794 5.5e-16
c21501 62 1 3.36e-15
c21502 56 26 1.03e-15
c21503 47 0 9.795e-15
c21504 617 3103 4.81e-16
c21505 922 752 5.14e-16
c21506 921 1083 1.58e-16
c21507 2305 2316 1.58e-16
c21508 1343 996 1.58e-16
c21509 4156 4158 2.254e-15
c21510 3008 3005 1.6e-16
c21511 595 881 2.22e-16
c21512 4327 4322 1.642e-15
c21513 3900 4506 1.58e-16
c21514 2469 868 1.813e-15
c21515 2682 677 4.81e-16
c21516 1801 1803 1.862e-15
c21517 4140 25 1.88e-16
c21518 3956 1 6.78e-16
c21519 4136 19 7.35e-16
c21520 601 4247 7.38e-16
c21521 2104 2070 1.75e-16
c21522 1161 0 3.7577e-14
c21523 507 509 1.58e-16
c21524 4582 3870 1.58e-16
c21525 1896 2405 1.58e-16
c21526 3202 707 1.58e-16
c21527 3585 722 4.81e-16
c21528 5039 1 4.669e-15
c21529 2328 2335 6.73e-16
c21530 3344 3411 1.58e-16
c21531 5409 5404 1.81e-15
c21532 2690 2299 4.11e-16
c21533 687 2557 3.15e-16
c21534 883 737 6.45e-16
c21535 909 1097 4.35e-16
c21536 907 1096 1.88e-16
c21537 890 1089 1.58e-16
c21538 2592 1 6.15e-16
c21539 5284 5345 1.6e-16
c21540 2214 2602 4.97e-16
c21541 1657 858 7.38e-16
c21542 1327 842 3.15e-16
c21543 1331 827 3.15e-16
c21544 2986 2984 1.167e-15
c21545 617 3440 5.03e-16
c21546 3158 1 1.716e-15
c21547 595 4234 1.58e-16
c21548 3599 4404 1.58e-16
c21549 3582 4421 2.386e-15
c21550 4430 4424 1.6e-16
c21551 4514 4582 5.5e-16
c21552 5585 5577 1.6e-16
c21553 3269 3260 3.46e-16
c21554 687 1803 1.58e-16
c21555 1625 1636 1.96e-16
c21556 4327 4689 1.58e-16
c21557 3083 3467 1.58e-16
c21558 1954 0 1.6491e-14
c21559 3409 3625 1.58e-16
c21560 5200 178 1.58e-16
c21561 596 835 2.45e-16
c21562 5317 5314 1.98e-16
c21563 2178 1953 1.58e-16
c21564 3898 827 4.46e-16
c21565 3882 868 4.03e-16
c21566 4536 852 2.4e-16
c21567 4545 858 6.67e-16
c21568 601 3434 7.38e-16
c21569 919 1203 1.58e-16
c21570 1777 662 3.15e-16
c21571 2010 868 1.58e-16
c21572 1345 1571 5.42e-16
c21573 1321 1559 1.58e-16
c21574 858 1 2.8086e-14
c21575 2583 3092 7.84e-16
c21576 2767 752 4.81e-16
c21577 1897 1888 3.92e-16
c21578 1505 1891 5.66e-16
c21579 1516 1883 1.58e-16
c21580 1784 1 1.716e-15
c21581 4786 4395 1.96e-16
c21582 9 187 5.8e-16
c21583 3411 3072 1.58e-16
c21584 2182 1953 1.58e-16
c21585 2386 1 9.28e-16
c21586 2356 0 3.6368e-14
c21587 5412 0 3.8102e-14
c21588 5134 5039 3.87e-16
c21589 1483 692 3.64e-16
c21590 5303 381 1.96e-16
c21591 2775 2776 1.6e-16
c21592 2856 2475 3.92e-16
c21593 3886 3616 5.5e-16
c21594 4509 4506 5.5e-16
c21595 2650 672 2.4e-16
c21596 4086 19 7.04e-16
c21597 1684 1624 1.58e-16
c21598 1690 1618 5.88e-16
c21599 1579 1 2.054e-15
c21600 1581 0 8e-16
c21601 1978 1975 3.01e-16
c21602 1974 1971 6.44e-16
c21603 37 436 1.88e-16
c21604 4582 4559 3.84e-16
c21605 4580 910 1.32e-16
c21606 5111 5114 3.92e-16
c21607 5116 5074 1.017e-15
c21608 5108 5101 9.81e-16
c21609 3497 702 1.58e-16
c21610 894 1038 3.54e-16
c21611 4152 4100 1.88e-16
c21612 1166 827 3.15e-16
c21613 1331 812 3.15e-16
c21614 2541 2735 1.96e-16
c21615 612 1331 7.99e-16
c21616 175 176 7.03e-16
c21617 5151 296 3.54e-16
c21618 3436 3022 1.532e-15
c21619 3442 3441 5.65e-16
c21620 1933 1 1.056e-15
c21621 4759 5174 3.92e-16
c21622 4793 236 1.88e-16
c21623 3876 3486 1.58e-16
c21624 3898 812 4.46e-16
c21625 2848 2841 1.96e-16
c21626 3876 4251 1.58e-16
c21627 3900 4263 5.42e-16
c21628 4317 3480 1.532e-15
c21629 910 1680 1.58e-16
c21630 1185 1 3.06e-16
c21631 602 3900 3.15e-16
c21632 612 3898 3.15e-16
c21633 4278 1 9.28e-16
c21634 4847 4849 2.15e-16
c21635 3034 3275 4.63e-16
c21636 4915 439 1.88e-16
c21637 2179 2197 1.94e-16
c21638 1718 0 3.3643e-14
c21639 4589 4590 9.93e-16
c21640 4567 4711 1.58e-16
c21641 4571 4327 5.5e-16
c21642 3393 3398 8.56e-16
c21643 1964 1953 1.58e-16
c21644 967 969 7.84e-16
c21645 4026 4024 7.1e-16
c21646 1462 677 1.09e-16
c21647 1208 1209 1.213e-15
c21648 3469 4302 7.84e-16
c21649 1518 1517 1.6e-16
c21650 1510 1508 2.15e-16
c21651 1327 1338 1.96e-16
c21652 4065 1 1.895e-14
c21653 2921 2933 5.37e-16
c21654 2923 2918 7.46e-16
c21655 2429 797 5.03e-16
c21656 1790 1788 1.6e-16
c21657 1785 1784 2.03e-16
c21658 4047 0 1.804e-14
c21659 1549 1 8.43e-16
c21660 4378 4728 2e-16
c21661 5158 5182 6.16e-16
c21662 0 342 1.4803e-14
c21663 37 349 1.88e-16
c21664 3508 3506 2.15e-16
c21665 3516 3515 1.6e-16
c21666 1794 0 6.914e-14
c21667 2375 1862 4.97e-16
c21668 2196 2235 5.42e-16
c21669 4708 5338 1.96e-16
c21670 282 286 1.372e-15
c21671 281 275 3.84e-16
c21672 107 305 1.88e-16
c21673 920 672 3.15e-16
c21674 3900 3896 3.92e-16
c21675 4122 4120 7.1e-16
c21676 2136 2072 1.58e-16
c21677 1166 812 3.15e-16
c21678 2736 0 3.5259e-14
c21679 2557 2683 1.58e-16
c21680 2541 2671 1.58e-16
c21681 3865 1 1.052e-15
c21682 2322 722 1.75e-16
c21683 3397 0 3.3139e-13
c21684 4413 1 1.868e-15
c21685 4665 4662 3.01e-16
c21686 508 368 1.88e-16
c21687 4403 0 2.93e-15
c21688 422 420 1.58e-16
c21689 4861 5114 3.92e-16
c21690 4844 5074 7.84e-16
c21691 4993 0 1.63e-15
c21692 1 458 1.44e-16
c21693 3397 3586 1.58e-16
c21694 3728 3729 5.67e-16
c21695 2549 2538 4.097e-15
c21696 4567 4860 3.92e-16
c21697 5538 5537 5.68e-16
c21698 5536 5535 1.96e-16
c21699 2566 1 4.41e-15
c21700 2820 2819 9.1e-16
c21701 1218 1299 1.96e-16
c21702 1300 1295 7.46e-16
c21703 3076 0 6.62e-16
c21704 2345 717 1.58e-16
c21705 1690 868 4.03e-16
c21706 1706 827 4.46e-16
c21707 1667 852 1.58e-16
c21708 919 1159 1.58e-16
c21709 1574 1576 1.862e-15
c21710 1121 1131 1.418e-15
c21711 506 15 5.8e-16
c21712 4276 4626 2e-16
c21713 4259 4643 1.36e-15
c21714 4652 4646 1.6e-16
c21715 3143 2628 2.386e-15
c21716 1690 1386 1.58e-16
c21717 3608 777 1.58e-16
c21718 1842 1839 3.01e-16
c21719 1838 1835 6.44e-16
c21720 4745 1 4.832e-15
c21721 3048 2719 1.58e-16
c21722 3046 2713 5.5e-16
c21723 3034 3240 1.58e-16
c21724 644 643 1.6e-16
c21725 273 274 1.482e-15
c21726 2469 0 6.9484e-14
c21727 752 743 1.078e-15
c21728 9 190 4.88e-16
c21729 1 158 2.946e-15
c21730 128 0 9.795e-15
c21731 5136 5031 1.58e-16
c21732 4861 323 1.88e-16
c21733 2451 2442 3.46e-16
c21734 1243 1231 2.238e-15
c21735 3836 3834 1.609e-15
c21736 5388 5391 3.54e-16
c21737 3002 2486 4.78e-16
c21738 506 507 5.8e-16
c21739 3609 0 6.62e-16
c21740 3419 1 1.716e-15
c21741 2316 702 3.79e-16
c21742 4008 1 5.1e-16
c21743 4182 26 4.48e-16
c21744 4457 4453 1.96e-16
c21745 1752 1761 3.92e-16
c21746 1380 1747 1.58e-16
c21747 1119 0 2.7376e-14
c21748 1708 1684 4.383e-15
c21749 1665 1663 2.61e-16
c21750 3594 3595 5.65e-16
c21751 889 901 5.8e-16
c21752 4730 4350 1.96e-16
c21753 1708 1935 3.92e-16
c21754 37 5 1.88e-16
c21755 4557 0 9.327e-15
c21756 3219 732 2.22e-16
c21757 3591 752 1.58e-16
c21758 632 2594 3.15e-16
c21759 2637 1 5.808e-15
c21760 1115 752 5.74e-16
c21761 4175 4166 1.88e-16
c21762 3027 3035 3.84e-16
c21763 2178 2528 2e-16
c21764 642 1389 1.58e-16
c21765 3400 0 6.35e-16
c21766 1146 1153 7.95e-16
c21767 3886 4370 1.58e-16
c21768 3876 3531 5.5e-16
c21769 2929 2934 1.96e-16
c21770 942 1 1.816e-15
c21771 2781 3305 4.36e-16
c21772 3990 26 4.48e-16
c21773 2696 3209 1.532e-15
c21774 3214 3215 5.65e-16
c21775 3034 3033 1.357e-15
c21776 1181 1647 2.38e-15
c21777 2628 662 3.15e-16
c21778 3882 0 3.63418e-13
c21779 1921 1539 2.48e-16
c21780 1293 1 1.594e-15
c21781 647 639 1.74e-16
c21782 2010 0 1.4092e-14
c21783 2647 1 9.28e-16
c21784 890 962 1.96e-16
c21785 233 1 4.22e-16
c21786 3706 827 1.58e-16
c21787 2802 2435 1.58e-16
c21788 3287 3654 1.58e-16
c21789 3276 3662 5.66e-16
c21790 3668 3659 3.92e-16
c21791 5484 410 7.46e-16
c21792 2721 2339 2.48e-16
c21793 2528 2182 6.18e-16
c21794 2041 2055 9.34e-16
c21795 1396 1389 1.96e-16
c21796 3049 1 2.86e-16
c21797 2194 2354 1.58e-16
c21798 2178 2342 1.58e-16
c21799 3531 3520 1.58e-16
c21800 721 1 4.03e-16
c21801 1800 692 1.75e-16
c21802 1706 812 4.46e-16
c21803 371 19 8.82e-16
c21804 2773 767 1.832e-15
c21805 3505 3117 4.97e-16
c21806 3589 762 1.58e-16
c21807 4548 3701 1.96e-16
c21808 2674 692 1.84e-16
c21809 612 1706 3.15e-16
c21810 602 1708 3.15e-16
c21811 573 580 3.54e-16
c21812 3502 672 2.4e-16
c21813 822 1956 1.58e-16
c21814 2702 737 1.75e-16
c21815 15 311 4.88e-16
c21816 1 305 1.9313e-14
c21817 2410 1 5.808e-15
c21818 2412 0 3.466e-15
c21819 595 2194 3.15e-16
c21820 602 2178 3.15e-16
c21821 762 25 1.58e-16
c21822 3662 812 1.84e-16
c21823 3918 3974 2.48e-16
c21824 5544 526 4.97e-16
c21825 777 1902 1.58e-16
c21826 2182 2342 1.58e-16
c21827 2799 2793 1.6e-16
c21828 378 360 1.58e-16
c21829 5407 5411 5.6e-16
c21830 5431 5409 9.18e-16
c21831 2545 2418 5.5e-16
c21832 2705 2712 1.96e-16
c21833 4267 3429 4.97e-16
c21834 601 1381 3.64e-16
c21835 1970 827 2.33e-16
c21836 3958 1 7.44e-16
c21837 762 1104 1.58e-16
c21838 3288 3289 1.6e-16
c21839 3279 3281 2.15e-16
c21840 3048 3173 3.92e-16
c21841 3644 3640 1.96e-16
c21842 4530 1 8.43e-16
c21843 602 2182 3.15e-16
c21844 747 1331 7.99e-16
c21845 19 535 3.84e-16
c21846 291 513 1.88e-16
c21847 470 441 3.75e-16
c21848 4582 3874 5.5e-16
c21849 1913 2393 1.58e-16
c21850 3270 2753 1.136e-15
c21851 3710 852 1.58e-16
c21852 894 1112 3.92e-16
c21853 909 1111 1.88e-16
c21854 883 1104 1.58e-16
c21855 981 984 1.58e-16
c21856 3397 3287 5.5e-16
c21857 4251 4263 2.32e-16
c21858 5262 5270 3.258e-15
c21859 3377 1 1.601e-15
c21860 1454 707 1.75e-16
c21861 1321 858 4.48e-16
c21862 617 3460 1.09e-16
c21863 3365 0 6.78e-16
c21864 3184 1 8.43e-16
c21865 1885 752 2.33e-16
c21866 4327 4706 1.58e-16
c21867 2822 827 1.339e-15
c21868 491 477 3.84e-16
c21869 3083 3472 2.386e-15
c21870 3481 3475 1.6e-16
c21871 3898 747 3.15e-16
c21872 5113 1 2.429e-15
c21873 3100 3455 1.58e-16
c21874 2327 1811 4.11e-16
c21875 4850 1 2.378e-15
c21876 3288 797 7.68e-16
c21877 1726 2239 4.97e-16
c21878 1087 732 1.58e-16
c21879 5262 5263 3.54e-16
c21880 5200 5205 3.84e-16
c21881 2194 1970 1.58e-16
c21882 105 104 6.67e-16
c21883 397 421 1.88e-16
c21884 4055 4054 1.58e-16
c21885 3876 852 3.15e-16
c21886 2903 2884 6.67e-16
c21887 1237 1238 1.96e-16
c21888 3909 37 1.88e-16
c21889 4343 4334 3.46e-16
c21890 5509 5511 1.609e-15
c21891 5417 5513 9.36e-16
c21892 2293 677 5.03e-16
c21893 1345 1576 1.58e-16
c21894 2594 3075 1.58e-16
c21895 1516 1888 1.58e-16
c21896 4847 4480 1.58e-16
c21897 1 340 1.607e-15
c21898 15 303 5.8e-16
c21899 3387 3083 5.5e-16
c21900 999 1006 2.27e-16
c21901 4048 4046 1.76e-16
c21902 2178 1777 5.88e-16
c21903 1046 692 3.15e-16
c21904 1203 894 3.54e-16
c21905 5514 5425 1.58e-16
c21906 5429 5426 4.41e-16
c21907 4725 5358 4.06e-16
c21908 146 218 1.88e-16
c21909 2683 2684 9.1e-16
c21910 659 26 2.65e-15
c21911 1539 767 2.33e-16
c21912 55 59 1.58e-16
c21913 3717 1 8.43e-16
c21914 2978 2969 3.92e-16
c21915 2282 692 1.58e-16
c21916 1038 1 1.56e-15
c21917 827 26 7.12e-16
c21918 3714 0 6.72e-16
c21919 3048 3138 5.42e-16
c21920 3024 3126 1.58e-16
c21921 4777 4780 6.67e-16
c21922 3409 3451 3.92e-16
c21923 3005 852 2.42e-16
c21924 632 2265 1.58e-16
c21925 5158 5220 6.67e-16
c21926 792 1121 1.813e-15
c21927 4861 265 1.88e-16
c21928 2391 1879 1.532e-15
c21929 2397 2396 5.65e-16
c21930 2182 1777 5.5e-16
c21931 5321 323 5.5e-16
c21932 2180 0 4.64e-16
c21933 4353 692 1.832e-15
c21934 1143 782 1.58e-16
c21935 4144 4142 1.76e-16
c21936 537 368 1.88e-16
c21937 2557 2752 3.92e-16
c21938 3773 1 1.021e-15
c21939 4403 4404 2.48e-16
c21940 2378 737 1.9e-16
c21941 1516 1071 1.136e-15
c21942 1615 1612 3.01e-16
c21943 1611 1608 6.44e-16
c21944 4696 4697 1.6e-16
c21945 4692 4310 1.443e-15
c21946 627 1331 7.99e-16
c21947 1690 0 3.63418e-13
c21948 1949 1 9.28e-16
c21949 5047 1 2.424e-15
c21950 2209 2206 5.5e-16
c21951 1080 707 6.48e-16
c21952 596 800 5.28e-16
c21953 4742 410 1.88e-16
c21954 602 3407 1.58e-16
c21955 3900 4268 1.58e-16
c21956 920 1205 3.92e-16
c21957 921 1204 2.54e-16
c21958 1999 842 7.68e-16
c21959 1992 827 1.9e-16
c21960 631 1 4.03e-16
c21961 3659 0 3.3633e-14
c21962 3073 2533 1.532e-15
c21963 3079 3078 5.65e-16
c21964 601 3900 3.15e-16
c21965 627 3898 3.15e-16
c21966 4291 1 6.15e-16
c21967 4395 3554 1.136e-15
c21968 1878 1482 1.96e-16
c21969 1873 1488 1.96e-16
c21970 4999 4978 5.92e-16
c21971 3347 3346 2.48e-16
c21972 3030 672 4.03e-16
c21973 3046 647 4.46e-16
c21974 1738 0 1.4092e-14
c21975 617 2616 1.58e-16
c21976 782 776 1.74e-16
c21977 1 440 4.92e-16
c21978 3393 767 3.15e-16
c21979 3710 3409 1.58e-16
c21980 4567 4728 1.58e-16
c21981 4571 4344 5.5e-16
c21982 4844 33 1.88e-16
c21983 1964 2487 4.36e-16
c21984 2485 2478 1.96e-16
c21985 3927 857 6.23e-16
c21986 4838 91 1.364e-15
c21987 2545 2339 1.58e-16
c21988 614 26 2.65e-15
c21989 3489 1 5.808e-15
c21990 910 3397 5.03e-16
c21991 3491 0 3.466e-15
c21992 4491 4489 2.15e-16
c21993 4499 4498 1.6e-16
c21994 2424 807 1.58e-16
c21995 2623 647 1.84e-16
c21996 2449 797 1.09e-16
c21997 1584 1579 1.642e-15
c21998 812 26 7.12e-16
c21999 2078 2049 1.37e-16
c22000 1635 2002 1.58e-16
c22001 100 117 1.138e-15
c22002 233 363 1.88e-16
c22003 612 26 1.58e-16
c22004 0 503 2.87e-16
c22005 5089 5064 5.87e-16
c22006 5066 5068 6.87e-16
c22007 2196 2240 1.58e-16
c22008 3910 3911 6.4e-16
c22009 1132 1133 7.46e-16
c22010 71 0 4.5712e-14
c22011 3900 3893 3.54e-16
c22012 2305 0 3.6368e-14
c22013 2166 2578 4.36e-16
c22014 2576 2569 1.96e-16
c22015 1427 1425 1.6e-16
c22016 1422 1421 2.03e-16
c22017 3882 4404 1.58e-16
c22018 3898 4416 1.58e-16
c22019 4484 4485 9.1e-16
c22020 82 81 1.58e-16
c22021 2535 2700 1.58e-16
c22022 2557 2688 1.58e-16
c22023 1007 0 1.0183e-14
c22024 657 1782 2.4e-16
c22025 3582 1 5.97e-15
c22026 3153 3152 1.6e-16
c22027 3145 3143 2.15e-16
c22028 4419 777 1.58e-16
c22029 3425 3423 1.6e-16
c22030 3420 3419 2.03e-16
c22031 2987 2955 1.58e-16
c22032 494 570 1.88e-16
c22033 5222 0 1.65e-16
c22034 1998 1607 1.136e-15
c22035 747 1706 3.15e-16
c22036 890 672 3.35e-16
c22037 907 647 4.8e-16
c22038 2549 2540 5.71e-16
c22039 4567 4877 3.92e-16
c22040 2673 0 3.466e-15
c22041 2542 2552 5.8e-16
c22042 596 755 5.28e-16
c22043 4007 4006 1.58e-16
c22044 3101 1 1.868e-15
c22045 1091 1094 6.13e-16
c22046 4736 5396 5.5e-16
c22047 2826 2822 1.96e-16
c22048 1684 852 3.15e-16
c22049 3890 0 8.1002e-14
c22050 1327 1504 1.96e-16
c22051 398 397 6.96e-16
c22052 4276 4643 1.58e-16
c22053 3138 3139 9.1e-16
c22054 1706 1403 1.58e-16
c22055 911 1331 3.45e-16
c22056 1357 0 3.466e-15
c22057 4572 4568 6.97e-16
c22058 4573 4566 1.71e-16
c22059 4561 4214 9.45e-16
c22060 3322 827 7.68e-16
c22061 4762 1 4.832e-15
c22062 1482 0 6.9481e-14
c22063 238 178 3.45e-16
c22064 612 2586 1.58e-16
c22065 5575 0 1.7164e-14
c22066 2457 2456 9.1e-16
c22067 2194 2388 1.58e-16
c22068 2178 2376 1.58e-16
c22069 2178 2171 1.58e-16
c22070 146 130 3.84e-16
c22071 3801 3806 1.291e-15
c22072 5464 5412 1.141e-15
c22073 5446 5449 3.54e-16
c22074 2509 2503 9.59e-16
c22075 920 797 3.69e-16
c22076 910 936 2.559e-15
c22077 3445 1 8.43e-16
c22078 911 3898 9.54e-16
c22079 910 3882 7.97e-16
c22080 1211 1345 3.92e-16
c22081 4208 0 2.2338e-14
c22082 2545 2854 4.63e-16
c22083 2423 782 7.38e-16
c22084 2172 702 3.15e-16
c22085 1752 1380 1.58e-16
c22086 3152 677 7.68e-16
c22087 3145 662 1.9e-16
c22088 2557 782 4.46e-16
c22089 2283 1 1.868e-15
c22090 2182 2376 1.58e-16
c22091 5447 439 5.5e-16
c22092 2273 0 2.93e-15
c22093 2182 2171 1.58e-16
c22094 986 672 1.58e-16
c22095 1434 647 4.81e-16
c22096 827 1187 1.58e-16
c22097 407 401 1.58e-16
c22098 4787 410 1.88e-16
c22099 2248 2635 1.532e-15
c22100 2640 2641 5.65e-16
c22101 543 535 2.218e-15
c22102 3029 3035 2.267e-15
c22103 642 1409 1.58e-16
c22104 4095 4086 1.96e-16
c22105 3415 0 1.23e-16
c22106 2196 692 3.15e-16
c22107 1750 1761 1.96e-16
c22108 2747 747 2.22e-16
c22109 953 0 1.9321e-14
c22110 3046 3031 1.632e-15
c22111 3030 3047 5.63e-16
c22112 4344 4724 1.96e-16
c22113 1708 1934 5.42e-16
c22114 1684 1922 1.58e-16
c22115 1694 1764 1.58e-16
c22116 2368 1851 1.96e-16
c22117 2369 2362 6.73e-16
c22118 2028 1 1.55e-16
c22119 2046 0 2.078e-15
c22120 2260 2261 5.65e-16
c22121 883 977 3.92e-16
c22122 890 976 1.88e-16
c22123 423 1 4.22e-16
c22124 227 233 1.58e-16
c22125 2810 2418 2.38e-15
c22126 3287 3659 1.58e-16
c22127 4685 33 1.88e-16
c22128 4072 4079 1.88e-16
c22129 3226 1 1.716e-15
c22130 2915 2913 5.66e-16
c22131 1771 647 5.03e-16
c22132 1274 1272 3.07e-16
c22133 4377 4370 1.96e-16
c22134 3531 4379 4.36e-16
c22135 2334 692 3.64e-16
c22136 3602 1 1.056e-15
c22137 1952 797 7.38e-16
c22138 1558 1116 2.48e-16
c22139 4628 4242 4.11e-16
c22140 4633 4624 3.46e-16
c22141 657 1794 2.22e-16
c22142 2508 842 1.58e-16
c22143 1437 1 4.41e-15
c22144 627 1706 3.15e-16
c22145 601 1708 3.15e-16
c22146 3322 812 3.64e-16
c22147 822 1976 1.58e-16
c22148 2787 3299 5.66e-16
c22149 2158 1635 1.96e-16
c22150 2156 2154 1.6e-16
c22151 1821 0 6.62e-16
c22152 1 30 8.8057e-14
c22153 24 22 7.1e-16
c22154 6 5 5.8e-16
c22155 9 49 5.8e-16
c22156 233 310 1.88e-16
c22157 3668 3657 1.96e-16
c22158 5165 5259 7.46e-16
c22159 2430 1 2.054e-15
c22160 1008 662 1.58e-16
c22161 642 3117 2.22e-16
c22162 2432 0 8e-16
c22163 601 2178 3.15e-16
c22164 3397 707 3.15e-16
c22165 3983 3976 1.88e-16
c22166 3041 1 7.228e-15
c22167 5378 1 3.36e-16
c22168 5514 5452 6.96e-16
c22169 3836 3840 1.202e-15
c22170 3032 0 4.64e-16
c22171 657 3397 7.99e-16
c22172 1556 807 5.73e-16
c22173 1331 1440 1.58e-16
c22174 3374 1 2.48e-16
c22175 4168 1 5.1e-16
c22176 3882 3684 5.88e-16
c22177 3876 3690 1.58e-16
c22178 4538 4539 1.6e-16
c22179 627 966 4e-16
c22180 617 1381 7.68e-16
c22181 4435 4811 3.92e-16
c22182 4548 1 1.106e-15
c22183 601 2182 3.15e-16
c22184 1 574 2.87e-16
c22185 310 305 1.88e-16
c22186 4582 4242 5.5e-16
c22187 2342 2349 1.96e-16
c22188 59 43 3.84e-16
c22189 3866 3858 7.29e-16
c22190 3856 3854 1.6e-16
c22191 4370 732 1.58e-16
c22192 4872 5104 2.037e-15
c22193 2712 2703 3.46e-16
c22194 1187 812 1.58e-16
c22195 921 918 3.84e-16
c22196 5324 5321 7.81e-16
c22197 1863 707 3.64e-16
c22198 2880 2893 1.96e-16
c22199 601 4251 1.832e-15
c22200 3281 3277 1.96e-16
c22201 4344 4706 1.58e-16
c22202 3192 3193 2.03e-16
c22203 2839 868 1.58e-16
c22204 1694 1505 1.58e-16
c22205 1468 1 1.056e-15
c22206 562 570 1.58e-16
c22207 4867 1 2.378e-15
c22208 5104 0 3.0503e-14
c22209 1089 737 1.58e-16
c22210 909 908 1.729e-15
c22211 5403 1 4.427e-15
c22212 2511 2510 1.6e-16
c22213 1576 782 1.832e-15
c22214 1374 1370 1.96e-16
c22215 3160 0 3.3874e-14
c22216 4349 4348 9.1e-16
c22217 2313 677 1.09e-16
c22218 667 1 5.62e-16
c22219 1203 1 1.704e-15
c22220 4322 1 2.054e-15
c22221 1516 1908 2.38e-15
c22222 1690 1689 3.15e-16
c22223 4324 0 8e-16
c22224 5038 5026 1.74e-16
c22225 4497 4847 2e-16
c22226 4864 4480 1.36e-15
c22227 4867 4873 1.6e-16
c22228 3411 3100 5.5e-16
c22229 2400 1 8.43e-16
c22230 1 546 2.87e-16
c22231 233 339 1.88e-16
c22232 4685 4680 1.536e-15
c22233 4776 4395 5.2e-16
c22234 4759 468 1.88e-16
c22235 2503 2498 1.642e-15
c22236 747 26 1.58e-16
c22237 3918 3935 8.1e-16
c22238 5450 0 4.0816e-14
c22239 3882 707 3.15e-16
c22240 2541 2373 1.58e-16
c22241 602 3409 4.46e-16
c22242 1533 782 1.58e-16
c22243 657 3882 4.03e-16
c22244 2518 2509 1.37e-16
c22245 2480 837 2.72e-16
c22246 3372 2849 1.96e-16
c22247 3369 3367 1.6e-16
c22248 910 1690 7.97e-16
c22249 911 1706 9.54e-16
c22250 3048 3143 1.58e-16
c22251 1786 0 3.3874e-14
c22252 1146 1 4.044e-15
c22253 4759 4761 4.93e-16
c22254 1594 0 6.62e-16
c22255 480 486 1.372e-15
c22256 302 320 1.58e-16
c22257 2189 1 7.228e-15
c22258 4793 178 5.8e-16
c22259 5133 5137 1.202e-15
c22260 2320 2321 9.1e-16
c22261 1147 797 6.38e-16
c22262 4241 4234 1.96e-16
c22263 3381 4243 4.36e-16
c22264 5270 149 7.16e-16
c22265 1647 842 1.58e-16
c22266 687 4319 1.58e-16
c22267 3876 4468 3.92e-16
c22268 702 0 2.86796e-13
c22269 4100 19 3.84e-16
c22270 1717 1719 2.03e-16
c22271 3169 3160 3.92e-16
c22272 2651 3163 5.66e-16
c22273 1590 1973 7.84e-16
c22274 1690 1833 1.96e-16
c22275 77 1 9.8e-16
c22276 5103 5074 1.58e-16
c22277 5127 5113 1.96e-16
c22278 3454 3455 2.48e-16
c22279 4458 792 1.58e-16
c22280 4470 0 1.6491e-14
c22281 332 342 8.86e-16
c22282 3557 717 1.58e-16
c22283 4969 4950 1.96e-16
c22284 792 1941 2.72e-16
c22285 5263 149 3.54e-16
c22286 2586 2593 1.96e-16
c22287 2558 1 2.471e-15
c22288 3310 3387 1.58e-16
c22289 4526 868 1.58e-16
c22290 5580 5579 9.13e-16
c22291 595 3021 1.58e-16
c22292 2804 0 3.5056e-14
c22293 2868 2867 1.6e-16
c22294 2860 2858 2.15e-16
c22295 3882 3452 1.58e-16
c22296 3124 0 1.6491e-14
c22297 1219 1220 7.51e-16
c22298 2541 2534 1.58e-16
c22299 2559 2554 1.58e-16
c22300 1801 1420 3.92e-16
c22301 839 0 7.709e-15
c22302 3160 3162 2.15e-16
c22303 3679 0 1.4092e-14
c22304 981 0 3.7577e-14
c22305 617 3900 3.15e-16
c22306 1667 1669 3.2e-16
c22307 595 911 1.58e-16
c22308 176 180 6.38e-16
c22309 164 163 2.84e-16
c22310 3030 3308 1.58e-16
c22311 3275 767 1.58e-16
c22312 3048 662 3.15e-16
c22313 2206 2213 1.96e-16
c22314 3397 3022 5.5e-16
c22315 2077 2078 2.123e-15
c22316 982 983 7.46e-16
c22317 4623 4242 5.2e-16
c22318 5562 497 3.54e-16
c22319 3886 677 3.15e-16
c22320 5478 5479 3.54e-16
c22321 4827 149 1.88e-16
c22322 3125 0 2.93e-15
c22323 2929 1 5.966e-15
c22324 1220 852 1.85e-16
c22325 1986 827 7.38e-16
c22326 919 1055 3.92e-16
c22327 922 1054 2.54e-16
c22328 3657 0 1.6491e-14
c22329 687 1420 5.73e-16
c22330 1523 1534 1.96e-16
c22331 1331 957 5.5e-16
c22332 1318 1316 3.54e-16
c22333 4078 1 6.76e-16
c22334 3024 2764 5.5e-16
c22335 4811 0 1.6462e-14
c22336 3393 3401 8.73e-16
c22337 2535 837 3.15e-16
c22338 1652 2020 1.96e-16
c22339 627 26 1.58e-16
c22340 339 340 6.96e-16
c22341 3521 3532 1.96e-16
c22342 5165 1 4.669e-15
c22343 2158 1 1.106e-15
c22344 2559 2350 5.5e-16
c22345 2170 2531 1.58e-16
c22346 3898 4421 1.58e-16
c22347 3876 4433 1.58e-16
c22348 1795 1786 3.92e-16
c22349 1403 1789 5.66e-16
c22350 2559 2717 5.42e-16
c22351 2535 2705 1.58e-16
c22352 3866 1 1.601e-15
c22353 4056 37 5.71e-16
c22354 3565 4383 1.96e-16
c22355 3373 0 2.7489e-14
c22356 4449 1 1.056e-15
c22357 4682 4679 3.01e-16
c22358 1690 1798 1.58e-16
c22359 1545 0 1.4092e-14
c22360 207 205 6.01e-16
c22361 2379 2376 5.5e-16
c22362 3521 702 1.58e-16
c22363 4982 4980 1.001e-15
c22364 4905 4930 1.96e-16
c22365 3030 797 3.15e-16
c22366 909 662 3.15e-16
c22367 4571 1 3.55e-15
c22368 4567 4894 3.92e-16
c22369 4770 468 1.88e-16
c22370 2866 3376 3.38e-16
c22371 2693 0 8e-16
c22372 2136 2106 6.53e-16
c22373 3673 3674 1.35e-16
c22374 4124 4126 2.254e-15
c22375 4623 497 1.88e-16
c22376 3266 0 6.72e-16
c22377 1324 1330 5.8e-16
c22378 5564 5422 2.12e-16
c22379 2764 762 2.22e-16
c22380 3869 0 2.0654e-14
c22381 2651 2645 1.418e-15
c22382 1343 1521 3.92e-16
c22383 4293 4643 2e-16
c22384 4276 4660 1.36e-15
c22385 4669 4663 1.6e-16
c22386 3062 3060 1.6e-16
c22387 3057 3056 2.03e-16
c22388 3225 3226 1.35e-16
c22389 1850 1465 1.96e-16
c22390 4549 3751 1.96e-16
c22391 2815 827 3.15e-16
c22392 4779 1 4.832e-15
c22393 1 465 4.22e-16
c22394 4580 4480 5.5e-16
c22395 4582 4486 1.58e-16
c22396 5278 5288 9.99e-16
c22397 627 2586 1.58e-16
c22398 456 0 1.0822e-14
c22399 5262 236 1.58e-16
c22400 4844 526 1.88e-16
c22401 2458 2452 1.418e-15
c22402 2441 2469 2.64e-16
c22403 2463 2459 1.96e-16
c22404 2194 1678 1.58e-16
c22405 4759 64 1.88e-16
c22406 1986 812 1.58e-16
c22407 1690 707 3.15e-16
c22408 1901 737 1.58e-16
c22409 1454 1837 7.84e-16
c22410 3392 3404 3.225e-15
c22411 2679 2288 1.136e-15
c22412 657 1690 4.03e-16
c22413 602 922 3.15e-16
c22414 595 919 4.37e-16
c22415 1693 0 1.5577e-14
c22416 822 25 1.58e-16
c22417 9 194 5.8e-16
c22418 3836 3841 9.94e-16
c22419 890 797 3.15e-16
c22420 907 1157 3.92e-16
c22421 2839 0 1.6491e-14
c22422 920 978 1.58e-16
c22423 3719 3710 3.92e-16
c22424 4223 3918 2.87e-16
c22425 3421 0 3.3643e-14
c22426 2545 2853 1.58e-16
c22427 3751 3734 1.541e-15
c22428 3323 3322 1.6e-16
c22429 1674 1206 1.96e-16
c22430 3139 662 7.38e-16
c22431 1708 1939 1.58e-16
c22432 642 1769 1.58e-16
c22433 632 1755 1.84e-16
c22434 3304 2787 1.136e-15
c22435 1938 1550 4.97e-16
c22436 1694 1769 1.58e-16
c22437 5058 5048 3.92e-16
c22438 612 1678 1.58e-16
c22439 3034 767 3.15e-16
c22440 2661 1 8.43e-16
c22441 883 991 1.88e-16
c22442 907 984 1.58e-16
c22443 877 878 3.62e-16
c22444 245 15 5.8e-16
c22445 284 19 8.82e-16
c22446 268 0 1.4515e-14
c22447 3287 3679 2.38e-15
c22448 5536 1 8.631e-15
c22449 657 3491 2.72e-16
c22450 1791 647 1.09e-16
c22451 1593 807 1.58e-16
c22452 1343 752 4.46e-16
c22453 1416 1415 1.6e-16
c22454 1408 1406 2.15e-16
c22455 2806 2808 2.03e-16
c22456 1828 692 3.15e-16
c22457 1465 1460 1.642e-15
c22458 1239 1 7.976e-15
c22459 1922 1934 2.32e-16
c22460 2305 707 1.75e-16
c22461 2815 812 3.15e-16
c22462 1846 1 1.868e-15
c22463 617 1708 3.15e-16
c22464 1836 0 2.93e-15
c22465 3239 737 4.81e-16
c22466 3387 3535 1.58e-16
c22467 2452 1 5.97e-15
c22468 837 844 1.6e-16
c22469 2448 0 6.72e-16
c22470 617 2178 3.15e-16
c22471 792 1913 1.813e-15
c22472 1930 777 2.22e-16
c22473 1511 722 1.58e-16
c22474 129 1 5.175e-15
c22475 160 13 1.88e-16
c22476 657 1007 2.68e-16
c22477 155 0 2.87e-16
c22478 2722 2724 2.15e-16
c22479 919 1113 1.58e-16
c22480 1694 677 3.15e-16
c22481 1490 1492 2.03e-16
c22482 3701 3898 5.5e-16
c22483 3707 3900 1.58e-16
c22484 4540 4552 3.13e-16
c22485 2753 2754 1.35e-16
c22486 1981 868 1.813e-15
c22487 687 2652 1.58e-16
c22488 2014 2005 3.46e-16
c22489 0 300 2.87e-16
c22490 3202 3570 1.96e-16
c22491 4582 4259 5.5e-16
c22492 5180 5162 6.67e-16
c22493 4674 439 1.88e-16
c22494 617 2182 3.15e-16
c22495 3976 3974 3.54e-16
c22496 5388 5326 6.96e-16
c22497 909 1098 3.54e-16
c22498 4271 4268 5.5e-16
c22499 238 239 3.84e-16
c22500 4606 1 7.849e-15
c22501 1482 707 3.15e-16
c22502 1472 1474 1.862e-15
c22503 1031 1041 1.418e-15
c22504 542 204 1.88e-16
c22505 3616 3588 2.64e-16
c22506 3972 1 2.259e-15
c22507 617 4251 1.58e-16
c22508 1740 1737 3.01e-16
c22509 1736 1733 6.44e-16
c22510 4815 4811 1.96e-16
c22511 2696 3190 1.96e-16
c22512 1618 2003 1.96e-16
c22513 601 1740 1.09e-16
c22514 1484 1 9.28e-16
c22515 4526 0 1.4092e-14
c22516 809 810 1.6e-16
c22517 204 188 3.84e-16
c22518 2349 2340 3.46e-16
c22519 14 1 1.607e-15
c22520 107 450 1.88e-16
c22521 3393 3688 1.58e-16
c22522 1083 1097 1.96e-16
c22523 2603 0 3.3717e-14
c22524 5229 5256 9.6e-16
c22525 4685 526 1.88e-16
c22526 2172 1981 5.5e-16
c22527 966 957 1.418e-15
c22528 3180 0 1.4092e-14
c22529 4355 4351 1.96e-16
c22530 4770 64 1.88e-16
c22531 2545 2616 4.63e-16
c22532 1321 1146 1.58e-16
c22533 1327 1136 5.88e-16
c22534 3393 3123 1.58e-16
c22535 4472 822 1.58e-16
c22536 4340 0 6.72e-16
c22537 4864 4497 1.58e-16
c22538 4871 1 8.43e-16
c22539 3046 3360 3.92e-16
c22540 3292 807 2.4e-16
c22541 797 813 1.621e-15
c22542 807 811 2.19e-16
c22543 9 507 6.48e-16
c22544 281 204 1.88e-16
c22545 5229 5231 5.25e-16
c22546 294 292 6.01e-16
c22547 4008 857 3.1e-16
c22548 3537 3538 1.35e-16
c22549 5484 5527 1.617e-15
c22550 921 1100 1.96e-16
c22551 601 3409 4.46e-16
c22552 1950 782 4.81e-16
c22553 1091 1545 2.38e-15
c22554 1327 1016 5.88e-16
c22555 3151 0 6.9481e-14
c22556 4599 4592 1.96e-16
c22557 3870 4601 1.914e-15
c22558 3701 4518 1.58e-16
c22559 2518 2521 1.138e-15
c22560 595 957 4.21e-16
c22561 1619 1 1.868e-15
c22562 4794 4797 6.67e-16
c22563 2104 2098 2.08e-16
c22564 4776 4783 1.81e-16
c22565 5227 5231 5.6e-16
c22566 1609 0 2.93e-15
c22567 520 522 7.1e-16
c22568 3185 3552 1.58e-16
c22569 3174 3560 5.66e-16
c22570 3566 3557 3.92e-16
c22571 4725 352 1.88e-16
c22572 5051 120 1.58e-16
c22573 3385 3381 1.58e-16
c22574 5296 5300 2.95e-16
c22575 4776 5207 6.9e-16
c22576 1084 1085 7.51e-16
c22577 52 53 1.58e-16
c22578 55 42 1.58e-16
c22579 2992 2982 1.98e-16
c22580 1833 702 2.4e-16
c22581 1642 852 1.58e-16
c22582 687 4339 1.58e-16
c22583 3900 4485 3.92e-16
c22584 4514 5588 4.69e-16
c22585 602 4236 1.9e-16
c22586 3261 3263 2.03e-16
c22587 2662 3160 1.58e-16
c22588 1601 1985 1.58e-16
c22589 1706 1850 3.92e-16
c22590 545 535 8.86e-16
c22591 1963 1 8.43e-16
c22592 5032 1 1.0083e-14
c22593 4949 4941 1.612e-15
c22594 3046 868 3.15e-16
c22595 3024 827 4.48e-16
c22596 3387 3236 5.5e-16
c22597 1072 1053 1.546e-15
c22598 2567 0 1.6491e-14
c22599 1116 1117 8.58e-16
c22600 4634 5412 2.675e-15
c22601 2559 2169 1.58e-16
c22602 2557 2166 1.58e-16
c22603 2545 2581 1.58e-16
c22604 922 1220 3.92e-16
c22605 1161 1610 7.84e-16
c22606 1690 1832 1.58e-16
c22607 1890 1499 4.11e-16
c22608 3046 3325 1.58e-16
c22609 3030 3313 1.58e-16
c22610 4855 439 1.88e-16
c22611 2196 2457 3.92e-16
c22612 3958 857 1.88e-16
c22613 3930 3928 7.1e-16
c22614 3605 767 2.33e-16
c22615 5511 381 5.5e-16
c22616 2777 2775 1.6e-16
c22617 2772 2771 2.03e-16
c22618 1238 858 3.15e-16
c22619 2003 868 2.4e-16
c22620 3873 911 1.88e-16
c22621 4504 4515 1.96e-16
c22622 2254 647 2.33e-16
c22623 1805 1414 4.11e-16
c22624 1798 1786 2.32e-16
c22625 2849 3343 1.96e-16
c22626 3048 2781 5.5e-16
c22627 2213 2204 3.46e-16
c22628 4828 0 1.6462e-14
c22629 2662 702 1.813e-15
c22630 1 450 4.2258e-14
c22631 15 419 5.8e-16
c22632 5039 5064 3.54e-16
c22633 2178 1743 5.88e-16
c22634 692 685 5.58e-16
c22635 3781 3868 1.6e-16
c22636 907 868 3.15e-16
c22637 883 827 6.45e-16
c22638 921 692 3.15e-16
c22639 957 960 2.03e-16
c22640 4338 692 5.03e-16
c22641 5396 5262 1.389e-15
c22642 542 175 1.88e-16
c22643 3684 3679 1.642e-15
c22644 3015 2929 4.06e-16
c22645 1447 1001 1.96e-16
c22646 1181 1158 6.54e-16
c22647 632 920 3.69e-16
c22648 3876 4438 1.58e-16
c22649 3900 4450 5.42e-16
c22650 2559 2722 1.58e-16
c22651 1689 1693 5.8e-16
c22652 2541 677 3.15e-16
c22653 2545 662 3.15e-16
c22654 1954 1567 1.532e-15
c22655 1960 1959 5.65e-16
c22656 2182 1743 5.5e-16
c22657 764 765 1.6e-16
c22658 3157 692 2.33e-16
c22659 4969 4531 7.01e-16
c22660 3024 812 4.48e-16
c22661 94 30 6.83e-16
c22662 88 37 1.88e-16
c22663 2709 0 6.72e-16
c22664 2581 2582 9.1e-16
c22665 1814 662 4.81e-16
c22666 1432 1423 3.92e-16
c22667 996 1426 5.66e-16
c22668 3119 1 9.28e-16
c22669 612 3024 3.15e-16
c22670 2194 762 3.15e-16
c22671 4508 827 1.9e-16
c22672 4515 842 7.68e-16
c22673 1845 732 1.813e-15
c22674 808 1 1.65e-16
c22675 657 1786 1.58e-16
c22676 3642 1 5.808e-15
c22677 911 1687 1.58e-16
c22678 4293 4660 1.58e-16
c22679 3242 792 5.73e-16
c22680 1369 0 3.6368e-14
c22681 263 265 6.01e-16
c22682 3430 3421 3.92e-16
c22683 3021 3424 5.66e-16
c22684 2832 868 1.813e-15
c22685 2186 2177 5.71e-16
c22686 4796 1 4.832e-15
c22687 1721 1 2.054e-15
c22688 4580 4497 5.5e-16
c22689 4582 4503 1.58e-16
c22690 707 702 2.77e-16
c22691 627 2606 1.58e-16
c22692 1981 0 6.9481e-14
c22693 281 175 1.88e-16
c22694 4725 294 5.8e-16
c22695 4804 352 1.88e-16
c22696 4674 5482 3.65e-16
c22697 2172 1682 5.5e-16
c22698 4423 752 1.9e-16
c22699 4770 5221 1.96e-16
c22700 2557 2503 3.92e-16
c22701 2518 2515 8.32e-16
c22702 921 1158 1.58e-16
c22703 4301 4302 2.48e-16
c22704 1343 1520 1.58e-16
c22705 1327 1508 1.58e-16
c22706 4214 3879 7.67e-16
c22707 1513 1510 3.01e-16
c22708 1509 1506 6.44e-16
c22709 2714 722 7.68e-16
c22710 1465 1849 1.58e-16
c22711 601 922 5.14e-16
c22712 4053 1 7.71e-16
c22713 4217 25 3.84e-16
c22714 4232 0 1.6491e-14
c22715 3330 3339 3.92e-16
c22716 3333 2821 5.66e-16
c22717 2832 3325 1.58e-16
c22718 1724 1 6.15e-16
c22719 3239 3237 1.6e-16
c22720 2045 2054 3.92e-16
c22721 1 337 3.6e-16
c22722 421 262 1.88e-16
c22723 3695 827 1.9e-16
c22724 5158 5171 1.96e-16
c22725 3370 2849 9.7e-16
c22726 2319 1 1.056e-15
c22727 3511 3508 3.01e-16
c22728 747 2357 1.58e-16
c22729 129 131 1.88e-16
c22730 3693 3393 1.58e-16
c22731 3705 3387 1.58e-16
c22732 1194 868 1.58e-16
c22733 883 812 6.45e-16
c22734 909 1172 4.35e-16
c22735 907 1171 1.88e-16
c22736 890 1164 1.58e-16
c22737 2288 1 4.41e-15
c22738 1113 1114 1.21e-16
c22739 2654 2282 1.58e-16
c22740 657 981 5.73e-16
c22741 3441 0 1.4092e-14
c22742 3254 1 1.868e-15
c22743 2545 2858 1.58e-16
c22744 612 883 3.15e-16
c22745 595 894 6.61e-16
c22746 2427 782 1.832e-15
c22747 1776 1380 1.96e-16
c22748 1771 1386 1.96e-16
c22749 3030 3070 1.58e-16
c22750 2026 2028 1.082e-15
c22751 2069 1 1.23e-16
c22752 3525 677 1.9e-16
c22753 890 978 3.54e-16
c22754 909 999 1.58e-16
c22755 3469 662 1.75e-16
c22756 3728 3736 3.54e-16
c22757 3784 3783 2.12e-16
c22758 1783 662 2.33e-16
c22759 1270 1300 2.93e-16
c22760 1331 1657 4.63e-16
c22761 763 1 1.65e-16
c22762 3410 3027 3.54e-16
c22763 3232 3230 1.6e-16
c22764 3227 3226 2.03e-16
c22765 3606 1 1.716e-15
c22766 1575 1121 4.97e-16
c22767 1347 1 2.86e-16
c22768 4645 4259 4.11e-16
c22769 4650 4641 3.46e-16
c22770 2799 782 3.64e-16
c22771 687 1794 1.813e-15
c22772 1326 0 4.3801e-14
c22773 3548 0 6.9481e-14
c22774 5007 1 6.03e-16
c22775 3390 3388 1.578e-15
c22776 3396 3403 7.06e-16
c22777 1465 1 5.97e-15
c22778 3387 3540 1.58e-16
c22779 3411 3552 5.42e-16
c22780 3393 3157 1.58e-16
c22781 3293 3678 1.96e-16
c22782 3287 3683 1.96e-16
c22783 279 291 1.58e-16
c22784 1 137 1.607e-15
c22785 410 30 3.84e-16
c22786 390 37 1.88e-16
c22787 426 27 1.88e-16
c22788 657 3485 2.4e-16
c22789 4087 4088 6.4e-16
c22790 2443 2445 2.03e-16
c22791 2265 1749 1.136e-15
c22792 4861 381 1.88e-16
c22793 687 3397 7.99e-16
c22794 1956 797 1.832e-15
c22795 1559 1571 2.32e-16
c22796 2498 858 1.84e-16
c22797 1818 1431 1.532e-15
c22798 1824 1823 5.65e-16
c22799 1331 1 4.57e-15
c22800 777 1117 1.58e-16
c22801 4452 4828 3.92e-16
c22802 4839 4840 1.6e-16
c22803 2151 2161 3.13e-16
c22804 1641 1708 1.58e-16
c22805 1635 1706 5.5e-16
c22806 81 71 8.86e-16
c22807 1659 0 1.7608e-14
c22808 41 43 2.84e-16
c22809 0 5 4.4191e-14
c22810 136 508 1.88e-16
c22811 3393 717 4.03e-16
c22812 4582 4276 5.5e-16
c22813 5397 1 3.36e-16
c22814 2425 2427 1.862e-15
c22815 1913 1919 1.418e-15
c22816 1930 1902 2.64e-16
c22817 3361 3809 4.06e-16
c22818 5366 0 2.9101e-14
c22819 2813 1 6.15e-16
c22820 894 1113 3.54e-16
c22821 996 997 8.58e-16
c22822 2724 2720 1.96e-16
c22823 5376 5353 2.12e-16
c22824 5360 5357 2.004e-15
c22825 2248 2616 1.96e-16
c22826 4175 4177 1.06e-16
c22827 3744 3748 3.01e-16
c22828 3046 0 3.5222e-13
c22829 617 4271 1.58e-16
c22830 3781 0 6.0757e-14
c22831 1651 1642 3.46e-16
c22832 3898 1 4.77e-16
c22833 3718 4552 3.38e-16
c22834 4709 4711 1.687e-15
c22835 4721 4714 6.73e-16
c22836 4720 4333 1.96e-16
c22837 627 1754 2.72e-16
c22838 1497 1 6.15e-16
c22839 4543 0 1.3715e-14
c22840 747 1527 2.72e-16
c22841 0 587 2.87e-16
c22842 19 576 3.45e-16
c22843 5185 1 3.36e-16
c22844 48 49 3.84e-16
c22845 42 43 5.8e-16
c22846 5025 122 3.54e-16
c22847 2011 0 6.72e-16
c22848 222 1 9.8e-16
c22849 4287 647 5.03e-16
c22850 1103 752 1.58e-16
c22851 4167 4166 1.58e-16
c22852 2623 0 1.4092e-14
c22853 3711 3709 2.03e-16
c22854 5403 410 3.54e-16
c22855 4804 294 1.88e-16
c22856 2041 2043 1.062e-15
c22857 1131 797 1.75e-16
c22858 4702 5388 1.58e-16
c22859 1218 919 1.58e-16
c22860 718 1 1.65e-16
c22861 3959 37 1.88e-16
c22862 1181 1640 1.96e-16
c22863 1345 1161 1.58e-16
c22864 1343 1151 5.5e-16
c22865 1331 1622 1.58e-16
c22866 3107 3109 1.862e-15
c22867 2594 2600 1.418e-15
c22868 2611 2583 2.64e-16
c22869 3501 3134 1.58e-16
c22870 3489 3488 2.48e-16
c22871 4492 822 1.58e-16
c22872 2778 767 1.09e-16
c22873 1533 1522 1.58e-16
c22874 5010 4920 1.58e-16
c22875 562 580 1.58e-16
c22876 3106 647 2.33e-16
c22877 4888 1 8.43e-16
c22878 4881 4497 1.365e-15
c22879 2601 0 1.6491e-14
c22880 4810 4435 4.9e-16
c22881 2178 2321 1.96e-16
c22882 1061 1038 6.54e-16
c22883 2995 0 1.5926e-14
c22884 617 3409 4.46e-16
c22885 2559 2390 1.58e-16
c22886 687 3882 4.03e-16
c22887 3109 3108 2.48e-16
c22888 601 971 3.57e-16
c22889 3684 4526 2.38e-15
c22890 2476 842 1.339e-15
c22891 907 0 3.45479e-13
c22892 3024 2651 1.58e-16
c22893 1166 1 5.821e-15
c22894 4793 4801 1.81e-16
c22895 0 559 2.87e-16
c22896 30 556 3.84e-16
c22897 37 548 1.88e-16
c22898 3185 3557 1.58e-16
c22899 3655 797 7.38e-16
c22900 4580 4605 3.92e-16
c22901 2396 0 1.4092e-14
c22902 2182 2321 4.63e-16
c22903 895 893 3.54e-16
c22904 1682 0 6.9718e-14
c22905 5300 0 2.8602e-14
c22906 78 305 1.88e-16
c22907 146 334 1.88e-16
c22908 3321 852 1.58e-16
c22909 4253 4251 2.15e-16
c22910 4261 4260 1.6e-16
c22911 2612 2603 3.92e-16
c22912 2220 2606 5.66e-16
c22913 2231 2598 1.58e-16
c22914 542 436 1.88e-16
c22915 3363 1 4.03e-16
c22916 1206 858 3.69e-16
c22917 1456 1026 2.48e-16
c22918 3932 1 4.64e-16
c22919 601 4236 5.03e-16
c22920 3024 747 3.15e-16
c22921 1718 1318 7.84e-16
c22922 870 1 7.18e-16
c22923 2662 3180 2.38e-15
c22924 1999 1993 1.6e-16
c22925 1601 1990 2.386e-15
c22926 1684 1867 3.92e-16
c22927 479 476 1.099e-15
c22928 308 320 1.58e-16
c22929 900 893 6.67e-16
c22930 2210 0 6.72e-16
c22931 485 494 1.58e-16
c22932 3174 732 5.73e-16
c22933 3048 852 3.58e-16
c22934 3411 3253 5.5e-16
c22935 5321 5332 9.85e-16
c22936 2786 2401 1.96e-16
c22937 1092 722 4.98e-16
c22938 601 3055 2.33e-16
c22939 595 3066 2.22e-16
c22940 2832 0 6.9481e-14
c22941 1561 782 5.03e-16
c22942 1121 1118 1.984e-15
c22943 3886 4314 1.58e-16
c22944 3898 3463 5.5e-16
c22945 3900 3469 1.58e-16
c22946 3707 852 1.58e-16
c22947 4668 381 7.84e-16
c22948 2894 2893 1.6e-16
c22949 1729 1727 1.6e-16
c22950 4335 4337 2.03e-16
c22951 2277 662 1.84e-16
c22952 2005 858 1.339e-15
c22953 1166 1622 1.58e-16
c22954 822 826 2.19e-16
c22955 1706 1849 1.58e-16
c22956 1690 1837 1.58e-16
c22957 85 26 1.03e-15
c22958 82 19 3.2e-16
c22959 4967 4946 5.14e-16
c22960 3083 3451 1.96e-16
c22961 3024 3342 1.58e-16
c22962 3046 3330 1.58e-16
c22963 2232 2233 1.6e-16
c22964 2223 2225 2.15e-16
c22965 675 674 1.6e-16
c22966 9 333 6.48e-16
c22967 3757 3732 7.65e-16
c22968 4168 857 3.1e-16
c22969 4657 4282 4.9e-16
c22970 632 3030 3.15e-16
c22971 1327 662 3.15e-16
c22972 2194 2269 1.58e-16
c22973 2178 2257 1.58e-16
c22974 2214 1681 1.136e-15
c22975 3599 782 1.58e-16
c22976 3321 3293 2.64e-16
c22977 4317 4319 1.862e-15
c22978 3515 1 1.868e-15
c22979 3090 3091 2.03e-16
c22980 2921 2977 9.34e-16
c22981 1194 0 2.7246e-14
c22982 2248 662 1.58e-16
c22983 747 883 3.15e-16
c22984 4845 0 1.6462e-14
c22985 2736 3245 7.84e-16
c22986 3180 707 1.84e-16
c22987 1771 0 3.466e-15
c22988 3393 3450 1.58e-16
c22989 632 2620 1.832e-15
c22990 5190 5197 8.94e-16
c22991 5192 5195 1.342e-15
c22992 2196 2456 5.42e-16
c22993 3542 3157 1.96e-16
c22994 3547 3151 1.96e-16
c22995 762 2384 3.79e-16
c22996 2182 2257 1.58e-16
c22997 5481 5491 2.114e-15
c22998 909 852 3.15e-16
c22999 5044 0 2.1607e-14
c23000 1160 782 1.58e-16
c23001 64 323 1.88e-16
c23002 4358 692 1.09e-16
c23003 1343 952 1.58e-16
c23004 542 349 1.88e-16
c23005 1459 1016 4.11e-16
c23006 3718 3754 2.31e-16
c23007 3046 3122 3.92e-16
c23008 1828 1823 1.642e-15
c23009 1116 0 3.7288e-14
c23010 4453 1 1.716e-15
c23011 4699 4696 3.01e-16
c23012 1706 1 4.77e-16
c23013 692 684 1.74e-16
c23014 325 321 6.38e-16
c23015 320 334 1.88e-16
c23016 310 450 1.88e-16
c23017 565 204 1.88e-16
c23018 3151 707 1.58e-16
c23019 5262 178 1.58e-16
c23020 5230 0 3.0503e-14
c23021 4944 4950 4.48e-16
c23022 3347 852 1.58e-16
c23023 2291 2289 1.862e-15
c23024 2154 0 1.3715e-14
c23025 1794 1766 2.64e-16
c23026 642 2559 3.58e-16
c23027 890 1052 1.96e-16
c23028 4571 4531 3.92e-16
c23029 632 890 3.15e-16
c23030 3297 0 6.62e-16
c23031 627 3024 3.15e-16
c23032 2172 777 3.15e-16
c23033 1106 1105 3.94e-16
c23034 3565 4387 1.58e-16
c23035 2350 752 1.58e-16
c23036 2628 2237 1.136e-15
c23037 2362 737 1.84e-16
c23038 672 25 1.58e-16
c23039 3662 1 2.054e-15
c23040 3853 0 1.7608e-14
c23041 1591 1136 1.532e-15
c23042 1597 1596 5.65e-16
c23043 966 1 4.044e-15
c23044 792 798 1.097e-15
c23045 3522 3524 2.03e-16
c23046 4310 4660 2e-16
c23047 4293 4677 1.36e-15
c23048 4686 4680 1.6e-16
c23049 2816 807 2.65e-16
c23050 3651 792 2.65e-16
c23051 1390 0 6.62e-16
c23052 4905 4960 1.139e-15
c23053 3022 3421 1.58e-16
c23054 642 1732 5.73e-16
c23055 3034 2770 1.58e-16
c23056 3409 3603 1.58e-16
c23057 4813 1 4.832e-15
c23058 1059 717 1.58e-16
c23059 858 867 1.74e-16
c23060 3606 3225 3.92e-16
c23061 4810 0 3.07588e-13
c23062 5136 5135 5.5e-16
c23063 2654 2271 7.84e-16
c23064 3321 3409 5.5e-16
c23065 4502 827 7.38e-16
c23066 5578 5576 1.6e-16
c23067 2907 1 7.51e-16
c23068 2756 2765 3.92e-16
c23069 3640 1 1.716e-15
c23070 1321 1537 1.58e-16
c23071 1343 1525 1.58e-16
c23072 537 136 1.88e-16
c23073 3067 3058 3.92e-16
c23074 2532 3061 5.66e-16
c23075 2333 722 3.15e-16
c23076 2724 732 2.72e-16
c23077 1863 1857 1.6e-16
c23078 1465 1854 2.386e-15
c23079 1482 1837 1.58e-16
c23080 687 1690 4.03e-16
c23081 617 922 5.14e-16
c23082 4490 4487 6.44e-16
c23083 4494 4491 3.01e-16
c23084 3330 2832 1.58e-16
c23085 2194 722 4.46e-16
c23086 792 797 2.77e-16
c23087 3243 767 1.339e-15
c23088 595 1 4.0331e-14
c23089 2031 2030 4.61e-16
c23090 1 499 5.698e-15
c23091 245 247 1.88e-16
c23092 3225 3607 2.48e-16
c23093 1947 822 1.813e-15
c23094 2335 1 9.28e-16
c23095 0 500 1.4515e-14
c23096 3497 3106 1.136e-15
c23097 3236 752 3.15e-16
c23098 3818 3819 1.6e-16
c23099 3916 3915 7.81e-16
c23100 5234 238 1.345e-15
c23101 1011 677 1.75e-16
c23102 1188 827 1.58e-16
c23103 894 1187 3.92e-16
c23104 909 1186 1.88e-16
c23105 883 1179 1.58e-16
c23106 103 9 4.88e-16
c23107 397 204 1.88e-16
c23108 4417 752 7.38e-16
c23109 4708 5286 2.45e-16
c23110 2766 2765 1.6e-16
c23111 922 1008 1.58e-16
c23112 4332 677 7.38e-16
c23113 2674 2282 2.38e-15
c23114 1891 752 1.84e-16
c23115 1331 1317 1.58e-16
c23116 600 19 1.96e-16
c23117 632 986 3.15e-16
c23118 2747 1 5.97e-15
c23119 627 883 3.15e-16
c23120 3886 3565 5.5e-16
c23121 3328 3339 1.96e-16
c23122 3046 3087 1.58e-16
c23123 3030 3075 1.58e-16
c23124 1684 1573 1.58e-16
c23125 1690 1567 5.88e-16
c23126 762 1551 2.65e-16
c23127 0 180 5.738e-14
c23128 339 450 1.88e-16
c23129 5034 5033 5.25e-16
c23130 2196 2219 3.92e-16
c23131 4954 1 5.28e-16
c23132 1126 1127 1.238e-15
c23133 883 993 3.54e-16
c23134 894 1014 1.58e-16
c23135 2557 2667 3.92e-16
c23136 1641 852 1.58e-16
c23137 1331 1321 4.116e-15
c23138 1661 1327 3.16e-16
c23139 3903 0 1.23e-16
c23140 1942 1939 5.5e-16
c23141 3519 677 7.38e-16
c23142 3390 3394 2.074e-15
c23143 1882 1 1.056e-15
c23144 5387 5385 1.167e-15
c23145 3411 3557 1.58e-16
c23146 3397 3570 4.63e-16
c23147 1970 1 4.41e-15
c23148 2178 1783 1.58e-16
c23149 842 835 5.58e-16
c23150 3344 852 1.58e-16
c23151 5586 1 1.23e-16
c23152 2538 2544 5.8e-16
c23153 5429 0 1.94e-14
c23154 2479 0 6.62e-16
c23155 3565 3560 1.642e-15
c23156 4502 812 1.58e-16
c23157 910 3046 1.014e-15
c23158 911 3024 1.88e-16
c23159 2818 2816 1.6e-16
c23160 1086 737 2.33e-16
c23161 3463 4281 1.96e-16
c23162 4216 1 7.71e-16
c23163 2515 858 1.58e-16
c23164 1113 1 1.56e-15
c23165 3677 3674 6.44e-16
c23166 3681 3678 3.01e-16
c23167 687 2673 2.72e-16
c23168 2182 1783 1.58e-16
c23169 4582 4293 5.5e-16
c23170 4844 207 1.88e-16
c23171 737 753 1.621e-15
c23172 3785 3783 7.3e-16
c23173 2822 1 1.716e-15
c23174 1001 672 1.813e-15
c23175 159 0 1.5696e-14
c23176 160 27 1.88e-16
c23177 5442 5453 6.73e-16
c23178 5446 5445 2.67e-16
c23179 617 633 1.621e-15
c23180 539 540 6.67e-16
c23181 1502 1500 1.6e-16
c23182 2944 2933 3.92e-16
c23183 1748 1363 1.96e-16
c23184 960 1 3.06e-16
c23185 943 0 2.6164e-14
c23186 4832 4828 1.96e-16
c23187 3129 647 1.58e-16
c23188 3126 672 1.58e-16
c23189 3034 3044 3.92e-16
c23190 3048 3020 3.54e-16
c23191 1660 0 3.26e-15
c23192 5182 5174 3.92e-16
c23193 440 437 6.67e-16
c23194 339 337 1.257e-15
c23195 565 175 1.88e-16
c23196 3604 737 1.58e-16
c23197 2339 2367 2.64e-16
c23198 2361 2357 1.96e-16
c23199 165 508 1.88e-16
c23200 64 265 1.88e-16
c23201 4068 4072 3.84e-16
c23202 4076 4075 4.41e-16
c23203 4719 0 3.9416e-13
c23204 2916 2917 2.67e-16
c23205 2924 2913 6.73e-16
c23206 910 907 6.76e-16
c23207 911 883 1.88e-16
c23208 2577 2169 1.136e-15
c23209 3973 19 9.67e-16
c23210 1321 1166 5.5e-16
c23211 1331 1627 1.58e-16
c23212 3537 1 4.41e-15
c23213 4371 0 6.62e-16
c23214 3100 662 1.58e-16
c23215 5288 352 3.54e-16
c23216 5188 207 3.54e-16
c23217 910 1682 3.45e-16
c23218 3387 3304 5.5e-16
c23219 5291 5318 4.01e-16
c23220 3397 3506 1.58e-16
c23221 3270 3655 1.96e-16
c23222 1 26 2.9261e-14
c23223 2155 2153 2.61e-16
c23224 1025 662 5.74e-16
c23225 642 3472 1.58e-16
c23226 3393 842 3.15e-16
c23227 5260 5165 3.87e-16
c23228 4915 149 1.88e-16
c23229 632 3458 1.84e-16
c23230 777 0 2.86343e-13
c23231 2194 2338 3.92e-16
c23232 3616 807 1.58e-16
c23233 1218 894 1.96e-16
c23234 1106 1101 1.58e-16
c23235 691 25 7.64e-16
c23236 4616 4609 1.96e-16
c23237 3874 4618 1.914e-15
c23238 1690 1318 1.58e-16
c23239 2535 2557 4.078e-15
c23240 2559 2541 4.312e-15
c23241 617 971 3.15e-16
c23242 711 700 7.23e-16
c23243 3048 2668 1.58e-16
c23244 3046 2662 5.5e-16
c23245 3034 3189 1.58e-16
c23246 3211 732 1.58e-16
c23247 2022 2133 1.58e-16
c23248 4810 4815 5.53e-16
c23249 1 571 1.607e-15
c23250 37 523 1.88e-16
c23251 27 513 1.88e-16
c23252 3185 3577 2.38e-15
c23253 4580 4622 3.92e-16
c23254 2409 1902 2.48e-16
c23255 48 15 6.58e-16
c23256 3851 2987 3.54e-16
c23257 60 63 6.67e-16
c23258 397 175 1.88e-16
c23259 642 3387 3.15e-16
c23260 3548 707 3.15e-16
c23261 2704 2706 2.03e-16
c23262 1363 1358 1.642e-15
c23263 2231 2603 1.58e-16
c23264 3558 0 6.62e-16
c23265 4826 797 1.23e-16
c23266 1806 1803 5.5e-16
c23267 822 827 2.77e-16
c23268 3748 0 2.703e-14
c23269 3947 1 6.66e-16
c23270 601 4256 1.09e-16
c23271 4437 3605 2.48e-16
c23272 1082 0 1.0044e-14
c23273 2559 732 3.58e-16
c23274 1708 1884 3.92e-16
c23275 37 317 5.71e-16
c23276 4563 4592 1.58e-16
c23277 2196 1800 1.58e-16
c23278 2866 2879 4.68e-16
c23279 3583 732 2.65e-16
c23280 3344 3409 1.58e-16
c23281 2249 2240 3.92e-16
c23282 1732 2243 5.66e-16
c23283 2612 2601 1.96e-16
c23284 2586 1 5.808e-15
c23285 907 906 8.88e-16
c23286 909 882 1.58e-16
c23287 890 895 3.54e-16
c23288 894 904 1.58e-16
c23289 883 879 3.84e-16
c23290 1837 702 1.58e-16
c23291 617 3055 1.75e-16
c23292 3163 1 2.054e-15
c23293 1581 782 1.09e-16
c23294 5587 4582 6.7e-16
c23295 4634 5450 3.54e-16
c23296 2702 747 5.73e-16
c23297 617 987 4.98e-16
c23298 669 1 5.57e-16
c23299 2668 3179 1.96e-16
c23300 1636 1630 1.6e-16
c23301 1166 1627 2.386e-15
c23302 1684 1866 1.58e-16
c23303 1706 1854 1.58e-16
c23304 4418 4419 1.35e-16
c23305 1912 1903 3.46e-16
c23306 1959 0 1.4092e-14
c23307 762 919 3.15e-16
c23308 3046 707 4.46e-16
c23309 3034 717 7.99e-16
c23310 3236 3625 2.386e-15
c23311 3634 3628 1.6e-16
c23312 657 3046 3.15e-16
c23313 2502 1981 1.96e-16
c23314 2497 1987 1.96e-16
c23315 2194 822 3.15e-16
c23316 2172 2286 1.58e-16
c23317 2194 2274 1.58e-16
c23318 3276 822 5.73e-16
c23319 2957 2921 1.58e-16
c23320 3368 3366 2.61e-16
c23321 1789 1 2.054e-15
c23322 2225 2221 1.96e-16
c23323 2747 3257 1.58e-16
c23324 2545 852 7.99e-16
c23325 2557 858 1.58e-16
c23326 1791 0 8e-16
c23327 462 465 3.54e-16
c23328 1 187 5.175e-15
c23329 3409 3072 1.58e-16
c23330 3628 3627 1.6e-16
c23331 3242 3623 3.92e-16
c23332 3393 3455 1.58e-16
c23333 2196 2461 1.58e-16
c23334 3781 3775 1.572e-15
c23335 3972 857 1.88e-16
c23336 3932 3934 2.254e-15
c23337 687 3160 1.58e-16
c23338 2782 2773 3.92e-16
c23339 601 3056 1.339e-15
c23340 2861 2475 5.66e-16
c23341 2680 2682 1.6e-16
c23342 1321 966 1.58e-16
c23343 2756 762 1.58e-16
c23344 3048 2538 3.54e-16
c23345 3898 3622 1.58e-16
c23346 2452 837 1.813e-15
c23347 2196 767 3.15e-16
c23348 822 812 3.28e-16
c23349 1042 0 1.8851e-14
c23350 2070 2069 1.96e-16
c23351 1694 2020 4.63e-16
c23352 3538 3541 6.44e-16
c23353 4479 1 8.43e-16
c23354 1972 1973 2.48e-16
c23355 19 432 3.45e-16
c23356 4567 4578 3.92e-16
c23357 5072 5125 3.18e-16
c23358 332 349 1.138e-15
c23359 3185 692 1.58e-16
c23360 3568 707 4.81e-16
c23361 4903 4944 5.5e-16
c23362 4954 4950 1.583e-15
c23363 113 100 1.58e-16
c23364 3696 3697 5.65e-16
c23365 907 707 4.8e-16
c23366 883 1067 3.92e-16
c23367 890 1066 1.88e-16
c23368 2740 0 6.62e-16
c23369 687 3532 2.65e-16
c23370 3322 1 1.868e-15
c23371 2756 2401 1.58e-16
c23372 1640 842 7.38e-16
c23373 657 907 3.15e-16
c23374 4033 4030 1.76e-16
c23375 3312 0 2.93e-15
c23376 3133 1 8.43e-16
c23377 361 9 5.8e-16
c23378 2863 2860 3.01e-16
c23379 2859 2856 6.44e-16
c23380 841 1 4.03e-16
c23381 3158 3161 6.44e-16
c23382 1415 1 1.868e-15
c23383 602 1343 4.46e-16
c23384 595 1321 1.511e-15
c23385 4310 4677 1.58e-16
c23386 2807 812 1.58e-16
c23387 3270 792 3.79e-16
c23388 1405 0 2.93e-15
c23389 4451 792 2.4e-16
c23390 3022 3441 2.38e-15
c23391 632 1726 1.58e-16
c23392 4830 1 4.832e-15
c23393 77 78 3.84e-16
c23394 3397 782 3.15e-16
c23395 2172 1902 1.58e-16
c23396 2178 1896 5.88e-16
c23397 4519 868 2.4e-16
c23398 2645 1 5.97e-15
c23399 2920 1 1.23e-16
c23400 3666 1 8.43e-16
c23401 4322 3480 2.38e-15
c23402 3159 3161 2.03e-16
c23403 1698 1324 1.121e-15
c23404 1687 1335 7.84e-16
c23405 1521 1076 1.96e-16
c23406 1331 1355 1.58e-16
c23407 2533 3058 1.58e-16
c23408 4819 1 6.42e-16
c23409 4480 4842 1.58e-16
c23410 4847 4856 3.92e-16
c23411 4600 4595 1.536e-15
c23412 4589 4592 6.02e-16
c23413 4563 4723 1.58e-16
c23414 3411 3386 2.38e-16
c23415 3387 3383 3.54e-16
c23416 617 2605 1.9e-16
c23417 2182 1896 5.5e-16
c23418 2348 1 6.15e-16
c23419 976 977 1.238e-15
c23420 3791 3773 1.23e-16
c23421 383 323 1.58e-16
c23422 747 2378 2.72e-16
c23423 1466 677 3.64e-16
c23424 858 1217 1.58e-16
c23425 1208 852 1.58e-16
c23426 5452 5447 7.37e-16
c23427 5486 5485 5.87e-16
c23428 3879 3887 3.84e-16
c23429 1071 1508 7.84e-16
c23430 2923 2928 3.54e-16
c23431 2951 2949 3.54e-16
c23432 1014 1 2.972e-15
c23433 537 165 1.88e-16
c23434 1919 797 1.75e-16
c23435 1788 1397 4.11e-16
c23436 4047 19 3.84e-16
c23437 4056 0 2.0707e-14
c23438 1015 0 6.29e-16
c23439 3873 1 4.076e-15
c23440 3024 3104 1.58e-16
c23441 3046 3092 1.58e-16
c23442 1708 1590 1.58e-16
c23443 1706 1584 5.5e-16
c23444 1694 1985 1.58e-16
c23445 1546 0 6.72e-16
c23446 4591 0 2.93e-15
c23447 777 1091 1.58e-16
c23448 19 342 8.82e-16
c23449 0 343 6.224e-15
c23450 209 205 6.38e-16
c23451 565 436 1.88e-16
c23452 5198 1 1.021e-15
c23453 2374 2385 1.96e-16
c23454 5241 0 2.078e-15
c23455 1766 2273 2.48e-16
c23456 272 273 6.67e-16
c23457 3497 647 1.58e-16
c23458 4330 662 4.81e-16
c23459 2850 2452 4.36e-16
c23460 2826 822 2.72e-16
c23461 2678 2282 1.96e-16
c23462 1134 767 8.3e-16
c23463 657 664 1.6e-16
c23464 4520 1 3.761e-15
c23465 4623 468 5.8e-16
c23466 2535 2684 3.92e-16
c23467 3871 1 1.96e-16
c23468 4389 3554 1.96e-16
c23469 4394 3548 1.96e-16
c23470 4662 4276 4.11e-16
c23471 4667 4658 3.46e-16
c23472 4421 762 1.58e-16
c23473 5022 5018 1.086e-15
c23474 1898 1 9.28e-16
c23475 426 427 6.96e-16
c23476 3393 3185 5.88e-16
c23477 2540 2544 5.8e-16
c23478 3882 782 3.15e-16
c23479 5558 5556 1.609e-15
c23480 5560 5543 9.36e-16
c23481 1076 752 1.58e-16
c23482 1579 1576 5.5e-16
c23483 758 0 1.1373e-14
c23484 594 1 5.57e-16
c23485 529 0 1.4515e-14
c23486 3608 0 3.3551e-14
c23487 1836 1837 2.48e-16
c23488 1687 1 8.766e-15
c23489 4367 0 3.6274e-14
c23490 1 190 1.65e-15
c23491 123 0 1.4515e-14
c23492 120 33 3.08e-16
c23493 3387 732 3.15e-16
c23494 3591 3603 2.32e-16
c23495 4582 4310 5.5e-16
c23496 4708 323 5.88e-16
c23497 2282 2271 1.58e-16
c23498 2455 2453 1.6e-16
c23499 3725 3844 1.52e-16
c23500 2848 1 8.43e-16
c23501 2172 2173 1.487e-15
c23502 59 479 1.88e-16
c23503 3463 4280 1.58e-16
c23504 3565 732 3.79e-16
c23505 5417 5404 1.96e-16
c23506 5388 5396 3.258e-15
c23507 920 995 3.92e-16
c23508 921 994 2.54e-16
c23509 3719 3321 4.36e-16
c23510 3424 1 2.054e-15
c23511 3426 0 8e-16
c23512 4027 1 6.78e-16
c23513 3876 4383 3.92e-16
c23514 4457 4458 1.6e-16
c23515 4453 3622 3.92e-16
c23516 2412 782 5.03e-16
c23517 974 1 3.06e-16
c23518 3318 3315 3.01e-16
c23519 3314 3311 6.44e-16
c23520 4016 0 6.8533e-14
c23521 4726 4728 1.687e-15
c23522 4738 4731 6.73e-16
c23523 4737 4350 1.96e-16
c23524 3338 2821 1.136e-15
c23525 3146 672 1.58e-16
c23526 565 349 1.88e-16
c23527 3808 3807 3.54e-16
c23528 59 189 1.88e-16
c23529 421 223 1.88e-16
c23530 5360 5291 3.54e-16
c23531 5355 5366 1.619e-15
c23532 1344 886 3.54e-16
c23533 2254 0 3.5926e-14
c23534 1604 797 4.81e-16
c23535 1411 1408 3.01e-16
c23536 1407 1404 6.44e-16
c23537 3882 4382 1.58e-16
c23538 2535 2649 1.58e-16
c23539 2557 2637 1.58e-16
c23540 3030 3035 8.56e-16
c23541 1932 1931 1.6e-16
c23542 1924 1922 2.15e-16
c23543 1694 1748 4.63e-16
c23544 1218 1 3.98e-16
c23545 5010 3744 1.14e-16
c23546 3034 3380 6.18e-16
c23547 4899 4897 8.88e-16
c23548 5277 5371 5.82e-16
c23549 596 685 2.45e-16
c23550 2172 2355 3.92e-16
c23551 926 929 1.928e-15
c23552 3799 3734 6.67e-16
c23553 3886 752 3.15e-16
c23554 4472 797 1.832e-15
c23555 3213 0 3.466e-15
c23556 919 1130 3.92e-16
c23557 922 1129 2.54e-16
c23558 1327 1453 1.96e-16
c23559 713 0 1.1384e-14
c23560 4553 3707 1.96e-16
c23561 2497 842 1.9e-16
c23562 4884 0 1.5788e-14
c23563 3024 2679 5.5e-16
c23564 3034 3194 1.58e-16
c23565 1684 1652 3.92e-16
c23566 1650 1 6.15e-16
c23567 4715 0 6.72e-16
c23568 1902 0 3.6368e-14
c23569 2006 2008 2.03e-16
c23570 3411 692 3.15e-16
c23571 3975 3972 1.58e-16
c23572 4580 4639 3.92e-16
c23573 5172 5171 1.6e-16
c23574 2407 2418 1.58e-16
c23575 378 362 3.84e-16
c23576 397 349 1.88e-16
c23577 4266 4277 1.96e-16
c23578 2231 2623 2.38e-15
c23579 3573 0 2.93e-15
c23580 2559 3003 3.25e-16
c23581 1473 1031 4.97e-16
c23582 627 4270 2.72e-16
c23583 2879 2900 4.41e-16
c23584 2907 2896 3.92e-16
c23585 3203 2685 1.96e-16
c23586 3204 3197 6.73e-16
c23587 3191 3576 1.96e-16
c23588 898 893 3.82e-16
c23589 291 508 1.88e-16
c23590 4527 0 6.72e-16
c23591 4563 4609 1.58e-16
c23592 4580 4621 1.58e-16
c23593 3574 737 1.58e-16
c23594 2341 2343 2.03e-16
c23595 2241 0 6.62e-16
c23596 4838 5074 1.53e-15
c23597 642 2577 1.58e-16
c23598 596 717 1.96e-16
c23599 2606 1 2.054e-15
c23600 7 13 1.88e-16
c23601 4855 4469 1.179e-15
c23602 1327 852 4.03e-16
c23603 1457 1469 2.32e-16
c23604 4158 3918 6.32e-16
c23605 617 3464 3.64e-16
c23606 601 3083 1.58e-16
c23607 3362 0 1.7608e-14
c23608 1388 957 4.97e-16
c23609 2832 2441 1.136e-15
c23610 4623 64 1.88e-16
c23611 2827 827 1.84e-16
c23612 1708 1883 5.42e-16
c23613 1684 1871 1.58e-16
c23614 1438 0 1.6491e-14
c23615 1241 1 1.23e-16
c23616 494 476 1.58e-16
c23617 1811 1817 1.418e-15
c23618 1828 1800 2.64e-16
c23619 2249 2238 1.96e-16
c23620 2790 2401 2.386e-15
c23621 2773 2418 1.58e-16
c23622 5229 5244 7.95e-16
c23623 4821 323 1.88e-16
c23624 2316 2311 1.642e-15
c23625 391 390 5.8e-16
c23626 381 412 1.88e-16
c23627 4060 4054 1.96e-16
c23628 1345 702 3.58e-16
c23629 3918 3948 2.87e-16
c23630 2976 1 7.49e-16
c23631 2172 2291 1.58e-16
c23632 4347 4345 1.6e-16
c23633 3182 3179 3.01e-16
c23634 1690 782 3.15e-16
c23635 1211 858 3.15e-16
c23636 3551 1 1.056e-15
c23637 2305 2688 7.84e-16
c23638 1549 1540 3.46e-16
c23639 3685 822 2.65e-16
c23640 642 1760 3.79e-16
c23641 595 1355 1.58e-16
c23642 4140 1 4.64e-16
c23643 3034 2838 1.58e-16
c23644 2657 677 1.84e-16
c23645 762 894 8.34e-16
c23646 4868 4866 1.6e-16
c23647 3271 3265 1.6e-16
c23648 2747 3262 2.386e-15
c23649 215 214 6.67e-16
c23650 3397 3134 5.5e-16
c23651 5247 5224 8.66e-16
c23652 3559 3168 4.11e-16
c23653 1678 1 5.329e-15
c23654 517 516 1.58e-16
c23655 762 2402 2.65e-16
c23656 894 883 4.116e-15
c23657 1232 890 1.96e-16
c23658 1234 909 1.58e-16
c23659 919 722 3.15e-16
c23660 920 1053 1.58e-16
c23661 1345 981 1.58e-16
c23662 1331 1418 1.58e-16
c23663 1196 1199 6.13e-16
c23664 602 1366 4.81e-16
c23665 3882 3633 5.88e-16
c23666 3876 3639 1.58e-16
c23667 4111 37 1.88e-16
c23668 2545 2768 1.58e-16
c23669 747 1089 1.58e-16
c23670 4401 4781 1.96e-16
c23671 2108 2105 1.931e-15
c23672 546 535 2.45e-16
c23673 1879 2396 2.38e-15
c23674 4954 4903 2.45e-16
c23675 5331 323 4.88e-16
c23676 3034 842 3.15e-16
c23677 2173 0 1.4835e-14
c23678 3411 3393 4.312e-15
c23679 2765 1 1.868e-15
c23680 2755 0 2.93e-15
c23681 2576 1 8.43e-16
c23682 687 3151 3.79e-16
c23683 3731 3762 6.73e-16
c23684 4520 4950 2.213e-15
c23685 5310 5299 1.96e-16
c23686 2815 1 5.97e-15
c23687 2559 2175 3.54e-16
c23688 1331 837 7.99e-16
c23689 4521 858 1.339e-15
c23690 3846 1 3.36e-16
c23691 4088 25 7.01e-16
c23692 4414 4407 6.73e-16
c23693 4413 3571 1.96e-16
c23694 1868 737 2.33e-16
c23695 1609 1610 2.48e-16
c23696 601 1343 4.46e-16
c23697 4310 4694 1.36e-15
c23698 4703 4697 1.6e-16
c23699 2827 812 1.58e-16
c23700 4455 0 3.3724e-14
c23701 2742 752 1.84e-16
c23702 4974 4975 3.54e-16
c23703 4993 4946 3.18e-16
c23704 2855 858 3.69e-16
c23705 3350 3347 5.5e-16
c23706 3271 782 7.68e-16
c23707 2546 1 3.009e-15
c23708 1082 707 1.58e-16
c23709 2547 0 5.86e-16
c23710 2194 1913 5.5e-16
c23711 3898 837 3.15e-16
c23712 4634 5461 1.96e-16
c23713 2645 2634 1.58e-16
c23714 1354 880 2.48e-16
c23715 919 1188 1.58e-16
c23716 2535 2536 1.487e-15
c23717 2545 2538 1.58e-16
c23718 1607 827 2.33e-16
c23719 1694 752 3.15e-16
c23720 1327 1101 1.58e-16
c23721 612 962 2.68e-16
c23722 623 0 1.1593e-14
c23723 4196 3879 9.33e-16
c23724 2533 3078 2.38e-15
c23725 4285 1 5.808e-15
c23726 4287 0 3.466e-15
c23727 3350 3357 6.73e-16
c23728 3030 3292 1.96e-16
c23729 4836 1 6.42e-16
c23730 3264 767 1.9e-16
c23731 2205 2207 2.03e-16
c23732 9 455 5.8e-16
c23733 4563 4740 1.58e-16
c23734 5165 5162 1.96e-16
c23735 4691 33 1.88e-16
c23736 2357 1 1.716e-15
c23737 782 775 5.58e-16
c23738 0 425 1.5723e-14
c23739 3781 3861 3.01e-16
c23740 5426 0 2.8602e-14
c23741 2937 1 1.257e-15
c23742 1031 677 3.15e-16
c23743 909 1173 3.54e-16
c23744 4708 5324 5.37e-16
c23745 2948 294 2.51e-16
c23746 1076 1520 1.58e-16
c23747 3106 0 3.5926e-14
c23748 3656 4489 7.84e-16
c23749 2453 797 3.64e-16
c23750 3354 2832 1.96e-16
c23751 3349 2838 1.96e-16
c23752 4231 1 4.442e-15
c23753 4745 4757 2.62e-16
c23754 1684 1601 5.5e-16
c23755 1694 1990 1.58e-16
c23756 4608 0 2.93e-15
c23757 677 693 1.621e-15
c23758 25 491 7.06e-16
c23759 3920 3917 1.76e-16
c23760 5068 5069 3.54e-16
c23761 2117 0 3.6242e-14
c23762 71 19 3.84e-16
c23763 78 450 1.88e-16
c23764 3514 672 2.22e-16
c23765 4336 677 1.832e-15
c23766 3327 3709 2.48e-16
c23767 1805 677 5.03e-16
c23768 1166 837 1.813e-15
c23769 1001 1435 1.58e-16
c23770 1016 1423 1.58e-16
c23771 1425 986 4.11e-16
c23772 3876 4417 3.92e-16
c23773 2559 2701 3.92e-16
c23774 787 1 5.62e-16
c23775 4038 19 7.04e-16
c23776 2361 722 1.9e-16
c23777 508 484 1.88e-16
c23778 4419 0 1.6491e-14
c23779 3423 3018 4.11e-16
c23780 2987 2518 7.46e-16
c23781 1911 1 6.15e-16
c23782 244 247 1.099e-15
c23783 3349 842 1.9e-16
c23784 2506 1 1.056e-15
c23785 1057 692 1.58e-16
c23786 1038 1044 1.58e-16
c23787 4005 4006 3.15e-16
c23788 2826 2827 1.6e-16
c23789 1322 1323 6.67e-16
c23790 921 1175 1.96e-16
c23791 1331 1061 5.5e-16
c23792 880 0 4.8002e-14
c23793 4241 1 8.43e-16
c23794 4215 4566 1.621e-15
c23795 4558 4559 4.57e-16
c23796 1781 1782 9.1e-16
c23797 3689 3304 1.96e-16
c23798 1704 0 1.2366e-14
c23799 4384 0 3.6274e-14
c23800 2045 2042 3.92e-16
c23801 4821 265 1.88e-16
c23802 2291 0 3.3692e-14
c23803 3801 3739 3.54e-16
c23804 3810 3811 5.07e-16
c23805 5170 0 2.1607e-14
c23806 3074 0 2.93e-15
c23807 2178 2186 8.73e-16
c23808 1436 672 2.4e-16
c23809 1192 1194 7.84e-16
c23810 1011 1018 7.95e-16
c23811 134 133 6.67e-16
c23812 3463 4285 1.58e-16
c23813 4407 737 1.58e-16
c23814 2637 2649 2.32e-16
c23815 537 291 1.88e-16
c23816 1890 737 1.9e-16
c23817 3442 0 6.72e-16
c23818 4208 19 3.84e-16
c23819 2518 2015 1.96e-16
c23820 2432 782 1.09e-16
c23821 4846 4463 4.97e-16
c23822 4849 4845 1.96e-16
c23823 942 889 1.185e-15
c23824 0 253 1.0822e-14
c23825 5457 439 4.88e-16
c23826 2196 2192 3.92e-16
c23827 2045 0 2.703e-14
c23828 2824 0 3.3717e-14
c23829 3417 0 3.22e-16
c23830 2136 2082 1.791e-15
c23831 1151 1149 1.931e-15
c23832 2713 0 6.9481e-14
c23833 742 1 5.62e-16
c23834 4398 1 1.056e-15
c23835 1339 1 1.002e-15
c23836 4980 1 4.081e-15
c23837 4902 4923 4.41e-16
c23838 4930 4919 3.92e-16
c23839 2260 1743 2.38e-15
c23840 229 216 1.58e-16
c23841 390 0 4.6653e-14
c23842 285 291 1.58e-16
c23843 4838 33 1.88e-16
c23844 1386 647 1.75e-16
c23845 902 926 3.54e-16
c23846 4719 5355 9.43e-16
c23847 3233 0 8e-16
c23848 1253 1243 1.318e-15
c23849 1076 1079 6.13e-16
c23850 1706 837 3.15e-16
c23851 1961 797 1.09e-16
c23852 1569 1568 1.6e-16
c23853 1561 1559 2.15e-16
c23854 1343 1470 3.92e-16
c23855 4633 4626 1.96e-16
c23856 4242 4635 1.914e-15
c23857 1708 1352 1.58e-16
c23858 1706 1319 5.5e-16
c23859 3327 1 4.41e-15
c23860 2688 702 1.58e-16
c23861 822 919 3.15e-16
c23862 721 719 5.88e-16
c23863 4920 0 1.63e-15
c23864 3048 2696 5.5e-16
c23865 2162 1641 1.96e-16
c23866 1 49 4.563e-15
c23867 3387 3519 3.92e-16
c23868 4563 4463 5.88e-16
c23869 5259 5263 1.202e-15
c23870 3202 3191 1.58e-16
c23871 0 37 3.65105e-13
c23872 4732 0 6.72e-16
c23873 926 928 1.61e-16
c23874 4580 4656 3.92e-16
c23875 5326 1 1.021e-15
c23876 2426 1913 4.97e-16
c23877 1243 1264 1.96e-16
c23878 3836 3842 6.23e-16
c23879 3804 3809 7.46e-16
c23880 3025 0 1.4835e-14
c23881 2541 2435 5.88e-16
c23882 921 767 3.15e-16
c23883 1001 978 6.54e-16
c23884 1327 1452 1.58e-16
c23885 3024 1 3.564e-15
c23886 3886 4536 4.63e-16
c23887 4543 4544 1.6e-16
c23888 4176 0 1.52701e-13
c23889 929 1 4.011e-15
c23890 2194 672 3.15e-16
c23891 2172 647 4.48e-16
c23892 3291 2781 1.58e-16
c23893 2696 2685 1.58e-16
c23894 1643 1645 2.03e-16
c23895 4710 4327 4.97e-16
c23896 4713 4709 1.96e-16
c23897 2541 752 3.15e-16
c23898 1 581 1.456e-15
c23899 4563 4626 1.58e-16
c23900 4580 4638 1.58e-16
c23901 2410 2422 2.32e-16
c23902 2196 1828 5.5e-16
c23903 2256 0 2.93e-15
c23904 3338 3857 3.92e-16
c23905 4872 5010 1.96e-16
c23906 2716 2714 1.6e-16
c23907 2788 0 1.6491e-14
c23908 2231 2627 1.96e-16
c23909 2237 2622 1.96e-16
c23910 2178 2508 1.96e-16
c23911 617 3083 3.15e-16
c23912 2880 2876 6.9e-16
c23913 2882 2897 1.96e-16
c23914 2545 2802 1.58e-16
c23915 4438 4450 2.32e-16
c23916 2545 2237 1.58e-16
c23917 697 1 5.62e-16
c23918 3725 468 1.952e-15
c23919 3944 37 5.71e-16
c23920 2679 3196 4.11e-16
c23921 595 1319 2.22e-16
c23922 3579 3576 3.01e-16
c23923 1708 1888 1.58e-16
c23924 3393 3672 1.96e-16
c23925 5010 0 2.81591e-13
c23926 2787 807 1.58e-16
c23927 2610 1 8.43e-16
c23928 890 898 8.05e-16
c23929 762 1 4.1542e-14
c23930 5483 410 3.54e-16
c23931 2514 2004 2.91e-16
c23932 2516 2515 1.6e-16
c23933 2508 2182 4.63e-16
c23934 3759 3734 1.96e-16
c23935 687 3046 3.15e-16
c23936 1370 952 3.92e-16
c23937 1374 1375 1.6e-16
c23938 3967 3918 8.1e-16
c23939 2317 677 3.64e-16
c23940 3567 1 9.28e-16
c23941 883 1 3.3e-15
c23942 4530 4521 3.46e-16
c23943 910 2173 7.06e-16
c23944 2764 797 1.58e-16
c23945 2679 722 1.58e-16
c23946 3409 3100 5.5e-16
c23947 2401 1 5.97e-15
c23948 657 2254 1.58e-16
c23949 592 655 6.34e-16
c23950 2397 0 6.72e-16
c23951 2234 1 1.056e-15
c23952 136 218 1.88e-16
c23953 3942 3951 1.88e-16
c23954 5411 468 3.54e-16
c23955 4844 497 1.88e-16
c23956 777 1879 1.58e-16
c23957 1046 717 1.813e-15
c23958 2305 2686 3.92e-16
c23959 2691 2690 1.6e-16
c23960 4252 4249 6.44e-16
c23961 4256 4253 3.01e-16
c23962 3886 4501 1.58e-16
c23963 3898 3650 5.5e-16
c23964 3900 3656 1.58e-16
c23965 3684 4519 1.96e-16
c23966 1970 837 1.58e-16
c23967 3377 2855 1.96e-16
c23968 3931 1 6.78e-16
c23969 2747 3260 1.532e-15
c23970 3265 3266 5.65e-16
c23971 1718 1717 2.48e-16
c23972 3184 3175 3.46e-16
c23973 3168 3553 1.96e-16
c23974 313 303 8.86e-16
c23975 311 320 1.58e-16
c23976 19 204 3.84e-16
c23977 3364 858 9.97e-16
c23978 2179 0 4.1004e-14
c23979 4353 717 1.58e-16
c23980 4776 5209 1.96e-16
c23981 894 722 3.15e-16
c23982 890 1053 3.54e-16
c23983 909 1074 1.58e-16
c23984 5284 5283 3.92e-16
c23985 3358 1 1.056e-15
c23986 2772 2390 2.48e-16
c23987 1431 692 1.58e-16
c23988 1447 1440 1.96e-16
c23989 595 604 1.6e-16
c23990 537 484 1.88e-16
c23991 687 907 3.15e-16
c23992 108 112 1.372e-15
c23993 2875 2874 5.87e-16
c23994 702 19 1.41e-15
c23995 542 88 1.88e-16
c23996 4102 37 1.88e-16
c23997 3898 3480 5.5e-16
c23998 3582 3571 1.58e-16
c23999 1862 752 1.58e-16
c24000 857 26 7.12e-16
c24001 2822 837 1.58e-16
c24002 1694 1448 5.5e-16
c24003 1433 1 9.28e-16
c24004 617 1343 4.46e-16
c24005 4100 3041 1.96e-16
c24006 4475 0 1.4092e-14
c24007 3464 3072 1.96e-16
c24008 3465 3458 6.73e-16
c24009 332 343 2.45e-16
c24010 4952 4946 3.54e-16
c24011 2307 1800 2.48e-16
c24012 4850 4847 5.5e-16
c24013 792 1556 1.58e-16
c24014 4657 4661 1.81e-16
c24015 2562 0 1.23e-16
c24016 2172 1930 5.5e-16
c24017 4126 3918 6.32e-16
c24018 3129 0 1.4092e-14
c24019 2545 2540 1.58e-16
c24020 2541 2549 8.73e-16
c24021 2270 647 7.38e-16
c24022 1806 1420 5.66e-16
c24023 4853 1 6.42e-16
c24024 3046 3309 3.92e-16
c24025 592 610 6.34e-16
c24026 5422 497 1.96e-16
c24027 5270 1 1.672e-15
c24028 894 1188 3.54e-16
c24029 1203 1217 1.96e-16
c24030 88 281 1.88e-16
c24031 5479 5481 1.387e-15
c24032 2946 0 2.28e-15
c24033 381 64 1.88e-16
c24034 1516 767 1.58e-16
c24035 1534 1528 1.6e-16
c24036 1076 1525 2.386e-15
c24037 1327 971 5.88e-16
c24038 4079 1 5.284e-15
c24039 3667 4501 1.58e-16
c24040 2265 677 1.58e-16
c24041 1947 797 3.15e-16
c24042 837 26 1.58e-16
c24043 4069 0 1.5061e-14
c24044 4071 19 3.45e-16
c24045 3030 2600 1.58e-16
c24046 1568 1 1.868e-15
c24047 4248 1 4.442e-15
c24048 3173 692 7.38e-16
c24049 2083 2029 1.191e-15
c24050 4625 0 2.93e-15
c24051 1558 0 2.93e-15
c24052 303 320 1.325e-15
c24053 3151 3506 1.58e-16
c24054 3532 3526 1.6e-16
c24055 5072 5088 1.23e-16
c24056 2156 0 8e-16
c24057 4520 4531 1.58e-16
c24058 1608 827 1.339e-15
c24059 3900 4434 3.92e-16
c24060 910 880 5.03e-16
c24061 647 0 2.80112e-13
c24062 1344 1328 3.54e-16
c24063 3886 4264 4.63e-16
c24064 3852 0 1.65e-16
c24065 4679 4293 4.11e-16
c24066 4684 4675 3.46e-16
c24067 1584 1951 1.58e-16
c24068 1706 1799 3.92e-16
c24069 910 1704 1.58e-16
c24070 117 252 1.88e-16
c24071 49 363 1.88e-16
c24072 5001 4992 3.92e-16
c24073 4982 4978 3.54e-16
c24074 2293 1777 4.11e-16
c24075 165 164 3.84e-16
c24076 407 479 1.88e-16
c24077 3411 3208 1.58e-16
c24078 4827 1 3.7282e-14
c24079 2866 3030 4.3e-16
c24080 2526 1 7.21e-16
c24081 1057 1059 7.84e-16
c24082 2492 0 3.7647e-14
c24083 4685 497 1.88e-16
c24084 5569 5422 1.666e-15
c24085 3882 3381 1.58e-16
c24086 3876 3384 1.58e-16
c24087 1992 837 2.72e-16
c24088 602 905 1.58e-16
c24089 3060 2529 4.11e-16
c24090 2987 2988 3.54e-16
c24091 5013 5011 3.92e-16
c24092 4546 3751 1.96e-16
c24093 4896 5007 1.58e-16
c24094 3258 752 1.58e-16
c24095 3024 3257 1.58e-16
c24096 3046 3245 1.58e-16
c24097 2177 2181 5.8e-16
c24098 5306 5288 6.67e-16
c24099 4401 0 3.5918e-14
c24100 462 26 1.03e-15
c24101 453 0 9.795e-15
c24102 136 130 3.84e-16
c24103 245 258 1.108e-15
c24104 5136 5034 1.58e-16
c24105 4691 526 1.88e-16
c24106 2459 1953 3.92e-16
c24107 2463 2464 1.6e-16
c24108 2311 0 1.4092e-14
c24109 2761 2758 3.01e-16
c24110 2757 2754 6.44e-16
c24111 1016 692 1.58e-16
c24112 1205 827 1.58e-16
c24113 922 1025 3.92e-16
c24114 632 1001 3.57e-16
c24115 1331 1330 1.357e-15
c24116 4476 4475 5.65e-16
c24117 4470 3633 1.532e-15
c24118 2541 2871 1.96e-16
c24119 1567 1116 1.136e-15
c24120 3326 2815 1.96e-16
c24121 4028 26 4.58e-16
c24122 3034 2533 5.5e-16
c24123 1 194 1.1938e-14
c24124 131 49 1.88e-16
c24125 4691 4697 5.87e-16
c24126 19 175 3.84e-16
c24127 2289 0 1.6491e-14
c24128 1423 662 1.58e-16
c24129 2844 0 1.4092e-14
c24130 2260 2257 5.5e-16
c24131 4193 4190 1.76e-16
c24132 160 161 1.079e-15
c24133 3310 3696 5.66e-16
c24134 1161 1163 7.72e-16
c24135 3839 3796 2.74e-16
c24136 3876 4387 1.58e-16
c24137 3900 4399 5.42e-16
c24138 2196 717 3.58e-16
c24139 3902 1 2.86e-16
c24140 4011 25 4.68e-16
c24141 2355 707 1.58e-16
c24142 1664 1661 5.5e-16
c24143 1206 1331 1.58e-16
c24144 3885 0 1.5577e-14
c24145 3148 662 1.09e-16
c24146 3124 2611 1.532e-15
c24147 1937 1948 1.96e-16
c24148 1690 1781 1.58e-16
c24149 3532 3134 4.36e-16
c24150 662 652 6.38e-16
c24151 595 2206 1.58e-16
c24152 910 3025 7.06e-16
c24153 421 233 1.88e-16
c24154 288 26 1.03e-15
c24155 277 0 1.051e-14
c24156 5514 1 5.868e-15
c24157 2658 0 6.72e-16
c24158 657 3106 1.58e-16
c24159 1403 672 5.73e-16
c24160 1795 647 3.64e-16
c24161 981 1406 7.84e-16
c24162 3068 1 9.28e-16
c24163 1270 1275 3.54e-16
c24164 4855 149 1.88e-16
c24165 1321 1487 3.92e-16
c24166 2611 3125 4.97e-16
c24167 2617 2628 1.58e-16
c24168 1684 1363 5.5e-16
c24169 3225 762 1.58e-16
c24170 2517 858 6.67e-16
c24171 2508 852 2.4e-16
c24172 3134 702 1.58e-16
c24173 4918 4920 3.92e-16
c24174 631 629 5.88e-16
c24175 3411 3536 3.92e-16
c24176 2748 2350 4.36e-16
c24177 837 841 2.19e-16
c24178 902 888 3.84e-16
c24179 595 2578 2.65e-16
c24180 602 2169 2.33e-16
c24181 1930 0 6.9481e-14
c24182 3781 3732 2.652e-15
c24183 4001 3998 1.76e-16
c24184 4580 4673 3.92e-16
c24185 5556 0 1.1948e-14
c24186 5498 470 5.93e-16
c24187 5066 91 3.54e-16
c24188 2196 2371 5.42e-16
c24189 2172 2359 1.58e-16
c24190 134 0 9.795e-15
c24191 146 25 5.71e-16
c24192 5410 5414 1.96e-16
c24193 3031 0 4.1004e-14
c24194 2557 2452 5.5e-16
c24195 1016 1020 2.03e-16
c24196 4287 3452 1.96e-16
c24197 4292 3446 1.96e-16
c24198 1343 1469 1.58e-16
c24199 1327 1457 1.58e-16
c24200 3412 1 2.86e-16
c24201 2248 2237 1.58e-16
c24202 4540 3882 3.16e-16
c24203 3886 3876 4.116e-15
c24204 3024 2634 1.58e-16
c24205 1448 1815 1.58e-16
c24206 822 894 8.34e-16
c24207 902 1 9.725e-15
c24208 3299 3305 1.6e-16
c24209 3296 2781 2.386e-15
c24210 2798 3279 1.58e-16
c24211 2696 3220 4.36e-16
c24212 2015 858 3.15e-16
c24213 2018 2016 1.6e-16
c24214 762 1321 3.15e-16
c24215 4563 4643 1.58e-16
c24216 4580 4655 1.58e-16
c24217 5171 5174 3.92e-16
c24218 5542 584 8.44e-16
c24219 824 825 1.6e-16
c24220 1187 837 2.68e-16
c24221 890 1127 1.96e-16
c24222 921 931 1.58e-16
c24223 230 232 7.1e-16
c24224 4702 1 2.3324e-14
c24225 1477 1474 5.5e-16
c24226 2702 1 4.41e-15
c24227 3886 3520 1.58e-16
c24228 915 0 2.94e-16
c24229 3122 647 7.38e-16
c24230 1690 1522 1.58e-16
c24231 601 1744 3.64e-16
c24232 602 1363 1.58e-16
c24233 204 195 1.58e-16
c24234 3489 3501 2.32e-16
c24235 5010 4918 1.715e-15
c24236 5036 5026 9.99e-16
c24237 2353 2351 1.6e-16
c24238 1 15 6.0789e-14
c24239 2625 2622 3.01e-16
c24240 2621 2618 6.44e-16
c24241 9 45 4.88e-16
c24242 7 27 1.88e-16
c24243 6 0 1.5696e-14
c24244 5200 5239 1.858e-15
c24245 4838 526 1.88e-16
c24246 2178 2507 1.58e-16
c24247 4076 4077 7.81e-16
c24248 1254 1255 3.92e-16
c24249 4355 4356 1.6e-16
c24250 4351 3520 3.92e-16
c24251 4457 797 5.03e-16
c24252 1811 677 3.15e-16
c24253 1331 1606 4.63e-16
c24254 689 0 7.709e-15
c24255 3580 1 6.15e-16
c24256 4161 1 3.3163e-14
c24257 3497 0 6.915e-14
c24258 2194 797 4.46e-16
c24259 4885 4883 1.6e-16
c24260 3364 3377 3.92e-16
c24261 3307 797 4.81e-16
c24262 4869 0 8e-16
c24263 3222 722 4.81e-16
c24264 2713 707 1.58e-16
c24265 2132 2131 1.08e-15
c24266 1 507 1.073e-15
c24267 13 508 1.88e-16
c24268 3642 3641 2.48e-16
c24269 5239 5251 1.96e-16
c24270 5230 5237 1.96e-16
c24271 5165 5224 3.54e-16
c24272 2196 1987 1.58e-16
c24273 2182 2507 1.58e-16
c24274 1013 647 3.57e-16
c24275 3581 3572 3.46e-16
c24276 3276 797 2.33e-16
c24277 3780 3770 1.668e-15
c24278 3971 3964 7.81e-16
c24279 5284 1 1.0125e-14
c24280 1245 1242 4.03e-16
c24281 5522 5388 1.389e-15
c24282 642 992 2.68e-16
c24283 65 0 1.4515e-14
c24284 3355 3397 3.92e-16
c24285 2968 0 3.6242e-14
c24286 922 1083 1.58e-16
c24287 4156 4163 7.81e-16
c24288 722 1 3.1284e-14
c24289 3886 4506 1.58e-16
c24290 3876 3667 5.5e-16
c24291 1801 1812 1.96e-16
c24292 4135 37 1.88e-16
c24293 3943 1 3.66e-16
c24294 4136 26 1.075e-15
c24295 4418 4798 1.96e-16
c24296 2104 2108 3.54e-16
c24297 523 514 1.58e-16
c24298 25 320 5.71e-16
c24299 3644 797 5.03e-16
c24300 4567 3870 3.54e-16
c24301 1896 1885 1.58e-16
c24302 2328 2327 1.6e-16
c24303 791 790 6.67e-16
c24304 165 218 1.88e-16
c24305 4373 717 1.58e-16
c24306 4838 5069 1.152e-15
c24307 2783 1 9.28e-16
c24308 2687 2299 4.97e-16
c24309 1162 807 1.58e-16
c24310 883 1068 3.54e-16
c24311 894 1089 1.58e-16
c24312 4150 4149 3.15e-16
c24313 2214 2599 1.96e-16
c24314 1848 692 4.81e-16
c24315 2982 2984 1.609e-15
c24316 2887 2986 9.36e-16
c24317 4520 5577 1.361e-15
c24318 4514 4567 5.5e-16
c24319 602 3384 2.33e-16
c24320 595 4243 2.65e-16
c24321 4428 4421 1.96e-16
c24322 3582 4430 4.36e-16
c24323 1690 1324 1.96e-16
c24324 3083 3072 1.58e-16
c24325 1904 1906 2.03e-16
c24326 5036 120 3.54e-16
c24327 1960 0 6.72e-16
c24328 777 1567 2.22e-16
c24329 1074 1081 2.27e-16
c24330 894 892 5.93e-16
c24331 2572 0 1.4092e-14
c24332 2287 672 2.4e-16
c24333 1618 868 1.813e-15
c24334 1166 1606 1.96e-16
c24335 1345 1116 1.58e-16
c24336 1343 1106 5.5e-16
c24337 1331 1571 1.58e-16
c24338 627 976 1.35e-16
c24339 3101 2583 1.96e-16
c24340 3102 3095 6.73e-16
c24341 1188 1 1.56e-15
c24342 1886 1888 1.862e-15
c24343 1499 1505 1.418e-15
c24344 1516 1488 2.64e-16
c24345 363 194 1.88e-16
c24346 4299 0 3.6274e-14
c24347 5226 178 3.54e-16
c24348 3024 3326 3.92e-16
c24349 978 991 1.58e-16
c24350 4651 4265 1.179e-15
c24351 4580 4745 1.58e-16
c24352 4571 4757 1.58e-16
c24353 1981 2490 1.58e-16
c24354 5470 0 1.23e-16
c24355 864 863 1.96e-16
c24356 3794 3770 6.73e-16
c24357 1041 1043 7.72e-16
c24358 2535 2356 1.58e-16
c24359 1550 752 1.58e-16
c24360 642 3876 3.15e-16
c24361 3758 1 3.36e-16
c24362 3667 4506 2.386e-15
c24363 4515 4509 1.6e-16
c24364 1050 1 3.06e-16
c24365 4086 26 4.48e-16
c24366 1712 1707 9.6e-16
c24367 1121 1 5.821e-15
c24368 4265 1 4.442e-15
c24369 4762 4774 2.62e-16
c24370 3393 3434 1.96e-16
c24371 4642 0 2.93e-15
c24372 792 1557 1.58e-16
c24373 0 445 2.87e-16
c24374 19 436 3.84e-16
c24375 4563 4215 1.96e-16
c24376 4567 4559 1.88e-16
c24377 2359 0 3.3692e-14
c24378 1155 782 6.48e-16
c24379 108 100 2.218e-15
c24380 101 117 3.84e-16
c24381 3503 692 1.75e-16
c24382 2170 2581 1.58e-16
c24383 1625 868 1.58e-16
c24384 1436 1435 9.1e-16
c24385 838 1 1.65e-16
c24386 1505 1506 1.35e-16
c24387 1567 1959 2.38e-15
c24388 3445 3436 3.46e-16
c24389 2144 0 1.5808e-14
c24390 186 189 1.099e-15
c24391 4878 236 1.88e-16
c24392 2316 0 6.9484e-14
c24393 4070 3918 2.48e-16
c24394 3886 4263 1.58e-16
c24395 3898 3385 5.5e-16
c24396 3900 3418 1.58e-16
c24397 3673 827 2.33e-16
c24398 2845 2844 5.65e-16
c24399 687 1042 1.58e-16
c24400 1151 1588 1.58e-16
c24401 3259 0 3.6368e-14
c24402 602 3886 3.15e-16
c24403 3048 3274 5.42e-16
c24404 3024 3262 1.58e-16
c24405 596 757 3.134e-15
c24406 4418 0 3.6274e-14
c24407 4589 4594 5.53e-16
c24408 4674 5388 1.96e-16
c24409 2178 2235 1.58e-16
c24410 3588 752 2.33e-16
c24411 5450 5446 5.32e-16
c24412 1207 1208 7.46e-16
c24413 383 381 3.84e-16
c24414 4312 4305 6.73e-16
c24415 4311 3469 1.96e-16
c24416 1986 837 2.4e-16
c24417 3089 1 4.41e-15
c24418 3310 3321 1.58e-16
c24419 911 3879 1.58e-16
c24420 1507 1508 2.48e-16
c24421 1343 1328 1.632e-15
c24422 1327 1344 5.63e-16
c24423 3473 0 6.62e-16
c24424 4237 0 1.4092e-14
c24425 4676 4299 2.48e-16
c24426 1157 0 1.0183e-14
c24427 1720 0 3.466e-15
c24428 4781 0 3.466e-15
c24429 2559 807 3.58e-16
c24430 5158 5154 7.1e-16
c24431 2196 2405 5.42e-16
c24432 19 349 3.84e-16
c24433 37 332 1.88e-16
c24434 2549 2175 1.121e-15
c24435 2538 2186 7.84e-16
c24436 2372 1862 1.96e-16
c24437 2196 1715 1.58e-16
c24438 2182 2235 1.58e-16
c24439 129 132 2.142e-15
c24440 657 3129 1.58e-16
c24441 1440 672 1.58e-16
c24442 919 672 3.15e-16
c24443 281 277 1.58e-16
c24444 3900 3872 3.54e-16
c24445 3886 3896 3.92e-16
c24446 4321 677 5.03e-16
c24447 5358 5366 1.725e-15
c24448 2824 2441 7.84e-16
c24449 2541 2870 1.58e-16
c24450 1166 1143 6.54e-16
c24451 4293 4288 1.642e-15
c24452 3245 777 1.58e-16
c24453 2557 2288 1.58e-16
c24454 984 0 2.7376e-14
c24455 3228 3235 1.96e-16
c24456 3046 3071 3.92e-16
c24457 2028 2059 6.73e-16
c24458 4402 1 1.716e-15
c24459 37 259 5.71e-16
c24460 3140 677 2.33e-16
c24461 3313 827 1.58e-16
c24462 3046 782 4.46e-16
c24463 1987 1988 1.35e-16
c24464 88 565 1.88e-16
c24465 4861 5103 6.5e-16
c24466 3397 3191 1.58e-16
c24467 4571 4847 1.58e-16
c24468 4582 4859 1.58e-16
c24469 2741 2356 1.96e-16
c24470 986 1389 1.58e-16
c24471 3246 0 6.62e-16
c24472 3081 1 6.15e-16
c24473 3548 4382 1.58e-16
c24474 1828 717 1.813e-15
c24475 642 1772 1.58e-16
c24476 539 1 4.22e-16
c24477 537 13 1.88e-16
c24478 3611 1 2.054e-15
c24479 3152 2628 4.36e-16
c24480 1574 1585 1.96e-16
c24481 4650 4643 1.96e-16
c24482 4259 4652 1.914e-15
c24483 1708 1380 5.5e-16
c24484 2172 868 3.15e-16
c24485 2815 837 1.813e-15
c24486 4754 1 1.749e-15
c24487 3744 0 2.1497e-14
c24488 3228 752 1.58e-16
c24489 3034 2719 1.58e-16
c24490 2730 732 2.22e-16
c24491 2165 1708 3.54e-16
c24492 1852 0 1.6491e-14
c24493 3409 3552 1.58e-16
c24494 822 1 4.1542e-14
c24495 596 712 3.134e-15
c24496 3601 3600 1.6e-16
c24497 601 2169 1.75e-16
c24498 2274 1 5.808e-15
c24499 4580 4690 3.92e-16
c24500 5044 5056 3.18e-16
c24501 1278 1226 7.4e-16
c24502 4736 5385 1.383e-15
c24503 4708 381 1.88e-16
c24504 657 647 3.28e-16
c24505 2535 2469 5.5e-16
c24506 1321 1486 1.58e-16
c24507 1343 1474 1.58e-16
c24508 542 523 1.88e-16
c24509 2697 707 7.68e-16
c24510 2196 842 3.15e-16
c24511 1431 1823 2.38e-15
c24512 642 1684 3.15e-16
c24513 1117 0 1.8851e-14
c24514 4188 26 4.58e-16
c24515 4020 1 6.78e-16
c24516 4454 4453 2.03e-16
c24517 4459 4457 1.6e-16
c24518 1752 1750 1.862e-15
c24519 1677 1 9.43e-16
c24520 1694 1684 4.116e-15
c24521 2151 1690 3.16e-16
c24522 81 88 3.54e-16
c24523 4561 1 3.132e-15
c24524 4727 4344 4.97e-16
c24525 4730 4726 1.96e-16
c24526 1694 1935 4.63e-16
c24527 777 1345 3.58e-16
c24528 19 5 3.84e-16
c24529 602 2574 1.09e-16
c24530 4563 4660 1.58e-16
c24531 4580 4672 1.58e-16
c24532 2430 2427 5.5e-16
c24533 3600 752 7.68e-16
c24534 5383 0 1.1948e-14
c24535 2021 236 8.6e-16
c24536 3820 3809 1.138e-15
c24537 4753 5157 9.82e-16
c24538 2807 1 5.808e-15
c24539 907 782 4.8e-16
c24540 883 1142 3.92e-16
c24541 890 1141 1.88e-16
c24542 2809 0 3.466e-15
c24543 2646 1 1.868e-15
c24544 3404 1 7.228e-15
c24545 5352 5355 3.54e-16
c24546 5378 5377 1.6e-16
c24547 1854 722 1.58e-16
c24548 397 88 1.88e-16
c24549 3395 0 4.64e-16
c24550 3294 2781 1.532e-15
c24551 3996 26 4.58e-16
c24552 2325 692 1.832e-15
c24553 1655 1653 1.6e-16
c24554 3718 3882 4.3e-16
c24555 617 1744 7.68e-16
c24556 601 1363 3.15e-16
c24557 1491 1 5.808e-15
c24558 1493 0 3.466e-15
c24559 2189 1698 5.8e-16
c24560 1927 1924 3.01e-16
c24561 1923 1920 6.44e-16
c24562 747 1086 4e-16
c24563 25 577 7.06e-16
c24564 3593 752 5.03e-16
c24565 4928 1 2.36e-16
c24566 5207 207 3.54e-16
c24567 3374 3364 1.65e-16
c24568 3313 812 1.832e-15
c24569 1618 0 6.9481e-14
c24570 236 1 3.36e-15
c24571 894 962 3.92e-16
c24572 909 961 1.58e-16
c24573 883 955 1.58e-16
c24574 4165 4166 3.15e-16
c24575 3452 647 1.75e-16
c24576 3270 3276 1.418e-15
c24577 3397 858 3.15e-16
c24578 3287 3259 2.64e-16
c24579 1321 722 4.48e-16
c24580 1393 1392 5.65e-16
c24581 3045 1 2.94e-16
c24582 146 9 5.8e-16
c24583 4477 797 1.09e-16
c24584 2559 2265 5.5e-16
c24585 2541 2633 1.96e-16
c24586 1448 1011 1.136e-15
c24587 3112 3109 5.5e-16
c24588 747 753 1.097e-15
c24589 3502 3117 1.96e-16
c24590 2782 767 3.64e-16
c24591 571 563 2.218e-15
c24592 2262 2259 3.01e-16
c24593 2258 2255 6.44e-16
c24594 602 1694 3.15e-16
c24595 4886 0 8e-16
c24596 2419 1 1.868e-15
c24597 1641 1652 1.58e-16
c24598 1027 672 1.58e-16
c24599 4088 4036 1.88e-16
c24600 3270 812 1.58e-16
c24601 5533 526 9.15e-16
c24602 5296 0 2.1607e-14
c24603 5153 5152 5.87e-16
c24604 2409 0 2.93e-15
c24605 3014 1 1.601e-15
c24606 1489 732 1.58e-16
c24607 3876 732 3.15e-16
c24608 2797 2790 1.96e-16
c24609 5414 5406 3.54e-16
c24610 3004 0 6.78e-16
c24611 2708 2709 5.65e-16
c24612 4264 3429 1.96e-16
c24613 4546 852 1.58e-16
c24614 2469 858 1.58e-16
c24615 2481 842 1.84e-16
c24616 1089 1 2.972e-15
c24617 1090 0 6.29e-16
c24618 3279 3278 2.48e-16
c24619 3034 3173 4.63e-16
c24620 762 1102 1.58e-16
c24621 3641 3640 2.03e-16
c24622 3646 3644 1.6e-16
c24623 1625 0 1.6491e-14
c24624 3393 662 3.15e-16
c24625 3664 797 1.09e-16
c24626 4567 3874 5.5e-16
c24627 1164 812 1.58e-16
c24628 981 982 8.58e-16
c24629 3418 4251 7.84e-16
c24630 1664 852 1.58e-16
c24631 1467 1466 1.6e-16
c24632 1459 1457 2.15e-16
c24633 1384 971 1.58e-16
c24634 595 3385 2.22e-16
c24635 601 3384 1.75e-16
c24636 3898 4315 3.92e-16
c24637 4327 4316 1.58e-16
c24638 1447 1 8.43e-16
c24639 3479 3472 1.96e-16
c24640 3083 3481 4.36e-16
c24641 495 499 6.38e-16
c24642 488 477 2.45e-16
c24643 2324 1811 4.97e-16
c24644 4867 4864 5.5e-16
c24645 1726 2236 1.96e-16
c24646 3409 3253 5.5e-16
c24647 5323 5316 8.94e-16
c24648 5321 5318 1.342e-15
c24649 5262 5261 5.5e-16
c24650 1068 722 1.58e-16
c24651 1116 782 1.75e-16
c24652 397 390 7.76e-16
c24653 107 103 1.58e-16
c24654 3882 858 3.15e-16
c24655 4821 381 1.88e-16
c24656 5403 5417 5.12e-16
c24657 3909 19 7.04e-16
c24658 2010 858 1.84e-16
c24659 1321 1121 5.5e-16
c24660 1331 1576 1.58e-16
c24661 601 963 1.58e-16
c24662 856 25 7.64e-16
c24663 1541 1543 2.03e-16
c24664 642 1777 2.22e-16
c24665 3048 3343 3.92e-16
c24666 2036 178 3.39e-16
c24667 3397 3484 1.58e-16
c24668 3253 3621 1.96e-16
c24669 998 999 1.213e-15
c24670 596 622 3.134e-15
c24671 1 333 1.073e-15
c24672 9 320 5.8e-16
c24673 223 204 1.88e-16
c24674 3387 807 3.15e-16
c24675 4580 4762 1.58e-16
c24676 4571 4774 1.58e-16
c24677 5105 62 3.54e-16
c24678 1998 2478 1.58e-16
c24679 2172 2270 3.92e-16
c24680 391 0 1.5696e-14
c24681 375 25 7.06e-16
c24682 3038 2538 1.121e-15
c24683 3937 3928 1.88e-16
c24684 3900 692 3.15e-16
c24685 5484 5450 1.58e-16
c24686 5514 5409 1.58e-16
c24687 3027 2549 7.84e-16
c24688 1046 1023 6.54e-16
c24689 4322 4319 5.5e-16
c24690 920 1070 3.92e-16
c24691 921 1069 2.54e-16
c24692 687 1438 1.58e-16
c24693 80 74 1.372e-15
c24694 4129 1 2.8425e-14
c24695 868 0 2.8609e-13
c24696 2921 2923 1.09e-15
c24697 1064 1 3.06e-16
c24698 4111 0 2.1639e-14
c24699 3048 2617 1.58e-16
c24700 3046 2611 5.5e-16
c24701 3034 3138 1.58e-16
c24702 1386 0 3.6368e-14
c24703 4282 1 4.442e-15
c24704 4659 0 2.93e-15
c24705 3638 782 7.38e-16
c24706 5106 5115 1.96e-16
c24707 2400 2391 3.46e-16
c24708 5136 31 6.06e-16
c24709 602 3061 1.58e-16
c24710 921 717 3.15e-16
c24711 971 969 1.931e-15
c24712 4362 692 3.64e-16
c24713 2214 2569 1.58e-16
c24714 1026 1016 1.418e-15
c24715 657 3497 2.22e-16
c24716 3839 3809 6.53e-16
c24717 4406 4402 1.96e-16
c24718 4458 1 2.054e-15
c24719 4696 4310 4.11e-16
c24720 4701 4692 3.46e-16
c24721 479 252 1.88e-16
c24722 4460 0 8e-16
c24723 3157 717 5.73e-16
c24724 3024 837 3.15e-16
c24725 5049 0 2.156e-15
c24726 2215 2209 1.6e-16
c24727 1678 2206 2.386e-15
c24728 107 247 1.88e-16
c24729 4821 4816 1.536e-15
c24730 5284 5295 1.37e-16
c24731 4827 410 1.88e-16
c24732 2172 0 3.14305e-13
c24733 1544 767 5.03e-16
c24734 1106 1103 1.984e-15
c24735 3886 4268 1.58e-16
c24736 3876 3429 5.5e-16
c24737 4617 5425 9.04e-16
c24738 2768 2769 9.1e-16
c24739 919 1205 3.92e-16
c24740 922 1204 2.54e-16
c24741 811 25 7.64e-16
c24742 1988 842 1.339e-15
c24743 1136 1596 2.38e-15
c24744 1684 1815 1.58e-16
c24745 1706 1803 1.58e-16
c24746 601 3886 3.15e-16
c24747 4564 4566 3.67e-16
c24748 3082 3073 3.46e-16
c24749 2735 737 7.38e-16
c24750 1870 1488 2.48e-16
c24751 771 760 7.23e-16
c24752 3048 3279 1.58e-16
c24753 5592 563 5.31e-16
c24754 4922 4920 1.072e-15
c24755 3236 3603 1.58e-16
c24756 3225 3611 5.66e-16
c24757 3617 3608 3.92e-16
c24758 4435 0 3.6274e-14
c24759 2512 0 3.8803e-14
c24760 1 447 4.59e-16
c24761 3411 767 3.15e-16
c24762 2476 1964 1.532e-15
c24763 2482 2481 5.65e-16
c24764 2015 2028 4.68e-16
c24765 5578 5575 6.67e-16
c24766 2194 2252 1.58e-16
c24767 2178 2240 1.58e-16
c24768 630 1 1.65e-16
c24769 1684 732 3.15e-16
c24770 3498 1 1.868e-15
c24771 3647 0 8e-16
c24772 1693 1324 1.176e-15
c24773 4488 4489 2.48e-16
c24774 2231 647 1.58e-16
c24775 4743 4367 3.92e-16
c24776 4755 4754 1.6e-16
c24777 4798 0 3.466e-15
c24778 2031 2049 4.06e-16
c24779 1635 1607 2.64e-16
c24780 3608 3610 2.15e-16
c24781 767 757 6.38e-16
c24782 1 496 4.92e-16
c24783 470 30 3.84e-16
c24784 2540 2186 9.72e-16
c24785 5080 5069 9.85e-16
c24786 2182 2240 1.58e-16
c24787 2118 1 2.397e-15
c24788 103 1 1.65e-15
c24789 883 837 3.15e-16
c24790 595 2557 3.15e-16
c24791 602 2541 3.15e-16
c24792 920 677 3.69e-16
c24793 110 0 1.4803e-14
c24794 4199 4208 1.88e-16
c24795 4341 677 1.09e-16
c24796 1327 1320 1.58e-16
c24797 1345 1340 1.58e-16
c24798 2567 2166 1.532e-15
c24799 3898 3571 1.58e-16
c24800 3265 777 1.58e-16
c24801 2535 2305 1.58e-16
c24802 2342 732 1.58e-16
c24803 789 1 5.57e-16
c24804 4367 4744 2.48e-16
c24805 3024 3088 3.92e-16
c24806 822 1321 3.15e-16
c24807 4428 1 8.43e-16
c24808 2128 1 3.36e-16
c24809 601 2223 1.832e-15
c24810 2120 0 1.65e-16
c24811 4905 1 2.341e-15
c24812 5195 0 3.1318e-14
c24813 3333 827 1.58e-16
c24814 3330 868 1.58e-16
c24815 894 672 8.34e-16
c24816 4922 5010 1.705e-15
c24817 4878 4915 1.96e-16
c24818 4571 4864 1.58e-16
c24819 4582 4876 1.58e-16
c24820 5514 410 1.58e-16
c24821 2475 1 4.41e-15
c24822 2751 2384 1.58e-16
c24823 2670 0 2.93e-15
c24824 2558 2542 3.54e-16
c24825 4111 4102 1.88e-16
c24826 3090 1 1.716e-15
c24827 1091 1090 3.94e-16
c24828 4508 837 2.72e-16
c24829 2828 2826 1.6e-16
c24830 2823 2822 2.03e-16
c24831 1690 858 3.15e-16
c24832 1321 1677 3.54e-16
c24833 1343 1327 4.274e-15
c24834 766 25 7.64e-16
c24835 1364 1 1.868e-15
c24836 4217 1 7.08e-16
c24837 1354 0 2.93e-15
c24838 3413 3394 9.83e-16
c24839 3311 827 1.339e-15
c24840 3409 3557 1.58e-16
c24841 4771 1 1.749e-15
c24842 223 175 1.88e-16
c24843 612 2595 2.65e-16
c24844 2294 1 2.054e-15
c24845 4079 857 1.88e-16
c24846 5403 470 3.54e-16
c24847 5396 1 1.672e-15
c24848 2194 1868 1.58e-16
c24849 5444 5449 7.25e-16
c24850 2559 2486 5.5e-16
c24851 2742 2748 1.6e-16
c24852 919 797 3.15e-16
c24853 920 1128 1.58e-16
c24854 3480 4285 1.58e-16
c24855 1708 692 3.15e-16
c24856 1345 1503 5.42e-16
c24857 1321 1491 1.58e-16
c24858 1061 1487 1.96e-16
c24859 4561 4560 6.67e-16
c24860 2316 707 3.15e-16
c24861 2707 717 2.72e-16
c24862 1211 1331 3.92e-16
c24863 2178 692 3.15e-16
c24864 777 782 2.77e-16
c24865 3141 677 1.339e-15
c24866 1 247 1.5625e-14
c24867 3695 837 2.72e-16
c24868 4674 4681 1.81e-16
c24869 4563 4677 1.58e-16
c24870 4580 4689 1.58e-16
c24871 612 2588 2.72e-16
c24872 2272 1 1.716e-15
c24873 632 2194 4.46e-16
c24874 941 939 5.88e-16
c24875 3219 737 3.15e-16
c24876 3801 3807 2.08e-16
c24877 2827 1 2.054e-15
c24878 1862 2342 1.58e-16
c24879 152 30 6.83e-16
c24880 407 404 3.54e-16
c24881 2829 0 8e-16
c24882 4702 410 1.88e-16
c24883 1874 722 1.58e-16
c24884 4092 4095 4.41e-16
c24885 3239 1 1.056e-15
c24886 2418 767 1.58e-16
c24887 2182 692 3.15e-16
c24888 3223 3224 9.1e-16
c24889 1708 1539 1.58e-16
c24890 1706 1533 5.5e-16
c24891 1694 1934 1.58e-16
c24892 617 1363 3.15e-16
c24893 3293 3294 1.35e-16
c24894 687 2291 1.58e-16
c24895 2055 1 3.36e-16
c24896 348 346 7.1e-16
c24897 331 349 1.58e-16
c24898 323 354 1.88e-16
c24899 642 2628 2.22e-16
c24900 2357 1851 3.92e-16
c24901 2361 2362 1.6e-16
c24902 2042 0 2.078e-15
c24903 420 9 6.48e-16
c24904 221 216 1.482e-15
c24905 894 976 1.58e-16
c24906 907 923 3.54e-16
c24907 3321 3705 1.58e-16
c24908 4078 4075 5.5e-16
c24909 4872 0 3.17264e-13
c24910 4600 33 1.88e-16
c24911 2911 2915 1.845e-15
c24912 642 4268 1.58e-16
c24913 3974 25 3.84e-16
c24914 4374 4373 5.65e-16
c24915 4368 3531 1.532e-15
c24916 1327 1639 1.58e-16
c24917 1564 1561 3.01e-16
c24918 1560 1557 6.44e-16
c24919 4174 1 6.76e-16
c24920 5199 207 3.54e-16
c24921 2987 2929 1.58e-16
c24922 822 1584 1.813e-15
c24923 1826 1 6.15e-16
c24924 601 1694 3.15e-16
c24925 726 715 7.23e-16
c24926 718 719 1.6e-16
c24927 1913 1 5.97e-15
c24928 2150 1641 1.96e-16
c24929 1029 677 1.58e-16
c24930 5200 5232 1.58e-16
c24931 792 2408 1.58e-16
c24932 777 19 1.41e-15
c24933 59 426 1.88e-16
c24934 4180 1 6.78e-16
c24935 617 1370 1.339e-15
c24936 4497 4884 1.188e-15
c24937 4152 37 5.71e-16
c24938 4435 4815 1.96e-16
c24939 1868 1869 1.35e-16
c24940 0 514 1.0822e-14
c24941 27 508 1.88e-16
c24942 136 334 1.88e-16
c24943 4567 4242 5.5e-16
c24944 2420 2419 1.6e-16
c24945 2412 2410 2.15e-16
c24946 0 564 1.5696e-14
c24947 3355 3869 1.58e-16
c24948 617 3105 1.58e-16
c24949 2797 1 8.43e-16
c24950 1158 1172 1.96e-16
c24951 3429 4263 1.58e-16
c24952 4793 5239 7.98e-16
c24953 922 918 1.88e-16
c24954 3015 3014 1.6e-16
c24955 3005 3003 1.96e-16
c24956 602 3429 1.58e-16
c24957 601 4260 3.64e-16
c24958 3876 4332 3.92e-16
c24959 4440 4438 2.15e-16
c24960 4448 4447 1.6e-16
c24961 3283 3281 1.6e-16
c24962 3278 3277 2.03e-16
c24963 3944 0 2.0499e-14
c24964 4344 4316 2.64e-16
c24965 1607 1 4.41e-15
c24966 3587 722 1.58e-16
c24967 4915 1 3.3585e-14
c24968 1991 0 6.62e-16
c24969 3387 3671 1.58e-16
c24970 1087 737 6.38e-16
c24971 909 905 3.92e-16
c24972 596 850 2.45e-16
c24973 1236 848 1.45e-16
c24974 2203 0 3.5936e-14
c24975 3752 3734 4.06e-16
c24976 1585 782 3.64e-16
c24977 1376 1374 1.6e-16
c24978 1371 1370 2.03e-16
c24979 4433 4434 9.1e-16
c24980 4571 4580 4.078e-15
c24981 4582 4563 4.312e-15
c24982 2535 2598 1.58e-16
c24983 2557 2586 1.58e-16
c24984 627 978 1.58e-16
c24985 617 963 1.58e-16
c24986 1229 1 3.64e-16
c24987 1916 1914 1.6e-16
c24988 4864 4871 1.96e-16
c24989 1947 1556 1.136e-15
c24990 5291 5280 7.92e-16
c24991 5339 5318 5.87e-16
c24992 3397 3489 1.58e-16
c24993 1 553 1.456e-15
c24994 4580 4779 1.58e-16
c24995 4571 4791 1.58e-16
c24996 5200 5190 1.021e-15
c24997 5104 62 4.44e-16
c24998 4844 468 1.88e-16
c24999 4838 207 1.88e-16
c25000 3029 2549 9.72e-16
c25001 3937 3942 4.33e-16
c25002 3162 0 3.466e-15
c25003 1493 707 1.9e-16
c25004 1159 1160 7.51e-16
c25005 3521 0 1.6491e-14
c25006 3574 747 1.58e-16
c25007 3839 3749 1.58e-16
c25008 3363 2855 1.96e-16
c25009 3034 3143 1.58e-16
c25010 1599 1 6.15e-16
c25011 4779 4791 2.62e-16
c25012 3194 717 1.58e-16
c25013 2072 2093 6.78e-16
c25014 420 419 5.8e-16
c25015 4676 0 2.93e-15
c25016 5198 5194 5.32e-16
c25017 481 482 6.67e-16
c25018 0 219 1.051e-14
c25019 316 303 1.108e-15
c25020 523 565 1.88e-16
c25021 5135 5133 1.167e-15
c25022 4878 178 1.88e-16
c25023 910 2172 5.22e-16
c25024 2195 1 2.471e-15
c25025 3723 3338 1.96e-16
c25026 3769 3767 6.87e-16
c25027 612 3075 1.58e-16
c25028 601 3061 1.84e-16
c25029 1147 1128 1.546e-15
c25030 4238 4237 5.65e-16
c25031 4232 3381 1.532e-15
c25032 3531 692 3.15e-16
c25033 1181 842 3.15e-16
c25034 1646 868 2.72e-16
c25035 1191 1194 1.58e-16
c25036 3330 0 3.3874e-14
c25037 3158 3160 1.862e-15
c25038 3540 3539 2.48e-16
c25039 2535 702 3.15e-16
c25040 1982 1590 1.96e-16
c25041 1983 1976 6.73e-16
c25042 4476 0 6.72e-16
c25043 5072 5114 3.15e-16
c25044 3633 777 2.22e-16
c25045 3616 792 1.813e-15
c25046 3457 3453 1.96e-16
c25047 360 359 6.67e-16
c25048 3566 717 2.65e-16
c25049 3696 3304 2.38e-15
c25050 3693 3691 1.862e-15
c25051 4905 4950 3.036e-15
c25052 4967 4944 1.96e-16
c25053 71 114 1.88e-16
c25054 3693 842 1.58e-16
c25055 5261 149 3.54e-16
c25056 2589 2590 5.65e-16
c25057 596 805 2.45e-16
c25058 612 3018 1.58e-16
c25059 361 1 5.175e-15
c25060 3900 3446 5.5e-16
c25061 3684 868 1.813e-15
c25062 4520 5576 1.96e-16
c25063 2857 2858 2.48e-16
c25064 2545 2554 1.58e-16
c25065 833 0 1.1593e-14
c25066 3160 3159 2.48e-16
c25067 3287 0 6.9481e-14
c25068 4480 4475 1.642e-15
c25069 617 3886 3.15e-16
c25070 3030 2787 1.58e-16
c25071 3030 677 3.15e-16
c25072 3034 662 3.15e-16
c25073 1678 2204 1.532e-15
c25074 2209 2210 5.65e-16
c25075 4452 0 3.6274e-14
c25076 5422 468 1.58e-16
c25077 5191 5188 1.98e-16
c25078 3943 857 6.23e-16
c25079 5560 497 3.54e-16
c25080 5476 5479 1.18e-15
c25081 4770 5200 1.53e-15
c25082 2882 1 3.016e-15
c25083 921 842 3.15e-16
c25084 3663 0 6.72e-16
c25085 2663 2654 3.92e-16
c25086 1327 1367 1.58e-16
c25087 4068 1 2.259e-15
c25088 2424 812 1.75e-16
c25089 4815 0 3.466e-15
c25090 2730 3228 1.58e-16
c25091 3158 702 1.58e-16
c25092 2068 2066 3.25e-16
c25093 4580 4724 3.92e-16
c25094 4708 4333 4.9e-16
c25095 3411 3401 5.5e-16
c25096 3409 3386 1.58e-16
c25097 3393 3407 3.92e-16
c25098 592 589 1.96e-16
c25099 2344 0 3.466e-15
c25100 777 1555 2.4e-16
c25101 339 333 3.84e-16
c25102 747 1868 1.58e-16
c25103 5452 5457 3.84e-16
c25104 5450 5489 3.18e-16
c25105 601 2541 3.15e-16
c25106 2545 2350 5.5e-16
c25107 2663 2664 1.6e-16
c25108 2654 2656 2.15e-16
c25109 1345 880 1.58e-16
c25110 1343 877 1.58e-16
c25111 672 1 4.1542e-14
c25112 2954 2949 1.291e-15
c25113 2951 2959 3.54e-16
c25114 3882 3582 5.88e-16
c25115 3876 3588 1.58e-16
c25116 2435 807 3.79e-16
c25117 1784 1786 1.862e-15
c25118 1397 1403 1.418e-15
c25119 3809 1 4.239e-15
c25120 4056 19 7.35e-16
c25121 2545 2717 1.58e-16
c25122 1013 0 1.4198e-14
c25123 3048 3105 3.92e-16
c25124 2029 2054 7.65e-16
c25125 1091 0 7.4292e-14
c25126 1732 1733 1.35e-16
c25127 19 343 3.2e-16
c25128 210 205 1.059e-15
c25129 201 204 3.54e-16
c25130 192 187 1.482e-15
c25131 2385 2379 1.6e-16
c25132 1862 2376 2.386e-15
c25133 1868 2384 1.136e-15
c25134 1879 2359 1.58e-16
c25135 3168 677 1.58e-16
c25136 4905 4904 4.61e-16
c25137 4903 4928 7.1e-16
c25138 2274 2276 2.15e-16
c25139 617 2223 1.58e-16
c25140 166 175 1.58e-16
c25141 2299 1 5.97e-15
c25142 2661 2652 3.46e-16
c25143 890 677 3.15e-16
c25144 907 1037 3.92e-16
c25145 657 661 2.19e-16
c25146 4571 4881 1.58e-16
c25147 4582 4893 1.58e-16
c25148 4685 468 1.88e-16
c25149 2136 2139 3.54e-16
c25150 4124 4131 7.81e-16
c25151 3273 1 1.056e-15
c25152 1538 752 7.38e-16
c25153 1326 1324 1.041e-15
c25154 2340 732 1.58e-16
c25155 657 1386 5.73e-16
c25156 3242 1 4.41e-15
c25157 3145 3147 1.6e-16
c25158 3141 3142 2.03e-16
c25159 4667 4660 1.96e-16
c25160 4276 4669 1.914e-15
c25161 2790 797 1.58e-16
c25162 4404 0 3.3608e-14
c25163 2705 722 1.58e-16
c25164 5350 354 9.1e-16
c25165 5387 265 3.54e-16
c25166 4549 5013 1.878e-15
c25167 3328 868 1.58e-16
c25168 4788 1 1.749e-15
c25169 4567 4486 1.58e-16
c25170 4861 4863 4.93e-16
c25171 5298 5297 1.6e-16
c25172 5177 5157 1.58e-16
c25173 118 120 6.01e-16
c25174 601 2597 4.81e-16
c25175 612 2214 3.79e-16
c25176 2465 2463 1.6e-16
c25177 2460 2459 2.03e-16
c25178 4502 837 2.4e-16
c25179 1239 1236 9.8e-16
c25180 1188 1189 1.21e-16
c25181 4844 64 1.88e-16
c25182 593 1 3.79e-16
c25183 1403 1404 1.35e-16
c25184 542 0 1.97336e-13
c25185 537 27 1.88e-16
c25186 1846 1454 1.96e-16
c25187 1847 1840 6.73e-16
c25188 3030 3241 1.96e-16
c25189 2172 707 4.48e-16
c25190 1710 1 2.86e-16
c25191 792 1141 1.35e-16
c25192 1689 0 4.3757e-14
c25193 1 178 3.36e-15
c25194 4691 4699 1.81e-16
c25195 4563 4694 1.58e-16
c25196 4580 4706 1.58e-16
c25197 5074 91 7.37e-16
c25198 2452 2447 1.642e-15
c25199 2298 1 8.43e-16
c25200 657 2172 3.15e-16
c25201 0 188 1.5696e-14
c25202 3834 3835 1.08e-15
c25203 3831 3775 9.34e-16
c25204 2178 2181 1.96e-16
c25205 1188 837 1.58e-16
c25206 894 797 3.15e-16
c25207 890 1128 3.54e-16
c25208 909 1149 1.58e-16
c25209 2845 0 6.72e-16
c25210 919 978 1.58e-16
c25211 4175 4182 2.45e-16
c25212 1061 1486 1.58e-16
c25213 4600 5564 5.5e-16
c25214 3622 4458 5.66e-16
c25215 4464 4455 3.92e-16
c25216 1902 782 1.75e-16
c25217 3879 1 8.766e-15
c25218 1659 1674 1.96e-16
c25219 972 0 6.29e-16
c25220 4546 4553 3.96e-16
c25221 1684 1550 5.5e-16
c25222 1694 1939 1.58e-16
c25223 627 1397 2.22e-16
c25224 910 0 4.47893e-13
c25225 687 2311 1.58e-16
c25226 1935 1550 1.96e-16
c25227 662 654 1.74e-16
c25228 2182 2181 1.357e-15
c25229 5300 352 7.94e-16
c25230 278 1 4.22e-16
c25231 4313 647 4.81e-16
c25232 3463 672 1.58e-16
c25233 909 963 3.54e-16
c25234 281 0 1.27746e-13
c25235 4086 4079 2.45e-16
c25236 1602 807 2.65e-16
c25237 1405 1406 2.48e-16
c25238 642 4288 1.58e-16
c25239 2559 2650 3.92e-16
c25240 4047 2189 2.697e-15
c25241 687 2289 1.58e-16
c25242 1539 1922 7.84e-16
c25243 632 627 2.77e-16
c25244 4407 747 1.58e-16
c25245 4902 4897 1.102e-15
c25246 1835 1 1.716e-15
c25247 617 1694 3.15e-16
c25248 636 625 7.23e-16
c25249 3387 3140 1.58e-16
c25250 2455 1 1.056e-15
c25251 747 1890 2.72e-16
c25252 217 0 1.5696e-14
c25253 3869 858 3.15e-16
c25254 3393 852 4.03e-16
c25255 3983 3990 2.45e-16
c25256 3047 1 2.471e-15
c25257 1061 722 3.15e-16
c25258 1510 732 2.72e-16
c25259 1071 1074 1.58e-16
c25260 632 993 1.58e-16
c25261 2722 2721 2.48e-16
c25262 719 26 2.65e-15
c25263 372 0 6.224e-15
c25264 4350 4351 1.35e-16
c25265 3707 3886 1.58e-16
c25266 4543 4540 5.5e-16
c25267 1987 842 2.33e-16
c25268 3030 3206 1.58e-16
c25269 1644 1 5.808e-15
c25270 625 626 6.67e-16
c25271 1646 0 3.466e-15
c25272 3409 692 4.46e-16
c25273 4567 4259 5.5e-16
c25274 4759 439 1.88e-16
c25275 595 2536 9.02e-16
c25276 891 917 1.067e-15
c25277 3972 3973 7.45e-16
c25278 3980 3982 2.239e-15
c25279 5366 294 7.62e-16
c25280 986 990 2.03e-16
c25281 361 363 1.88e-16
c25282 3446 4251 1.58e-16
c25283 3429 4268 2.386e-15
c25284 4277 4271 1.6e-16
c25285 5436 5425 1.96e-16
c25286 160 59 1.88e-16
c25287 1472 1483 1.96e-16
c25288 3987 1 6.78e-16
c25289 601 3429 3.15e-16
c25290 617 4260 7.68e-16
c25291 627 3435 1.58e-16
c25292 3900 4349 3.92e-16
c25293 2395 767 5.03e-16
c25294 2781 3275 1.96e-16
c25295 2293 1783 1.96e-16
c25296 3491 3489 2.15e-16
c25297 3499 3498 1.6e-16
c25298 3684 0 6.9481e-14
c25299 165 334 1.88e-16
c25300 14 20 1.372e-15
c25301 3387 3676 1.58e-16
c25302 3411 3688 5.42e-16
c25303 3393 3293 1.58e-16
c25304 921 925 5.35e-16
c25305 920 924 3.54e-16
c25306 1024 1025 7.51e-16
c25307 4600 526 1.88e-16
c25308 1136 767 3.57e-16
c25309 3898 4319 1.58e-16
c25310 3876 4331 1.58e-16
c25311 4685 64 1.88e-16
c25312 2662 0 6.9481e-14
c25313 2559 2615 5.42e-16
c25314 2535 2603 1.58e-16
c25315 884 0 1.4741e-14
c25316 691 1 4.03e-16
c25317 3926 37 1.88e-16
c25318 3935 25 4.68e-16
c25319 4352 4351 2.03e-16
c25320 4357 4355 1.6e-16
c25321 4347 1 1.056e-15
c25322 1708 1691 3.62e-16
c25323 1706 1698 4.63e-16
c25324 1443 0 1.4092e-14
c25325 477 484 7.76e-16
c25326 3484 3485 9.1e-16
c25327 3411 3123 1.58e-16
c25328 657 2270 2.4e-16
c25329 3364 3363 2.49e-16
c25330 1743 2223 1.58e-16
c25331 1658 2118 5.71e-16
c25332 1012 993 1.546e-15
c25333 4580 4796 1.58e-16
c25334 4571 4808 1.58e-16
c25335 91 89 6.01e-16
c25336 3918 3950 6.32e-16
c25337 4455 782 1.832e-15
c25338 2969 1 2.397e-15
c25339 922 1100 3.92e-16
c25340 1553 1551 1.6e-16
c25341 1343 1419 3.92e-16
c25342 2995 2518 5.5e-16
c25343 3701 3673 2.64e-16
c25344 4142 1 6.76e-16
c25345 2654 662 1.832e-15
c25346 4863 4486 2.48e-16
c25347 4316 1 4.442e-15
c25348 2118 2070 3.15e-16
c25349 1608 1 1.716e-15
c25350 1 351 4.92e-16
c25351 217 219 1.58e-16
c25352 5249 5227 1.74e-16
c25353 5234 5226 3.54e-16
c25354 3168 3174 1.418e-15
c25355 3555 3557 1.862e-15
c25356 4693 0 2.93e-15
c25357 3185 3157 2.64e-16
c25358 4563 4564 1.239e-15
c25359 4810 352 1.88e-16
c25360 3338 3855 1.885e-15
c25361 627 3075 1.58e-16
c25362 1167 797 4.98e-16
c25363 59 513 1.88e-16
c25364 5303 5311 9.34e-16
c25365 5388 5310 1.58e-16
c25366 687 689 5.59e-16
c25367 74 73 7.08e-16
c25368 65 60 1.059e-15
c25369 2983 2982 1.08e-15
c25370 687 3497 1.813e-15
c25371 3886 4485 4.63e-16
c25372 3839 3836 7.46e-16
c25373 4120 37 5.71e-16
c25374 707 0 2.8008e-13
c25375 2126 2125 1.6e-16
c25376 657 0 2.86553e-13
c25377 1601 1590 1.58e-16
c25378 305 204 1.88e-16
c25379 5106 5074 1.58e-16
c25380 3185 717 3.79e-16
c25381 4940 4936 3.82e-16
c25382 5071 1 1.23e-16
c25383 4954 4967 3.92e-16
c25384 4903 4905 1.96e-16
c25385 3865 3869 1.96e-16
c25386 3393 3409 4.274e-15
c25387 3397 3637 1.58e-16
c25388 3722 3355 1.58e-16
c25389 3328 0 1.6491e-14
c25390 2178 2457 1.96e-16
c25391 1355 1364 3.92e-16
c25392 1116 1123 7.95e-16
c25393 4526 858 1.84e-16
c25394 4640 5459 6.9e-16
c25395 2545 2169 1.58e-16
c25396 3775 0 4.4655e-14
c25397 1766 647 2.33e-16
c25398 2009 842 1.9e-16
c25399 1619 1161 1.96e-16
c25400 1620 1613 6.73e-16
c25401 1690 1437 1.58e-16
c25402 3094 3090 1.96e-16
c25403 1887 1499 4.97e-16
c25404 3367 852 1.58e-16
c25405 781 779 5.88e-16
c25406 3393 3621 1.96e-16
c25407 13 218 1.88e-16
c25408 4770 439 1.88e-16
c25409 4861 120 1.88e-16
c25410 2182 2457 4.63e-16
c25411 642 3048 3.58e-16
c25412 1321 672 3.15e-16
c25413 1345 647 3.15e-16
c25414 1365 1364 1.6e-16
c25415 2541 2544 1.96e-16
c25416 1343 1384 1.58e-16
c25417 629 26 2.65e-15
c25418 4877 842 1.23e-16
c25419 1871 1883 2.32e-16
c25420 642 1743 1.813e-15
c25421 3452 0 3.6368e-14
c25422 3034 2781 5.5e-16
c25423 1802 1414 4.97e-16
c25424 4760 4384 3.92e-16
c25425 4772 4771 1.6e-16
c25426 4832 0 3.466e-15
c25427 2668 692 2.33e-16
c25428 1753 0 6.62e-16
c25429 534 536 2.84e-16
c25430 1 455 3.0375e-14
c25431 4580 4741 3.92e-16
c25432 3387 3433 1.58e-16
c25433 632 2220 1.75e-16
c25434 2362 1 2.054e-15
c25435 0 441 5.5238e-14
c25436 2364 0 8e-16
c25437 3628 767 1.58e-16
c25438 2917 1 2.53e-16
c25439 890 1202 1.96e-16
c25440 5422 5424 1.062e-15
c25441 5400 5262 3.54e-16
c25442 617 2541 3.15e-16
c25443 922 692 5.14e-16
c25444 921 1023 1.58e-16
c25445 2702 2703 1.35e-16
c25446 1181 1184 6.13e-16
c25447 632 919 3.15e-16
c25448 4310 3469 1.136e-15
c25449 3886 4450 1.58e-16
c25450 3898 3599 5.5e-16
c25451 3900 3605 1.58e-16
c25452 3667 4485 1.96e-16
c25453 2634 672 1.58e-16
c25454 2545 2722 1.58e-16
c25455 1690 2002 1.58e-16
c25456 1963 1954 3.46e-16
c25457 5032 5094 6.67e-16
c25458 158 175 1.138e-15
c25459 5356 265 1.58e-16
c25460 3437 3439 2.03e-16
c25461 617 2243 1.58e-16
c25462 2022 0 5.5809e-14
c25463 88 19 3.84e-16
c25464 91 33 1.88e-16
c25465 2716 1 1.056e-15
c25466 3731 3729 1.082e-15
c25467 3289 1 9.28e-16
c25468 1421 1423 1.862e-15
c25469 986 996 1.418e-15
c25470 642 909 3.15e-16
c25471 4504 842 1.339e-15
c25472 1851 722 2.33e-16
c25473 1257 1255 1.186e-15
c25474 657 1795 2.65e-16
c25475 3651 1 1.868e-15
c25476 1382 1 9.28e-16
c25477 4424 0 1.4092e-14
c25478 2725 722 1.58e-16
c25479 262 253 1.58e-16
c25480 246 252 3.84e-16
c25481 3419 3421 1.862e-15
c25482 3018 3021 1.576e-15
c25483 2838 842 2.33e-16
c25484 2276 2272 1.96e-16
c25485 617 2221 1.339e-15
c25486 1905 1 5.808e-15
c25487 1907 0 3.466e-15
c25488 4805 1 1.749e-15
c25489 777 1522 5.73e-16
c25490 1038 702 1.05e-15
c25491 4567 4503 1.58e-16
c25492 4810 294 1.88e-16
c25493 4719 352 1.88e-16
c25494 627 2214 1.813e-15
c25495 1964 2457 1.96e-16
c25496 2172 1879 5.5e-16
c25497 2833 2824 3.92e-16
c25498 3092 0 3.3874e-14
c25499 922 1158 1.58e-16
c25500 4304 4300 1.96e-16
c25501 3001 2492 3.92e-16
c25502 2518 2527 1.6e-16
c25503 1343 1071 1.58e-16
c25504 392 393 1.079e-15
c25505 397 391 3.84e-16
c25506 797 1 3.1284e-14
c25507 2703 722 1.339e-15
c25508 1465 1454 1.58e-16
c25509 3394 3417 1.003e-15
c25510 4223 25 1.88e-16
c25511 4238 0 6.72e-16
c25512 3330 3328 1.862e-15
c25513 687 2316 2.22e-16
c25514 1896 1891 1.642e-15
c25515 9 368 5.8e-16
c25516 3691 842 1.339e-15
c25517 3370 3371 3.01e-16
c25518 822 2442 1.58e-16
c25519 0 332 4.5547e-14
c25520 3693 3411 1.58e-16
c25521 4520 4521 1.35e-16
c25522 1201 1202 1.238e-15
c25523 1200 827 6.48e-16
c25524 1192 868 1.58e-16
c25525 883 1143 3.54e-16
c25526 894 1164 1.58e-16
c25527 129 128 1.482e-15
c25528 5474 5412 6.67e-16
c25529 5356 5324 1.75e-16
c25530 1505 737 2.33e-16
c25531 1061 1491 1.58e-16
c25532 3022 0 6.9483e-14
c25533 3633 4455 1.58e-16
c25534 2436 782 3.64e-16
c25535 1706 1420 1.58e-16
c25536 1768 1386 2.48e-16
c25537 4845 4856 1.96e-16
c25538 3030 2532 1.58e-16
c25539 1086 1 4.044e-15
c25540 1526 0 6.62e-16
c25541 37 262 1.88e-16
c25542 305 175 1.88e-16
c25543 657 3122 2.4e-16
c25544 4992 4991 1.353e-15
c25545 407 426 1.88e-16
c25546 894 978 3.54e-16
c25547 1593 812 1.58e-16
c25548 1151 807 3.79e-16
c25549 2958 2959 5.07e-16
c25550 1281 1300 1.54e-16
c25551 2344 707 1.9e-16
c25552 1345 1656 5.42e-16
c25553 1321 1644 1.58e-16
c25554 1550 1934 1.58e-16
c25555 1690 1765 1.96e-16
c25556 419 424 1.482e-15
c25557 4978 1 3.56e-15
c25558 1861 1 8.43e-16
c25559 736 734 5.88e-16
c25560 3411 3157 1.58e-16
c25561 3293 3675 2.48e-16
c25562 4910 0 5.9239e-14
c25563 2471 1 9.28e-16
c25564 1043 677 3.57e-16
c25565 1023 1036 1.58e-16
c25566 390 19 3.84e-16
c25567 3338 827 1.58e-16
c25568 5051 5274 9.75e-16
c25569 5044 5045 3.18e-16
c25570 2441 0 3.5724e-14
c25571 5537 5535 5.25e-16
c25572 1287 1275 6.73e-16
c25573 1284 1243 7.55e-16
c25574 1280 1226 1.96e-16
c25575 1965 797 3.64e-16
c25576 1116 1559 7.84e-16
c25577 1226 0 6.0838e-14
c25578 1125 1 3.06e-16
c25579 3713 1 2.054e-15
c25580 1981 858 1.58e-16
c25581 1827 1818 3.46e-16
c25582 4452 4832 1.96e-16
c25583 3046 3223 1.58e-16
c25584 3030 3211 1.58e-16
c25585 2154 2151 5.5e-16
c25586 1641 1694 1.58e-16
c25587 77 71 5.8e-16
c25588 17 18 1.58e-16
c25589 19 37 2.8387e-14
c25590 0 34 1.4515e-14
c25591 28 33 6.38e-16
c25592 3411 717 3.58e-16
c25593 4567 4276 5.5e-16
c25594 2425 2436 1.96e-16
c25595 3480 3089 1.136e-15
c25596 5355 0 3.6193e-14
c25597 996 1003 7.95e-16
c25598 4390 722 1.58e-16
c25599 2726 2724 1.6e-16
c25600 2721 2720 2.03e-16
c25601 910 884 9.54e-16
c25602 5375 5360 6.67e-16
c25603 920 964 3.98e-16
c25604 632 957 1.58e-16
c25605 617 3429 3.15e-16
c25606 2882 2896 2.217e-15
c25607 2557 2803 3.92e-16
c25608 4713 4711 2.15e-16
c25609 4709 4720 1.96e-16
c25610 822 1612 2.72e-16
c25611 15 563 3.92e-16
c25612 4915 410 1.88e-16
c25613 2018 1 1.056e-15
c25614 3857 3859 2.61e-16
c25615 3853 3854 1.6e-16
c25616 4793 5232 4.06e-16
c25617 239 1 5.62e-16
c25618 5326 5333 3.54e-16
c25619 5324 5364 1.062e-15
c25620 2793 0 1.4092e-14
c25621 2231 0 6.9484e-14
c25622 4217 857 1.88e-16
c25623 4719 294 7.67e-16
c25624 1413 971 1.96e-16
c25625 1136 1134 1.931e-15
c25626 3876 4336 1.58e-16
c25627 3900 4348 5.42e-16
c25628 2559 2620 1.58e-16
c25629 2566 2567 1.35e-16
c25630 3959 19 3.45e-16
c25631 3531 4349 1.96e-16
c25632 1331 1161 1.58e-16
c25633 4363 1 9.28e-16
c25634 3107 3118 1.96e-16
c25635 3650 822 1.813e-15
c25636 3106 3134 2.64e-16
c25637 2987 2907 1.58e-16
c25638 4881 4888 1.96e-16
c25639 3048 732 3.58e-16
c25640 1 324 4.92e-16
c25641 3642 3654 2.32e-16
c25642 4580 4813 1.58e-16
c25643 4571 4825 1.58e-16
c25644 5522 1 1.672e-15
c25645 2607 0 6.72e-16
c25646 2520 2512 2.15e-16
c25647 1998 2004 1.545e-15
c25648 642 3072 5.73e-16
c25649 1381 1372 3.92e-16
c25650 952 1375 5.66e-16
c25651 777 2406 2.4e-16
c25652 3002 1 4.03e-16
c25653 1061 1064 6.13e-16
c25654 2955 0 2.9272e-14
c25655 2545 2390 1.58e-16
c25656 2557 762 3.15e-16
c25657 1706 1680 1.58e-16
c25658 1684 1683 1.58e-16
c25659 1224 0 2.8146e-14
c25660 4534 4532 1.6e-16
c25661 2474 827 7.38e-16
c25662 1721 1718 5.5e-16
c25663 4796 4808 2.62e-16
c25664 2685 732 5.73e-16
c25665 1634 1 8.43e-16
c25666 15 535 5.8e-16
c25667 3387 3502 3.92e-16
c25668 1879 0 6.9481e-14
c25669 0 565 1.56098e-13
c25670 19 548 3.45e-16
c25671 3957 3951 7.45e-16
c25672 4691 497 1.88e-16
c25673 2196 2320 5.42e-16
c25674 627 3095 1.58e-16
c25675 2557 2401 5.5e-16
c25676 2688 2697 3.92e-16
c25677 2316 2683 1.58e-16
c25678 4250 4251 2.48e-16
c25679 2214 2220 1.418e-15
c25680 2231 2203 2.64e-16
c25681 2041 2990 2.12e-16
c25682 1462 1459 3.01e-16
c25683 1458 1455 6.44e-16
c25684 2389 752 7.38e-16
c25685 1721 1728 6.73e-16
c25686 1319 1703 2.79e-16
c25687 3188 3186 1.6e-16
c25688 3673 1 4.41e-15
c25689 1601 1999 4.36e-16
c25690 1997 1990 1.96e-16
c25691 1760 1755 1.642e-15
c25692 291 334 1.88e-16
c25693 4507 0 6.62e-16
c25694 5148 5010 8.12e-16
c25695 565 564 1.88e-16
c25696 3034 852 7.99e-16
c25697 3046 858 1.58e-16
c25698 909 732 3.15e-16
c25699 3397 3642 1.58e-16
c25700 1085 722 5.74e-16
c25701 3781 858 1.58e-16
c25702 5286 5299 1.138e-15
c25703 5262 5239 1.58e-16
c25704 1437 702 5.73e-16
c25705 595 600 2.19e-16
c25706 2194 2474 3.92e-16
c25707 107 105 1.257e-15
c25708 4053 4047 7.45e-16
c25709 4543 858 1.58e-16
c25710 3886 3469 1.58e-16
c25711 1725 1315 1.96e-16
c25712 1720 1318 1.96e-16
c25713 601 980 1.58e-16
c25714 854 0 7.709e-15
c25715 1166 1161 1.58e-16
c25716 1706 1454 1.58e-16
c25717 355 354 3.84e-16
c25718 81 0 1.4803e-14
c25719 2866 2861 1.642e-15
c25720 2318 2317 1.6e-16
c25721 642 2257 1.58e-16
c25722 2223 2222 2.48e-16
c25723 2552 0 5.5167e-14
c25724 4657 4658 9.93e-16
c25725 2178 2456 1.58e-16
c25726 396 1 9.8e-16
c25727 2194 1749 1.58e-16
c25728 397 0 1.62163e-13
c25729 4317 4328 1.96e-16
c25730 4804 5270 5.5e-16
c25731 2279 647 1.09e-16
c25732 3504 1 1.716e-15
c25733 3694 0 6.62e-16
c25734 1918 767 7.38e-16
c25735 2713 2708 1.642e-15
c25736 1192 0 1.8851e-14
c25737 4117 1 7.71e-16
c25738 2474 812 1.58e-16
c25739 1778 1 1.868e-15
c25740 4849 0 3.466e-15
c25741 3254 2736 1.96e-16
c25742 2662 707 1.58e-16
c25743 1768 0 2.93e-15
c25744 5209 5158 1.191e-15
c25745 3393 3055 1.58e-16
c25746 3411 3450 5.42e-16
c25747 3387 3438 1.58e-16
c25748 632 2629 3.64e-16
c25749 2196 1936 1.58e-16
c25750 2182 2456 1.58e-16
c25751 556 553 6.38e-16
c25752 2392 2394 2.03e-16
c25753 1457 692 1.58e-16
c25754 883 1217 3.92e-16
c25755 907 858 1.58e-16
c25756 890 1216 1.88e-16
c25757 5481 5508 9.6e-16
c25758 5506 5452 9.34e-16
c25759 5503 5492 3.92e-16
c25760 4804 5263 2.137e-15
c25761 2871 2486 1.96e-16
c25762 3313 1 5.808e-15
c25763 1456 1016 4.97e-16
c25764 4088 1 5.1e-16
c25765 5419 528 5.93e-16
c25766 2282 662 3.15e-16
c25767 2849 2821 2.64e-16
c25768 3836 1 1.81e-16
c25769 1698 1687 4.097e-15
c25770 4069 19 9.67e-16
c25771 1691 1701 5.8e-16
c25772 4378 4761 4.97e-16
c25773 2730 3252 1.96e-16
c25774 2736 3247 1.96e-16
c25775 3182 692 1.09e-16
c25776 2069 2071 9.16e-16
c25777 642 2622 2.72e-16
c25778 1969 1968 9.1e-16
c25779 777 1559 1.58e-16
c25780 330 331 6.67e-16
c25781 4982 4977 3.73e-16
c25782 2732 1 9.28e-16
c25783 642 2545 7.99e-16
c25784 894 1052 3.92e-16
c25785 909 1051 1.88e-16
c25786 883 1044 1.58e-16
c25787 5262 5173 1.58e-16
c25788 3302 1 6.15e-16
c25789 1613 827 1.84e-16
c25790 1321 797 4.48e-16
c25791 4872 4922 3.41e-16
c25792 632 894 3.15e-16
c25793 3281 792 2.72e-16
c25794 647 19 1.676e-15
c25795 1845 737 1.58e-16
c25796 3270 1 5.97e-15
c25797 1600 1591 3.46e-16
c25798 809 0 7.709e-15
c25799 4684 4677 1.96e-16
c25800 4293 4686 1.914e-15
c25801 1395 1 6.15e-16
c25802 1652 1647 1.642e-15
c25803 2832 858 1.58e-16
c25804 3393 3591 1.58e-16
c25805 3409 3208 1.58e-16
c25806 4822 1 1.749e-15
c25807 2522 1 2.48e-16
c25808 2200 2195 9.6e-16
c25809 762 1533 3.79e-16
c25810 1066 1067 1.238e-15
c25811 1057 717 1.58e-16
c25812 3748 3745 3.92e-16
c25813 4674 1 1.4793e-14
c25814 4922 0 2.37076e-13
c25815 4838 497 1.88e-16
c25816 2663 2271 1.96e-16
c25817 3876 807 3.15e-16
c25818 910 3022 3.45e-16
c25819 1542 752 1.832e-15
c25820 2756 2754 1.862e-15
c25821 1607 837 1.58e-16
c25822 1136 1589 1.96e-16
c25823 1321 1086 1.58e-16
c25824 1327 1076 5.88e-16
c25825 3056 3058 1.862e-15
c25826 2529 2532 1.576e-15
c25827 1164 1 2.972e-15
c25828 1465 1863 4.36e-16
c25829 1861 1854 1.96e-16
c25830 5007 5020 9.41e-16
c25831 1165 0 6.29e-16
c25832 792 1128 1.05e-15
c25833 3048 3258 3.92e-16
c25834 3606 3609 6.44e-16
c25835 2656 2271 1.96e-16
c25836 2470 2461 3.92e-16
c25837 1953 2464 5.66e-16
c25838 1964 2456 1.58e-16
c25839 687 2172 3.15e-16
c25840 767 759 1.74e-16
c25841 851 850 6.67e-16
c25842 0 478 1.5696e-14
c25843 5246 238 5.93e-16
c25844 5160 236 7.46e-16
c25845 2178 2219 1.96e-16
c25846 1209 842 8.3e-16
c25847 106 15 6.58e-16
c25848 105 1 3.6e-16
c25849 99 0 9.795e-15
c25850 1499 752 1.58e-16
c25851 1343 1342 1.009e-15
c25852 1327 1332 8.56e-16
c25853 4048 1 2.3688e-14
c25854 3633 4475 2.38e-15
c25855 1930 782 3.15e-16
c25856 978 1 1.56e-15
c25857 87 85 7.1e-16
c25858 3046 2566 1.58e-16
c25859 3607 3609 2.03e-16
c25860 5032 5029 3.54e-16
c25861 2544 2175 1.176e-15
c25862 2182 2219 4.63e-16
c25863 3830 3820 1.96e-16
c25864 3702 3693 3.92e-16
c25865 4111 4113 1.06e-16
c25866 2554 2555 1.736e-15
c25867 1613 812 1.58e-16
c25868 657 3452 5.73e-16
c25869 3875 1 2.259e-15
c25870 4023 37 1.88e-16
c25871 2154 858 1.58e-16
c25872 764 0 7.709e-15
c25873 2611 3129 2.38e-15
c25874 1948 1942 1.6e-16
c25875 1550 1939 2.386e-15
c25876 1706 1782 3.92e-16
c25877 5010 4946 1.58e-16
c25878 3571 762 5.73e-16
c25879 5277 5385 1.58e-16
c25880 646 644 5.88e-16
c25881 271 0 2.87e-16
c25882 268 30 6.83e-16
c25883 3387 3168 5.5e-16
c25884 2484 1 6.15e-16
c25885 4068 857 1.88e-16
c25886 3900 767 3.15e-16
c25887 1270 1291 3.04e-16
c25888 920 1145 3.92e-16
c25889 921 1144 2.54e-16
c25890 1584 797 3.15e-16
c25891 1121 1571 1.58e-16
c25892 1139 1 3.06e-16
c25893 2527 858 7.12e-16
c25894 1833 1832 9.1e-16
c25895 5039 180 1.76e-16
c25896 3241 737 1.58e-16
c25897 1837 0 3.3874e-14
c25898 3409 3536 3.92e-16
c25899 929 889 3.84e-16
c25900 948 936 7.81e-16
c25901 4567 4293 5.5e-16
c25902 5069 91 5.5e-16
c25903 143 25 7.06e-16
c25904 5444 5445 8.03e-16
c25905 542 565 1.88e-16
c25906 1498 1046 1.96e-16
c25907 1493 1056 1.96e-16
c25908 3898 3882 4.274e-15
c25909 3876 4556 3.54e-16
c25910 2918 2928 1.668e-15
c25911 2535 2820 3.92e-16
c25912 3134 3129 1.642e-15
c25913 3034 3020 1.58e-16
c25914 2611 647 3.15e-16
c25915 5185 5184 1.6e-16
c25916 340 349 1.58e-16
c25917 5162 236 3.54e-16
c25918 2363 2361 1.6e-16
c25919 2358 2357 2.03e-16
c25920 647 637 6.38e-16
c25921 5388 5385 7.46e-16
c25922 642 3109 1.58e-16
c25923 1406 647 1.58e-16
c25924 438 1 4.92e-16
c25925 78 247 1.88e-16
c25926 4855 1 3.1272e-14
c25927 2633 2265 1.96e-16
c25928 4634 0 4.72366e-13
c25929 4259 3418 1.136e-15
c25930 3900 4353 1.58e-16
c25931 2916 2915 8.03e-16
c25932 2196 662 3.15e-16
c25933 1744 1352 1.96e-16
c25934 901 0 5.1519e-14
c25935 2747 2356 1.136e-15
c25936 1221 1253 1.014e-15
c25937 822 1606 2.4e-16
c25938 4376 1 6.15e-16
c25939 4544 0 6.72e-16
c25940 1684 1730 1.58e-16
c25941 1706 1718 1.58e-16
c25942 192 194 1.257e-15
c25943 2350 2345 1.642e-15
c25944 5167 296 5.93e-16
c25945 2150 2152 1.6e-16
c25946 1 45 1.65e-15
c25947 407 513 1.88e-16
c25948 281 565 1.88e-16
c25949 3411 842 3.15e-16
c25950 4580 4830 1.58e-16
c25951 4571 4842 1.58e-16
c25952 812 828 1.621e-15
c25953 642 3481 2.65e-16
c25954 632 3066 1.58e-16
c25955 3195 0 6.62e-16
c25956 1253 1262 1.96e-16
c25957 3531 4348 1.58e-16
c25958 3520 4356 5.66e-16
c25959 4362 4353 3.92e-16
c25960 3622 797 1.75e-16
c25961 4702 5333 7.87e-16
c25962 1684 807 3.15e-16
c25963 2535 777 3.15e-16
c25964 3574 1 5.808e-15
c25965 1708 1315 1.58e-16
c25966 2545 2541 4.431e-15
c25967 3013 3017 1.96e-16
c25968 627 1385 2.4e-16
c25969 3024 2855 1.58e-16
c25970 3030 2849 5.88e-16
c25971 3134 647 1.58e-16
c25972 4152 0 2.0707e-14
c25973 4880 4503 2.48e-16
c25974 3305 807 2.65e-16
c25975 4480 0 6.8832e-14
c25976 3279 3291 2.32e-16
c25977 3220 732 2.65e-16
c25978 3034 2668 1.58e-16
c25979 1801 0 1.6491e-14
c25980 1 504 4.22e-16
c25981 3585 3583 1.6e-16
c25982 19 523 3.84e-16
c25983 2415 2412 3.01e-16
c25984 2411 2408 6.44e-16
c25985 2196 2325 1.58e-16
c25986 2178 1800 1.58e-16
c25987 2237 2238 1.35e-16
c25988 596 852 1.96e-16
c25989 59 50 1.58e-16
c25990 2873 0 5.5809e-14
c25991 2688 2316 1.58e-16
c25992 920 752 3.69e-16
c25993 1321 1435 1.58e-16
c25994 1343 1423 1.58e-16
c25995 4159 4158 5.5e-16
c25996 3882 4518 1.58e-16
c25997 3004 3001 6.71e-16
c25998 1812 1806 1.6e-16
c25999 2535 2785 1.58e-16
c26000 3941 1 7.71e-16
c26001 4439 4436 6.44e-16
c26002 4443 4440 3.01e-16
c26003 595 1718 1.58e-16
c26004 1610 0 3.3846e-14
c26005 687 0 2.85914e-13
c26006 2557 722 4.46e-16
c26007 2545 732 7.99e-16
c26008 2233 1 9.28e-16
c26009 1694 1884 4.63e-16
c26010 19 317 8.4e-16
c26011 4580 3873 1.58e-16
c26012 2182 1800 1.58e-16
c26013 2325 2334 3.92e-16
c26014 2328 1817 5.66e-16
c26015 1828 2320 1.58e-16
c26016 795 794 1.6e-16
c26017 4838 5079 5.91e-16
c26018 3446 3055 1.136e-15
c26019 2686 2697 1.96e-16
c26020 2595 1 1.868e-15
c26021 1726 1732 1.418e-15
c26022 894 895 6.91e-16
c26023 3710 3708 1.862e-15
c26024 1846 702 2.65e-16
c26025 1345 868 3.58e-16
c26026 73 70 1.099e-15
c26027 2984 2990 6.23e-16
c26028 4520 4580 1.58e-16
c26029 3839 3830 8.15e-16
c26030 1166 1636 4.36e-16
c26031 1634 1627 1.96e-16
c26032 617 980 5.74e-16
c26033 2668 3176 2.48e-16
c26034 1684 1471 1.58e-16
c26035 1690 1465 5.88e-16
c26036 602 1729 4.81e-16
c26037 1694 1692 5.93e-16
c26038 1567 0 6.9481e-14
c26039 5095 0 2.285e-15
c26040 1081 732 1.35e-16
c26041 596 832 3.134e-15
c26042 9 566 4.88e-16
c26043 3236 3634 4.36e-16
c26044 2494 1987 2.48e-16
c26045 2194 2473 1.58e-16
c26046 2178 2461 1.58e-16
c26047 2172 1766 1.58e-16
c26048 2271 662 2.33e-16
c26049 2541 2582 1.96e-16
c26050 1708 767 3.15e-16
c26051 642 1327 4.03e-16
c26052 3530 1 8.43e-16
c26053 595 3397 9.84e-16
c26054 1891 1888 5.5e-16
c26055 2955 2952 5.5e-16
c26056 2178 767 3.15e-16
c26057 3363 3365 1.6e-16
c26058 1397 1 5.97e-15
c26059 3290 782 4.81e-16
c26060 2781 767 1.58e-16
c26061 2227 2225 1.6e-16
c26062 2222 2221 2.03e-16
c26063 4777 4401 3.92e-16
c26064 4789 4788 1.6e-16
c26065 2747 2736 1.58e-16
c26066 3205 707 4.81e-16
c26067 2696 692 1.58e-16
c26068 456 465 1.58e-16
c26069 1 220 4.22e-16
c26070 3397 3468 4.63e-16
c26071 3236 3627 4.11e-16
c26072 4582 4758 3.92e-16
c26073 4742 4367 4.9e-16
c26074 3411 3455 1.58e-16
c26075 657 2231 1.58e-16
c26076 642 2248 3.79e-16
c26077 2182 2461 1.58e-16
c26078 1868 1 4.41e-15
c26079 2377 0 6.62e-16
c26080 27 218 1.88e-16
c26081 3514 3509 1.642e-15
c26082 3259 782 2.33e-16
c26083 3706 3397 4.63e-16
c26084 3781 3773 4.48e-16
c26085 3932 3940 7.81e-16
c26086 687 3169 2.65e-16
c26087 1477 692 1.58e-16
c26088 3033 2538 1.176e-15
c26089 2771 2773 1.862e-15
c26090 2288 2673 1.96e-16
c26091 3333 1 2.054e-15
c26092 2182 767 3.15e-16
c26093 3626 3623 6.44e-16
c26094 3630 3627 3.01e-16
c26095 632 1 3.1284e-14
c26096 2070 2088 1.23e-16
c26097 1708 2019 5.42e-16
c26098 1684 2007 1.58e-16
c26099 1975 1971 1.96e-16
c26100 1574 0 1.6491e-14
c26101 5115 5074 3.18e-16
c26102 5101 5105 5.6e-16
c26103 687 3162 2.72e-16
c26104 4952 4944 1.58e-16
c26105 116 114 7.1e-16
c26106 2870 2486 1.58e-16
c26107 2745 1 6.15e-16
c26108 1157 782 1.58e-16
c26109 894 1066 1.58e-16
c26110 907 1038 3.54e-16
c26111 3311 1 1.716e-15
c26112 2758 762 2.72e-16
c26113 1831 677 4.81e-16
c26114 4525 842 1.9e-16
c26115 3882 4281 1.96e-16
c26116 2816 812 7.68e-16
c26117 1404 1 1.716e-15
c26118 3449 3447 1.6e-16
c26119 4839 1 1.749e-15
c26120 5283 5281 1.441e-15
c26121 5299 5301 3.92e-16
c26122 4922 4918 1.58e-16
c26123 2775 2384 4.11e-16
c26124 5417 5444 4.01e-16
c26125 595 3882 4.03e-16
c26126 3435 1 4.41e-15
c26127 2724 737 5.03e-16
c26128 4269 0 6.62e-16
c26129 4480 4452 2.64e-16
c26130 4847 4853 7.25e-16
c26131 4469 4463 9.42e-16
c26132 4015 4024 3.84e-16
c26133 4563 4333 1.58e-16
c26134 4708 4712 1.81e-16
c26135 5136 5114 1.58e-16
c26136 1964 2461 1.58e-16
c26137 2194 2236 3.92e-16
c26138 88 223 1.88e-16
c26139 1026 1028 7.72e-16
c26140 5476 5477 5.87e-16
c26141 2559 2322 1.58e-16
c26142 1916 752 4.81e-16
c26143 1517 1071 1.96e-16
c26144 1518 1511 6.73e-16
c26145 4062 1 6.76e-16
c26146 2923 2944 6.78e-16
c26147 1785 1397 4.97e-16
c26148 1414 1403 1.58e-16
c26149 1012 1 3.54e-16
c26150 1009 0 9.602e-15
c26151 3024 2583 1.58e-16
c26152 3030 2577 5.88e-16
c26153 1318 0 4.4783e-14
c26154 1553 1 1.056e-15
c26155 4590 1 1.806e-15
c26156 2029 2042 1.96e-16
c26157 1694 1590 1.58e-16
c26158 5158 5157 3.92e-16
c26159 0 364 1.051e-14
c26160 3516 3509 6.73e-16
c26161 5237 0 2.078e-15
c26162 1132 767 1.58e-16
c26163 1113 1119 1.58e-16
c26164 159 158 5.8e-16
c26165 129 175 1.88e-16
c26166 3898 3890 4.63e-16
c26167 3900 3895 1.58e-16
c26168 5356 5395 1.738e-15
c26169 2839 2452 1.532e-15
c26170 2653 2655 2.03e-16
c26171 2735 747 2.4e-16
c26172 4111 4120 3.84e-16
c26173 4125 4124 6.67e-16
c26174 1799 672 2.4e-16
c26175 1608 837 1.58e-16
c26176 632 3463 3.15e-16
c26177 4775 752 1.23e-16
c26178 3245 0 3.3551e-14
c26179 2594 2589 1.642e-15
c26180 4386 3554 2.48e-16
c26181 4407 1 2.054e-15
c26182 204 450 1.88e-16
c26183 4409 0 8e-16
c26184 4430 762 2.65e-16
c26185 2029 0 2.8699e-14
c26186 5015 5005 1.98e-16
c26187 420 418 2.84e-16
c26188 3411 3185 5.5e-16
c26189 5279 5278 5.87e-16
c26190 5262 5175 4.2e-16
c26191 4103 4104 6.4e-16
c26192 3075 1 5.808e-15
c26193 5558 5563 9.94e-16
c26194 5538 5544 1.203e-15
c26195 2764 2373 1.136e-15
c26196 3077 0 3.466e-15
c26197 1585 1579 1.6e-16
c26198 1121 1576 2.386e-15
c26199 534 1 4.59e-16
c26200 1839 1835 1.96e-16
c26201 5010 352 1.88e-16
c26202 3048 3228 1.58e-16
c26203 1857 0 1.4092e-14
c26204 1702 1 1.002e-15
c26205 421 49 1.88e-16
c26206 3208 3591 7.84e-16
c26207 902 889 4.481e-15
c26208 4743 0 1.6462e-14
c26209 4567 4310 5.5e-16
c26210 5136 5048 1.237e-15
c26211 5044 5047 1.817e-15
c26212 4793 323 1.88e-16
c26213 2451 1930 1.96e-16
c26214 2446 1936 1.96e-16
c26215 1766 0 3.5926e-14
c26216 3725 3834 6.31e-16
c26217 3833 3806 9.6e-16
c26218 3005 2486 3.92e-16
c26219 2557 822 3.15e-16
c26220 1001 677 1.58e-16
c26221 911 898 1.829e-15
c26222 3463 3435 2.64e-16
c26223 919 995 3.92e-16
c26224 922 994 2.54e-16
c26225 3610 0 3.466e-15
c26226 4175 4183 3.45e-16
c26227 3018 1 5.329e-15
c26228 3052 3047 9.6e-16
c26229 4011 1 6.66e-16
c26230 4184 25 7.01e-16
c26231 4457 3616 4.11e-16
c26232 2559 2837 3.92e-16
c26233 4463 4826 1.96e-16
c26234 1706 1690 4.274e-15
c26235 92 89 6.67e-16
c26236 1345 0 3.46872e-13
c26237 4579 1 2.94e-16
c26238 4730 4728 2.15e-16
c26239 4726 4737 1.96e-16
c26240 4744 0 2.93e-15
c26241 22 36 1.88e-16
c26242 5028 5029 3.54e-16
c26243 3806 3807 5.88e-16
c26244 280 1 9.8e-16
c26245 3480 672 1.813e-15
c26246 5324 5365 1.817e-15
c26247 4804 236 1.88e-16
c26248 2048 2044 1.64e-16
c26249 4589 5544 3.92e-16
c26250 3388 0 1.4835e-14
c26251 2535 2819 1.58e-16
c26252 2557 2807 1.58e-16
c26253 3882 3537 1.58e-16
c26254 1363 1352 1.58e-16
c26255 3732 0 2.8687e-14
c26256 3992 25 7.01e-16
c26257 2535 2254 1.58e-16
c26258 2541 2248 5.88e-16
c26259 3123 662 2.33e-16
c26260 1794 1789 1.642e-15
c26261 1921 1922 2.48e-16
c26262 1708 1747 5.42e-16
c26263 1684 1735 1.58e-16
c26264 1056 0 3.7097e-14
c26265 33 584 3.75e-16
c26266 831 820 7.23e-16
c26267 3376 3048 6.7e-16
c26268 4919 1 5.21e-16
c26269 3030 752 3.15e-16
c26270 2165 1652 1.58e-16
c26271 241 0 2.87e-16
c26272 3662 3659 5.5e-16
c26273 2424 1 4.41e-15
c26274 2734 2350 1.58e-16
c26275 2638 0 6.62e-16
c26276 2178 2196 4.312e-15
c26277 2136 2056 1.58e-16
c26278 642 3100 3.79e-16
c26279 632 3483 4.81e-16
c26280 1327 732 4.03e-16
c26281 3983 3991 3.45e-16
c26282 3210 0 2.93e-15
c26283 2248 2243 1.642e-15
c26284 1239 1240 1.03e-16
c26285 1236 1241 1.81e-16
c26286 146 1 4.22e-16
c26287 3960 36 1.88e-16
c26288 3531 4353 1.58e-16
c26289 4481 797 3.64e-16
c26290 1327 1623 1.96e-16
c26291 632 1010 1.58e-16
c26292 366 1 3.6e-16
c26293 2559 792 3.58e-16
c26294 3219 747 3.79e-16
c26295 3202 762 1.58e-16
c26296 4538 4553 1.96e-16
c26297 2288 702 5.73e-16
c26298 595 1690 4.03e-16
c26299 2798 807 3.79e-16
c26300 4721 1 8.85e-16
c26301 4813 4825 2.62e-16
c26302 4497 0 6.9455e-14
c26303 3211 737 1.58e-16
c26304 1670 1249 6.17e-16
c26305 1 313 1.44e-16
c26306 4827 4831 1.81e-16
c26307 2182 2196 4.274e-15
c26308 2333 1817 1.136e-15
c26309 662 1022 1.58e-16
c26310 895 888 2.335e-15
c26311 3702 3691 1.96e-16
c26312 777 2410 1.58e-16
c26313 2194 1817 1.58e-16
c26314 1226 1224 1.963e-15
c26315 5352 294 3.54e-16
c26316 378 369 1.58e-16
c26317 3702 842 7.68e-16
c26318 5414 5409 3.73e-16
c26319 601 2594 1.58e-16
c26320 3001 0 1.7608e-14
c26321 2946 2503 9.1e-16
c26322 2708 2316 2.38e-15
c26323 2631 2629 1.6e-16
c26324 1470 1031 1.96e-16
c26325 2478 827 1.832e-15
c26326 601 1375 1.58e-16
c26327 1088 0 1.4198e-14
c26328 895 1 2.048e-15
c26329 3282 3289 6.73e-16
c26330 4534 1 1.056e-15
c26331 3192 2685 3.92e-16
c26332 2854 842 7.38e-16
c26333 2559 737 3.15e-16
c26334 1630 0 1.4092e-14
c26335 3191 3573 2.48e-16
c26336 2246 1 6.15e-16
c26337 891 893 1.58e-16
c26338 4580 4231 1.58e-16
c26339 3490 3487 6.44e-16
c26340 3494 3491 3.01e-16
c26341 3583 737 7.68e-16
c26342 2325 1828 1.58e-16
c26343 890 752 3.15e-16
c26344 907 1112 3.92e-16
c26345 2214 1 5.97e-15
c26346 7 8 7.08e-16
c26347 1837 707 1.58e-16
c26348 1465 702 3.79e-16
c26349 1026 1457 7.84e-16
c26350 3188 1 1.056e-15
c26351 2879 2884 3.73e-16
c26352 1385 957 1.96e-16
c26353 2393 752 1.832e-15
c26354 3927 37 1.88e-16
c26355 2308 677 1.832e-15
c26356 2002 2003 9.1e-16
c26357 1708 1488 1.58e-16
c26358 1706 1482 5.5e-16
c26359 1694 1883 1.58e-16
c26360 1444 0 6.72e-16
c26361 482 484 1.257e-15
c26362 494 483 3.84e-16
c26363 450 175 1.88e-16
c26364 3576 722 1.9e-16
c26365 2323 2334 1.96e-16
c26366 3387 3655 3.92e-16
c26367 5010 294 1.88e-16
c26368 3282 797 1.84e-16
c26369 5262 5232 1.604e-15
c26370 2799 2401 4.36e-16
c26371 4736 323 1.88e-16
c26372 2492 2503 1.58e-16
c26373 2172 2490 1.58e-16
c26374 2194 2478 1.58e-16
c26375 3315 822 2.72e-16
c26376 2884 2877 8.3e-16
c26377 1343 692 4.46e-16
c26378 1331 702 7.99e-16
c26379 74 9 4.88e-16
c26380 4338 3503 1.96e-16
c26381 4343 3497 1.96e-16
c26382 4460 782 1.09e-16
c26383 1327 1588 1.58e-16
c26384 1211 1188 6.54e-16
c26385 632 1321 4.48e-16
c26386 4596 4594 1.6e-16
c26387 2172 782 4.48e-16
c26388 4865 4863 2.03e-16
c26389 2747 3271 4.36e-16
c26390 3393 3083 5.88e-16
c26391 1 320 4.22e-16
c26392 13 334 1.88e-16
c26393 4582 4775 3.92e-16
c26394 2196 1964 5.5e-16
c26395 512 523 3.84e-16
c26396 3948 3949 7.81e-16
c26397 687 2662 3.79e-16
c26398 1472 717 1.58e-16
c26399 1203 907 3.54e-16
c26400 3898 702 3.15e-16
c26401 4742 5170 6.17e-16
c26402 919 1053 1.58e-16
c26403 661 19 1.96e-16
c26404 1922 767 1.832e-15
c26405 1331 981 1.58e-16
c26406 3506 0 3.3874e-14
c26407 1196 1195 3.94e-16
c26408 3030 2549 3.15e-16
c26409 2951 2887 2.249e-15
c26410 2509 2969 5.71e-16
c26411 595 1357 2.72e-16
c26412 612 1353 1.58e-16
c26413 822 1177 1.58e-16
c26414 868 19 1.41e-15
c26415 1062 0 6.29e-16
c26416 4111 19 3.84e-16
c26417 4120 0 2.0707e-14
c26418 3083 3078 1.642e-15
c26419 747 1087 1.58e-16
c26420 4395 4778 4.97e-16
c26421 4777 4781 1.96e-16
c26422 2115 2070 3.18e-16
c26423 2123 2108 6.67e-16
c26424 3540 3552 2.32e-16
c26425 3647 782 1.09e-16
c26426 5104 5101 3.54e-16
c26427 4793 265 1.88e-16
c26428 2404 2402 1.6e-16
c26429 2183 1 3.009e-15
c26430 707 699 1.74e-16
c26431 2184 0 5.86e-16
c26432 4954 4952 7.26e-16
c26433 2754 1 1.716e-15
c26434 2676 2673 3.01e-16
c26435 2672 2669 6.44e-16
c26436 3337 1 8.43e-16
c26437 4634 5464 1.96e-16
c26438 3830 1 7.87e-16
c26439 4406 4407 1.6e-16
c26440 4402 3571 3.92e-16
c26441 1612 1608 1.96e-16
c26442 4701 4694 1.96e-16
c26443 4310 4703 1.914e-15
c26444 371 361 8.86e-16
c26445 1556 1 4.41e-15
c26446 786 775 7.23e-16
c26447 778 779 1.6e-16
c26448 4944 4990 9.29e-16
c26449 1940 0 6.62e-16
c26450 3387 3620 1.58e-16
c26451 5284 5288 1.96e-16
c26452 4674 410 1.88e-16
c26453 1053 1067 1.96e-16
c26454 2539 0 6.78e-16
c26455 5463 1 3.36e-16
c26456 1101 767 1.75e-16
c26457 1360 1357 3.01e-16
c26458 1356 1353 6.44e-16
c26459 3882 4280 1.58e-16
c26460 1993 842 1.84e-16
c26461 1345 1091 5.5e-16
c26462 595 953 1.58e-16
c26463 602 954 1.222e-15
c26464 910 1318 3.75e-16
c26465 3086 3084 1.6e-16
c26466 4294 1 1.868e-15
c26467 2744 737 1.09e-16
c26468 1881 1880 1.6e-16
c26469 1873 1871 2.15e-16
c26470 4284 0 2.93e-15
c26471 3350 3349 1.6e-16
c26472 538 537 7.08e-16
c26473 2080 2081 2.12e-16
c26474 963 969 1.58e-16
c26475 1 446 4.22e-16
c26476 3409 767 4.46e-16
c26477 4563 4350 1.58e-16
c26478 4725 4727 4.93e-16
c26479 4776 33 1.88e-16
c26480 1964 2481 2.38e-15
c26481 5151 238 3.54e-16
c26482 2172 2253 3.92e-16
c26483 397 565 1.88e-16
c26484 3781 3866 3.96e-16
c26485 3919 3910 9.33e-16
c26486 1031 1008 6.54e-16
c26487 921 1040 1.96e-16
c26488 5391 5389 3.92e-16
c26489 1076 1071 1.58e-16
c26490 616 19 1.96e-16
c26491 4499 4492 6.73e-16
c26492 4498 3656 1.96e-16
c26493 3346 2838 2.48e-16
c26494 4607 1 1.806e-15
c26495 4367 4745 7.84e-16
c26496 421 194 1.88e-16
c26497 1955 1957 2.03e-16
c26498 30 500 6.83e-16
c26499 37 490 1.88e-16
c26500 3621 767 7.38e-16
c26501 5064 5071 8.94e-16
c26502 5066 5069 1.342e-15
c26503 2131 1 1.88e-16
c26504 93 0 5.7351e-14
c26505 1132 1134 7.84e-16
c26506 921 662 3.15e-16
c26507 110 19 8.82e-16
c26508 146 363 1.88e-16
c26509 4216 4208 7.45e-16
c26510 4345 677 3.64e-16
c26511 2688 0 3.3717e-14
c26512 2166 2572 2.38e-15
c26513 3731 3736 3.73e-16
c26514 2923 2913 1.021e-15
c26515 1422 986 4.97e-16
c26516 1001 996 1.58e-16
c26517 3265 0 1.4092e-14
c26518 84 85 6.4e-16
c26519 2545 2701 4.63e-16
c26520 4038 26 4.48e-16
c26521 3387 792 3.15e-16
c26522 3153 3146 6.73e-16
c26523 30 180 3.84e-16
c26524 3599 762 3.79e-16
c26525 4425 0 6.72e-16
c26526 3582 777 1.58e-16
c26527 3420 3018 4.97e-16
c26528 627 2236 2.4e-16
c26529 2168 2167 4.57e-16
c26530 1055 702 1.85e-16
c26531 4012 4006 1.96e-16
c26532 3095 1 2.054e-15
c26533 1091 1088 1.984e-15
c26534 3673 837 1.58e-16
c26535 4770 5262 1.58e-16
c26536 3097 0 8e-16
c26537 2557 2475 1.58e-16
c26538 922 1175 3.92e-16
c26539 910 1345 5.03e-16
c26540 777 783 1.097e-15
c26541 1706 1786 1.58e-16
c26542 4561 4197 1.886e-15
c26543 4214 4215 3.225e-15
c26544 4760 0 1.6462e-14
c26545 752 768 1.621e-15
c26546 1 380 4.92e-16
c26547 3387 737 4.48e-16
c26548 4088 857 3.1e-16
c26549 4736 265 7.84e-16
c26550 910 3388 7.06e-16
c26551 5358 0 3.974e-14
c26552 2178 2192 3.92e-16
c26553 146 131 1.88e-16
c26554 151 120 1.88e-16
c26555 3565 737 3.15e-16
c26556 5449 5447 1.373e-15
c26557 2968 2503 8.82e-16
c26558 1706 702 3.15e-16
c26559 3449 1 1.056e-15
c26560 2254 2637 7.84e-16
c26561 2196 852 3.58e-16
c26562 1211 1677 1.58e-16
c26563 782 0 2.79792e-13
c26564 4199 37 1.88e-16
c26565 4843 4463 1.96e-16
c26566 2713 3223 1.58e-16
c26567 3146 677 1.84e-16
c26568 1 267 5.698e-15
c26569 2356 2357 1.35e-16
c26570 2279 0 8e-16
c26571 2182 2192 3.92e-16
c26572 2196 2168 3.54e-16
c26573 4855 410 1.88e-16
c26574 642 644 5.59e-16
c26575 2764 2759 1.642e-15
c26576 2041 2031 1.58e-16
c26577 3394 0 4.1004e-14
c26578 2559 2836 5.42e-16
c26579 2535 2824 1.58e-16
c26580 1151 1147 3.78e-16
c26581 1363 1761 4.36e-16
c26582 2325 717 1.58e-16
c26583 1708 1752 1.58e-16
c26584 436 450 1.88e-16
c26585 320 363 1.88e-16
c26586 5543 584 3.19e-16
c26587 2368 2359 3.92e-16
c26588 1851 2362 5.66e-16
c26589 741 730 7.23e-16
c26590 733 734 1.6e-16
c26591 3508 672 2.72e-16
c26592 3313 837 1.58e-16
c26593 2266 2268 1.6e-16
c26594 420 1 1.073e-15
c26595 4537 0 1.7584e-14
c26596 632 624 1.74e-16
c26597 9 136 5.8e-16
c26598 4753 33 1.88e-16
c26599 2739 2350 2.386e-15
c26600 2722 2367 1.58e-16
c26601 4012 3918 2.87e-16
c26602 1076 1075 3.94e-16
c26603 3531 4373 2.38e-15
c26604 3650 797 3.15e-16
c26605 4656 647 1.23e-16
c26606 5514 5417 6.72e-16
c26607 1343 1640 3.92e-16
c26608 746 1 5.57e-16
c26609 2722 2734 2.32e-16
c26610 1558 1559 2.48e-16
c26611 1231 1 2.808e-15
c26612 3505 3507 2.03e-16
c26613 1694 1352 1.58e-16
c26614 4175 1 5.284e-15
c26615 1819 1821 2.03e-16
c26616 4889 4503 1.812e-15
c26617 1820 1 5.808e-15
c26618 3299 3296 5.5e-16
c26619 3034 2696 5.5e-16
c26620 1822 0 3.466e-15
c26621 3659 3666 1.96e-16
c26622 4738 1 8.85e-16
c26623 4916 0 1.63e-15
c26624 2149 2162 1.96e-16
c26625 14 5 2.218e-15
c26626 4844 4846 4.93e-16
c26627 5261 5259 1.167e-15
c26628 0 19 7.1256e-13
c26629 2425 0 1.6491e-14
c26630 3035 1 3.009e-15
c26631 2423 1913 1.96e-16
c26632 2172 1834 1.58e-16
c26633 2178 1828 5.88e-16
c26634 1243 1242 5.64e-16
c26635 64 120 1.88e-16
c26636 146 310 1.88e-16
c26637 617 2594 3.15e-16
c26638 3036 0 5.86e-16
c26639 922 767 5.14e-16
c26640 921 1098 1.58e-16
c26641 1001 1004 6.13e-16
c26642 1939 807 1.58e-16
c26643 1327 1011 1.58e-16
c26644 3876 4523 1.58e-16
c26645 3900 4535 5.42e-16
c26646 627 1389 1.58e-16
c26647 617 1375 1.84e-16
c26648 3983 1 5.284e-15
c26649 2770 2781 1.58e-16
c26650 3030 3190 1.96e-16
c26651 1735 1737 2.15e-16
c26652 4813 4811 1.687e-15
c26653 3209 737 1.339e-15
c26654 4554 1 7.21e-16
c26655 601 1735 1.832e-15
c26656 4580 4248 1.58e-16
c26657 1902 2410 7.84e-16
c26658 2182 1828 5.5e-16
c26659 2255 1 1.716e-15
c26660 732 734 5.59e-16
c26661 3202 722 3.15e-16
c26662 2892 3850 1.33e-16
c26663 3866 3853 1.96e-16
c26664 3338 3858 5.69e-16
c26665 632 3094 5.03e-16
c26666 42 50 2.218e-15
c26667 47 49 1.257e-15
c26668 2712 2316 1.96e-16
c26669 2794 0 6.72e-16
c26670 2631 1 1.056e-15
c26671 5324 5345 1.96e-16
c26672 2792 2407 1.96e-16
c26673 2237 2619 2.48e-16
c26674 1857 707 1.58e-16
c26675 1031 1469 1.58e-16
c26676 3204 1 9.28e-16
c26677 3605 4438 7.84e-16
c26678 3281 2764 4.11e-16
c26679 3948 25 1.88e-16
c26680 3944 19 7.35e-16
c26681 2679 3193 4.97e-16
c26682 2852 827 4.81e-16
c26683 1684 1499 5.5e-16
c26684 1694 1888 1.58e-16
c26685 526 584 3.45e-16
c26686 657 1766 1.58e-16
c26687 1533 1901 1.96e-16
c26688 450 349 1.88e-16
c26689 571 575 1.372e-15
c26690 5148 0 1.376e-15
c26691 5133 31 5.5e-16
c26692 3411 3672 3.92e-16
c26693 1083 732 1.58e-16
c26694 890 891 1.343e-15
c26695 3652 3651 1.6e-16
c26696 2514 2510 1.96e-16
c26697 1345 707 3.15e-16
c26698 971 1372 1.58e-16
c26699 1374 881 4.11e-16
c26700 1221 1222 2.377e-15
c26701 2559 2599 3.92e-16
c26702 1639 1640 9.1e-16
c26703 657 1345 3.58e-16
c26704 1232 1 3.24e-16
c26705 1690 1687 1.123e-15
c26706 4317 0 1.6491e-14
c26707 5042 5026 7.48e-16
c26708 1227 0 6.29e-16
c26709 689 688 1.6e-16
c26710 3637 3638 9.1e-16
c26711 4794 4418 3.92e-16
c26712 4806 4805 1.6e-16
c26713 2404 1 1.056e-15
c26714 1635 2078 9.7e-16
c26715 4582 4792 3.92e-16
c26716 5165 5192 4.01e-16
c26717 4691 468 1.88e-16
c26718 5010 62 1.88e-16
c26719 2495 2507 2.32e-16
c26720 0 557 1.4515e-14
c26721 3287 782 1.58e-16
c26722 5310 1 7.87e-16
c26723 3900 717 3.58e-16
c26724 1056 707 2.33e-16
c26725 146 339 1.88e-16
c26726 3526 0 1.4092e-14
c26727 3886 3656 1.58e-16
c26728 3362 3377 1.96e-16
c26729 3813 410 9.02e-16
c26730 3030 3155 1.58e-16
c26731 1593 1 5.808e-15
c26732 1595 0 3.466e-15
c26733 310 320 3.75e-16
c26734 26 204 8.41e-16
c26735 37 201 5.71e-16
c26736 3732 3775 2.15e-16
c26737 2199 0 1.23e-16
c26738 1149 1156 2.27e-16
c26739 894 1053 3.54e-16
c26740 3381 4237 2.38e-15
c26741 2586 2598 2.32e-16
c26742 2541 2186 3.15e-16
c26743 1191 868 4e-16
c26744 1444 1443 5.65e-16
c26745 394 395 6.67e-16
c26746 856 1 4.03e-16
c26747 702 26 1.58e-16
c26748 3920 1 9.475e-15
c26749 4102 19 7.04e-16
c26750 3900 4298 3.92e-16
c26751 3163 3160 5.5e-16
c26752 3633 0 6.9481e-14
c26753 3453 3072 3.92e-16
c26754 3457 3458 1.6e-16
c26755 349 337 1.58e-16
c26756 3570 707 1.58e-16
c26757 5316 323 3.15e-16
c26758 2313 2310 3.01e-16
c26759 2309 2306 6.44e-16
c26760 5424 5423 1.6e-16
c26761 5232 149 1.58e-16
c26762 3310 3393 1.58e-16
c26763 595 3421 1.58e-16
c26764 398 15 4.88e-16
c26765 3882 4285 1.58e-16
c26766 3898 4297 1.58e-16
c26767 5588 5589 1.6e-16
c26768 4514 5590 1.23e-16
c26769 4520 5575 3.92e-16
c26770 5577 5579 1.96e-16
c26771 2868 2861 6.73e-16
c26772 2611 0 6.9481e-14
c26773 2541 2555 3.92e-16
c26774 2559 2563 1.6e-16
c26775 601 954 1.58e-16
c26776 839 26 2.65e-15
c26777 656 1 5.57e-16
c26778 1406 0 3.3656e-14
c26779 1200 1 3.06e-16
c26780 1667 1675 4.06e-16
c26781 2098 178 1.108e-15
c26782 982 984 7.84e-16
c26783 5196 5194 3.25e-16
c26784 762 2356 5.73e-16
c26785 5493 5491 3.92e-16
c26786 2880 0 2.8687e-14
c26787 920 1054 1.58e-16
c26788 1076 1534 4.36e-16
c26789 1532 1525 1.96e-16
c26790 1343 1368 3.92e-16
c26791 2566 3074 2.48e-16
c26792 3667 3656 1.58e-16
c26793 3048 2594 5.5e-16
c26794 1557 1 1.716e-15
c26795 4624 1 1.806e-15
c26796 3409 3401 4.63e-16
c26797 2087 2064 5.87e-16
c26798 339 320 1.88e-16
c26799 3530 3523 1.96e-16
c26800 2373 2384 1.58e-16
c26801 1834 0 3.583e-14
c26802 2163 1 7.21e-16
c26803 3767 3739 4.39e-16
c26804 3514 677 3.15e-16
c26805 2708 0 1.4092e-14
c26806 2170 2554 2.79e-16
c26807 542 262 1.88e-16
c26808 3134 0 6.921e-14
c26809 2968 2966 3.92e-16
c26810 2954 2959 3.73e-16
c26811 3886 4434 4.63e-16
c26812 1789 1786 5.5e-16
c26813 3338 1 5.343e-15
c26814 811 1 4.03e-16
c26815 1690 1986 1.96e-16
c26816 3851 0 1.376e-15
c26817 1592 1594 2.03e-16
c26818 2557 672 3.15e-16
c26819 2535 647 4.48e-16
c26820 1584 1556 2.64e-16
c26821 187 204 1.325e-15
c26822 4993 4980 1.96e-16
c26823 3048 807 3.58e-16
c26824 2290 1777 4.97e-16
c26825 162 163 6.67e-16
c26826 88 305 1.88e-16
c26827 2171 2191 2.07e-16
c26828 4787 4401 1.179e-15
c26829 4838 468 1.88e-16
c26830 2686 0 1.6491e-14
c26831 2169 2571 1.96e-16
c26832 3708 3712 1.96e-16
c26833 4127 4126 5.5e-16
c26834 1803 672 1.58e-16
c26835 3327 3397 1.58e-16
c26836 4600 497 7.84e-16
c26837 1547 752 1.09e-16
c26838 4387 4399 2.32e-16
c26839 5573 5514 3.54e-16
c26840 2557 2299 5.5e-16
c26841 2535 2492 1.58e-16
c26842 611 1 5.57e-16
c26843 3878 0 5.96e-16
c26844 3160 2645 2.386e-15
c26845 3057 2529 4.97e-16
c26846 5005 5007 1.417e-15
c26847 5013 4546 5.5e-16
c26848 2987 2986 5.5e-16
c26849 3024 2736 1.58e-16
c26850 3030 2730 5.88e-16
c26851 792 1145 1.85e-16
c26852 4946 0 4.4619e-14
c26853 1 459 2.87e-16
c26854 4777 0 1.6462e-14
c26855 122 120 1.96e-16
c26856 281 262 1.88e-16
c26857 5160 5155 7.46e-16
c26858 5044 5032 1.75e-16
c26859 4804 178 1.88e-16
c26860 4776 526 1.88e-16
c26861 2463 1947 4.11e-16
c26862 4691 64 1.88e-16
c26863 1708 717 3.58e-16
c26864 3465 1 9.28e-16
c26865 1331 1326 1.58e-16
c26866 543 0 1.0822e-14
c26867 529 30 6.83e-16
c26868 528 33 1.88e-16
c26869 602 920 9.47e-16
c26870 4479 4470 3.46e-16
c26871 2178 717 4.03e-16
c26872 1684 1952 3.92e-16
c26873 1 163 3.6e-16
c26874 123 30 6.83e-16
c26875 114 37 5.71e-16
c26876 4691 4310 5.2e-16
c26877 4571 4707 3.92e-16
c26878 2295 0 6.72e-16
c26879 2078 1 5.966e-15
c26880 0 195 1.0822e-14
c26881 26 175 8.41e-16
c26882 37 158 1.88e-16
c26883 5296 352 1.58e-16
c26884 5210 1 3.36e-16
c26885 3806 3821 1.739e-15
c26886 3822 3820 3.92e-16
c26887 1432 662 7.68e-16
c26888 909 807 3.15e-16
c26889 2266 2260 1.6e-16
c26890 1335 898 3.84e-16
c26891 4184 4182 3.54e-16
c26892 4315 672 2.4e-16
c26893 2820 2452 1.96e-16
c26894 4226 3918 8.1e-16
c26895 4600 5569 5.5e-16
c26896 4606 5429 1.96e-16
c26897 2559 2841 1.58e-16
c26898 3886 4399 1.58e-16
c26899 3898 3548 5.5e-16
c26900 3900 3554 1.58e-16
c26901 3322 2804 1.96e-16
c26902 2182 717 7.99e-16
c26903 4008 37 5.71e-16
c26904 2736 762 1.58e-16
c26905 2156 858 6.67e-16
c26906 923 0 5.6106e-14
c26907 766 1 4.03e-16
c26908 2645 702 1.58e-16
c26909 1690 1951 1.58e-16
c26910 3397 762 7.99e-16
c26911 3133 3124 3.46e-16
c26912 3521 3134 1.532e-15
c26913 910 19 2.105e-15
c26914 841 839 5.88e-16
c26915 3333 837 1.58e-16
c26916 595 2215 2.65e-16
c26917 602 1681 2.33e-16
c26918 4844 5093 3.92e-16
c26919 2665 1 1.056e-15
c26920 890 992 1.96e-16
c26921 642 649 1.6e-16
c26922 5561 1 5.04e-16
c26923 4086 4088 3.54e-16
c26924 1606 797 1.58e-16
c26925 1415 981 1.96e-16
c26926 1416 1409 6.73e-16
c26927 2178 2371 1.58e-16
c26928 1521 737 7.38e-16
c26929 1270 1273 1.021e-15
c26930 2323 717 1.58e-16
c26931 3725 439 1.707e-15
c26932 2611 3122 1.96e-16
c26933 3763 1 1.88e-16
c26934 2492 858 3.69e-16
c26935 2688 707 1.58e-16
c26936 4918 4916 3.92e-16
c26937 3311 837 1.58e-16
c26938 1840 1 2.054e-15
c26939 1842 0 8e-16
c26940 3393 3535 1.58e-16
c26941 4830 4842 2.62e-16
c26942 747 1505 1.58e-16
c26943 233 37 1.88e-16
c26944 2737 2350 1.532e-15
c26945 792 2435 2.22e-16
c26946 2194 1845 5.5e-16
c26947 2182 2371 1.58e-16
c26948 1749 1 4.41e-15
c26949 932 918 5.74e-16
c26950 165 9 5.8e-16
c26951 3992 3990 3.54e-16
c26952 1071 732 4e-16
c26953 3051 0 1.23e-16
c26954 2725 2732 6.73e-16
c26955 372 19 3.2e-16
c26956 4284 3452 2.48e-16
c26957 1343 1026 1.58e-16
c26958 3408 1 2.94e-16
c26959 537 552 1.88e-16
c26960 3020 3019 4.57e-16
c26961 2503 868 2.22e-16
c26962 2920 2922 9.16e-16
c26963 3296 3303 1.96e-16
c26964 3046 3207 3.92e-16
c26965 2194 677 4.46e-16
c26966 629 630 1.6e-16
c26967 3666 3657 3.46e-16
c26968 2014 1618 1.96e-16
c26969 2009 1624 1.96e-16
c26970 617 1735 1.58e-16
c26971 1191 0 3.7577e-14
c26972 25 291 5.71e-16
c26973 4580 4265 1.58e-16
c26974 5162 5155 9.38e-16
c26975 1913 2422 1.58e-16
c26976 898 888 3.54e-16
c26977 3974 3979 1.96e-16
c26978 894 1127 3.92e-16
c26979 909 1126 1.88e-16
c26980 883 1119 1.58e-16
c26981 234 237 6.67e-16
c26982 4617 1 8.21e-15
c26983 922 931 1.58e-16
c26984 1483 1477 1.6e-16
c26985 1031 1474 2.386e-15
c26986 1046 1457 1.58e-16
c26987 898 1 7.867e-15
c26988 3217 1 6.15e-16
c26989 3974 1 7.08e-16
c26990 3616 4421 1.58e-16
c26991 1885 767 1.75e-16
c26992 1706 1369 1.58e-16
c26993 1737 1733 1.96e-16
c26994 3958 37 1.88e-16
c26995 3967 25 4.68e-16
c26996 2858 842 1.832e-15
c26997 1708 1516 5.5e-16
c26998 1041 1 4.044e-15
c26999 1475 0 6.62e-16
c27000 3106 3489 7.84e-16
c27001 3882 762 4.03e-16
c27002 204 190 1.58e-16
c27003 2349 1828 1.96e-16
c27004 2344 1834 1.96e-16
c27005 5098 122 9.1e-16
c27006 2787 812 1.75e-16
c27007 29 1 4.92e-16
c27008 13 11 1.257e-15
c27009 3409 3688 1.58e-16
c27010 5324 5316 3.54e-16
c27011 4172 3918 2.87e-16
c27012 5229 5240 1.619e-15
c27013 4753 526 1.88e-16
c27014 2178 1987 1.58e-16
c27015 1389 957 2.386e-15
c27016 4838 64 1.88e-16
c27017 1254 1250 3.92e-16
c27018 4355 3514 4.11e-16
c27019 1345 1605 5.42e-16
c27020 1321 1593 1.58e-16
c27021 1437 1438 1.35e-16
c27022 683 0 1.1593e-14
c27023 1106 1538 1.96e-16
c27024 3409 3123 1.58e-16
c27025 4613 4611 1.6e-16
c27026 1533 1900 1.58e-16
c27027 1237 0 1.1576e-14
c27028 4875 1 1.013e-15
c27029 4882 4880 2.03e-16
c27030 1810 1 8.43e-16
c27031 1014 1021 2.27e-16
c27032 4793 4799 5.87e-16
c27033 4582 4809 3.92e-16
c27034 5151 5245 5.82e-16
c27035 2182 1987 1.58e-16
c27036 0 512 1.5723e-14
c27037 5323 1 1.23e-16
c27038 53 1 2.87e-16
c27039 73 13 1.88e-16
c27040 3958 3959 1.58e-16
c27041 5514 5412 1.58e-16
c27042 5526 5388 3.54e-16
c27043 2982 1 1.88e-16
c27044 3870 4595 2.196e-15
c27045 612 1374 2.72e-16
c27046 1053 1 1.56e-15
c27047 4143 1 5.284e-15
c27048 2463 827 5.03e-16
c27049 4875 4873 1.6e-16
c27050 4133 0 1.5061e-14
c27051 4135 19 3.45e-16
c27052 3274 3275 9.1e-16
c27053 1613 1 2.054e-15
c27054 4412 4795 4.97e-16
c27055 4794 4798 1.96e-16
c27056 5198 5252 9.34e-16
c27057 1615 0 8e-16
c27058 512 514 1.58e-16
c27059 511 510 6.67e-16
c27060 523 505 1.58e-16
c27061 0 331 9.795e-15
c27062 27 334 1.88e-16
c27063 33 325 4.12e-16
c27064 3560 3557 5.5e-16
c27065 2196 2304 3.92e-16
c27066 2209 0 1.4092e-14
c27067 1143 797 1.58e-16
c27068 59 508 1.88e-16
c27069 3531 717 1.813e-15
c27070 2684 2299 1.96e-16
c27071 5320 5321 3.54e-16
c27072 65 62 4.6e-16
c27073 3321 3708 1.532e-15
c27074 2989 2984 9.94e-16
c27075 1181 852 1.58e-16
c27076 1196 827 3.57e-16
c27077 3744 3745 3.18e-16
c27078 1367 1368 9.1e-16
c27079 3839 3822 8.15e-16
c27080 4425 4424 5.65e-16
c27081 4419 3582 1.532e-15
c27082 5588 5580 7.29e-16
c27083 2541 2769 1.96e-16
c27084 707 19 1.676e-15
c27085 687 1801 1.58e-16
c27086 657 19 1.41e-15
c27087 1967 1 1.056e-15
c27088 4965 4941 5.87e-16
c27089 5034 1 3.944e-15
c27090 2223 2235 2.32e-16
c27091 3393 3236 5.88e-16
c27092 1073 1074 1.213e-15
c27093 4143 4151 3.45e-16
c27094 2166 0 4.79e-14
c27095 1570 767 4.81e-16
c27096 3900 842 3.15e-16
c27097 2559 2569 1.58e-16
c27098 920 1220 3.92e-16
c27099 921 1219 2.54e-16
c27100 601 975 6.48e-16
c27101 627 968 1.58e-16
c27102 3707 3708 1.35e-16
c27103 1624 842 2.33e-16
c27104 1331 1116 1.58e-16
c27105 4706 4707 8.22e-16
c27106 4312 1 9.28e-16
c27107 3090 2583 3.92e-16
c27108 3094 3095 1.6e-16
c27109 1886 1897 1.96e-16
c27110 1214 1 3.06e-16
c27111 1414 1 5.97e-15
c27112 5224 178 3.54e-16
c27113 466 465 7.03e-16
c27114 4640 4646 5.87e-16
c27115 4563 4361 5.88e-16
c27116 4571 4367 1.58e-16
c27117 1981 1970 1.58e-16
c27118 3919 3928 3.84e-16
c27119 3933 3932 6.67e-16
c27120 4438 767 1.832e-15
c27121 5482 381 1.58e-16
c27122 921 852 3.15e-16
c27123 1321 1385 3.92e-16
c27124 4513 4506 1.96e-16
c27125 3667 4515 4.36e-16
c27126 2637 647 1.832e-15
c27127 2463 812 1.9e-16
c27128 4092 26 4.58e-16
c27129 4641 1 1.806e-15
c27130 4384 4762 7.84e-16
c27131 2082 2093 3.92e-16
c27132 1583 1 8.43e-16
c27133 542 543 6.96e-16
c27134 1 424 3.6e-16
c27135 479 117 1.88e-16
c27136 3411 3434 3.92e-16
c27137 26 436 8.41e-16
c27138 4567 4566 1.357e-15
c27139 5121 5098 8.66e-16
c27140 692 682 6.38e-16
c27141 3723 3387 3.92e-16
c27142 2541 2367 5.88e-16
c27143 2756 2373 7.84e-16
c27144 2170 2169 1.58e-16
c27145 2541 2734 1.58e-16
c27146 1687 1693 5.8e-16
c27147 1257 1254 5.47e-16
c27148 1249 1253 1.836e-15
c27149 1037 0 1.0065e-14
c27150 1706 2003 3.92e-16
c27151 1967 1965 1.6e-16
c27152 117 189 1.88e-16
c27153 3540 692 1.832e-15
c27154 5262 265 1.96e-16
c27155 2104 0 2.9272e-14
c27156 762 1690 4.03e-16
c27157 1426 1423 5.5e-16
c27158 2600 1 4.41e-15
c27159 595 3046 3.15e-16
c27160 602 3030 3.15e-16
c27161 2172 2406 3.92e-16
c27162 4015 1701 2.697e-15
c27163 3886 3418 1.58e-16
c27164 4509 842 1.84e-16
c27165 2848 2839 3.46e-16
c27166 2367 732 2.22e-16
c27167 2535 2316 5.5e-16
c27168 602 935 1.11e-16
c27169 3625 792 1.58e-16
c27170 262 259 3.54e-16
c27171 3424 3421 5.5e-16
c27172 3048 2753 1.58e-16
c27173 3046 2747 5.5e-16
c27174 3034 3274 1.58e-16
c27175 1522 0 3.6012e-14
c27176 2186 2175 4.097e-15
c27177 592 760 6.34e-16
c27178 4794 0 1.6462e-14
c27179 2574 2571 3.01e-16
c27180 4872 352 1.88e-16
c27181 2503 0 5.6922e-14
c27182 2178 2405 1.58e-16
c27183 2178 1715 1.58e-16
c27184 2518 2512 9.61e-16
c27185 379 381 6.01e-16
c27186 4304 4305 1.6e-16
c27187 4300 3469 3.92e-16
c27188 3478 1 6.15e-16
c27189 4197 3879 1.96e-16
c27190 1510 1506 1.96e-16
c27191 3839 3786 9.01e-16
c27192 2921 2918 9.58e-16
c27193 601 920 5.92e-16
c27194 3381 0 4.7676e-14
c27195 2866 1 1.492e-15
c27196 1727 1 1.868e-15
c27197 2651 677 2.33e-16
c27198 2557 797 4.46e-16
c27199 2545 807 7.99e-16
c27200 2045 2028 1.287e-15
c27201 1708 1969 3.92e-16
c27202 1717 0 2.93e-15
c27203 1 368 2.3e-14
c27204 3370 3367 8.32e-16
c27205 2196 1885 1.58e-16
c27206 2182 2405 1.58e-16
c27207 3508 3504 1.96e-16
c27208 0 352 1.24903e-13
c27209 26 349 8.41e-16
c27210 19 332 3.84e-16
c27211 3705 3393 1.58e-16
c27212 3693 3409 1.58e-16
c27213 657 2611 1.813e-15
c27214 747 1845 1.58e-16
c27215 2182 1715 1.58e-16
c27216 1449 672 2.65e-16
c27217 1202 827 1.58e-16
c27218 5358 5355 7.84e-16
c27219 2833 2441 1.96e-16
c27220 2671 1 5.808e-15
c27221 3886 3872 1.58e-16
c27222 4205 4206 7.81e-16
c27223 657 1406 1.58e-16
c27224 3248 1 2.054e-15
c27225 1166 1169 6.13e-16
c27226 595 907 3.15e-16
c27227 602 890 3.15e-16
c27228 632 3480 1.58e-16
c27229 2815 2804 1.58e-16
c27230 1779 1778 1.6e-16
c27231 982 0 1.8851e-14
c27232 2713 3226 1.532e-15
c27233 3231 3232 5.65e-16
c27234 19 259 8.4e-16
c27235 601 1681 1.75e-16
c27236 595 1682 2.22e-16
c27237 4302 662 1.58e-16
c27238 4844 5072 5.37e-16
c27239 2819 2452 1.58e-16
c27240 883 1007 3.92e-16
c27241 890 1006 1.88e-16
c27242 3355 868 2.22e-16
c27243 3757 3758 1.6e-16
c27244 4109 4108 7.81e-16
c27245 4567 4859 1.58e-16
c27246 4582 4469 1.58e-16
c27247 4821 120 6.4e-16
c27248 3251 1 6.15e-16
c27249 2738 2356 2.48e-16
c27250 2971 2970 1.6e-16
c27251 3548 3537 1.58e-16
c27252 1834 707 2.33e-16
c27253 1708 842 3.15e-16
c27254 2742 2739 5.5e-16
c27255 642 1380 1.813e-15
c27256 3219 1 5.97e-15
c27257 3141 2628 1.532e-15
c27258 2793 782 1.58e-16
c27259 1694 1380 5.5e-16
c27260 3606 777 1.58e-16
c27261 1324 0 8.2949e-14
c27262 2708 707 1.58e-16
c27263 2178 842 3.15e-16
c27264 3390 3404 6.4e-16
c27265 602 2211 1.09e-16
c27266 1858 0 6.72e-16
c27267 3393 3540 1.58e-16
c27268 3409 3157 1.58e-16
c27269 3676 3678 2.15e-16
c27270 3685 3686 1.6e-16
c27271 4751 1 6.42e-16
c27272 3237 752 7.68e-16
c27273 2165 1694 6.18e-16
c27274 1023 662 1.58e-16
c27275 592 715 6.34e-16
c27276 279 274 1.482e-15
c27277 1 127 4.22e-16
c27278 245 291 1.88e-16
c27279 657 3134 2.22e-16
c27280 3397 722 3.15e-16
c27281 4793 381 1.88e-16
c27282 3838 3836 1.167e-15
c27283 1321 1041 1.58e-16
c27284 1327 1031 5.88e-16
c27285 506 516 8.86e-16
c27286 528 526 1.96e-16
c27287 3049 3031 1.94e-16
c27288 3023 3043 2.07e-16
c27289 2686 707 1.339e-15
c27290 2182 842 3.15e-16
c27291 1987 852 5.73e-16
c27292 1831 1829 1.6e-16
c27293 1211 1644 1.58e-16
c27294 537 59 1.88e-16
c27295 4007 1 6.03e-16
c27296 3024 3224 3.92e-16
c27297 4830 4828 1.687e-15
c27298 4833 4840 6.73e-16
c27299 3230 752 5.03e-16
c27300 77 88 3.84e-16
c27301 617 1755 1.58e-16
c27302 777 1331 7.99e-16
c27303 27 18 1.58e-16
c27304 3409 717 3.15e-16
c27305 4580 4282 1.58e-16
c27306 5385 1 1.81e-16
c27307 2436 2430 1.6e-16
c27308 1913 2427 2.386e-15
c27309 1919 2435 1.136e-15
c27310 1930 2410 1.58e-16
c27311 3589 752 1.339e-15
c27312 2816 1 1.868e-15
c27313 894 1141 1.58e-16
c27314 907 1113 3.54e-16
c27315 2724 2333 4.11e-16
c27316 2806 0 2.93e-15
c27317 1863 722 7.68e-16
c27318 642 1387 1.58e-16
c27319 3751 3747 1.64e-16
c27320 4168 37 5.71e-16
c27321 3303 3294 3.46e-16
c27322 1651 1181 1.96e-16
c27323 1646 1191 1.96e-16
c27324 4333 4714 5.66e-16
c27325 4720 4711 3.92e-16
c27326 617 1733 1.339e-15
c27327 822 1161 4e-16
c27328 1500 1 1.868e-15
c27329 1490 0 2.93e-15
c27330 3898 777 3.15e-16
c27331 4540 0 3.8805e-14
c27332 565 262 1.88e-16
c27333 4899 1 1.23e-16
c27334 5353 5350 1.18e-15
c27335 1104 752 1.58e-16
c27336 4172 4166 1.96e-16
c27337 223 0 1.09879e-13
c27338 4872 294 1.88e-16
c27339 2194 2004 1.58e-16
c27340 1576 797 1.58e-16
c27341 1396 1387 3.46e-16
c27342 2545 2265 5.5e-16
c27343 367 1 9.8e-16
c27344 1345 1610 1.58e-16
c27345 687 1345 3.58e-16
c27346 3118 3112 1.6e-16
c27347 2594 3109 2.386e-15
c27348 2611 3092 1.58e-16
c27349 1533 1905 1.58e-16
c27350 3489 647 1.832e-15
c27351 4892 1 9.72e-16
c27352 822 1954 1.58e-16
c27353 4823 4822 1.6e-16
c27354 2408 1 1.716e-15
c27355 9 291 5.8e-16
c27356 4810 4813 6.02e-16
c27357 4582 4826 3.92e-16
c27358 0 294 1.24426e-13
c27359 5484 0 3.974e-14
c27360 3882 722 3.15e-16
c27361 4702 5335 1.96e-16
c27362 2794 2793 5.65e-16
c27363 632 983 1.58e-16
c27364 2518 0 5.4517e-14
c27365 1087 1 3.54e-16
c27366 1964 842 1.58e-16
c27367 2483 827 1.09e-16
c27368 1084 0 9.602e-15
c27369 3048 3172 5.42e-16
c27370 3024 3160 1.58e-16
c27371 1631 0 6.72e-16
c27372 792 1151 4.21e-16
c27373 0 545 1.4803e-14
c27374 448 451 2.142e-15
c27375 461 419 9.5e-16
c27376 3411 662 3.15e-16
c27377 5338 1 1.257e-15
c27378 910 2166 1.58e-16
c27379 1162 812 6.38e-16
c27380 981 988 7.95e-16
c27381 397 262 1.88e-16
c27382 4261 4254 6.73e-16
c27383 4260 3418 1.96e-16
c27384 5388 5286 1.58e-16
c27385 4861 91 1.88e-16
c27386 2606 2603 5.5e-16
c27387 612 610 3.327e-15
c27388 1456 1457 2.48e-16
c27389 3882 4502 1.96e-16
c27390 3935 1 6.66e-16
c27391 2398 752 1.09e-16
c27392 1533 1086 1.136e-15
c27393 886 893 5.5e-16
c27394 480 484 1.58e-16
c27395 485 477 2.218e-15
c27396 500 499 3.84e-16
c27397 3476 3475 5.65e-16
c27398 3470 3083 1.532e-15
c27399 3557 732 1.58e-16
c27400 5125 1 7.49e-16
c27401 2321 1811 1.96e-16
c27402 1983 1 9.28e-16
c27403 4776 5158 2.69e-16
c27404 5284 5335 1.191e-15
c27405 2773 2390 7.84e-16
c27406 4175 857 1.88e-16
c27407 4134 3918 2.48e-16
c27408 601 3438 1.832e-15
c27409 1121 1119 1.931e-15
c27410 106 105 2.84e-16
c27411 107 102 1.88e-16
c27412 3900 4302 1.58e-16
c27413 4736 381 1.88e-16
c27414 1241 1240 1.65e-16
c27415 922 921 4.274e-15
c27416 3909 26 4.48e-16
c27417 1618 858 1.58e-16
c27418 81 19 8.82e-16
c27419 368 363 1.88e-16
c27420 3034 3343 4.63e-16
c27421 3024 702 3.15e-16
c27422 2226 2233 6.73e-16
c27423 1936 1937 1.35e-16
c27424 2072 2077 3.54e-16
c27425 223 219 1.58e-16
c27426 3397 3089 1.58e-16
c27427 4657 4660 6.02e-16
c27428 4563 4378 5.88e-16
c27429 4571 4384 1.58e-16
c27430 997 998 7.46e-16
c27431 592 625 6.34e-16
c27432 3385 3875 1.62e-16
c27433 4044 4052 6.67e-16
c27434 4050 4040 7.1e-16
c27435 3983 857 1.88e-16
c27436 3321 3676 1.58e-16
c27437 3886 692 3.15e-16
c27438 5484 5486 1.001e-15
c27439 5482 5479 3.54e-16
c27440 5422 5434 3.18e-16
c27441 3144 0 6.62e-16
c27442 1046 1049 6.13e-16
c27443 4328 4322 1.6e-16
c27444 2283 647 3.64e-16
c27445 919 1070 3.92e-16
c27446 922 1069 2.54e-16
c27447 3509 1 2.054e-15
c27448 1927 767 1.09e-16
c27449 1345 1402 3.92e-16
c27450 3718 868 2.22e-16
c27451 2577 3091 4.97e-16
c27452 3511 0 8e-16
c27453 2956 2954 3.73e-16
c27454 3721 1 1.056e-15
c27455 3024 2804 1.58e-16
c27456 3030 2798 5.88e-16
c27457 1601 1596 1.642e-15
c27458 4658 1 1.806e-15
c27459 2668 717 5.73e-16
c27460 3034 2617 1.58e-16
c27461 2535 868 3.15e-16
c27462 2559 827 3.15e-16
c27463 2078 2070 4.48e-16
c27464 5197 5199 9.16e-16
c27465 3409 3450 1.58e-16
c27466 3542 3540 2.15e-16
c27467 3550 3549 1.6e-16
c27468 5025 5108 1.67e-16
c27469 5452 5491 1.858e-15
c27470 602 2529 1.58e-16
c27471 612 2532 5.73e-16
c27472 2966 0 2.078e-15
c27473 922 717 3.15e-16
c27474 971 967 3.78e-16
c27475 1343 1372 1.58e-16
c27476 4140 4148 6.67e-16
c27477 4146 4136 7.1e-16
c27478 2635 662 1.339e-15
c27479 3745 0 2.078e-15
c27480 4070 25 3.84e-16
c27481 4403 4402 2.03e-16
c27482 4408 4406 1.6e-16
c27483 2557 2751 1.58e-16
c27484 2541 2739 1.58e-16
c27485 2372 737 7.38e-16
c27486 3046 2645 5.5e-16
c27487 3030 2628 5.88e-16
c27488 3355 0 5.7036e-14
c27489 1559 0 3.3846e-14
c27490 3535 3536 9.1e-16
c27491 3616 1 5.97e-15
c27492 5074 5069 7.37e-16
c27493 5108 5107 5.87e-16
c27494 5057 1 3.36e-16
c27495 4982 4972 8.28e-16
c27496 4993 4994 1.6e-16
c27497 3360 858 7.38e-16
c27498 2294 2300 1.6e-16
c27499 1794 2274 1.58e-16
c27500 2151 0 3.8836e-14
c27501 777 1706 3.15e-16
c27502 883 702 3.15e-16
c27503 5045 0 2.156e-15
c27504 1678 2215 4.36e-16
c27505 687 3506 1.58e-16
c27506 1327 807 4.03e-16
c27507 3298 0 3.466e-15
c27508 601 3030 3.15e-16
c27509 910 3381 1.58e-16
c27510 4617 5409 9.82e-16
c27511 4623 5425 8.41e-16
c27512 2854 2853 9.1e-16
c27513 2559 2333 5.5e-16
c27514 3397 822 7.99e-16
c27515 3854 0 3.26e-15
c27516 1604 1602 1.6e-16
c27517 1327 1538 1.96e-16
c27518 1389 1 5.808e-15
c27519 2810 807 1.58e-16
c27520 3645 792 1.58e-16
c27521 4196 4215 1.922e-15
c27522 4564 4214 8.97e-16
c27523 1876 1873 3.01e-16
c27524 1872 1869 6.44e-16
c27525 1391 0 3.466e-15
c27526 2838 852 5.73e-16
c27527 642 2240 1.58e-16
c27528 3034 3279 1.58e-16
c27529 2179 2189 5.8e-16
c27530 2031 2044 1.138e-15
c27531 3219 3225 1.418e-15
c27532 3606 3608 1.862e-15
c27533 4606 4608 4.93e-16
c27534 5436 1 7.87e-16
c27535 4742 0 3.2607e-13
c27536 5136 5139 3.54e-16
c27537 4878 31 5.88e-16
c27538 3236 3208 2.64e-16
c27539 2485 2476 3.46e-16
c27540 2900 1 8.09e-16
c27541 2194 1732 1.58e-16
c27542 2756 2759 5.5e-16
c27543 1690 722 3.15e-16
c27544 3487 1 1.716e-15
c27545 1689 1324 7.67e-16
c27546 3061 3058 5.5e-16
c27547 1163 0 1.4198e-14
c27548 617 920 3.69e-16
c27549 4491 4487 1.96e-16
c27550 4747 4367 1.96e-16
c27551 2559 812 3.15e-16
c27552 138 132 1.372e-15
c27553 465 37 1.88e-16
c27554 9 484 5.8e-16
c27555 3608 3607 2.48e-16
c27556 2469 822 2.22e-16
c27557 1817 1 4.41e-15
c27558 2326 0 6.62e-16
c27559 855 854 1.6e-16
c27560 1440 677 1.58e-16
c27561 907 1187 3.92e-16
c27562 858 868 2.77e-16
c27563 102 1 1.0533e-14
c27564 71 15 5.8e-16
c27565 2766 2759 6.73e-16
c27566 2894 0 1.65e-16
c27567 2691 1 2.054e-15
c27568 612 2559 3.58e-16
c27569 919 677 3.15e-16
c27570 920 1008 1.58e-16
c27571 1331 1340 1.58e-16
c27572 3731 3733 3.54e-16
c27573 2576 2567 3.46e-16
c27574 601 890 3.15e-16
c27575 2815 3339 4.36e-16
c27576 2747 777 1.813e-15
c27577 4743 4744 2.03e-16
c27578 1708 1968 5.42e-16
c27579 1684 1956 1.58e-16
c27580 3145 3141 1.96e-16
c27581 762 1545 1.58e-16
c27582 601 2232 3.64e-16
c27583 602 1726 1.58e-16
c27584 4319 672 1.58e-16
c27585 4861 5106 4.06e-16
c27586 4922 5148 5.74e-16
c27587 2824 2452 1.58e-16
c27588 2669 1 1.716e-15
c27589 883 1021 1.88e-16
c27590 907 1014 1.58e-16
c27591 4567 4876 1.58e-16
c27592 4514 4877 1.96e-16
c27593 1343 767 4.46e-16
c27594 1353 1 1.716e-15
c27595 3882 822 4.03e-16
c27596 4223 1 4.64e-16
c27597 2172 858 4.48e-16
c27598 612 2225 2.72e-16
c27599 4768 1 6.42e-16
c27600 2730 737 3.15e-16
c27601 2478 1 5.808e-15
c27602 842 832 6.38e-16
c27603 3868 858 7.12e-16
c27604 5578 0 7.67e-16
c27605 2480 0 3.466e-15
c27606 1525 737 1.832e-15
c27607 919 1128 1.58e-16
c27608 5440 5442 1.77e-15
c27609 2545 2486 5.5e-16
c27610 2739 2746 1.96e-16
c27611 1694 692 3.15e-16
c27612 1345 1056 1.58e-16
c27613 1343 1046 5.5e-16
c27614 1331 1503 1.58e-16
c27615 3786 1 1.257e-15
c27616 4361 4356 1.642e-15
c27617 2512 858 9.97e-16
c27618 2525 852 3.64e-16
c27619 1137 0 6.29e-16
c27620 777 1113 1.05e-15
c27621 3313 3315 2.15e-16
c27622 3678 3674 1.96e-16
c27623 4776 207 5.88e-16
c27624 5079 91 4.88e-16
c27625 0 270 2.87e-16
c27626 1420 672 1.58e-16
c27627 166 0 1.0822e-14
c27628 129 37 1.88e-16
c27629 4285 4297 2.32e-16
c27630 5449 5454 3.07e-16
c27631 534 535 1.482e-15
c27632 3038 3027 4.097e-15
c27633 3410 1 2.471e-15
c27634 3031 3041 5.8e-16
c27635 1482 722 3.15e-16
c27636 1873 732 2.72e-16
c27637 2946 2929 1.96e-16
c27638 2931 2933 7.3e-16
c27639 2421 767 4.81e-16
c27640 3030 3023 1.58e-16
c27641 3048 3043 1.58e-16
c27642 4344 4723 1.58e-16
c27643 1694 1539 1.58e-16
c27644 1811 1783 2.64e-16
c27645 5157 5174 1.443e-15
c27646 449 451 1.58e-16
c27647 430 419 2.45e-16
c27648 331 332 1.482e-15
c27649 3876 792 3.15e-16
c27650 2361 1845 4.11e-16
c27651 400 1 1.44e-16
c27652 223 217 3.84e-16
c27653 2814 2418 1.96e-16
c27654 4071 4079 9.33e-16
c27655 4072 4070 3.54e-16
c27656 4787 0 3.5424e-13
c27657 4640 33 1.88e-16
c27658 1402 1401 9.1e-16
c27659 3972 37 1.88e-16
c27660 4377 4368 3.46e-16
c27661 1327 1176 1.58e-16
c27662 4370 1 5.808e-15
c27663 4630 4628 1.6e-16
c27664 1708 1731 3.92e-16
c27665 204 194 3.75e-16
c27666 4372 0 3.466e-15
c27667 2987 2882 1.58e-16
c27668 3393 3304 5.88e-16
c27669 4889 4882 2.67e-16
c27670 5285 352 3.54e-16
c27671 88 450 1.88e-16
c27672 3718 0 6.0716e-14
c27673 2150 2149 1.6e-16
c27674 11 27 1.58e-16
c27675 1 31 3.53e-16
c27676 407 508 1.88e-16
c27677 2434 1 8.43e-16
c27678 1027 677 6.38e-16
c27679 3338 837 2.22e-16
c27680 3387 827 4.48e-16
c27681 3409 842 4.46e-16
c27682 4582 4843 3.92e-16
c27683 2718 2350 1.96e-16
c27684 777 26 1.58e-16
c27685 378 479 1.88e-16
c27686 3983 3975 9.33e-16
c27687 3876 737 4.48e-16
c27688 4872 62 1.88e-16
c27689 1251 1250 1.96e-16
c27690 1218 907 1.96e-16
c27691 632 1005 6.48e-16
c27692 2535 0 3.17834e-13
c27693 921 1115 1.96e-16
c27694 2929 2492 1.958e-15
c27695 2541 2407 1.58e-16
c27696 2717 2718 9.1e-16
c27697 1567 782 3.15e-16
c27698 1754 1369 1.96e-16
c27699 1106 1542 1.58e-16
c27700 3874 4612 2.196e-15
c27701 3191 0 3.6368e-14
c27702 2541 3017 2e-16
c27703 4167 1 6.03e-16
c27704 4152 19 7.35e-16
c27705 4892 4890 1.6e-16
c27706 4429 4812 4.97e-16
c27707 3224 722 1.58e-16
c27708 3048 3177 1.58e-16
c27709 2145 2133 8.94e-16
c27710 1806 0 1.4092e-14
c27711 5230 5198 1.75e-16
c27712 1 582 4.92e-16
c27713 0 505 9.795e-15
c27714 306 304 1.58e-16
c27715 37 519 1.88e-16
c27716 33 526 2.52e-16
c27717 2409 2410 2.48e-16
c27718 5347 0 2.285e-15
c27719 62 0 1.30646e-13
c27720 65 30 6.83e-16
c27721 73 27 1.88e-16
c27722 642 3393 4.03e-16
c27723 3429 3418 1.58e-16
c27724 4368 732 1.58e-16
c27725 1099 1100 7.51e-16
c27726 3008 3006 1.6e-16
c27727 3898 4519 3.92e-16
c27728 4437 4438 2.48e-16
c27729 2559 2786 3.92e-16
c27730 4571 647 1.33e-16
c27731 687 1822 2.72e-16
c27732 2843 842 5.03e-16
c27733 687 19 1.41e-15
c27734 3577 732 1.58e-16
c27735 5277 323 3.54e-16
c27736 1996 1 6.15e-16
c27737 3387 3276 1.58e-16
c27738 5039 0 5.8525e-14
c27739 2243 2240 5.5e-16
c27740 1087 1068 1.546e-15
c27741 907 904 1.58e-16
c27742 2603 2610 1.96e-16
c27743 3616 3225 1.136e-15
c27744 617 3438 1.58e-16
c27745 1131 1133 7.72e-16
c27746 4231 4232 1.35e-16
c27747 5587 5591 1.96e-16
c27748 4567 4563 4.431e-15
c27749 4657 5491 7.98e-16
c27750 2541 2773 1.58e-16
c27751 3211 747 1.58e-16
c27752 3158 0 1.6491e-14
c27753 2535 2203 1.58e-16
c27754 2541 2170 5.5e-16
c27755 3177 3179 2.15e-16
c27756 4326 1 8.43e-16
c27757 4505 0 2.93e-15
c27758 1912 1516 1.96e-16
c27759 1907 1522 1.96e-16
c27760 822 1690 4.03e-16
c27761 890 886 8.76e-16
c27762 1 566 1.65e-15
c27763 3387 812 4.48e-16
c27764 4563 4395 5.88e-16
c27765 4571 4401 1.58e-16
c27766 5506 1 3.36e-16
c27767 2373 1 4.41e-15
c27768 2587 0 6.62e-16
c27769 2505 2504 1.6e-16
c27770 2497 2495 2.15e-16
c27771 3159 0 2.93e-15
c27772 2300 672 2.65e-16
c27773 1327 1572 1.96e-16
c27774 822 820 3.327e-15
c27775 612 3387 3.15e-16
c27776 2559 747 3.58e-16
c27777 3659 822 1.58e-16
c27778 3527 0 6.72e-16
c27779 858 0 2.79654e-13
c27780 2957 2978 1.96e-16
c27781 3363 3362 1.6e-16
c27782 3048 2821 1.58e-16
c27783 3046 2815 5.5e-16
c27784 2474 837 2.4e-16
c27785 4675 1 1.806e-15
c27786 4401 4779 7.84e-16
c27787 3203 717 2.65e-16
c27788 1784 0 1.6491e-14
c27789 453 465 1.58e-16
c27790 15 204 5.8e-16
c27791 3625 3623 1.862e-15
c27792 3409 3455 1.58e-16
c27793 3769 3772 3.54e-16
c27794 3974 857 1.88e-16
c27795 3935 3934 5.5e-16
c27796 5489 0 2.078e-15
c27797 5388 323 1.58e-16
c27798 5025 5133 1.58e-16
c27799 2776 2773 5.5e-16
c27800 612 3084 2.65e-16
c27801 601 2529 1.58e-16
c27802 2559 2384 5.5e-16
c27803 4241 4232 3.46e-16
c27804 1345 1401 5.42e-16
c27805 1321 1389 1.58e-16
c27806 2596 2595 1.6e-16
c27807 1191 1192 8.58e-16
c27808 687 4317 1.58e-16
c27809 3898 4455 1.58e-16
c27810 3876 4467 1.58e-16
c27811 4518 4519 9.1e-16
c27812 602 1341 1.58e-16
c27813 3582 4400 1.96e-16
c27814 853 1 1.65e-16
c27815 590 589 1.96e-16
c27816 3158 3169 1.96e-16
c27817 1579 0 1.4092e-14
c27818 4483 1 1.056e-15
c27819 2541 692 3.15e-16
c27820 1971 1590 3.92e-16
c27821 1975 1976 1.6e-16
c27822 4571 4570 2.14e-16
c27823 4582 4577 1.58e-16
c27824 5072 5103 1.58e-16
c27825 3459 3457 1.6e-16
c27826 3454 3453 2.03e-16
c27827 792 1684 3.15e-16
c27828 113 117 1.58e-16
c27829 5405 5404 5.87e-16
c27830 5388 5301 4.2e-16
c27831 632 2557 4.46e-16
c27832 2741 0 3.466e-15
c27833 2534 1 2.259e-15
c27834 1682 1678 1.58e-16
c27835 792 1935 2.4e-16
c27836 687 3526 1.58e-16
c27837 3690 3691 1.35e-16
c27838 5151 149 5.11e-16
c27839 2584 2593 3.46e-16
c27840 1431 662 3.15e-16
c27841 3690 842 2.33e-16
c27842 602 3423 1.9e-16
c27843 3318 0 8e-16
c27844 3137 1 1.056e-15
c27845 617 3030 3.15e-16
c27846 2860 2856 1.96e-16
c27847 3886 3446 5.5e-16
c27848 3158 3162 1.96e-16
c27849 1409 1 2.054e-15
c27850 1411 0 8e-16
c27851 175 194 1.88e-16
c27852 2849 827 1.58e-16
c27853 4143 857 1.88e-16
c27854 4623 4630 1.81e-16
c27855 2475 2469 1.418e-15
c27856 2172 2410 1.58e-16
c27857 922 842 5.14e-16
c27858 921 1173 1.58e-16
c27859 4423 767 5.03e-16
c27860 1684 737 4.48e-16
c27861 642 2238 1.58e-16
c27862 4083 1 6.78e-16
c27863 1745 1 9.28e-16
c27864 2764 752 1.58e-16
c27865 2679 677 1.58e-16
c27866 1652 2019 1.58e-16
c27867 4708 4709 9.93e-16
c27868 3387 3406 1.58e-16
c27869 3393 3383 3.54e-16
c27870 3411 3407 3.92e-16
c27871 2351 1 1.868e-15
c27872 596 605 5.28e-16
c27873 2341 0 2.93e-15
c27874 1670 1 1.286e-15
c27875 5239 1 2.429e-15
c27876 1460 677 1.58e-16
c27877 1209 852 1.58e-16
c27878 5452 5471 4.78e-16
c27879 3879 3881 1.041e-15
c27880 2654 2653 2.48e-16
c27881 627 2559 3.58e-16
c27882 3117 1 5.97e-15
c27883 1331 880 1.58e-16
c27884 2427 797 1.58e-16
c27885 1784 1795 1.96e-16
c27886 617 890 3.15e-16
c27887 4065 0 7.8627e-14
c27888 4056 26 1.075e-15
c27889 3034 3105 4.63e-16
c27890 4592 1 4.832e-15
c27891 2029 2025 6.9e-16
c27892 1708 1973 1.58e-16
c27893 1862 2385 4.36e-16
c27894 2383 2376 1.96e-16
c27895 3525 692 5.03e-16
c27896 5360 354 1.345e-15
c27897 4903 4899 6.9e-16
c27898 4977 4531 9.58e-16
c27899 2274 2273 2.48e-16
c27900 627 1732 1.58e-16
c27901 617 2232 7.68e-16
c27902 601 1726 3.15e-16
c27903 2844 2452 2.38e-15
c27904 2695 1 8.43e-16
c27905 911 2532 1.88e-16
c27906 894 677 3.15e-16
c27907 890 1008 3.54e-16
c27908 909 1029 1.58e-16
c27909 4119 4118 1.58e-16
c27910 4567 4893 1.58e-16
c27911 4514 4894 1.96e-16
c27912 1345 782 3.15e-16
c27913 1333 1332 6.97e-16
c27914 1334 1330 1.71e-16
c27915 4389 4387 2.15e-16
c27916 4397 4396 1.6e-16
c27917 3631 1 6.15e-16
c27918 3865 0 1.1956e-14
c27919 537 407 1.88e-16
c27920 2799 797 7.68e-16
c27921 2987 2969 1.58e-16
c27922 1505 1 4.41e-15
c27923 5277 265 5.11e-16
c27924 3839 5018 9.36e-16
c27925 1889 0 6.62e-16
c27926 3409 3185 5.5e-16
c27927 4785 1 6.42e-16
c27928 1 481 4.22e-16
c27929 15 456 4.88e-16
c27930 687 3134 1.813e-15
c27931 4112 4110 1.76e-16
c27932 458 0 1.4803e-14
c27933 3879 3390 1.96e-16
c27934 627 2584 1.58e-16
c27935 1309 1236 5.5e-16
c27936 2566 0 3.5325e-14
c27937 911 945 2.135e-15
c27938 2770 2771 1.35e-16
c27939 617 986 3.57e-16
c27940 1835 1454 3.92e-16
c27941 1839 1840 1.6e-16
c27942 4471 4473 2.03e-16
c27943 792 1133 1.58e-16
c27944 3219 3587 1.96e-16
c27945 4745 0 3.4656e-14
c27946 15 175 5.8e-16
c27947 3393 732 4.03e-16
c27948 4580 4316 1.58e-16
c27949 0 158 4.512e-14
c27950 3355 3775 1.19e-16
c27951 5173 1 2.424e-15
c27952 2852 1 1.056e-15
c27953 2178 2177 3.15e-16
c27954 1016 662 3.15e-16
c27955 894 1128 3.54e-16
c27956 2746 2737 3.46e-16
c27957 911 924 4.5e-16
c27958 134 129 1.482e-15
c27959 3038 3029 5.71e-16
c27960 4183 4184 6.4e-16
c27961 632 1408 1.9e-16
c27962 3419 0 1.6491e-14
c27963 3616 3622 1.418e-15
c27964 4453 4455 1.862e-15
c27965 968 1 4.59e-16
c27966 3315 3311 1.96e-16
c27967 965 0 1.2487e-14
c27968 4008 0 2.0592e-14
c27969 3396 3038 5.8e-16
c27970 2713 3207 1.96e-16
c27971 1663 1206 2.91e-16
c27972 1665 1664 1.6e-16
c27973 1518 1 9.28e-16
c27974 4350 4731 5.66e-16
c27975 4737 4728 3.92e-16
c27976 5388 265 6.06e-16
c27977 5029 5031 1.441e-15
c27978 5049 5047 3.92e-16
c27979 2182 2177 1.58e-16
c27980 846 835 7.23e-16
c27981 838 839 1.6e-16
c27982 911 2559 3.45e-16
c27983 910 2535 5.22e-16
c27984 1118 752 3.57e-16
c27985 1098 1111 1.58e-16
c27986 5326 5366 4.39e-16
c27987 2637 0 3.3485e-14
c27988 1408 1404 1.96e-16
c27989 642 3446 1.813e-15
c27990 2545 2650 4.63e-16
c27991 3387 747 3.15e-16
c27992 1931 1539 1.96e-16
c27993 1932 1925 6.73e-16
c27994 5010 5007 5.5e-16
c27995 3565 747 1.813e-15
c27996 3024 3046 4.078e-15
c27997 3048 3030 4.312e-15
c27998 595 2173 9.02e-16
c27999 4571 4299 1.58e-16
c28000 5277 5350 1.03e-16
c28001 3411 852 3.58e-16
c28002 2731 2339 1.96e-16
c28003 596 682 3.134e-15
c28004 3554 3555 1.35e-16
c28005 3798 3781 1.96e-16
c28006 3991 3992 6.4e-16
c28007 1071 1072 8.58e-16
c28008 920 1129 1.58e-16
c28009 2557 2424 1.58e-16
c28010 3030 2685 1.58e-16
c28011 1653 1 1.868e-15
c28012 3658 3660 2.03e-16
c28013 4827 4828 9.93e-16
c28014 1643 0 2.93e-15
c28015 3202 3569 1.58e-16
c28016 2410 0 3.3692e-14
c28017 0 305 9.4544e-14
c28018 3975 3974 1.58e-16
c28019 5543 526 4.02e-16
c28020 4844 439 1.88e-16
c28021 5355 294 5.5e-16
c28022 2354 2355 9.1e-16
c28023 4275 4268 1.96e-16
c28024 3429 4277 4.36e-16
c28025 3579 0 8e-16
c28026 617 4249 1.339e-15
c28027 3886 4349 4.63e-16
c28028 3046 762 3.15e-16
c28029 2900 2896 6.35e-16
c28030 912 1 2.86e-16
c28031 3203 3194 3.92e-16
c28032 2685 3197 5.66e-16
c28033 2696 3189 1.58e-16
c28034 3574 3576 2.15e-16
c28035 2863 842 1.09e-16
c28036 2290 1783 2.48e-16
c28037 1618 2002 1.58e-16
c28038 1690 1901 1.96e-16
c28039 199 195 1.372e-15
c28040 2242 0 3.466e-15
c28041 3411 3293 1.58e-16
c28042 1107 737 4.98e-16
c28043 919 924 3.54e-16
c28044 922 925 1.96e-16
c28045 3 1 4.22e-16
c28046 9 13 5.8e-16
c28047 4640 526 1.88e-16
c28048 617 3458 1.58e-16
c28049 3926 19 7.04e-16
c28050 4600 64 1.88e-16
c28051 2559 2220 1.58e-16
c28052 2557 2214 5.5e-16
c28053 2545 2615 1.58e-16
c28054 896 0 5.86e-16
c28055 872 25 7.64e-16
c28056 4429 3588 1.136e-15
c28057 1706 1704 1.96e-16
c28058 1690 1703 1.58e-16
c28059 1708 1711 1.6e-16
c28060 477 476 1.482e-15
c28061 535 577 1.88e-16
c28062 4470 822 1.58e-16
c28063 3046 3359 1.58e-16
c28064 3030 3347 1.58e-16
c28065 3185 2668 1.136e-15
c28066 3474 647 5.03e-16
c28067 5113 0 3.4847e-14
c28068 2240 2247 1.96e-16
c28069 4850 0 1.4233e-14
c28070 2610 2601 3.46e-16
c28071 2103 1658 6.55e-16
c28072 2127 2072 3.18e-16
c28073 223 565 1.88e-16
c28074 4563 4412 5.88e-16
c28075 4571 4418 1.58e-16
c28076 2196 2491 3.92e-16
c28077 4063 4054 1.96e-16
c28078 2804 822 1.58e-16
c28079 4007 857 6.23e-16
c28080 74 1 1.65e-15
c28081 4464 782 3.64e-16
c28082 5517 5515 3.92e-16
c28083 3209 747 1.58e-16
c28084 1794 672 3.79e-16
c28085 1343 1589 3.92e-16
c28086 627 3387 3.15e-16
c28087 3679 822 1.58e-16
c28088 1549 1091 1.96e-16
c28089 1544 1101 1.96e-16
c28090 4591 3873 2.48e-16
c28091 2999 2136 3.54e-16
c28092 2955 2518 2.037e-15
c28093 4132 1 2.259e-15
c28094 3024 2832 5.5e-16
c28095 2663 662 3.64e-16
c28096 762 907 3.15e-16
c28097 4863 4862 2.03e-16
c28098 4692 1 1.806e-15
c28099 2696 717 3.79e-16
c28100 2103 2070 1.58e-16
c28101 1 326 5.62e-16
c28102 233 219 1.58e-16
c28103 5224 5234 1.125e-15
c28104 3555 3566 1.96e-16
c28105 523 519 1.58e-16
c28106 0 340 1.0822e-14
c28107 3397 672 7.99e-16
c28108 3992 3907 1.88e-16
c28109 4582 4196 5.5e-16
c28110 5293 412 5.93e-16
c28111 4922 352 1.88e-16
c28112 762 2396 1.58e-16
c28113 1896 2389 1.96e-16
c28114 2194 1760 5.5e-16
c28115 883 907 4.078e-15
c28116 909 890 4.312e-15
c28117 1234 1235 1.96e-16
c28118 5514 5461 9.01e-16
c28119 3719 842 3.64e-16
c28120 4372 707 1.9e-16
c28121 601 3086 4.81e-16
c28122 612 2577 3.79e-16
c28123 1160 797 5.74e-16
c28124 3657 822 1.58e-16
c28125 4247 4246 9.1e-16
c28126 1345 1406 1.58e-16
c28127 1646 858 5.03e-16
c28128 1196 1193 1.984e-15
c28129 59 52 3.54e-16
c28130 3876 4472 1.58e-16
c28131 3900 4484 5.42e-16
c28132 2435 827 1.58e-16
c28133 2656 662 1.9e-16
c28134 595 880 1.58e-16
c28135 2559 2756 1.58e-16
c28136 1038 0 4.6723e-14
c28137 4120 19 7.35e-16
c28138 3030 3139 1.96e-16
c28139 4779 4781 2.15e-16
c28140 3006 852 1.58e-16
c28141 595 1704 2.13e-16
c28142 4111 3041 2.697e-15
c28143 4499 1 9.28e-16
c28144 2535 707 4.48e-16
c28145 2401 2396 1.642e-15
c28146 4938 4941 1.316e-15
c28147 4945 4936 1.873e-15
c28148 3411 3409 4.506e-15
c28149 2759 1 2.054e-15
c28150 657 2535 3.15e-16
c28151 3397 3242 1.58e-16
c28152 2761 0 8e-16
c28153 2580 1 1.056e-15
c28154 4136 4143 1.88e-16
c28155 3684 858 1.58e-16
c28156 601 3423 5.03e-16
c28157 3334 0 6.72e-16
c28158 2798 792 2.22e-16
c28159 3153 1 9.28e-16
c28160 2645 2254 1.136e-15
c28161 1355 1353 1.862e-15
c28162 3571 4407 5.66e-16
c28163 4413 4404 3.92e-16
c28164 2376 737 1.832e-15
c28165 3773 0 4.1103e-14
c28166 1608 1161 3.92e-16
c28167 1612 1613 1.6e-16
c28168 1345 1555 3.92e-16
c28169 1708 1431 5.5e-16
c28170 3096 3094 1.6e-16
c28171 1884 1499 1.96e-16
c28172 1769 1 5.808e-15
c28173 3411 3621 3.92e-16
c28174 5047 0 3.5057e-14
c28175 3265 782 1.84e-16
c28176 2218 2219 9.1e-16
c28177 4640 4648 1.81e-16
c28178 4685 439 1.88e-16
c28179 2551 0 5.86e-16
c28180 2288 2289 1.35e-16
c28181 978 979 1.21e-16
c28182 642 3034 7.99e-16
c28183 1331 647 3.15e-16
c28184 3686 1 9.28e-16
c28185 4443 767 1.09e-16
c28186 1990 827 1.832e-15
c28187 1343 1554 1.58e-16
c28188 1327 1542 1.58e-16
c28189 645 1 1.65e-16
c28190 2748 737 3.64e-16
c28191 1488 1871 7.84e-16
c28192 2194 752 4.46e-16
c28193 1799 1414 1.96e-16
c28194 3347 3356 3.92e-16
c28195 3350 2838 5.66e-16
c28196 2849 3342 1.58e-16
c28197 1758 1 6.15e-16
c28198 4764 4384 1.96e-16
c28199 3387 3021 1.58e-16
c28200 1845 1 5.97e-15
c28201 782 772 6.38e-16
c28202 15 436 5.8e-16
c28203 3236 767 3.15e-16
c28204 1203 868 1.58e-16
c28205 894 1202 3.92e-16
c28206 909 1201 1.88e-16
c28207 883 1194 1.58e-16
c28208 3898 647 4.46e-16
c28209 3882 672 4.03e-16
c28210 121 118 6.67e-16
c28211 59 218 1.88e-16
c28212 5391 5170 2.12e-16
c28213 922 1023 1.58e-16
c28214 4217 4208 2.45e-16
c28215 911 3387 1.88e-16
c28216 3489 0 3.3874e-14
c28217 2787 1 4.41e-15
c28218 1181 1180 3.94e-16
c28219 677 1 3.1284e-14
c28220 3886 3605 1.58e-16
c28221 2955 2966 1.96e-16
c28222 2435 812 3.15e-16
c28223 2447 797 1.58e-16
c28224 3357 3356 1.6e-16
c28225 4609 1 4.832e-15
c28226 1690 1607 1.58e-16
c28227 3630 767 1.09e-16
c28228 617 1726 3.15e-16
c28229 3545 692 1.09e-16
c28230 3350 842 1.58e-16
c28231 595 3025 9.02e-16
c28232 1141 1142 1.238e-15
c28233 88 26 8.41e-16
c28234 1421 1432 1.96e-16
c28235 2887 2915 4.39e-16
c28236 4004 1701 1.96e-16
c28237 2840 2842 2.03e-16
c28238 4040 25 7.01e-16
c28239 3900 4247 3.92e-16
c28240 1499 1494 1.642e-15
c28241 3582 0 6.9481e-14
c28242 3419 3430 1.96e-16
c28243 1914 1 1.868e-15
c28244 248 252 1.58e-16
c28245 2278 2276 1.6e-16
c28246 2273 2272 2.03e-16
c28247 4802 1 6.42e-16
c28248 4969 0 1.666e-15
c28249 1904 0 2.93e-15
c28250 4054 3918 2.48e-16
c28251 4922 294 1.88e-16
c28252 2822 2824 1.862e-15
c28253 687 1037 2.68e-16
c28254 4301 4300 2.03e-16
c28255 4306 4304 1.6e-16
c28256 5417 5414 1.96e-16
c28257 2518 2520 3.2e-16
c28258 783 0 7.86e-15
c28259 398 396 1.58e-16
c28260 384 383 3.84e-16
c28261 542 233 1.88e-16
c28262 2533 3020 1.58e-16
c28263 1128 1 1.56e-15
c28264 4245 1 1.056e-15
c28265 4566 4568 3.84e-16
c28266 4762 0 3.485e-14
c28267 1 365 4.22e-16
c28268 15 349 5.8e-16
c28269 3689 827 7.38e-16
c28270 146 132 1.58e-16
c28271 5410 5471 1.6e-16
c28272 2868 1 9.28e-16
c28273 5356 5360 1.96e-16
c28274 3882 3879 1.123e-15
c28275 1774 1771 3.01e-16
c28276 1770 1767 6.44e-16
c28277 990 1 3.06e-16
c28278 782 19 1.676e-15
c28279 3048 2529 1.58e-16
c28280 1531 1 6.15e-16
c28281 3143 662 1.832e-15
c28282 2053 2026 1.79e-16
c28283 2033 2030 2.208e-15
c28284 19 262 3.84e-16
c28285 5010 4954 1.826e-15
c28286 2086 1 1.257e-15
c28287 2873 352 1.952e-15
c28288 1330 898 5.8e-16
c28289 403 390 1.58e-16
c28290 281 233 1.88e-16
c28291 2826 2435 4.11e-16
c28292 5270 5044 1.666e-15
c28293 3789 3785 1.96e-16
c28294 1602 812 7.68e-16
c28295 1281 1303 7.53e-16
c28296 1293 1294 2.023e-15
c28297 1196 1657 1.96e-16
c28298 1345 1191 1.58e-16
c28299 1343 1181 5.5e-16
c28300 1331 1656 1.58e-16
c28301 4647 4645 1.6e-16
c28302 1550 1539 1.58e-16
c28303 508 252 1.88e-16
c28304 3506 3134 1.58e-16
c28305 4923 4889 1.301e-15
c28306 233 217 3.84e-16
c28307 285 274 2.45e-16
c28308 1 136 8.25e-15
c28309 403 37 1.88e-16
c28310 281 305 1.88e-16
c28311 4736 4350 1.179e-15
c28312 1040 662 1.58e-16
c28313 943 929 2.679e-15
c28314 3726 3739 5.78e-16
c28315 4014 3918 6.32e-16
c28316 3226 0 1.6491e-14
c28317 1510 737 5.03e-16
c28318 1076 1073 1.984e-15
c28319 5532 5533 3.54e-16
c28320 5514 5515 3.54e-16
c28321 2535 2441 1.58e-16
c28322 738 0 7.86e-15
c28323 1568 1116 1.96e-16
c28324 1569 1562 6.73e-16
c28325 4242 4629 2.196e-15
c28326 1289 0 2.285e-15
c28327 4184 1 5.1e-16
c28328 2987 2970 8.15e-16
c28329 2701 692 1.58e-16
c28330 4446 4829 4.97e-16
c28331 3046 2702 1.58e-16
c28332 1437 0 3.6368e-14
c28333 1196 1 5.194e-15
c28334 1 46 4.22e-16
c28335 15 5 5.8e-16
c28336 3393 3519 1.96e-16
c28337 3202 3574 1.58e-16
c28338 2430 0 1.4092e-14
c28339 26 37 3.001e-15
c28340 889 895 7.94e-16
c28341 0 30 2.66612e-13
c28342 27 25 5.71e-16
c28343 3689 812 1.58e-16
c28344 3041 0 5.5167e-14
c28345 4389 732 2.72e-16
c28346 3548 722 3.15e-16
c28347 4810 5270 5.5e-16
c28348 4844 5136 1.606e-15
c28349 1690 672 4.03e-16
c28350 1706 647 4.46e-16
c28351 919 964 1.58e-16
c28352 3595 0 6.72e-16
c28353 2248 2615 1.58e-16
c28354 3024 777 3.15e-16
c28355 2882 2909 2.84e-16
c28356 1112 0 1.0183e-14
c28357 938 1 1.65e-16
c28358 3992 1 5.1e-16
c28359 4168 0 2.0592e-14
c28360 3295 3297 2.03e-16
c28361 1735 1352 7.84e-16
c28362 1249 1667 4.79e-16
c28363 2696 3194 1.58e-16
c28364 627 1748 2.4e-16
c28365 4550 1 2.48e-16
c28366 309 308 2.84e-16
c28367 1678 1679 1.76e-16
c28368 747 1521 2.4e-16
c28369 0 574 6.224e-15
c28370 2262 0 8e-16
c28371 2892 3807 2.24e-16
c28372 3858 3859 1.6e-16
c28373 3866 3868 1.6e-16
c28374 3344 3857 2.91e-16
c28375 632 2583 1.75e-16
c28376 596 866 2.45e-16
c28377 4872 4867 1.536e-15
c28378 2620 2622 2.15e-16
c28379 2559 2790 1.58e-16
c28380 1388 1390 2.03e-16
c28381 1136 1132 3.78e-16
c28382 3886 4348 1.58e-16
c28383 3898 3497 5.5e-16
c28384 3900 3503 1.58e-16
c28385 2535 2231 5.5e-16
c28386 2545 2620 1.58e-16
c28387 1181 1639 1.58e-16
c28388 1690 1900 1.58e-16
c28389 3487 3488 2.03e-16
c28390 204 247 1.88e-16
c28391 2892 2905 3.18e-16
c28392 704 703 1.6e-16
c28393 570 568 1.257e-15
c28394 3494 647 1.09e-16
c28395 3409 3672 3.92e-16
c28396 3296 807 1.58e-16
c28397 3046 722 4.46e-16
c28398 3034 732 7.99e-16
c28399 4867 0 1.4233e-14
c28400 5351 5350 5.87e-16
c28401 3259 3642 7.84e-16
c28402 4563 4429 5.88e-16
c28403 4571 4435 1.58e-16
c28404 2510 1998 1.477e-15
c28405 1343 717 3.15e-16
c28406 1370 1372 1.862e-15
c28407 881 952 1.418e-15
c28408 5403 0 5.7679e-14
c28409 2048 1 1.031e-15
c28410 2178 2320 1.58e-16
c28411 1061 1060 3.94e-16
c28412 3633 782 3.15e-16
c28413 4685 5299 9.04e-16
c28414 686 1 5.57e-16
c28415 3174 1 4.41e-15
c28416 3107 3108 2.03e-16
c28417 4322 0 1.4092e-14
c28418 4525 3690 1.96e-16
c28419 4530 3684 1.96e-16
c28420 1203 0 4.6617e-14
c28421 777 883 3.15e-16
c28422 2247 2238 3.46e-16
c28423 4418 4796 7.84e-16
c28424 1 555 4.92e-16
c28425 657 2637 1.58e-16
c28426 592 652 1.96e-16
c28427 0 546 6.224e-15
c28428 3253 807 1.58e-16
c28429 4580 4604 1.58e-16
c28430 4776 497 1.88e-16
c28431 777 2401 3.79e-16
c28432 2182 2320 1.58e-16
c28433 627 2577 1.813e-15
c28434 2873 294 7.57e-16
c28435 2688 2686 1.862e-15
c28436 2305 2299 1.418e-15
c28437 2316 2288 2.64e-16
c28438 4253 4249 1.96e-16
c28439 3900 4489 1.58e-16
c28440 2452 868 1.58e-16
c28441 2478 837 1.58e-16
c28442 3271 3273 1.6e-16
c28443 3046 3156 3.92e-16
c28444 1721 1720 1.6e-16
c28445 747 752 2.77e-16
c28446 4512 1 6.15e-16
c28447 3184 2662 1.96e-16
c28448 1988 1601 1.532e-15
c28449 1994 1993 5.65e-16
c28450 1146 0 3.7577e-14
c28451 479 494 1.88e-16
c28452 33 207 1.88e-16
c28453 37 187 1.88e-16
c28454 2189 0 5.4993e-14
c28455 3435 3436 1.35e-16
c28456 1156 807 1.35e-16
c28457 907 722 4.8e-16
c28458 883 1082 3.92e-16
c28459 890 1081 1.88e-16
c28460 5286 5283 7.84e-16
c28461 5320 5322 3.25e-16
c28462 2785 2401 1.58e-16
c28463 642 596 1.96e-16
c28464 4555 858 7.12e-16
c28465 601 3443 1.09e-16
c28466 2886 2874 1.74e-16
c28467 3582 4404 1.58e-16
c28468 2384 752 3.15e-16
c28469 1717 1318 2.48e-16
c28470 848 0 1.1394e-14
c28471 996 1 4.044e-15
c28472 1424 0 6.62e-16
c28473 4196 4564 7.37e-16
c28474 3464 3455 3.92e-16
c28475 3072 3458 5.66e-16
c28476 3083 3450 1.58e-16
c28477 642 2266 2.65e-16
c28478 627 1760 2.22e-16
c28479 77 0 1.5723e-14
c28480 4943 4946 9.03e-16
c28481 792 1939 1.58e-16
c28482 2558 0 1.4914e-14
c28483 3397 797 3.15e-16
c28484 4167 857 6.23e-16
c28485 4657 4662 5.53e-16
c28486 2178 1936 1.58e-16
c28487 1321 677 4.48e-16
c28488 3699 1 6.15e-16
c28489 5403 5486 1.67e-16
c28490 655 1 3.79e-16
c28491 648 0 7.86e-15
c28492 632 2259 1.9e-16
c28493 1499 1883 1.58e-16
c28494 4463 1 6.275e-15
c28495 2108 178 1.038e-15
c28496 1767 1 1.716e-15
c28497 3411 3055 1.58e-16
c28498 991 992 1.238e-15
c28499 592 607 1.96e-16
c28500 5213 5192 5.87e-16
c28501 1981 822 2.22e-16
c28502 2182 1936 1.58e-16
c28503 3545 3542 3.01e-16
c28504 3900 662 3.15e-16
c28505 1466 692 7.68e-16
c28506 1224 858 5.75e-16
c28507 894 1216 1.58e-16
c28508 907 1188 3.54e-16
c28509 2929 0 6.1551e-14
c28510 1453 1016 1.96e-16
c28511 4507 4505 2.03e-16
c28512 2634 677 1.75e-16
c28513 2736 3244 2.48e-16
c28514 3046 3121 1.58e-16
c28515 3030 3109 1.58e-16
c28516 3066 2532 1.136e-15
c28517 1562 1 2.054e-15
c28518 4626 1 4.832e-15
c28519 4378 4758 1.96e-16
c28520 2062 2066 3.82e-16
c28521 1564 0 8e-16
c28522 777 1568 2.65e-16
c28523 335 334 1.079e-15
c28524 136 363 1.88e-16
c28525 5232 1 3.914e-15
c28526 5072 5068 5.32e-16
c28527 2159 1 2.48e-16
c28528 3774 3775 6.26e-16
c28529 3879 3890 4.097e-15
c28530 5165 0 5.8577e-14
c28531 151 91 1.58e-16
c28532 537 252 1.88e-16
c28533 1151 827 1.58e-16
c28534 2541 2718 1.96e-16
c28535 1344 1338 1.988e-15
c28536 647 26 7.12e-16
c28537 803 0 1.1456e-14
c28538 175 247 1.88e-16
c28539 4999 4991 1.96e-16
c28540 4989 4992 3.92e-16
c28541 4938 4934 1.845e-15
c28542 3411 3591 1.58e-16
c28543 3397 3604 4.63e-16
c28544 4759 1 2.0331e-14
c28545 2004 1 4.946e-15
c28546 852 850 3.327e-15
c28547 2516 0 6.72e-16
c28548 4753 497 1.88e-16
c28549 2477 2479 2.03e-16
c28550 1551 752 3.64e-16
c28551 3876 4234 1.58e-16
c28552 3900 4246 5.42e-16
c28553 3882 797 3.15e-16
c28554 5514 5429 8.28e-16
c28555 610 1 3.79e-16
c28556 603 0 7.86e-15
c28557 3056 3067 1.96e-16
c28558 1162 1 3.54e-16
c28559 4261 1 9.28e-16
c28560 3393 3027 1.96e-16
c28561 2718 732 2.4e-16
c28562 1852 1465 1.532e-15
c28563 1858 1857 5.65e-16
c28564 1159 0 9.602e-15
c28565 3034 3258 4.63e-16
c28566 2175 2181 5.8e-16
c28567 426 117 1.88e-16
c28568 5288 5281 9.38e-16
c28569 4779 0 3.4504e-14
c28570 601 2599 1.58e-16
c28571 1 488 2.87e-16
c28572 118 117 7.03e-16
c28573 136 131 1.88e-16
c28574 2653 2271 2.48e-16
c28575 2459 2461 1.862e-15
c28576 1947 1953 1.418e-15
c28577 1964 1936 2.64e-16
c28578 2169 2167 3.54e-16
c28579 4770 5212 1.96e-16
c28580 4922 62 1.88e-16
c28581 2758 2754 1.96e-16
c28582 1207 842 1.58e-16
c28583 1188 1194 1.58e-16
c28584 920 1025 3.92e-16
c28585 921 1024 2.54e-16
c28586 1004 1 3.06e-16
c28587 3898 4400 3.92e-16
c28588 4483 4481 1.6e-16
c28589 520 477 1.88e-16
c28590 2196 2218 5.42e-16
c28591 3773 3775 1.09e-15
c28592 2095 0 1.666e-15
c28593 160 157 1.099e-15
c28594 64 91 1.88e-16
c28595 78 102 1.88e-16
c28596 3310 3693 7.84e-16
c28597 3046 822 3.15e-16
c28598 1151 812 3.15e-16
c28599 1161 1164 1.58e-16
c28600 4023 19 3.45e-16
c28601 2557 2666 1.58e-16
c28602 2541 2654 1.58e-16
c28603 2164 858 7.12e-16
c28604 1196 1321 5.5e-16
c28605 3137 3135 1.6e-16
c28606 1550 1948 4.36e-16
c28607 1946 1939 1.96e-16
c28608 3526 3134 2.38e-15
c28609 3517 662 4.81e-16
c28610 3397 3569 1.58e-16
c28611 2547 2546 6.97e-16
c28612 2548 2544 1.71e-16
c28613 2136 2093 2.74e-16
c28614 842 834 1.74e-16
c28615 657 3489 1.58e-16
c28616 1789 647 1.58e-16
c28617 1786 672 1.58e-16
c28618 902 943 3.92e-16
c28619 2532 1 4.044e-15
c28620 2194 2372 3.92e-16
c28621 1530 737 1.09e-16
c28622 1270 1251 1.58e-16
c28623 146 421 1.88e-16
c28624 3886 767 3.15e-16
c28625 3059 0 6.62e-16
c28626 2559 2458 1.58e-16
c28627 919 1145 3.92e-16
c28628 922 1144 2.54e-16
c28629 3126 2628 1.58e-16
c28630 1121 1116 1.58e-16
c28631 3608 762 1.58e-16
c28632 1239 0 3.6229e-14
c28633 777 1130 1.85e-16
c28634 687 2667 2.4e-16
c28635 2452 0 6.9025e-14
c28636 595 2572 1.58e-16
c28637 602 2569 1.832e-15
c28638 3781 3796 1.96e-16
c28639 165 1 1.1938e-14
c28640 129 0 4.3431e-14
c28641 5412 5414 1.001e-15
c28642 4287 4285 2.15e-16
c28643 4295 4294 1.6e-16
c28644 1708 662 3.15e-16
c28645 1380 1375 1.642e-15
c28646 3763 3764 2.67e-16
c28647 2248 2620 1.58e-16
c28648 1490 1056 2.48e-16
c28649 2299 702 1.813e-15
c28650 822 907 3.15e-16
c28651 3048 792 3.58e-16
c28652 2390 767 2.33e-16
c28653 2178 662 3.15e-16
c28654 1747 1363 1.58e-16
c28655 2696 3214 2.38e-15
c28656 3124 672 1.58e-16
c28657 3046 3045 1.009e-15
c28658 1708 1918 3.92e-16
c28659 33 296 1.88e-16
c28660 340 332 2.218e-15
c28661 333 349 3.84e-16
c28662 642 3118 2.65e-16
c28663 1415 647 7.68e-16
c28664 596 732 1.96e-16
c28665 395 1 3.6e-16
c28666 4770 1 2.7499e-14
c28667 4606 0 3.61969e-13
c28668 4071 4068 1.58e-16
c28669 3211 1 5.808e-15
c28670 924 1 8.63e-16
c28671 3886 4353 1.58e-16
c28672 3876 3514 5.5e-16
c28673 2182 662 3.15e-16
c28674 1733 1352 3.92e-16
c28675 3980 26 4.58e-16
c28676 3972 0 2.0172e-14
c28677 4369 4371 2.03e-16
c28678 1196 1627 1.58e-16
c28679 916 0 3.8e-16
c28680 2645 647 1.58e-16
c28681 1706 1917 1.58e-16
c28682 1690 1905 1.58e-16
c28683 1253 1 2.223e-15
c28684 2179 1687 1.939e-15
c28685 2183 1698 1.018e-15
c28686 3486 662 2.33e-16
c28687 5278 352 3.54e-16
c28688 3048 737 3.15e-16
c28689 1 17 1.44e-16
c28690 12 11 2.84e-16
c28691 2802 2418 1.58e-16
c28692 2622 2618 1.96e-16
c28693 14 0 1.0822e-14
c28694 9 27 5.8e-16
c28695 3270 3654 1.58e-16
c28696 4563 4446 5.88e-16
c28697 4571 4452 1.58e-16
c28698 2832 822 2.22e-16
c28699 2559 1 2.222e-15
c28700 2194 2337 1.58e-16
c28701 2178 2325 1.58e-16
c28702 3531 3503 2.64e-16
c28703 3514 3520 1.418e-15
c28704 4351 4353 1.862e-15
c28705 1690 797 3.15e-16
c28706 689 26 2.65e-15
c28707 3583 1 1.868e-15
c28708 1264 1 7.87e-16
c28709 4608 4231 2.48e-16
c28710 657 2283 2.65e-16
c28711 1694 1315 3.54e-16
c28712 4158 1 6.76e-16
c28713 792 909 3.15e-16
c28714 4880 4879 2.03e-16
c28715 2770 3279 7.84e-16
c28716 1807 0 6.72e-16
c28717 3645 3644 1.6e-16
c28718 3259 3640 3.92e-16
c28719 2127 2106 1.96e-16
c28720 1014 647 8.3e-16
c28721 1021 672 1.35e-16
c28722 812 806 1.74e-16
c28723 1 510 4.22e-16
c28724 233 565 1.88e-16
c28725 421 320 1.88e-16
c28726 2196 2495 1.58e-16
c28727 26 523 8.41e-16
c28728 9 570 3.92e-16
c28729 3581 3185 1.96e-16
c28730 3659 797 1.832e-15
c28731 5286 1 3.986e-15
c28732 2182 2325 1.58e-16
c28733 1732 1 4.41e-15
c28734 70 1 4.59e-16
c28735 3958 3964 1.96e-16
c28736 3373 3809 2.107e-15
c28737 919 752 3.15e-16
c28738 920 1083 1.58e-16
c28739 1321 996 1.58e-16
c28740 1327 986 5.88e-16
c28741 4156 4150 1.96e-16
c28742 3882 3673 1.58e-16
c28743 3007 3005 2.61e-16
c28744 1953 827 1.75e-16
c28745 1810 1803 1.96e-16
c28746 612 952 1.58e-16
c28747 602 881 1.58e-16
c28748 3948 1 4.64e-16
c28749 4133 19 9.67e-16
c28750 4796 4798 2.15e-16
c28751 2104 2105 3.54e-16
c28752 26 317 1.03e-15
c28753 911 2549 1.829e-15
c28754 1896 2393 1.58e-16
c28755 5025 1 4.55e-15
c28756 687 2535 3.15e-16
c28757 2325 2323 1.862e-15
c28758 909 737 3.15e-16
c28759 883 1096 1.88e-16
c28760 907 1089 1.58e-16
c28761 4838 5093 1.96e-16
c28762 3397 3270 5.5e-16
c28763 5284 5346 6.67e-16
c28764 2774 0 6.62e-16
c28765 2584 1 1.716e-15
c28766 601 590 1.078e-15
c28767 52 42 8.86e-16
c28768 60 62 6.01e-16
c28769 3713 3714 5.65e-16
c28770 1343 842 4.46e-16
c28771 1331 868 7.99e-16
c28772 627 3457 2.72e-16
c28773 3167 1 8.43e-16
c28774 602 4234 1.832e-15
c28775 595 4237 1.58e-16
c28776 3582 4424 2.38e-15
c28777 1625 1166 1.532e-15
c28778 1631 1630 5.65e-16
c28779 4503 4504 1.35e-16
c28780 4327 4677 2e-16
c28781 3175 3178 6.44e-16
c28782 595 1720 2.72e-16
c28783 612 1716 1.58e-16
c28784 3556 3558 2.03e-16
c28785 3083 3455 1.58e-16
c28786 2756 752 1.832e-15
c28787 5032 0 3.0289e-14
c28788 5033 120 3.54e-16
c28789 5315 5314 2.67e-16
c28790 722 1082 1.58e-16
c28791 1073 732 1.58e-16
c28792 592 835 6.34e-16
c28793 3759 3747 1.96e-16
c28794 2500 2497 3.01e-16
c28795 2496 2493 6.44e-16
c28796 2194 1953 1.58e-16
c28797 397 233 1.88e-16
c28798 3876 827 4.48e-16
c28799 3898 868 3.15e-16
c28800 3142 2634 2.48e-16
c28801 601 977 1.58e-16
c28802 1694 767 3.15e-16
c28803 1345 1559 1.58e-16
c28804 3101 3092 3.92e-16
c28805 2583 3095 5.66e-16
c28806 1897 1891 1.6e-16
c28807 1499 1888 2.386e-15
c28808 1516 1871 1.58e-16
c28809 1212 0 6.29e-16
c28810 1793 1 8.43e-16
c28811 3236 3624 4.97e-16
c28812 3387 3066 5.5e-16
c28813 2382 1 6.15e-16
c28814 448 454 5.8e-16
c28815 1 197 1.44e-16
c28816 3745 3732 1.96e-16
c28817 4567 4758 3.92e-16
c28818 4742 4743 9.93e-16
c28819 5474 0 1.65e-16
c28820 3765 3769 3.82e-16
c28821 3927 3926 1.58e-16
c28822 5388 381 1.96e-16
c28823 2771 2782 1.96e-16
c28824 1031 692 3.15e-16
c28825 1476 702 2.72e-16
c28826 1041 1044 1.58e-16
c28827 4233 4235 2.03e-16
c28828 2288 2670 2.48e-16
c28829 542 465 1.88e-16
c28830 528 497 1.88e-16
c28831 4112 1 3.3163e-14
c28832 1953 812 2.33e-16
c28833 1803 1414 2.386e-15
c28834 1707 1691 3.54e-16
c28835 4643 1 4.832e-15
c28836 4395 4758 1.96e-16
c28837 3409 3434 3.92e-16
c28838 1635 2020 1.96e-16
c28839 1708 1624 1.58e-16
c28840 1706 1618 5.5e-16
c28841 1694 2019 1.58e-16
c28842 4742 4744 4.93e-16
c28843 1977 1975 1.6e-16
c28844 1972 1971 2.03e-16
c28845 1580 0 6.72e-16
c28846 792 1106 1.58e-16
c28847 777 1121 3.79e-16
c28848 0 450 1.24687e-13
c28849 25 433 7.06e-16
c28850 30 441 3.84e-16
c28851 4580 4579 1.009e-15
c28852 4563 4568 9.81e-16
c28853 5123 5101 1.74e-16
c28854 5108 5100 3.54e-16
c28855 1128 1142 1.96e-16
c28856 108 117 1.58e-16
c28857 91 122 1.88e-16
c28858 4336 692 1.58e-16
c28859 1166 868 1.58e-16
c28860 1638 827 4.81e-16
c28861 1452 1016 1.58e-16
c28862 3882 4451 1.96e-16
c28863 2557 2735 3.92e-16
c28864 2805 812 1.339e-15
c28865 3445 3022 1.96e-16
c28866 3440 3055 1.96e-16
c28867 1932 1 9.28e-16
c28868 165 363 1.88e-16
c28869 5299 5297 3.92e-16
c28870 4810 236 1.88e-16
c28871 2772 2384 4.97e-16
c28872 868 870 5.59e-16
c28873 4132 857 1.88e-16
c28874 3900 3486 1.58e-16
c28875 1106 737 3.57e-16
c28876 3900 4251 1.58e-16
c28877 3876 812 4.48e-16
c28878 4506 827 1.832e-15
c28879 2852 2850 1.6e-16
c28880 921 1190 1.96e-16
c28881 4326 3480 1.96e-16
c28882 1975 827 5.03e-16
c28883 3642 0 3.3874e-14
c28884 612 3876 3.15e-16
c28885 4274 1 6.15e-16
c28886 4850 4849 1.6e-16
c28887 1721 0 1.4092e-14
c28888 4796 0 3.4717e-14
c28889 3393 3396 1.96e-16
c28890 617 2599 7.38e-16
c28891 4582 4327 5.5e-16
c28892 5136 5103 1.58e-16
c28893 747 2372 2.4e-16
c28894 4421 752 1.832e-15
c28895 5450 5447 7.81e-16
c28896 1453 662 1.58e-16
c28897 1207 1209 7.84e-16
c28898 3469 4305 5.66e-16
c28899 4311 4302 3.92e-16
c28900 3472 1 5.808e-15
c28901 2545 2322 1.58e-16
c28902 1506 1071 3.92e-16
c28903 1510 1511 1.6e-16
c28904 3474 0 3.466e-15
c28905 2407 807 5.73e-16
c28906 1782 1397 1.96e-16
c28907 4053 0 1.5176e-14
c28908 3228 3240 2.32e-16
c28909 4587 0 2.96e-16
c28910 0 337 9.795e-15
c28911 3508 3509 1.6e-16
c28912 2196 2223 1.58e-16
c28913 160 117 1.88e-16
c28914 3882 3875 1.58e-16
c28915 3886 3895 1.58e-16
c28916 2820 822 2.4e-16
c28917 2288 0 3.6368e-14
c28918 4388 4385 6.44e-16
c28919 4392 4389 3.01e-16
c28920 3387 1 3.564e-15
c28921 2535 2683 1.58e-16
c28922 2557 2671 1.58e-16
c28923 632 1782 1.58e-16
c28924 3880 0 6.78e-16
c28925 3565 1 5.97e-15
c28926 4664 4662 1.6e-16
c28927 204 455 1.88e-16
c28928 3151 672 2.22e-16
c28929 3523 677 1.832e-15
c28930 5006 5005 1.08e-15
c28931 422 428 1.372e-15
c28932 421 420 1.88e-16
c28933 417 418 6.67e-16
c28934 4944 0 4.0267e-14
c28935 3397 3574 1.58e-16
c28936 4844 4469 4.9e-16
c28937 3247 0 3.466e-15
c28938 3084 1 1.868e-15
c28939 1270 1295 1.25e-15
c28940 5538 5533 7.46e-16
c28941 2350 717 2.22e-16
c28942 1706 868 3.15e-16
c28943 1684 827 4.48e-16
c28944 533 1 4.22e-16
c28945 3146 2628 2.38e-15
c28946 1975 812 1.9e-16
c28947 1121 1585 4.36e-16
c28948 1583 1576 1.96e-16
c28949 3606 0 1.6491e-14
c28950 4463 3622 1.136e-15
c28951 4259 4646 2.196e-15
c28952 1706 1386 1.58e-16
c28953 1841 1839 1.6e-16
c28954 1836 1835 2.03e-16
c28955 4935 4934 2.67e-16
c28956 3024 2713 5.5e-16
c28957 3034 3228 1.58e-16
c28958 1465 0 6.9481e-14
c28959 4748 1 2.378e-15
c28960 4747 0 3.466e-15
c28961 137 0 1.0822e-14
c28962 3601 3594 6.73e-16
c28963 3600 3208 1.96e-16
c28964 5044 5031 1.58e-16
c28965 5051 5058 3.18e-16
c28966 4878 323 1.88e-16
c28967 601 2569 1.58e-16
c28968 2443 1936 2.48e-16
c28969 3886 3401 1.58e-16
c28970 1243 1291 1.6e-16
c28971 1289 1226 1.96e-16
c28972 5358 294 7.46e-16
c28973 2738 2740 2.03e-16
c28974 3607 0 2.93e-15
c28975 3428 1 8.43e-16
c28976 2545 2837 4.63e-16
c28977 4005 1 7.71e-16
c28978 4454 3616 4.97e-16
c28979 4571 707 1.33e-16
c28980 1755 1761 1.6e-16
c28981 1752 1363 2.386e-15
c28982 1380 1735 1.58e-16
c28983 4215 1 7.228e-15
c28984 3128 662 5.03e-16
c28985 2541 767 3.15e-16
c28986 1331 0 3.26142e-13
c28987 30 34 6.83e-16
c28988 117 513 1.88e-16
c28989 3208 3593 1.96e-16
c28990 889 898 1.872e-15
c28991 3594 752 1.84e-16
c28992 632 3120 4.81e-16
c28993 5380 5379 1.6e-16
c28994 2640 1 2.054e-15
c28995 3027 3033 5.8e-16
c28996 2194 2528 4.22e-16
c28997 3399 0 5.86e-16
c28998 2933 2934 1.96e-16
c28999 2918 2913 3.54e-16
c29000 2849 2458 1.136e-15
c29001 3505 3123 2.48e-16
c29002 3900 3531 5.5e-16
c29003 3307 3305 1.6e-16
c29004 3797 0 1.65e-16
c29005 2713 762 1.58e-16
c29006 2730 747 3.79e-16
c29007 1652 842 1.58e-16
c29008 2696 3218 1.96e-16
c29009 2702 3213 1.96e-16
c29010 3024 3025 1.487e-15
c29011 3034 3027 1.58e-16
c29012 2858 852 1.58e-16
c29013 642 2196 3.58e-16
c29014 3898 0 3.47397e-13
c29015 1924 1920 1.96e-16
c29016 1694 1747 1.58e-16
c29017 747 1525 1.58e-16
c29018 25 580 3.84e-16
c29019 5010 4980 6.15e-16
c29020 3706 868 2.4e-16
c29021 4285 647 1.58e-16
c29022 5365 5367 3.92e-16
c29023 2790 2435 1.58e-16
c29024 2643 1 6.15e-16
c29025 907 962 3.92e-16
c29026 3287 3642 1.58e-16
c29027 3270 3659 2.386e-15
c29028 3668 3662 1.6e-16
c29029 222 0 1.5723e-14
c29030 3736 3735 5.87e-16
c29031 3209 1 1.716e-15
c29032 2178 2182 4.431e-15
c29033 2528 2524 1.96e-16
c29034 1400 1398 1.6e-16
c29035 2172 2354 1.58e-16
c29036 2194 2342 1.58e-16
c29037 2541 2282 5.88e-16
c29038 2317 692 7.68e-16
c29039 1684 812 4.48e-16
c29040 2545 792 7.99e-16
c29041 4622 4621 8.22e-16
c29042 2776 767 1.58e-16
c29043 4542 3707 2.91e-16
c29044 2491 842 7.38e-16
c29045 568 580 1.58e-16
c29046 576 577 6.4e-16
c29047 3305 812 7.68e-16
c29048 2259 2255 1.96e-16
c29049 612 1684 3.15e-16
c29050 4435 4813 7.84e-16
c29051 3220 737 7.68e-16
c29052 2413 1 2.054e-15
c29053 1 291 4.22e-16
c29054 5164 5152 1.74e-16
c29055 2415 0 8e-16
c29056 777 2419 2.65e-16
c29057 602 2194 4.46e-16
c29058 595 2172 1.511e-15
c29059 3310 3691 3.92e-16
c29060 3693 3705 2.32e-16
c29061 1046 732 1.58e-16
c29062 632 3397 3.15e-16
c29063 3310 842 1.75e-16
c29064 2832 2827 1.642e-15
c29065 1970 868 5.73e-16
c29066 2487 827 3.64e-16
c29067 601 881 3.15e-16
c29068 627 952 5.73e-16
c29069 3967 1 6.66e-16
c29070 627 4264 2.4e-16
c29071 2770 3277 3.92e-16
c29072 3282 3281 1.6e-16
c29073 3213 722 1.9e-16
c29074 2545 737 3.15e-16
c29075 1166 0 7.407e-14
c29076 19 545 8.82e-16
c29077 456 455 6.96e-16
c29078 3409 662 4.46e-16
c29079 3572 3575 6.44e-16
c29080 722 713 1.078e-15
c29081 3572 737 1.339e-15
c29082 1158 807 1.58e-16
c29083 894 752 3.15e-16
c29084 890 1083 3.54e-16
c29085 909 1104 1.58e-16
c29086 4838 5072 3.54e-16
c29087 2849 1 5.343e-15
c29088 1846 707 7.68e-16
c29089 1661 852 2.8e-16
c29090 1345 858 3.15e-16
c29091 1466 1026 1.96e-16
c29092 1467 1460 6.73e-16
c29093 3363 0 3.26e-15
c29094 601 4234 1.58e-16
c29095 2402 752 3.64e-16
c29096 870 0 7.709e-15
c29097 3927 19 3.45e-16
c29098 4327 4694 1.58e-16
c29099 1694 1488 1.58e-16
c29100 1451 1 1.056e-15
c29101 3083 3475 2.38e-15
c29102 3876 747 3.15e-16
c29103 566 563 2.142e-15
c29104 488 487 1.58e-16
c29105 455 175 1.88e-16
c29106 5114 1 2.424e-15
c29107 5262 5265 3.54e-16
c29108 2788 2401 1.532e-15
c29109 2602 2604 2.03e-16
c29110 4184 857 3.1e-16
c29111 5200 5207 3.54e-16
c29112 627 3451 2.4e-16
c29113 2172 1970 1.58e-16
c29114 2178 1964 5.88e-16
c29115 1559 782 1.58e-16
c29116 393 407 1.58e-16
c29117 378 426 1.88e-16
c29118 3900 852 3.58e-16
c29119 4724 707 1.23e-16
c29120 5403 5513 1.58e-16
c29121 2529 2530 1.76e-16
c29122 617 977 1.58e-16
c29123 3911 25 7.01e-16
c29124 4335 3503 2.48e-16
c29125 1624 852 5.73e-16
c29126 1327 1131 1.58e-16
c29127 1211 1214 6.13e-16
c29128 4593 4591 2.03e-16
c29129 676 674 5.88e-16
c29130 88 194 1.88e-16
c29131 3411 3083 5.5e-16
c29132 2103 2098 1.291e-15
c29133 1 323 3.36e-15
c29134 281 450 1.88e-16
c29135 3393 807 4.03e-16
c29136 4036 4040 3.84e-16
c29137 4044 4043 4.41e-16
c29138 4668 4663 1.536e-15
c29139 4567 4775 3.92e-16
c29140 5233 5234 5.87e-16
c29141 2182 1964 5.5e-16
c29142 3992 857 3.1e-16
c29143 2194 1777 5.5e-16
c29144 5514 5426 1.237e-15
c29145 5403 5519 1.52e-16
c29146 5484 5505 1.96e-16
c29147 5422 5425 1.817e-15
c29148 4742 5358 1.344e-15
c29149 1931 767 3.64e-16
c29150 1091 1537 1.58e-16
c29151 632 3882 3.15e-16
c29152 74 78 1.58e-16
c29153 2978 2923 3.18e-16
c29154 2976 2968 1.96e-16
c29155 2954 2509 6.55e-16
c29156 1058 1 4.59e-16
c29157 868 26 1.58e-16
c29158 4126 1 6.76e-16
c29159 3711 0 6.62e-16
c29160 1055 0 1.0077e-14
c29161 4660 1 4.832e-15
c29162 4395 4775 1.96e-16
c29163 3048 3126 1.58e-16
c29164 2098 2101 1.099e-15
c29165 1601 1969 1.96e-16
c29166 3157 3540 7.84e-16
c29167 5104 5122 1.37e-16
c29168 4878 265 1.88e-16
c29169 2400 1879 1.96e-16
c29170 2395 1885 1.96e-16
c29171 702 708 1.097e-15
c29172 2176 0 6.78e-16
c29173 59 334 1.88e-16
c29174 4356 692 1.58e-16
c29175 4132 4136 3.84e-16
c29176 4140 4139 4.41e-16
c29177 1196 837 4.21e-16
c29178 1457 1016 2.386e-15
c29179 4079 37 1.88e-16
c29180 4406 3565 4.11e-16
c29181 2535 2752 3.92e-16
c29182 2381 737 1.09e-16
c29183 1614 1612 1.6e-16
c29184 1609 1608 2.03e-16
c29185 1690 1816 1.96e-16
c29186 4453 0 1.6491e-14
c29187 5074 5079 3.84e-16
c29188 1945 1 6.15e-16
c29189 1706 0 3.5222e-13
c29190 3540 717 1.58e-16
c29191 5048 1 2.386e-15
c29192 3387 3225 1.58e-16
c29193 4759 410 1.88e-16
c29194 5160 5173 1.138e-15
c29195 1106 1104 1.931e-15
c29196 3882 3435 1.58e-16
c29197 687 1038 1.58e-16
c29198 920 1204 1.58e-16
c29199 1601 842 1.58e-16
c29200 1995 827 1.09e-16
c29201 1331 1091 5.5e-16
c29202 3662 0 1.4092e-14
c29203 627 3876 3.15e-16
c29204 4283 1 1.716e-15
c29205 3082 2533 1.96e-16
c29206 3077 2566 1.96e-16
c29207 1870 1871 2.48e-16
c29208 966 0 3.7577e-14
c29209 3030 3291 1.58e-16
c29210 3258 767 7.38e-16
c29211 3046 672 3.15e-16
c29212 3024 647 4.48e-16
c29213 426 479 1.88e-16
c29214 4813 0 3.4075e-14
c29215 1 430 2.87e-16
c29216 15 425 6.58e-16
c29217 3611 3608 5.5e-16
c29218 3397 3018 3.54e-16
c29219 782 774 1.74e-16
c29220 4582 4344 5.5e-16
c29221 5165 5152 1.96e-16
c29222 5136 5144 3.258e-15
c29223 4861 33 1.88e-16
c29224 2489 2487 1.6e-16
c29225 5579 5575 1.96e-16
c29226 1031 1034 6.13e-16
c29227 922 1040 3.92e-16
c29228 3492 1 2.054e-15
c29229 3640 0 1.6491e-14
c29230 911 3877 2.09e-16
c29231 3494 0 8e-16
c29232 4491 4492 1.6e-16
c29233 4487 3656 3.92e-16
c29234 3352 3349 3.01e-16
c29235 3348 3345 6.44e-16
c29236 4743 4745 1.687e-15
c29237 4755 4748 6.73e-16
c29238 4754 4367 1.96e-16
c29239 1635 1990 1.58e-16
c29240 1 484 3.0375e-14
c29241 595 0 3.03776e-13
c29242 19 490 3.45e-16
c29243 0 499 5.6218e-14
c29244 33 497 1.88e-16
c29245 3922 3911 7.1e-16
c29246 3915 3924 6.67e-16
c29247 5083 5032 1.191e-15
c29248 88 15 5.8e-16
c29249 2274 2286 2.32e-16
c29250 97 0 2.87e-16
c29251 922 662 5.14e-16
c29252 1327 1341 3.92e-16
c29253 2580 2578 1.6e-16
c29254 1419 986 1.96e-16
c29255 3898 4404 1.58e-16
c29256 3876 4416 1.58e-16
c29257 2747 0 6.9041e-14
c29258 2196 732 3.58e-16
c29259 2559 2700 5.42e-16
c29260 2535 2688 1.58e-16
c29261 2355 722 7.38e-16
c29262 4745 4744 2.48e-16
c29263 3145 3146 1.6e-16
c29264 4432 1 1.056e-15
c29265 291 363 1.88e-16
c29266 248 254 1.372e-15
c29267 5219 0 1.963e-15
c29268 4941 1 1.18e-16
c29269 3343 842 7.38e-16
c29270 747 1684 3.15e-16
c29271 907 672 3.15e-16
c29272 883 647 6.45e-16
c29273 4954 0 2.8939e-14
c29274 2676 0 8e-16
c29275 2558 2552 1.988e-15
c29276 62 93 1.88e-16
c29277 2577 1 5.97e-15
c29278 1708 852 3.58e-16
c29279 1343 1504 3.92e-16
c29280 1358 1 2.054e-15
c29281 910 1331 5.03e-16
c29282 1684 1403 1.58e-16
c29283 1690 1397 5.88e-16
c29284 2178 852 4.03e-16
c29285 1465 1833 1.96e-16
c29286 1360 0 8e-16
c29287 2798 827 1.58e-16
c29288 3688 3304 1.58e-16
c29289 4765 1 2.378e-15
c29290 2866 2855 1.58e-16
c29291 4764 0 3.466e-15
c29292 2441 2452 1.58e-16
c29293 612 2589 1.58e-16
c29294 1970 0 3.6368e-14
c29295 2172 2388 1.58e-16
c29296 2194 2376 1.58e-16
c29297 2807 2819 2.32e-16
c29298 2178 2168 3.54e-16
c29299 2194 2171 1.58e-16
c29300 146 128 1.58e-16
c29301 5442 5451 2.177e-15
c29302 2646 2254 1.96e-16
c29303 1884 737 7.38e-16
c29304 911 3876 1.88e-16
c29305 910 3898 1.014e-15
c29306 2182 852 7.99e-16
c29307 632 1690 3.15e-16
c29308 1113 0 4.6566e-14
c29309 4199 19 7.04e-16
c29310 4216 0 1.5176e-14
c29311 3313 2804 7.84e-16
c29312 2713 2702 1.58e-16
c29313 2535 782 4.48e-16
c29314 2023 2033 9.99e-16
c29315 792 1327 4.03e-16
c29316 15 253 4.88e-16
c29317 1 265 3.36e-15
c29318 465 565 1.88e-16
c29319 2196 1862 5.5e-16
c29320 1760 1 5.97e-15
c29321 4514 4509 1.642e-15
c29322 2182 2168 1.58e-16
c29323 3480 677 1.58e-16
c29324 4770 410 1.88e-16
c29325 2822 0 1.6491e-14
c29326 2541 2271 1.58e-16
c29327 2248 2644 1.96e-16
c29328 2254 2639 1.96e-16
c29329 921 963 1.58e-16
c29330 3029 3033 5.8e-16
c29331 1488 732 1.58e-16
c29332 1491 1503 2.32e-16
c29333 3789 3734 1.141e-15
c29334 4097 4094 1.76e-16
c29335 3414 0 1.23e-16
c29336 2545 2836 1.58e-16
c29337 1750 1363 1.532e-15
c29338 3034 3029 1.58e-16
c29339 3030 3038 8.73e-16
c29340 1708 1922 1.58e-16
c29341 642 1752 1.58e-16
c29342 3508 3117 4.11e-16
c29343 4452 4453 1.35e-16
c29344 1694 1752 1.58e-16
c29345 433 419 3.84e-16
c29346 436 455 1.88e-16
c29347 2357 2359 1.862e-15
c29348 1845 1851 1.418e-15
c29349 4904 4902 3.54e-16
c29350 1749 2259 1.96e-16
c29351 417 1 4.22e-16
c29352 390 15 5.8e-16
c29353 909 977 4.35e-16
c29354 907 976 1.88e-16
c29355 890 969 1.58e-16
c29356 1023 1024 1.21e-16
c29357 4668 33 1.88e-16
c29358 3235 1 8.43e-16
c29359 1327 737 3.15e-16
c29360 4381 4379 1.6e-16
c29361 3216 3213 3.01e-16
c29362 3212 3209 6.44e-16
c29363 1811 692 3.15e-16
c29364 2327 702 2.72e-16
c29365 3601 1 9.28e-16
c29366 1561 1557 1.96e-16
c29367 4625 4248 2.48e-16
c29368 3537 0 3.583e-14
c29369 4889 4879 8.06e-16
c29370 5158 207 1.58e-16
c29371 2798 812 3.15e-16
c29372 1829 1 1.868e-15
c29373 627 1684 3.15e-16
c29374 1819 0 2.93e-15
c29375 3387 3518 1.58e-16
c29376 3662 3663 5.65e-16
c29377 3270 3657 1.532e-15
c29378 2713 722 3.15e-16
c29379 2435 1 5.97e-15
c29380 2153 1641 2.91e-16
c29381 2155 2154 1.6e-16
c29382 1028 662 3.57e-16
c29383 1 44 4.096e-15
c29384 0 26 4.89201e-13
c29385 5151 5259 1.58e-16
c29386 5324 1 1.021e-15
c29387 2431 0 6.72e-16
c29388 792 1896 1.58e-16
c29389 777 1913 3.79e-16
c29390 601 2194 4.46e-16
c29391 1076 717 4.21e-16
c29392 1243 1255 1.96e-16
c29393 632 1007 1.58e-16
c29394 3028 0 6.78e-16
c29395 922 1098 1.58e-16
c29396 1001 1000 3.94e-16
c29397 392 107 1.88e-16
c29398 752 1 3.1284e-14
c29399 627 1398 2.65e-16
c29400 617 881 1.58e-16
c29401 4165 1 7.71e-16
c29402 3886 4535 1.58e-16
c29403 3898 3684 5.5e-16
c29404 3900 3690 1.58e-16
c29405 3701 4536 1.96e-16
c29406 1735 1734 2.48e-16
c29407 4813 4815 2.15e-16
c29408 4822 4811 1.96e-16
c29409 9 580 3.92e-16
c29410 309 311 1.58e-16
c29411 310 291 1.88e-16
c29412 2419 1902 1.96e-16
c29413 2420 2413 6.73e-16
c29414 0 571 1.0822e-14
c29415 2892 3847 1.666e-15
c29416 2801 1 1.056e-15
c29417 4872 5137 2.137e-15
c29418 2789 2407 2.48e-16
c29419 920 918 5.74e-16
c29420 1465 707 3.15e-16
c29421 1856 717 2.72e-16
c29422 1031 1026 1.58e-16
c29423 601 4254 1.58e-16
c29424 4448 4441 6.73e-16
c29425 4447 3605 1.96e-16
c29426 1896 737 1.58e-16
c29427 3278 2764 4.97e-16
c29428 687 1437 1.58e-16
c29429 3943 37 1.88e-16
c29430 3944 26 1.06e-15
c29431 2679 3190 1.96e-16
c29432 612 1737 2.72e-16
c29433 1467 1 9.28e-16
c29434 4344 4694 2e-16
c29435 1618 1986 1.96e-16
c29436 601 612 3.28e-16
c29437 455 349 1.88e-16
c29438 1990 1 5.808e-15
c29439 1992 0 3.466e-15
c29440 64 584 4.48e-16
c29441 3393 3671 1.58e-16
c29442 1089 1096 2.27e-16
c29443 894 891 5.52e-16
c29444 596 847 3.134e-15
c29445 2586 0 3.3717e-14
c29446 5509 1 1.88e-16
c29447 2508 1998 1.96e-16
c29448 1579 782 1.58e-16
c29449 1331 707 3.15e-16
c29450 1371 881 4.97e-16
c29451 957 952 1.58e-16
c29452 4563 5591 2e-16
c29453 4651 5491 9.98e-16
c29454 3163 0 1.4092e-14
c29455 2545 2599 4.63e-16
c29456 1221 1228 1.078e-15
c29457 2304 662 1.58e-16
c29458 657 1331 7.99e-16
c29459 1708 1701 3.54e-16
c29460 1690 1702 6.67e-16
c29461 1222 1 5.63e-16
c29462 4323 0 6.72e-16
c29463 4867 4480 2.196e-15
c29464 5230 178 4.44e-16
c29465 2239 2241 2.03e-16
c29466 5318 5316 8.35e-16
c29467 2157 2078 3.01e-16
c29468 993 1006 1.58e-16
c29469 4567 4792 3.92e-16
c29470 5491 1 2.429e-15
c29471 5200 5199 5.01e-16
c29472 4776 468 1.88e-16
c29473 1987 2495 7.84e-16
c29474 3886 717 7.99e-16
c29475 3898 707 4.46e-16
c29476 2557 2373 1.58e-16
c29477 1550 767 3.15e-16
c29478 657 3898 3.15e-16
c29479 858 19 1.676e-15
c29480 3684 4518 1.58e-16
c29481 3366 2855 2.91e-16
c29482 3368 3367 1.6e-16
c29483 910 1706 1.014e-15
c29484 911 1684 1.88e-16
c29485 4677 1 4.832e-15
c29486 4412 4775 1.96e-16
c29487 3207 707 1.58e-16
c29488 1789 0 1.4092e-14
c29489 1602 1 1.868e-15
c29490 427 419 2.218e-15
c29491 4759 4763 1.81e-16
c29492 5198 5195 7.81e-16
c29493 1592 0 2.93e-15
c29494 3168 3552 1.58e-16
c29495 309 303 5.8e-16
c29496 0 187 4.6772e-14
c29497 19 201 8.4e-16
c29498 291 339 1.88e-16
c29499 33 209 2.92e-16
c29500 3732 3773 5.71e-16
c29501 3772 3767 7.25e-16
c29502 5133 5139 6.23e-16
c29503 4810 178 1.88e-16
c29504 1148 1149 1.213e-15
c29505 4245 4243 1.6e-16
c29506 4351 717 1.58e-16
c29507 2203 2586 7.84e-16
c29508 1447 1438 3.46e-16
c29509 3900 4468 3.92e-16
c29510 4102 26 4.48e-16
c29511 3886 4298 4.63e-16
c29512 3169 3163 1.6e-16
c29513 1982 1973 3.92e-16
c29514 1590 1976 5.66e-16
c29515 1601 1968 1.58e-16
c29516 1706 1833 3.92e-16
c29517 5127 5114 3.92e-16
c29518 350 354 6.38e-16
c29519 332 337 1.482e-15
c29520 3560 717 1.58e-16
c29521 5314 323 3.54e-16
c29522 4941 4950 1.193e-15
c29523 3457 3066 4.11e-16
c29524 3693 3304 2.386e-15
c29525 2549 1 8.822e-15
c29526 596 802 3.134e-15
c29527 3696 827 1.58e-16
c29528 5265 149 3.54e-16
c29529 3310 3411 1.58e-16
c29530 595 3430 2.65e-16
c29531 602 3021 2.33e-16
c29532 392 1 3.6971e-14
c29533 3898 3452 1.58e-16
c29534 4514 5584 1.96e-16
c29535 5580 5582 1.6e-16
c29536 2860 2861 1.6e-16
c29537 2541 2531 3.54e-16
c29538 2557 2534 1.58e-16
c29539 3163 3162 1.6e-16
c29540 602 911 1.58e-16
c29541 595 910 1.58e-16
c29542 178 180 1.96e-16
c29543 3046 3308 1.58e-16
c29544 3030 3296 1.58e-16
c29545 2110 178 9.02e-16
c29546 4830 0 3.485e-14
c29547 2080 2078 7.82e-16
c29548 2196 2440 3.92e-16
c29549 5564 497 3.54e-16
c29550 2645 0 6.9063e-14
c29551 2933 1 2.224e-15
c29552 1227 858 6.47e-16
c29553 378 513 1.88e-16
c29554 107 276 1.88e-16
c29555 3588 767 1.75e-16
c29556 5502 5479 2.12e-16
c29557 5486 5483 2.004e-15
c29558 4844 149 1.88e-16
c29559 919 1054 1.58e-16
c29560 2657 2654 5.5e-16
c29561 1523 1076 1.532e-15
c29562 1529 1528 5.65e-16
c29563 1187 0 1.0183e-14
c29564 4070 1 7.08e-16
c29565 3048 2764 5.5e-16
c29566 3034 2594 5.5e-16
c29567 2559 837 3.58e-16
c29568 421 368 1.88e-16
c29569 4708 4711 6.02e-16
c29570 3409 3407 1.96e-16
c29571 3527 3526 5.65e-16
c29572 5543 497 7.46e-16
c29573 5151 1 4.427e-15
c29574 747 2376 1.58e-16
c29575 5592 0 2.537e-15
c29576 2657 2664 6.73e-16
c29577 642 921 3.15e-16
c29578 3876 4421 1.58e-16
c29579 3900 4433 5.42e-16
c29580 1795 1789 1.6e-16
c29581 1397 1786 2.386e-15
c29582 2559 2705 1.58e-16
c29583 1014 0 2.7256e-14
c29584 2029 2028 3.92e-16
c29585 4448 1 9.28e-16
c29586 3873 0 4.4689e-14
c29587 4681 4679 1.6e-16
c29588 1706 1798 1.58e-16
c29589 3140 692 1.75e-16
c29590 5198 0 4.0816e-14
c29591 4938 4939 8.03e-16
c29592 4903 4902 3.92e-16
c29593 3046 797 4.46e-16
c29594 3034 807 7.99e-16
c29595 2287 1777 1.96e-16
c29596 1766 2283 1.96e-16
c29597 2277 2284 6.73e-16
c29598 2824 822 1.58e-16
c29599 2866 3364 1.66e-16
c29600 2692 0 6.72e-16
c29601 4124 4118 1.96e-16
c29602 4582 1 1.795e-15
c29603 4753 468 1.88e-16
c29604 2748 747 2.65e-16
c29605 2169 2568 2.48e-16
c29606 1812 672 2.65e-16
c29607 4520 0 3.7003e-14
c29608 4640 497 1.88e-16
c29609 4491 827 5.03e-16
c29610 5538 5574 1.617e-15
c29611 5572 5422 1.33e-16
c29612 3554 4387 7.84e-16
c29613 1828 732 1.58e-16
c29614 3625 1 5.808e-15
c29615 1414 1420 1.418e-15
c29616 1321 1521 3.92e-16
c29617 3169 2645 4.36e-16
c29618 4276 4663 2.196e-15
c29619 3242 777 1.58e-16
c29620 4910 5007 9.2e-16
c29621 2815 868 1.58e-16
c29622 3341 827 4.81e-16
c29623 3387 3587 3.92e-16
c29624 4782 1 2.378e-15
c29625 1052 702 2.68e-16
c29626 4571 4480 5.5e-16
c29627 5177 5174 4.41e-16
c29628 458 19 8.82e-16
c29629 5160 5175 1.96e-16
c29630 5170 236 1.58e-16
c29631 4861 526 1.88e-16
c29632 2460 1947 4.97e-16
c29633 4043 3918 8.1e-16
c29634 592 596 6.485e-15
c29635 2172 1678 3.54e-16
c29636 4406 752 5.03e-16
c29637 4776 64 1.88e-16
c29638 1706 707 4.46e-16
c29639 1694 717 7.99e-16
c29640 1588 1589 9.1e-16
c29641 595 884 1.201e-15
c29642 589 1 5.62e-16
c29643 3162 2645 4.11e-16
c29644 1846 1837 3.92e-16
c29645 1454 1840 5.66e-16
c29646 1465 1832 1.58e-16
c29647 657 1706 3.15e-16
c29648 602 919 3.15e-16
c29649 3325 2815 1.58e-16
c29650 1687 0 8.2949e-14
c29651 1 168 1.44e-16
c29652 114 19 8.4e-16
c29653 3678 827 5.03e-16
c29654 2444 2456 2.32e-16
c29655 2302 1 1.056e-15
c29656 2031 1 3.016e-15
c29657 0 190 1.051e-14
c29658 19 158 3.84e-16
c29659 3225 752 2.33e-16
c29660 3828 3773 3.18e-16
c29661 1421 662 1.339e-15
c29662 907 797 4.8e-16
c29663 883 1157 3.92e-16
c29664 890 1156 1.88e-16
c29665 397 450 1.88e-16
c29666 2750 2748 1.6e-16
c29667 632 981 2.33e-16
c29668 3424 0 1.4092e-14
c29669 3839 3785 1.791e-15
c29670 3886 3554 1.58e-16
c29671 4458 4455 5.5e-16
c29672 4600 5538 2.039e-15
c29673 2545 2841 1.58e-16
c29674 2410 782 1.58e-16
c29675 3311 2804 3.92e-16
c29676 3883 1 3.358e-15
c29677 4012 25 1.88e-16
c29678 4008 19 7.35e-16
c29679 1669 1661 2.15e-16
c29680 1196 1206 1.545e-15
c29681 1690 1556 1.58e-16
c29682 910 26 1.58e-16
c29683 305 262 1.88e-16
c29684 5031 5061 9.6e-16
c29685 5056 5047 1.96e-16
c29686 3508 677 5.03e-16
c29687 3396 3398 3.84e-16
c29688 276 1 2.6396e-14
c29689 894 992 3.92e-16
c29690 909 991 1.88e-16
c29691 883 984 1.58e-16
c29692 2537 2536 6.67e-16
c29693 1596 807 1.58e-16
c29694 1321 752 4.48e-16
c29695 1404 981 3.92e-16
c29696 1408 1409 1.6e-16
c29697 4491 812 1.9e-16
c29698 939 25 1.163e-15
c29699 642 1750 1.58e-16
c29700 4639 4638 8.22e-16
c29701 1218 0 5.303e-14
c29702 1448 1 5.97e-15
c29703 4934 1 1.88e-16
c29704 3387 3523 1.58e-16
c29705 3411 3535 5.42e-16
c29706 3393 3140 1.58e-16
c29707 4452 4830 7.84e-16
c29708 233 19 3.84e-16
c29709 632 3485 1.58e-16
c29710 3790 3767 5.87e-16
c29711 3409 852 3.15e-16
c29712 5568 1 1.65e-16
c29713 617 2194 4.46e-16
c29714 161 9 4.88e-16
c29715 139 1 1.44e-16
c29716 3781 3780 2.123e-15
c29717 4286 4283 6.44e-16
c29718 4290 4287 3.01e-16
c29719 2725 2724 1.6e-16
c29720 721 19 1.96e-16
c29721 4589 4600 4.67e-16
c29722 617 1400 4.81e-16
c29723 3701 3876 5.5e-16
c29724 2690 692 1.9e-16
c29725 2495 842 1.832e-15
c29726 584 585 3.84e-16
c29727 762 1117 1.58e-16
c29728 3299 3300 5.65e-16
c29729 2006 1624 2.48e-16
c29730 891 888 8.95e-16
c29731 0 299 2.87e-16
c29732 3678 812 1.9e-16
c29733 4691 439 1.88e-16
c29734 1913 1902 1.58e-16
c29735 3973 3974 3.15e-16
c29736 4623 1 7.831e-15
c29737 1031 1483 4.36e-16
c29738 1481 1474 1.96e-16
c29739 617 4254 1.84e-16
c29740 627 4268 1.58e-16
c29741 1739 1737 1.6e-16
c29742 1734 1733 2.03e-16
c29743 891 1 3.901e-15
c29744 904 0 9.683e-15
c29745 3958 19 7.04e-16
c29746 1480 1 6.15e-16
c29747 2867 842 3.64e-16
c29748 1694 1516 5.5e-16
c29749 617 612 2.77e-16
c29750 187 188 5.8e-16
c29751 3499 3492 6.73e-16
c29752 3498 3106 1.96e-16
c29753 5010 236 1.88e-16
c29754 2341 1834 2.48e-16
c29755 809 808 1.6e-16
c29756 3393 3676 1.58e-16
c29757 3409 3293 1.58e-16
c29758 1083 737 1.58e-16
c29759 13 1 8.75e-16
c29760 2606 0 1.4092e-14
c29761 4668 526 1.88e-16
c29762 1398 957 4.36e-16
c29763 4753 64 1.88e-16
c29764 4352 3514 4.97e-16
c29765 1181 1623 1.96e-16
c29766 1345 1146 1.58e-16
c29767 1343 1136 5.5e-16
c29768 1331 1605 1.58e-16
c29769 4610 4608 2.03e-16
c29770 1533 1505 2.64e-16
c29771 3364 3366 1.96e-16
c29772 3024 3360 3.92e-16
c29773 3089 647 1.75e-16
c29774 2118 2117 1.353e-15
c29775 15 523 5.8e-16
c29776 1 516 1.44e-16
c29777 3387 837 3.15e-16
c29778 4793 4412 5.2e-16
c29779 4567 4809 3.92e-16
c29780 5229 5227 1.387e-15
c29781 1998 2507 1.58e-16
c29782 1013 1014 1.213e-15
c29783 2178 2304 1.96e-16
c29784 5517 5296 2.12e-16
c29785 5422 5410 1.75e-16
c29786 4336 4348 2.32e-16
c29787 920 1100 3.92e-16
c29788 921 1099 2.54e-16
c29789 4215 857 1.96e-16
c29790 1343 1016 5.5e-16
c29791 1327 1001 5.88e-16
c29792 4603 4601 1.6e-16
c29793 2048 2521 1.96e-16
c29794 602 957 3.57e-16
c29795 1079 1 3.06e-16
c29796 3701 4506 1.58e-16
c29797 4871 4480 1.96e-16
c29798 4694 1 4.832e-15
c29799 4412 4792 1.96e-16
c29800 1151 1 5.821e-15
c29801 4776 4778 4.93e-16
c29802 3185 3540 1.58e-16
c29803 3168 3557 2.386e-15
c29804 3566 3560 1.6e-16
c29805 523 507 3.84e-16
c29806 4742 352 1.88e-16
c29807 2182 2304 4.63e-16
c29808 5136 120 1.58e-16
c29809 1678 0 4.7708e-14
c29810 3321 827 3.15e-16
c29811 3327 868 1.58e-16
c29812 3338 3397 5.5e-16
c29813 3344 3855 1.361e-15
c29814 3537 707 2.33e-16
c29815 4776 5221 3.92e-16
c29816 4759 5160 5.87e-16
c29817 921 732 3.15e-16
c29818 2214 2598 1.58e-16
c29819 78 70 1.58e-16
c29820 59 73 1.88e-16
c29821 4152 4154 7.1e-16
c29822 1191 858 1.75e-16
c29823 1453 1452 9.1e-16
c29824 602 4239 1.09e-16
c29825 4428 4419 3.46e-16
c29826 707 26 7.12e-16
c29827 2541 717 4.03e-16
c29828 1601 1973 1.58e-16
c29829 1684 1850 3.92e-16
c29830 657 26 1.58e-16
c29831 541 540 2.84e-16
c29832 3024 868 3.15e-16
c29833 3048 827 3.15e-16
c29834 3411 3236 5.5e-16
c29835 1715 2223 7.84e-16
c29836 1072 1073 7.46e-16
c29837 3752 3747 7.46e-16
c29838 3690 852 5.73e-16
c29839 3886 842 3.15e-16
c29840 601 3021 1.75e-16
c29841 595 3022 2.22e-16
c29842 2815 0 6.8914e-14
c29843 1355 1358 5.5e-16
c29844 919 1220 3.92e-16
c29845 922 1219 2.54e-16
c29846 2535 2166 3.54e-16
c29847 2545 2569 1.58e-16
c29848 2274 647 1.832e-15
c29849 1619 1610 3.92e-16
c29850 1161 1613 5.66e-16
c29851 1166 1605 1.58e-16
c29852 1706 1832 1.58e-16
c29853 1690 1820 1.58e-16
c29854 4401 4402 1.35e-16
c29855 3094 2577 4.11e-16
c29856 5002 5001 1.6e-16
c29857 3066 3451 1.96e-16
c29858 3359 3360 9.1e-16
c29859 3024 3325 1.58e-16
c29860 3046 3313 1.58e-16
c29861 3409 3621 3.92e-16
c29862 88 247 1.88e-16
c29863 461 462 6.4e-16
c29864 1 193 9.8e-16
c29865 4640 4259 5.2e-16
c29866 4838 439 1.88e-16
c29867 2546 0 1.157e-14
c29868 1364 880 1.96e-16
c29869 1365 1358 6.73e-16
c29870 922 852 3.15e-16
c29871 392 310 1.88e-16
c29872 4447 767 3.64e-16
c29873 528 468 3.45e-16
c29874 631 19 1.96e-16
c29875 3310 3702 1.96e-16
c29876 3873 910 3.75e-16
c29877 3870 4559 6.19e-16
c29878 4285 0 3.3589e-14
c29879 4510 4509 5.65e-16
c29880 4504 3667 1.532e-15
c29881 2254 672 5.73e-16
c29882 2646 647 3.64e-16
c29883 1703 1704 1.736e-15
c29884 4760 4762 1.687e-15
c29885 4772 4765 6.73e-16
c29886 4771 4384 1.96e-16
c29887 3177 692 1.832e-15
c29888 1670 1211 1.96e-16
c29889 2077 2067 1.668e-15
c29890 1754 0 3.466e-15
c29891 1 452 4.22e-16
c29892 3393 3433 1.58e-16
c29893 632 2603 1.58e-16
c29894 2196 2439 5.42e-16
c29895 2357 0 1.6491e-14
c29896 4567 4214 1.58e-16
c29897 2194 1743 5.5e-16
c29898 883 868 3.15e-16
c29899 909 827 3.15e-16
c29900 596 807 1.96e-16
c29901 5429 5428 1.062e-15
c29902 2294 2291 5.5e-16
c29903 3321 812 1.58e-16
c29904 5396 5170 1.666e-15
c29905 920 692 3.69e-16
c29906 1629 842 5.03e-16
c29907 1181 1178 1.984e-15
c29908 3900 4438 1.58e-16
c29909 3001 2929 5.95e-16
c29910 2957 2959 1.001e-15
c29911 2639 647 1.9e-16
c29912 1689 1687 1.041e-15
c29913 4231 0 3.5842e-14
c29914 2820 797 1.58e-16
c29915 2557 677 4.46e-16
c29916 1667 1 5.051e-15
c29917 1963 1567 1.96e-16
c29918 1958 1573 1.96e-16
c29919 5069 5079 1.462e-15
c29920 188 190 1.58e-16
c29921 3549 692 3.64e-16
c29922 3048 812 3.15e-16
c29923 2004 2005 1.35e-16
c29924 764 763 1.6e-16
c29925 93 30 3.84e-16
c29926 3710 3709 2.48e-16
c29927 3748 3749 3.92e-16
c29928 2758 2373 1.96e-16
c29929 1803 677 1.58e-16
c29930 1432 1426 1.6e-16
c29931 986 1423 2.386e-15
c29932 2172 762 3.15e-16
c29933 4511 827 1.09e-16
c29934 3667 842 1.58e-16
c29935 3280 0 6.62e-16
c29936 3115 1 6.15e-16
c29937 612 3048 3.58e-16
c29938 806 1 5.57e-16
c29939 2359 722 1.832e-15
c29940 1862 717 2.22e-16
c29941 657 1789 1.58e-16
c29942 3645 1 2.054e-15
c29943 952 1 4.044e-15
c29944 1373 0 6.62e-16
c29945 3430 3424 1.6e-16
c29946 3018 3421 2.386e-15
c29947 612 1743 2.22e-16
c29948 250 252 1.257e-15
c29949 4905 4920 1.96e-16
c29950 2849 837 2.22e-16
c29951 2276 1760 4.11e-16
c29952 3034 2753 1.58e-16
c29953 4799 1 2.378e-15
c29954 777 1905 1.58e-16
c29955 4571 4497 5.5e-16
c29956 4787 352 1.88e-16
c29957 4742 294 1.88e-16
c29958 2178 1885 1.58e-16
c29959 4006 4015 1.88e-16
c29960 2827 2824 5.5e-16
c29961 920 1158 1.58e-16
c29962 392 339 1.88e-16
c29963 4304 3463 4.11e-16
c29964 3480 4314 1.58e-16
c29965 4426 752 1.09e-16
c29966 4770 5160 2.675e-15
c29967 3014 2492 1.96e-16
c29968 2535 2503 3.92e-16
c29969 1321 1520 1.58e-16
c29970 1343 1508 1.58e-16
c29971 779 25 1.13e-15
c29972 783 19 1.58e-16
c29973 1512 1510 1.6e-16
c29974 1507 1506 2.03e-16
c29975 2316 722 1.58e-16
c29976 1465 1837 1.58e-16
c29977 4217 37 1.88e-16
c29978 4226 25 4.68e-16
c29979 4061 1 6.78e-16
c29980 1782 1414 1.96e-16
c29981 601 919 3.15e-16
c29982 3333 3339 1.6e-16
c29983 3330 2815 2.386e-15
c29984 2832 3313 1.58e-16
c29985 1716 1 1.716e-15
c29986 3691 3304 1.532e-15
c29987 3238 3237 1.6e-16
c29988 4564 1 3.358e-15
c29989 3370 3379 1.6e-16
c29990 1694 1969 4.63e-16
c29991 1 355 5.62e-16
c29992 13 363 1.88e-16
c29993 3698 827 1.09e-16
c29994 3304 842 1.58e-16
c29995 822 1930 1.58e-16
c29996 2182 1885 1.58e-16
c29997 2318 1 9.28e-16
c29998 3510 3508 1.6e-16
c29999 3705 3411 5.42e-16
c30000 2371 1862 1.58e-16
c30001 909 812 3.15e-16
c30002 883 1171 1.88e-16
c30003 907 1164 1.58e-16
c30004 4691 5299 8.41e-16
c30005 2822 2441 3.92e-16
c30006 2680 1 1.868e-15
c30007 2654 2265 2.386e-15
c30008 1888 737 1.832e-15
c30009 1516 732 2.22e-16
c30010 2730 1 5.97e-15
c30011 1166 1165 3.94e-16
c30012 2430 782 1.58e-16
c30013 612 909 3.15e-16
c30014 602 894 3.15e-16
c30015 3877 1 2.606e-15
c30016 3046 3070 1.58e-16
c30017 3030 3058 1.58e-16
c30018 1525 1 5.808e-15
c30019 2055 2054 1.6e-16
c30020 2025 2028 3.54e-16
c30021 1527 0 3.466e-15
c30022 26 259 1.03e-15
c30023 5010 4905 1.58e-16
c30024 2066 1 2.53e-16
c30025 657 2645 2.22e-16
c30026 3528 677 1.09e-16
c30027 4311 662 7.68e-16
c30028 894 1006 1.58e-16
c30029 907 978 3.54e-16
c30030 4567 4469 1.58e-16
c30031 761 1 5.57e-16
c30032 3401 3027 1.121e-15
c30033 1694 842 3.15e-16
c30034 538 9 4.88e-16
c30035 4642 4265 2.48e-16
c30036 1346 1 2.86e-16
c30037 3396 3402 1.6e-16
c30038 1865 1 1.056e-15
c30039 288 291 3.54e-16
c30040 9 100 5.8e-16
c30041 13 131 1.88e-16
c30042 412 33 1.88e-16
c30043 3411 3540 1.58e-16
c30044 3397 3553 4.63e-16
c30045 3676 3675 2.48e-16
c30046 687 2288 1.58e-16
c30047 1953 1 4.41e-15
c30048 1044 677 8.3e-16
c30049 2462 0 6.62e-16
c30050 4485 812 7.38e-16
c30051 5535 5544 4.95e-16
c30052 5514 5296 4.35e-16
c30053 4878 381 1.88e-16
c30054 1071 737 1.75e-16
c30055 1275 1276 1.649e-15
c30056 4400 722 1.58e-16
c30057 1959 797 1.58e-16
c30058 1397 1369 2.64e-16
c30059 734 25 1.13e-15
c30060 738 19 1.58e-16
c30061 506 520 3.84e-16
c30062 4174 4171 5.5e-16
c30063 3710 1 5.808e-15
c30064 2503 858 3.15e-16
c30065 1827 1431 1.96e-16
c30066 1822 1437 1.96e-16
c30067 3327 0 3.6368e-14
c30068 528 64 3.08e-16
c30069 4830 4832 2.15e-16
c30070 4839 4828 1.96e-16
c30071 1635 1684 5.5e-16
c30072 1673 1 1.052e-15
c30073 84 71 1.108e-15
c30074 0 49 5.4059e-14
c30075 5395 1 3.36e-16
c30076 1913 2436 4.36e-16
c30077 2434 2427 1.96e-16
c30078 5326 0 4.4446e-14
c30079 3811 3809 1.001e-15
c30080 3554 732 1.58e-16
c30081 2805 1 1.716e-15
c30082 2721 2333 4.97e-16
c30083 911 886 1.58e-16
c30084 5360 5353 9.81e-16
c30085 4174 4176 1.76e-16
c30086 1852 722 1.339e-15
c30087 632 1369 1.75e-16
c30088 3751 3759 1.077e-15
c30089 3024 0 3.17834e-13
c30090 3785 1 2.224e-15
c30091 4172 25 1.88e-16
c30092 4168 19 7.35e-16
c30093 3882 4366 1.96e-16
c30094 1363 1731 1.96e-16
c30095 687 1465 2.22e-16
c30096 929 0 2.4086e-14
c30097 3798 0 2.28e-15
c30098 1643 1191 2.48e-16
c30099 1489 1 1.716e-15
c30100 3876 1 3.564e-15
c30101 3718 4540 1.66e-16
c30102 4717 4711 7.25e-16
c30103 4327 4333 9.42e-16
c30104 617 627 3.28e-16
c30105 19 574 3.2e-16
c30106 5182 1 7.49e-16
c30107 2339 2350 1.58e-16
c30108 5176 0 1.65e-16
c30109 1102 752 6.38e-16
c30110 221 1 3.6e-16
c30111 4787 294 1.88e-16
c30112 4668 5303 1.96e-16
c30113 1585 797 7.68e-16
c30114 2541 2632 1.58e-16
c30115 716 1 5.57e-16
c30116 3964 26 4.58e-16
c30117 1321 1151 5.5e-16
c30118 1331 1610 1.58e-16
c30119 687 1331 7.99e-16
c30120 3520 1 4.41e-15
c30121 2594 3118 4.36e-16
c30122 3116 3109 1.96e-16
c30123 3489 3134 1.58e-16
c30124 3501 3117 1.58e-16
c30125 4354 0 6.62e-16
c30126 2892 2895 1.887e-15
c30127 910 1678 1.58e-16
c30128 569 568 2.84e-16
c30129 3498 647 3.64e-16
c30130 3106 672 5.73e-16
c30131 3270 3638 1.96e-16
c30132 4567 4826 3.92e-16
c30133 5491 410 9.42e-16
c30134 2004 2515 8.31e-16
c30135 762 0 2.8669e-13
c30136 642 3455 1.58e-16
c30137 1375 1372 5.5e-16
c30138 2194 2321 3.92e-16
c30139 1493 722 5.03e-16
c30140 1061 1058 1.984e-15
c30141 2797 2788 3.46e-16
c30142 3000 0 1.65e-16
c30143 1174 1175 7.51e-16
c30144 678 0 7.86e-15
c30145 687 3898 3.15e-16
c30146 3874 3870 1.58e-16
c30147 601 957 3.15e-16
c30148 883 0 3.11441e-13
c30149 2684 677 1.58e-16
c30150 4429 4792 1.96e-16
c30151 3194 732 1.58e-16
c30152 3048 2651 1.58e-16
c30153 3034 3172 1.58e-16
c30154 1638 1 1.056e-15
c30155 3393 3502 1.96e-16
c30156 4793 4800 1.81e-16
c30157 2401 0 6.908e-14
c30158 19 546 3.2e-16
c30159 30 557 6.83e-16
c30160 25 552 5.71e-16
c30161 4571 4605 3.92e-16
c30162 5296 5284 1.75e-16
c30163 1162 1143 1.546e-15
c30164 4253 4254 1.6e-16
c30165 4249 3418 3.92e-16
c30166 3541 0 6.62e-16
c30167 2612 2606 1.6e-16
c30168 2214 2603 2.386e-15
c30169 2231 2586 1.58e-16
c30170 1674 858 1.58e-16
c30171 1459 1455 1.96e-16
c30172 3744 3758 9.34e-16
c30173 2518 2988 2.241e-15
c30174 2521 2990 1.722e-15
c30175 3048 747 3.58e-16
c30176 872 1 4.03e-16
c30177 612 4253 2.72e-16
c30178 1718 1727 3.92e-16
c30179 1721 1318 5.66e-16
c30180 3560 3561 5.65e-16
c30181 4506 1 5.808e-15
c30182 1601 1993 2.38e-15
c30183 1708 1867 3.92e-16
c30184 899 893 1.6e-16
c30185 4508 0 3.466e-15
c30186 3479 3470 3.46e-16
c30187 1726 2235 1.58e-16
c30188 2782 2390 1.96e-16
c30189 1820 702 1.58e-16
c30190 4553 852 3.64e-16
c30191 4540 858 9.97e-16
c30192 601 3447 3.64e-16
c30193 602 3066 1.58e-16
c30194 1121 1117 3.78e-16
c30195 3886 4302 1.58e-16
c30196 3876 3463 5.5e-16
c30197 1728 1727 1.6e-16
c30198 3823 0 1.65e-16
c30199 2291 672 1.58e-16
c30200 1166 1610 1.58e-16
c30201 854 26 2.65e-15
c30202 1684 1849 1.58e-16
c30203 1706 1837 1.58e-16
c30204 4969 4946 1.96e-16
c30205 2317 1800 1.96e-16
c30206 3048 3342 5.42e-16
c30207 3024 3330 1.58e-16
c30208 681 670 7.23e-16
c30209 673 674 1.6e-16
c30210 4859 4860 8.22e-16
c30211 3030 692 3.15e-16
c30212 1715 2221 3.92e-16
c30213 2226 2225 1.6e-16
c30214 9 335 4.88e-16
c30215 3253 3620 1.58e-16
c30216 381 1 3.36e-15
c30217 632 3046 4.46e-16
c30218 1343 662 4.46e-16
c30219 2172 2269 1.58e-16
c30220 2194 2257 1.58e-16
c30221 1046 1045 3.94e-16
c30222 361 37 1.88e-16
c30223 4326 4319 1.96e-16
c30224 5482 5500 1.37e-16
c30225 4838 5136 1.58e-16
c30226 644 25 1.13e-15
c30227 648 19 1.58e-16
c30228 3695 0 3.466e-15
c30229 2577 3088 1.96e-16
c30230 1331 1402 4.63e-16
c30231 3874 4559 1.88e-16
c30232 747 909 3.15e-16
c30233 4571 782 1.33e-16
c30234 1772 1 2.054e-15
c30235 3254 3245 3.92e-16
c30236 2736 3248 5.66e-16
c30237 1774 0 8e-16
c30238 2541 842 3.15e-16
c30239 2545 827 3.15e-16
c30240 2518 858 1.58e-16
c30241 5190 5194 3.54e-16
c30242 3409 3055 1.58e-16
c30243 3393 3438 1.58e-16
c30244 632 2623 1.58e-16
c30245 2196 2444 1.58e-16
c30246 5481 5492 1.619e-15
c30247 4804 5232 2.039e-15
c30248 5270 0 1.5838e-14
c30249 64 325 1.88e-16
c30250 1321 952 1.58e-16
c30251 1327 881 5.5e-16
c30252 2435 837 1.58e-16
c30253 3725 1 4.493e-15
c30254 4068 37 1.88e-16
c30255 4079 0 2.1071e-14
c30256 3254 3255 1.6e-16
c30257 3245 3247 2.15e-16
c30258 3024 3122 3.92e-16
c30259 632 2601 1.339e-15
c30260 2091 2067 6.73e-16
c30261 4462 1 8.43e-16
c30262 4248 0 3.6274e-14
c30263 4698 4696 1.6e-16
c30264 5098 5099 5.87e-16
c30265 1879 2388 1.58e-16
c30266 1684 1 3.564e-15
c30267 3236 2719 1.136e-15
c30268 3168 692 3.15e-16
c30269 4982 4997 6.67e-16
c30270 2291 2298 1.96e-16
c30271 890 692 3.15e-16
c30272 907 1052 3.92e-16
c30273 3397 3219 5.5e-16
c30274 2723 0 6.62e-16
c30275 2528 1 9.43e-16
c30276 4140 4141 7.81e-16
c30277 4582 4531 3.92e-16
c30278 3305 1 1.868e-15
c30279 632 907 4.8e-16
c30280 4623 5409 6.58e-16
c30281 3295 0 2.93e-15
c30282 627 3048 3.58e-16
c30283 2545 2333 5.5e-16
c30284 3252 3243 3.46e-16
c30285 2367 737 3.15e-16
c30286 1600 1136 1.96e-16
c30287 1595 1146 1.96e-16
c30288 809 26 2.65e-15
c30289 4293 4680 2.196e-15
c30290 1398 1 1.868e-15
c30291 3270 777 2.22e-16
c30292 3253 792 1.813e-15
c30293 1388 0 2.93e-15
c30294 617 2251 4.81e-16
c30295 627 1743 3.79e-16
c30296 4816 1 2.378e-15
c30297 2195 2179 3.54e-16
c30298 3409 3591 1.58e-16
c30299 858 865 1.74e-16
c30300 3606 3617 1.96e-16
c30301 617 2220 2.33e-16
c30302 4827 0 2.82384e-13
c30303 2657 2271 5.66e-16
c30304 2342 1 5.808e-15
c30305 2908 1 2.94e-16
c30306 3649 1 8.43e-16
c30307 1990 837 1.58e-16
c30308 1345 1537 5.42e-16
c30309 1321 1525 1.58e-16
c30310 603 19 1.58e-16
c30311 3067 3061 1.6e-16
c30312 2529 3058 2.386e-15
c30313 1076 1504 1.96e-16
c30314 2733 722 4.81e-16
c30315 1465 1857 2.38e-15
c30316 687 1706 3.15e-16
c30317 4488 4487 2.03e-16
c30318 4493 4491 1.6e-16
c30319 2172 722 4.48e-16
c30320 617 919 3.15e-16
c30321 4803 1 8.43e-16
c30322 3606 3610 1.96e-16
c30323 602 1 3.3074e-14
c30324 4747 4743 1.96e-16
c30325 2545 812 3.15e-16
c30326 2331 1 6.15e-16
c30327 2031 2026 7.46e-16
c30328 465 19 3.84e-16
c30329 268 267 3.84e-16
c30330 137 141 1.372e-15
c30331 128 127 6.67e-16
c30332 136 132 1.58e-16
c30333 468 33 3.08e-16
c30334 2464 2461 5.5e-16
c30335 5078 5066 1.37e-16
c30336 1449 677 7.68e-16
c30337 1442 662 1.9e-16
c30338 1188 868 1.05e-15
c30339 890 1158 3.54e-16
c30340 909 1179 1.58e-16
c30341 2758 2759 1.6e-16
c30342 107 27 1.88e-16
c30343 612 2545 7.99e-16
c30344 919 1008 1.58e-16
c30345 1419 1001 1.96e-16
c30346 4040 1 5.1e-16
c30347 911 1322 2.09e-16
c30348 627 909 3.15e-16
c30349 601 894 3.15e-16
c30350 3328 2815 1.532e-15
c30351 1002 0 6.29e-16
c30352 3024 3087 1.58e-16
c30353 3046 3075 1.58e-16
c30354 1708 1573 1.58e-16
c30355 1706 1567 5.5e-16
c30356 1694 1968 1.58e-16
c30357 762 1091 1.813e-15
c30358 747 1106 4.21e-16
c30359 0 194 9.3355e-14
c30360 513 494 1.88e-16
c30361 5032 5056 6.16e-16
c30362 5034 5029 7.46e-16
c30363 672 670 3.327e-15
c30364 2269 2270 9.1e-16
c30365 909 993 3.54e-16
c30366 4328 672 2.65e-16
c30367 4878 5139 1.628e-15
c30368 3355 858 3.15e-16
c30369 657 4285 1.58e-16
c30370 2887 2884 1.96e-16
c30371 2535 2667 3.92e-16
c30372 3392 3038 9.72e-16
c30373 2151 858 9.97e-16
c30374 2162 852 3.64e-16
c30375 632 1771 1.9e-16
c30376 1331 1345 4.274e-15
c30377 1671 1327 1.96e-16
c30378 1482 1041 1.136e-15
c30379 764 26 2.65e-15
c30380 4656 4655 8.22e-16
c30381 1690 1414 5.88e-16
c30382 1350 0 2.96e-16
c30383 4404 762 1.58e-16
c30384 3396 3401 4.17e-16
c30385 1881 1 9.28e-16
c30386 822 1618 2.22e-16
c30387 2194 1783 1.58e-16
c30388 3393 3168 5.88e-16
c30389 5583 1 5.01e-16
c30390 2487 1 1.868e-15
c30391 2477 0 2.93e-15
c30392 4070 857 1.88e-16
c30393 5514 0 5.8355e-14
c30394 911 3048 3.45e-16
c30395 910 3024 5.22e-16
c30396 1534 737 3.64e-16
c30397 2817 2816 1.6e-16
c30398 2809 2807 2.15e-16
c30399 2742 2743 5.65e-16
c30400 1331 1056 1.58e-16
c30401 1329 0 4.64e-16
c30402 1133 1 4.59e-16
c30403 4224 1 6.78e-16
c30404 2701 717 2.4e-16
c30405 1130 0 1.0077e-14
c30406 5010 178 1.88e-16
c30407 3313 3312 2.48e-16
c30408 1885 1886 1.35e-16
c30409 3675 3674 2.03e-16
c30410 3680 3678 1.6e-16
c30411 612 2582 2.4e-16
c30412 1777 1 5.97e-15
c30413 3689 837 2.4e-16
c30414 3797 3732 6.67e-16
c30415 4861 207 1.88e-16
c30416 129 19 3.84e-16
c30417 151 33 3e-16
c30418 5412 5436 1.96e-16
c30419 5440 5456 7.38e-16
c30420 2831 1 8.43e-16
c30421 1173 1186 1.58e-16
c30422 3452 4285 7.84e-16
c30423 921 980 1.96e-16
c30424 1501 1500 1.6e-16
c30425 1493 1491 2.15e-16
c30426 506 549 1.88e-16
c30427 2882 2946 1.6e-16
c30428 2880 2929 2.652e-15
c30429 902 0 7.2392e-14
c30430 3034 3043 1.58e-16
c30431 4344 4333 1.58e-16
c30432 2007 2019 2.32e-16
c30433 5159 236 3.54e-16
c30434 2358 1845 4.97e-16
c30435 223 233 1.88e-16
c30436 230 216 3.84e-16
c30437 4702 0 4.30397e-13
c30438 2722 2339 7.84e-16
c30439 4068 4069 7.45e-16
c30440 4076 4078 2.239e-15
c30441 910 883 5.54e-16
c30442 911 909 3.45e-16
c30443 642 4266 1.58e-16
c30444 3882 4365 1.58e-16
c30445 2702 0 3.5142e-14
c30446 3972 19 3.84e-16
c30447 1345 1166 5.5e-16
c30448 928 0 3.79e-16
c30449 4379 1 1.868e-15
c30450 4627 4625 2.03e-16
c30451 1694 1731 4.63e-16
c30452 1284 1 1.257e-15
c30453 334 252 1.88e-16
c30454 4369 0 2.93e-15
c30455 3411 3304 5.5e-16
c30456 1964 1573 1.136e-15
c30457 88 455 1.88e-16
c30458 15 0 2.10863e-13
c30459 1 27 4.22e-16
c30460 223 305 1.88e-16
c30461 4567 4843 3.92e-16
c30462 4827 4452 4.9e-16
c30463 1027 1008 1.546e-15
c30464 642 3475 1.58e-16
c30465 3196 0 3.466e-15
c30466 2172 2338 3.92e-16
c30467 1253 1248 2.067e-15
c30468 1218 1224 1.58e-16
c30469 4356 4353 5.5e-16
c30470 4455 797 1.58e-16
c30471 922 1115 3.92e-16
c30472 3701 3696 1.642e-15
c30473 1751 1369 2.48e-16
c30474 1327 1436 1.96e-16
c30475 4620 4618 1.6e-16
c30476 1706 1318 1.58e-16
c30477 2559 2557 4.506e-15
c30478 617 957 3.15e-16
c30479 4888 4497 1.96e-16
c30480 4161 0 1.28788e-13
c30481 4152 26 1.075e-15
c30482 4429 4809 1.96e-16
c30483 3214 732 1.58e-16
c30484 3024 2662 5.5e-16
c30485 3034 3177 1.58e-16
c30486 2131 2133 1.609e-15
c30487 2036 2135 9.36e-16
c30488 1658 1667 1.37e-16
c30489 15 514 4.88e-16
c30490 4810 4818 1.81e-16
c30491 5230 5234 1.96e-16
c30492 1 570 3.775e-14
c30493 25 520 7.06e-16
c30494 19 519 3.45e-16
c30495 0 507 1.5696e-14
c30496 292 291 7.03e-16
c30497 4571 4622 3.92e-16
c30498 4907 64 8.88e-16
c30499 2390 2418 2.64e-16
c30500 2412 2408 1.96e-16
c30501 5284 0 3.0268e-14
c30502 59 25 5.71e-16
c30503 64 33 1.88e-16
c30504 3370 2892 4.79e-16
c30505 3809 3852 1.489e-15
c30506 3355 3865 3.38e-16
c30507 1182 812 4.98e-16
c30508 642 3411 3.58e-16
c30509 922 927 2.598e-15
c30510 3556 0 2.93e-15
c30511 2196 807 3.58e-16
c30512 722 0 2.8022e-13
c30513 2545 2786 4.63e-16
c30514 3950 1 6.76e-16
c30515 4134 25 3.84e-16
c30516 4440 4436 1.96e-16
c30517 687 26 1.58e-16
c30518 4580 4592 1.58e-16
c30519 3185 732 1.813e-15
c30520 2224 0 6.62e-16
c30521 5425 5423 3.92e-16
c30522 2299 2697 4.36e-16
c30523 2589 1 2.054e-15
c30524 2249 2243 1.6e-16
c30525 1726 2240 2.386e-15
c30526 909 879 4.9e-16
c30527 3719 3720 1.6e-16
c30528 2214 2601 1.532e-15
c30529 2606 2607 5.65e-16
c30530 1840 702 1.58e-16
c30531 1327 827 3.15e-16
c30532 3731 3734 7.84e-16
c30533 5577 4582 5.76e-16
c30534 627 3072 1.58e-16
c30535 617 3447 7.68e-16
c30536 601 3066 3.15e-16
c30537 1166 1630 2.38e-15
c30538 3177 3176 2.48e-16
c30539 1708 1866 5.42e-16
c30540 1684 1854 1.58e-16
c30541 595 1318 1.58e-16
c30542 1904 1522 2.48e-16
c30543 450 262 1.88e-16
c30544 1811 1800 1.58e-16
c30545 3024 707 4.48e-16
c30546 3174 3175 1.35e-16
c30547 3327 3328 1.35e-16
c30548 894 886 1.58e-16
c30549 883 884 1.534e-15
c30550 5327 5316 6.73e-16
c30551 9 552 5.8e-16
c30552 3236 3628 2.38e-15
c30553 5039 62 4.02e-16
c30554 2494 2495 2.48e-16
c30555 2172 822 3.15e-16
c30556 797 791 1.74e-16
c30557 657 3024 3.15e-16
c30558 1572 767 1.58e-16
c30559 881 877 1.58e-16
c30560 3943 3944 6.4e-16
c30561 2172 2274 1.58e-16
c30562 1487 707 7.38e-16
c30563 2545 747 7.99e-16
c30564 3534 1 1.056e-15
c30565 3718 858 3.15e-16
c30566 3572 747 1.58e-16
c30567 2957 2956 1.624e-15
c30568 2955 2976 6.16e-16
c30569 1188 0 4.6723e-14
c30570 3034 2821 1.58e-16
c30571 2747 3245 1.58e-16
c30572 1790 0 6.72e-16
c30573 3634 3623 1.96e-16
c30574 4777 4779 1.687e-15
c30575 4789 4782 6.73e-16
c30576 4788 4401 1.96e-16
c30577 2535 858 4.48e-16
c30578 2376 1 5.808e-15
c30579 2072 2062 1.021e-15
c30580 420 436 3.84e-16
c30581 1 205 1.456e-15
c30582 4742 4745 6.02e-16
c30583 3642 782 1.832e-15
c30584 2378 0 3.466e-15
c30585 2171 1 2.259e-15
c30586 707 697 6.38e-16
c30587 3798 3775 1.96e-16
c30588 3765 3767 5.66e-16
c30589 3918 3914 8.1e-16
c30590 3932 3926 1.96e-16
c30591 687 3163 1.58e-16
c30592 1041 702 4e-16
c30593 2782 2776 1.6e-16
c30594 2545 2384 5.5e-16
c30595 2680 2681 1.6e-16
c30596 2671 2673 2.15e-16
c30597 1345 966 1.58e-16
c30598 1331 1401 1.58e-16
c30599 1439 1441 2.03e-16
c30600 1191 1198 7.95e-16
c30601 3882 3616 5.88e-16
c30602 3876 3622 1.58e-16
c30603 822 1171 1.35e-16
c30604 3627 3623 1.96e-16
c30605 2070 2066 5.32e-16
c30606 4265 0 3.6274e-14
c30607 1975 1584 4.11e-16
c30608 1121 0 7.4124e-14
c30609 3538 3539 2.03e-16
c30610 3542 3544 1.6e-16
c30611 3907 886 2.538e-15
c30612 4567 4577 1.58e-16
c30613 5108 5103 5.63e-16
c30614 5072 5126 9.34e-16
c30615 4943 4944 1.96e-16
c30616 2748 1 1.868e-15
c30617 883 707 6.45e-16
c30618 909 1067 4.35e-16
c30619 907 1066 1.88e-16
c30620 890 1059 1.58e-16
c30621 952 955 1.58e-16
c30622 111 100 2.45e-16
c30623 2738 0 2.93e-15
c30624 2798 1 5.97e-15
c30625 1327 812 3.15e-16
c30626 657 883 3.15e-16
c30627 2862 2860 1.6e-16
c30628 2857 2856 2.03e-16
c30629 3158 3159 2.03e-16
c30630 2810 812 1.84e-16
c30631 612 1327 4.03e-16
c30632 595 1345 3.15e-16
c30633 602 1321 3.46e-16
c30634 2739 737 1.832e-15
c30635 190 196 1.372e-15
c30636 175 163 1.58e-16
c30637 178 176 6.01e-16
c30638 188 194 3.84e-16
c30639 2298 2289 3.46e-16
c30640 4833 1 2.378e-15
c30641 2753 767 2.33e-16
c30642 5583 4950 3.01e-16
c30643 1053 702 1.58e-16
c30644 595 3388 9.02e-16
c30645 2628 1 5.97e-15
c30646 2194 1896 5.5e-16
c30647 922 1173 1.58e-16
c30648 4315 4314 9.1e-16
c30649 1590 827 1.75e-16
c30650 392 78 1.88e-16
c30651 4268 1 5.808e-15
c30652 4270 0 3.466e-15
c30653 4820 1 8.43e-16
c30654 4480 4830 2e-16
c30655 4847 4463 1.36e-15
c30656 4850 4856 1.6e-16
c30657 3030 3275 1.96e-16
c30658 601 1 3.0651e-14
c30659 3411 3383 3.54e-16
c30660 617 2608 1.09e-16
c30661 2340 1 1.716e-15
c30662 2061 2060 2.67e-16
c30663 1652 1624 2.64e-16
c30664 4589 4595 5.87e-16
c30665 4563 4711 1.58e-16
c30666 4580 4723 1.58e-16
c30667 4708 4713 5.53e-16
c30668 3765 3739 3.54e-16
c30669 1216 1217 1.238e-15
c30670 1207 852 1.58e-16
c30671 1026 1029 1.58e-16
c30672 3879 3885 5.8e-16
c30673 627 2545 7.99e-16
c30674 1517 1508 3.92e-16
c30675 1071 1511 5.66e-16
c30676 3089 0 3.6368e-14
c30677 2923 2931 3.54e-16
c30678 2436 797 7.68e-16
c30679 1414 1786 1.58e-16
c30680 617 894 3.15e-16
c30681 4053 19 9.67e-16
c30682 3048 3104 5.42e-16
c30683 3024 3092 1.58e-16
c30684 4601 1 1.749e-15
c30685 1684 1584 5.5e-16
c30686 1694 1973 1.58e-16
c30687 4593 0 7.67e-16
c30688 0 358 2.87e-16
c30689 209 207 3.84e-16
c30690 30 352 3.84e-16
c30691 27 363 1.88e-16
c30692 3515 3506 3.92e-16
c30693 2374 1862 1.532e-15
c30694 2380 2379 5.65e-16
c30695 3823 3775 1.062e-15
c30696 687 2645 1.813e-15
c30697 894 1008 3.54e-16
c30698 166 158 2.218e-15
c30699 3497 672 3.79e-16
c30700 4319 677 1.58e-16
c30701 5389 5385 1.202e-15
c30702 5588 1 1.601e-15
c30703 4640 468 1.88e-16
c30704 1151 837 1.58e-16
c30705 1331 782 3.15e-16
c30706 3893 1 7.228e-15
c30707 4386 4387 2.48e-16
c30708 5571 5558 8.94e-16
c30709 2559 2684 3.92e-16
c30710 2344 722 5.03e-16
c30711 4659 4282 2.48e-16
c30712 2788 797 1.339e-15
c30713 4402 0 1.6491e-14
c30714 4424 762 1.58e-16
c30715 2987 2954 1.58e-16
c30716 1894 1 6.15e-16
c30717 5001 1 2.73e-16
c30718 3839 4549 1.96e-16
c30719 3332 842 5.03e-16
c30720 762 1907 2.72e-16
c30721 1 467 4.92e-16
c30722 421 136 1.88e-16
c30723 4514 4486 2.64e-16
c30724 4563 4860 1.96e-16
c30725 5290 5278 1.74e-16
c30726 2540 2538 1.041e-15
c30727 1043 692 1.58e-16
c30728 1091 722 3.57e-16
c30729 1309 1307 3.92e-16
c30730 3898 782 4.46e-16
c30731 5560 5529 1.58e-16
c30732 591 1 5.57e-16
c30733 1590 812 2.33e-16
c30734 1414 981 1.136e-15
c30735 3611 0 1.4092e-14
c30736 1839 1448 4.11e-16
c30737 3030 3240 1.58e-16
c30738 3304 3672 1.96e-16
c30739 822 0 2.86609e-13
c30740 122 33 1.88e-16
c30741 131 27 1.88e-16
c30742 3411 732 3.58e-16
c30743 5291 412 1.76e-16
c30744 5072 91 5.5e-16
c30745 4725 323 1.88e-16
c30746 2265 2271 1.418e-15
c30747 2454 2453 1.6e-16
c30748 2446 2444 2.15e-16
c30749 5566 5529 1.52e-16
c30750 2274 0 3.3474e-14
c30751 3804 3808 5.6e-16
c30752 1420 677 1.75e-16
c30753 3463 4268 1.58e-16
c30754 920 994 1.58e-16
c30755 1873 737 5.03e-16
c30756 151 147 6.38e-16
c30757 3047 3031 3.54e-16
c30758 3425 0 6.72e-16
c30759 3839 3734 1.58e-16
c30760 3900 4383 3.92e-16
c30761 4453 4464 1.96e-16
c30762 3317 3315 1.6e-16
c30763 3312 3311 2.03e-16
c30764 1663 1659 1.96e-16
c30765 4734 4728 7.25e-16
c30766 4344 4350 9.42e-16
c30767 2617 662 1.75e-16
c30768 1677 0 2.0654e-14
c30769 117 508 1.88e-16
c30770 4561 0 1.4175e-14
c30771 5045 5047 3.92e-16
c30772 1335 886 1.121e-15
c30773 2807 0 3.3544e-14
c30774 911 2545 3.45e-16
c30775 282 1 1.607e-15
c30776 5379 5365 1.96e-16
c30777 5360 5277 1.67e-16
c30778 5355 5326 1.58e-16
c30779 4872 236 1.88e-16
c30780 3404 0 5.4893e-14
c30781 1410 1408 1.6e-16
c30782 1405 1404 2.03e-16
c30783 3882 4370 1.58e-16
c30784 3898 4382 1.58e-16
c30785 3796 0 2.28e-15
c30786 2559 2649 5.42e-16
c30787 2535 2637 1.58e-16
c30788 1644 1656 2.32e-16
c30789 1211 1253 8.49e-16
c30790 3030 3033 1.96e-16
c30791 1491 0 3.3846e-14
c30792 1920 1539 3.92e-16
c30793 1924 1925 1.6e-16
c30794 204 368 1.88e-16
c30795 5010 4978 1.58e-16
c30796 3034 3030 4.431e-15
c30797 3376 3380 1.96e-16
c30798 236 0 1.25288e-13
c30799 747 1884 2.4e-16
c30800 5544 1 3.85e-16
c30801 2720 2339 3.92e-16
c30802 2639 0 3.466e-15
c30803 592 685 6.34e-16
c30804 1589 807 2.4e-16
c30805 3216 0 8e-16
c30806 3023 1 2.259e-15
c30807 792 2407 1.58e-16
c30808 1504 732 2.4e-16
c30809 1071 1078 7.95e-16
c30810 140 1 2.87e-16
c30811 78 276 1.88e-16
c30812 4475 797 1.58e-16
c30813 919 1129 1.58e-16
c30814 3121 3122 9.1e-16
c30815 1343 1453 3.92e-16
c30816 3701 3707 1.545e-15
c30817 4548 4540 2.15e-16
c30818 2475 868 1.58e-16
c30819 2671 702 1.58e-16
c30820 2500 842 1.09e-16
c30821 3048 2679 5.5e-16
c30822 1735 1747 2.32e-16
c30823 1642 1 1.716e-15
c30824 4333 1 4.442e-15
c30825 4446 4809 1.96e-16
c30826 1708 1652 3.92e-16
c30827 4710 0 2.93e-15
c30828 4827 4832 5.53e-16
c30829 30 294 3.84e-16
c30830 27 310 1.88e-16
c30831 3202 3174 2.64e-16
c30832 3702 3304 4.36e-16
c30833 4571 4639 3.92e-16
c30834 5411 5409 5.25e-16
c30835 2541 2418 5.88e-16
c30836 4272 4271 5.65e-16
c30837 4266 3429 1.532e-15
c30838 919 944 1.687e-15
c30839 2559 3011 1.96e-16
c30840 2905 2895 1.96e-16
c30841 2879 2910 6.73e-16
c30842 1089 0 2.6946e-14
c30843 3696 1 2.054e-15
c30844 2781 3274 1.58e-16
c30845 3192 3194 1.862e-15
c30846 2679 2685 1.418e-15
c30847 3111 647 5.03e-16
c30848 2696 2668 2.64e-16
c30849 1618 1607 1.58e-16
c30850 747 1327 4.03e-16
c30851 25 549 7.06e-16
c30852 453 455 1.257e-15
c30853 49 565 1.88e-16
c30854 3574 3573 2.48e-16
c30855 4580 4609 1.58e-16
c30856 4571 4621 1.58e-16
c30857 2196 1811 5.5e-16
c30858 888 886 2.144e-15
c30859 3491 3487 1.96e-16
c30860 2239 0 2.93e-15
c30861 201 158 1.88e-16
c30862 3577 737 1.84e-16
c30863 592 717 5.8e-16
c30864 5388 5367 2.85e-16
c30865 8 9 4.88e-16
c30866 7 4 1.284e-15
c30867 4132 3390 2.573e-15
c30868 1100 737 5.74e-16
c30869 2773 792 1.58e-16
c30870 1343 852 3.15e-16
c30871 2178 2491 1.96e-16
c30872 3726 3738 1.74e-16
c30873 886 1 9.051e-15
c30874 4150 3918 2.48e-16
c30875 617 3066 3.15e-16
c30876 2879 2881 3.54e-16
c30877 3926 26 4.48e-16
c30878 4640 64 1.88e-16
c30879 2545 2220 1.58e-16
c30880 892 0 4.64e-16
c30881 1708 1871 1.58e-16
c30882 477 483 5.8e-16
c30883 1811 2334 4.36e-16
c30884 4876 4877 8.22e-16
c30885 2770 807 5.73e-16
c30886 1726 2238 1.532e-15
c30887 2243 2244 5.65e-16
c30888 691 689 5.88e-16
c30889 3393 3655 1.96e-16
c30890 2793 2401 2.38e-15
c30891 4060 4063 4.41e-16
c30892 4804 323 1.88e-16
c30893 2182 2491 4.63e-16
c30894 396 390 5.8e-16
c30895 2877 2881 5.6e-16
c30896 59 9 5.8e-16
c30897 2866 3373 1.96e-16
c30898 2977 1 3.36e-16
c30899 4338 4336 2.15e-16
c30900 4346 4345 1.6e-16
c30901 2300 677 7.68e-16
c30902 2293 662 1.9e-16
c30903 1706 782 4.46e-16
c30904 1431 1426 1.642e-15
c30905 3181 3179 1.6e-16
c30906 2305 2691 5.66e-16
c30907 3550 1 9.28e-16
c30908 3287 822 1.813e-15
c30909 1541 1101 2.48e-16
c30910 4591 4590 2.03e-16
c30911 4147 1 6.78e-16
c30912 602 1355 1.832e-15
c30913 2747 3265 2.38e-15
c30914 3409 3083 5.5e-16
c30915 3397 3117 5.5e-16
c30916 2117 2115 3.92e-16
c30917 2103 2108 3.73e-16
c30918 4046 4043 5.5e-16
c30919 5237 5198 3.18e-16
c30920 5113 62 9.42e-16
c30921 0 333 1.5696e-14
c30922 27 339 1.88e-16
c30923 762 1879 1.813e-15
c30924 1896 747 2.22e-16
c30925 2217 1 1.056e-15
c30926 383 33 3e-16
c30927 1031 717 1.58e-16
c30928 894 909 4.274e-15
c30929 627 3073 1.58e-16
c30930 64 526 1.88e-16
c30931 1331 1406 1.58e-16
c30932 687 694 1.6e-16
c30933 59 56 3.54e-16
c30934 3886 4484 1.58e-16
c30935 3898 3633 5.5e-16
c30936 3900 3639 1.58e-16
c30937 3684 4502 1.96e-16
c30938 2969 2968 1.353e-15
c30939 2719 2720 1.35e-16
c30940 2652 677 1.339e-15
c30941 1953 837 5.73e-16
c30942 612 877 1.58e-16
c30943 2545 2756 1.58e-16
c30944 3725 410 7.57e-16
c30945 4129 0 1.11604e-13
c30946 4120 26 1.075e-15
c30947 4420 4422 2.03e-16
c30948 3196 707 1.9e-16
c30949 2108 2101 8.96e-16
c30950 1845 1454 1.136e-15
c30951 4282 0 3.5831e-14
c30952 546 545 1.58e-16
c30953 552 540 1.58e-16
c30954 3168 3536 1.96e-16
c30955 5104 5125 6.16e-16
c30956 5106 5072 1.58e-16
c30957 2188 0 5.86e-16
c30958 5302 0 1.65e-16
c30959 5333 323 3.54e-16
c30960 5086 1 1.257e-15
c30961 2308 2310 2.15e-16
c30962 2673 2669 1.96e-16
c30963 5588 4950 3.96e-16
c30964 5310 5300 3.92e-16
c30965 2754 777 1.58e-16
c30966 4142 4139 5.5e-16
c30967 3341 1 1.056e-15
c30968 3848 1 3.36e-16
c30969 4088 37 5.71e-16
c30970 3565 3571 1.418e-15
c30971 4402 4404 1.862e-15
c30972 2385 737 3.64e-16
c30973 1612 1151 4.11e-16
c30974 1331 1555 4.63e-16
c30975 4310 4697 2.196e-15
c30976 2662 3156 1.96e-16
c30977 1694 1431 5.5e-16
c30978 627 1327 4.03e-16
c30979 601 1321 4.48e-16
c30980 374 378 1.58e-16
c30981 4458 0 1.4092e-14
c30982 1939 1 5.808e-15
c30983 368 175 1.88e-16
c30984 4944 4946 1.035e-15
c30985 3377 858 1.58e-16
c30986 5031 0 3.6422e-14
c30987 2747 782 1.58e-16
c30988 1941 0 3.466e-15
c30989 792 1539 5.73e-16
c30990 3393 3620 1.58e-16
c30991 5286 5288 1.001e-15
c30992 2544 1 2.56e-15
c30993 1072 717 1.58e-16
c30994 627 2248 2.22e-16
c30995 3722 3338 1.58e-16
c30996 1981 2474 1.96e-16
c30997 2172 1913 5.5e-16
c30998 1542 767 1.58e-16
c30999 1357 1353 1.96e-16
c31000 3876 837 3.15e-16
c31001 2628 2634 1.418e-15
c31002 602 955 3e-16
c31003 1607 868 5.73e-16
c31004 1999 827 3.64e-16
c31005 1343 1101 1.58e-16
c31006 4564 4584 9.83e-16
c31007 4288 1 2.054e-15
c31008 1880 1488 1.96e-16
c31009 1881 1874 6.73e-16
c31010 4290 0 8e-16
c31011 4837 1 8.43e-16
c31012 3347 3345 1.862e-15
c31013 3046 3292 3.92e-16
c31014 3267 767 1.09e-16
c31015 538 536 1.58e-16
c31016 617 1 3.1284e-14
c31017 4764 4760 1.96e-16
c31018 2366 1 8.43e-16
c31019 2078 2083 1.96e-16
c31020 4563 4728 1.58e-16
c31021 4580 4740 1.58e-16
c31022 4708 33 1.88e-16
c31023 2486 2481 1.642e-15
c31024 0 447 9.795e-15
c31025 3781 3338 9.7e-16
c31026 2936 1 3.36e-16
c31027 4219 4218 6.4e-16
c31028 2541 2339 1.58e-16
c31029 1076 1508 1.58e-16
c31030 537 117 1.88e-16
c31031 1008 1 1.56e-15
c31032 3667 4484 1.58e-16
c31033 3656 4492 5.66e-16
c31034 4498 4489 3.92e-16
c31035 1930 797 3.15e-16
c31036 2446 807 2.72e-16
c31037 3055 3056 1.35e-16
c31038 4618 1 1.749e-15
c31039 1708 1601 5.5e-16
c31040 4610 0 7.67e-16
c31041 595 19 1.41e-15
c31042 37 491 5.71e-16
c31043 5071 5073 9.16e-16
c31044 3907 3911 3.84e-16
c31045 3915 3914 4.41e-16
c31046 2118 0 2.6642e-14
c31047 103 0 1.051e-14
c31048 4339 677 1.58e-16
c31049 3321 3709 4.97e-16
c31050 1001 1423 1.58e-16
c31051 3900 4417 3.92e-16
c31052 3886 4247 4.63e-16
c31053 2339 732 1.58e-16
c31054 2364 722 1.09e-16
c31055 3393 792 4.03e-16
c31056 3152 3143 3.92e-16
c31057 4673 4672 8.22e-16
c31058 1567 1951 1.58e-16
c31059 251 252 3.84e-16
c31060 1903 1 1.716e-15
c31061 3352 842 1.09e-16
c31062 4563 4877 1.96e-16
c31063 4514 4503 1.58e-16
c31064 2505 1 9.28e-16
c31065 1065 692 6.48e-16
c31066 2475 0 3.6368e-14
c31067 3582 3191 1.136e-15
c31068 4017 4015 1.06e-16
c31069 4004 4006 4.33e-16
c31070 4060 3918 2.87e-16
c31071 1091 1089 1.931e-15
c31072 4506 837 1.58e-16
c31073 2822 2833 1.96e-16
c31074 3090 0 1.6491e-14
c31075 3002 2492 1.96e-16
c31076 920 1175 3.92e-16
c31077 921 1174 2.54e-16
c31078 384 379 1.059e-15
c31079 911 1327 7.6e-16
c31080 4215 4197 6.4e-16
c31081 4214 4568 2.268e-15
c31082 1154 1 3.06e-16
c31083 4896 4934 8.35e-16
c31084 3415 3410 9.6e-16
c31085 9 362 6.48e-16
c31086 1 360 4.59e-16
c31087 15 332 5.8e-16
c31088 3393 737 3.15e-16
c31089 5173 5184 1.96e-16
c31090 4804 265 1.88e-16
c31091 2196 2389 3.92e-16
c31092 165 421 1.88e-16
c31093 5396 0 1.5838e-14
c31094 2294 0 1.4092e-14
c31095 2194 2186 4.63e-16
c31096 921 807 3.15e-16
c31097 1893 737 1.09e-16
c31098 2541 2854 1.96e-16
c31099 782 26 7.12e-16
c31100 4079 2552 2.697e-15
c31101 4216 19 9.67e-16
c31102 617 3463 1.58e-16
c31103 2815 3309 1.96e-16
c31104 3152 662 3.64e-16
c31105 3034 2529 3.54e-16
c31106 2052 2033 6.67e-16
c31107 3344 3345 1.35e-16
c31108 2272 0 1.6491e-14
c31109 0 247 7.7468e-14
c31110 26 262 8.41e-16
c31111 37 258 1.88e-16
c31112 3818 3807 1.96e-16
c31113 5459 439 3.54e-16
c31114 2196 2191 1.58e-16
c31115 1326 898 9.72e-16
c31116 2827 0 1.4092e-14
c31117 3972 1324 2.573e-15
c31118 5356 5363 1.96e-16
c31119 2823 2435 4.97e-16
c31120 2650 2282 1.96e-16
c31121 632 623 1.078e-15
c31122 3650 3645 1.642e-15
c31123 2953 2949 5.87e-16
c31124 1591 812 1.339e-15
c31125 4276 4271 1.642e-15
c31126 632 4287 1.9e-16
c31127 3548 4366 1.96e-16
c31128 2583 2584 1.35e-16
c31129 2338 707 7.38e-16
c31130 1652 852 3.15e-16
c31131 1331 1191 1.58e-16
c31132 962 0 1.018e-14
c31133 1322 1 2.606e-15
c31134 762 764 5.59e-16
c31135 4397 1 9.28e-16
c31136 3684 822 2.22e-16
c31137 4644 4642 2.03e-16
c31138 1690 1764 1.58e-16
c31139 436 424 1.58e-16
c31140 565 194 1.88e-16
c31141 2362 2359 5.5e-16
c31142 4928 4918 1.96e-16
c31143 4549 1 2.54e-16
c31144 427 1 1.607e-15
c31145 215 216 1.482e-15
c31146 403 19 3.45e-16
c31147 407 25 5.71e-16
c31148 284 291 3.54e-16
c31149 657 3089 5.73e-16
c31150 4821 33 1.88e-16
c31151 1778 647 7.68e-16
c31152 3232 0 6.72e-16
c31153 1254 1243 1.58e-15
c31154 1285 1273 5.87e-16
c31155 5530 5533 1.18e-15
c31156 5514 5513 5.5e-16
c31157 1817 702 1.58e-16
c31158 1684 837 3.15e-16
c31159 1557 1116 3.92e-16
c31160 1561 1562 1.6e-16
c31161 1321 1470 3.92e-16
c31162 4637 4635 1.6e-16
c31163 1684 1319 5.5e-16
c31164 3321 1 5.97e-15
c31165 2691 702 1.58e-16
c31166 1668 1 5.01e-16
c31167 3411 3519 3.92e-16
c31168 4350 1 4.442e-15
c31169 4446 4826 1.96e-16
c31170 2158 2151 2.15e-16
c31171 1635 1641 1.545e-15
c31172 233 305 1.88e-16
c31173 4727 0 2.93e-15
c31174 4580 4463 5.5e-16
c31175 5259 5265 6.23e-16
c31176 4040 857 3.1e-16
c31177 4571 4656 3.92e-16
c31178 1913 0 6.9108e-14
c31179 3040 0 5.86e-16
c31180 920 767 3.69e-16
c31181 1001 998 1.984e-15
c31182 2557 2435 5.5e-16
c31183 1343 1452 1.58e-16
c31184 1327 1440 1.58e-16
c31185 3048 1 2.222e-15
c31186 2248 2220 2.64e-16
c31187 627 625 3.327e-15
c31188 2669 702 1.58e-16
c31189 1431 1815 1.58e-16
c31190 3734 1 3.016e-15
c31191 3279 2781 1.58e-16
c31192 2172 672 3.15e-16
c31193 1738 1745 6.73e-16
c31194 3707 1 4.946e-15
c31195 2557 752 4.46e-16
c31196 1 580 4.22e-16
c31197 4580 4626 1.58e-16
c31198 4571 4638 1.58e-16
c31199 1743 1 5.97e-15
c31200 3370 3807 2.037e-15
c31201 3858 3344 8.31e-16
c31202 3338 3853 1.477e-15
c31203 47 46 6.67e-16
c31204 62 30 3.84e-16
c31205 5410 5423 1.96e-16
c31206 4872 4915 1.96e-16
c31207 2715 2714 1.6e-16
c31208 5324 5333 1.58e-16
c31209 5326 5325 5.01e-16
c31210 2620 2619 2.48e-16
c31211 3006 3003 5.5e-16
c31212 1471 717 1.58e-16
c31213 627 3100 2.22e-16
c31214 2685 1 4.41e-15
c31215 2194 2508 3.92e-16
c31216 4668 5511 1.383e-15
c31217 2545 2790 1.58e-16
c31218 3886 3503 1.58e-16
c31219 1181 1176 1.58e-16
c31220 1690 1505 1.58e-16
c31221 612 1352 1.58e-16
c31222 602 1319 1.58e-16
c31223 3578 3576 1.6e-16
c31224 657 2274 1.58e-16
c31225 4915 0 2.39764e-13
c31226 5104 31 1.58e-16
c31227 1607 0 3.6368e-14
c31228 5364 5363 1.6e-16
c31229 907 898 3.98e-16
c31230 3652 3645 6.73e-16
c31231 3651 3259 1.96e-16
c31232 5479 410 9.15e-16
c31233 687 3024 3.15e-16
c31234 1370 1381 1.96e-16
c31235 3967 3966 5.5e-16
c31236 4685 5283 9.82e-16
c31237 2957 1 4.239e-15
c31238 2789 2791 2.03e-16
c31239 1794 677 3.15e-16
c31240 3563 1 6.15e-16
c31241 909 1 2.305e-15
c31242 1905 1917 2.32e-16
c31243 2730 2725 1.642e-15
c31244 601 1355 1.58e-16
c31245 3387 3501 1.58e-16
c31246 4794 4796 1.687e-15
c31247 4806 4799 6.73e-16
c31248 4805 4418 1.96e-16
c31249 657 2646 2.65e-16
c31250 2154 2078 8.32e-16
c31251 596 665 5.28e-16
c31252 1 541 9.8e-16
c31253 3397 677 3.15e-16
c31254 3259 797 1.75e-16
c31255 5407 468 9.68e-16
c31256 4861 497 1.88e-16
c31257 1491 707 1.832e-15
c31258 4250 4249 2.03e-16
c31259 4255 4253 1.6e-16
c31260 2015 2004 1.58e-16
c31261 3347 1 5.808e-15
c31262 3886 4489 1.58e-16
c31263 3876 3650 5.5e-16
c31264 2849 2855 1.545e-15
c31265 2487 837 2.65e-16
c31266 2747 3269 1.96e-16
c31267 2753 3264 1.96e-16
c31268 747 1083 1.05e-15
c31269 657 2639 2.72e-16
c31270 1997 1988 3.46e-16
c31271 19 187 3.84e-16
c31272 3471 3473 2.03e-16
c31273 3796 3775 6.78e-16
c31274 2195 0 1.4914e-14
c31275 797 1157 1.58e-16
c31276 1148 807 1.58e-16
c31277 894 1081 1.58e-16
c31278 907 1053 3.54e-16
c31279 3357 1 9.28e-16
c31280 1644 868 1.58e-16
c31281 1451 1449 1.6e-16
c31282 687 883 3.15e-16
c31283 3911 1 5.1e-16
c31284 4104 25 7.01e-16
c31285 3876 3480 5.5e-16
c31286 3145 2634 1.96e-16
c31287 1879 722 1.58e-16
c31288 1723 1720 3.01e-16
c31289 1719 1716 6.44e-16
c31290 4784 4781 3.01e-16
c31291 1429 1 6.15e-16
c31292 617 1321 4.48e-16
c31293 3453 3455 1.862e-15
c31294 3066 3072 1.418e-15
c31295 3083 3055 2.64e-16
c31296 360 363 1.099e-15
c31297 349 368 1.88e-16
c31298 4954 4946 7.84e-16
c31299 2310 2306 1.96e-16
c31300 792 1948 2.65e-16
c31301 3310 3409 1.58e-16
c31302 4118 3918 2.48e-16
c31303 389 1 4.59e-16
c31304 2867 2858 3.92e-16
c31305 361 0 4.5712e-14
c31306 2559 2542 3.62e-16
c31307 2557 2549 4.63e-16
c31308 601 955 1.58e-16
c31309 595 923 1.58e-16
c31310 841 19 1.96e-16
c31311 1151 1606 1.96e-16
c31312 1499 1488 1.58e-16
c31313 1667 1206 1.958e-15
c31314 3024 3309 3.92e-16
c31315 4854 1 8.43e-16
c31316 596 620 5.28e-16
c31317 223 450 1.88e-16
c31318 4634 4248 1.179e-15
c31319 1981 2473 1.58e-16
c31320 5569 497 7.16e-16
c31321 378 508 1.88e-16
c31322 3886 662 3.15e-16
c31323 3882 677 3.15e-16
c31324 5478 5481 3.54e-16
c31325 5504 5503 1.6e-16
c31326 1455 692 1.339e-15
c31327 1203 858 1.58e-16
c31328 2882 0 3.8149e-14
c31329 1533 752 3.15e-16
c31330 1076 1528 2.38e-15
c31331 1343 971 5.5e-16
c31332 1327 957 5.88e-16
c31333 3075 3074 2.48e-16
c31334 4085 1 7.71e-16
c31335 3667 4489 1.58e-16
c31336 4076 26 4.58e-16
c31337 4068 0 2.3316e-14
c31338 4635 1 1.749e-15
c31339 3046 2600 1.58e-16
c31340 2064 2062 5.66e-16
c31341 1106 1 5.821e-15
c31342 3393 3392 3.15e-16
c31343 642 2616 2.4e-16
c31344 4627 0 7.67e-16
c31345 1641 1 4.946e-15
c31346 2022 236 1.952e-15
c31347 2155 0 6.72e-16
c31348 3883 3899 3.54e-16
c31349 2968 2970 3.92e-16
c31350 1335 1328 7.37e-16
c31351 3344 1 4.946e-15
c31352 4054 25 3.84e-16
c31353 672 0 2.8647e-13
c31354 3275 792 2.4e-16
c31355 3244 3246 2.03e-16
c31356 3809 0 4.0391e-14
c31357 2809 797 1.9e-16
c31358 1584 1939 1.58e-16
c31359 1684 1799 3.92e-16
c31360 4905 4918 1.138e-15
c31361 3384 3382 3.54e-16
c31362 3387 3202 5.5e-16
c31363 2866 3046 3.92e-16
c31364 2299 0 6.9484e-14
c31365 2510 1 1.886e-15
c31366 2191 2192 1.736e-15
c31367 4563 4894 1.96e-16
c31368 4844 1 3.2245e-14
c31369 2569 2571 2.15e-16
c31370 4668 497 1.88e-16
c31371 1101 1103 7.72e-16
c31372 3886 4246 1.58e-16
c31373 3898 3381 1.58e-16
c31374 3900 3384 1.58e-16
c31375 3656 827 1.75e-16
c31376 2600 2601 1.35e-16
c31377 1136 1588 1.58e-16
c31378 3242 0 3.6368e-14
c31379 1861 1852 3.46e-16
c31380 4978 3744 1.33e-16
c31381 3411 3027 3.54e-16
c31382 2987 2990 3.54e-16
c31383 3048 3257 5.42e-16
c31384 3024 3245 1.58e-16
c31385 2177 2175 1.041e-15
c31386 4861 4486 4.9e-16
c31387 1 485 1.607e-15
c31388 136 128 1.58e-16
c31389 5044 5034 1.58e-16
c31390 4872 178 1.88e-16
c31391 4708 526 1.88e-16
c31392 2441 822 1.58e-16
c31393 2459 2470 1.96e-16
c31394 5236 238 8.44e-16
c31395 2178 2218 1.58e-16
c31396 1205 868 1.85e-16
c31397 3571 752 1.75e-16
c31398 2760 2758 1.6e-16
c31399 2755 2754 2.03e-16
c31400 919 1025 3.92e-16
c31401 922 1024 2.54e-16
c31402 4200 4201 6.4e-16
c31403 3072 1 4.41e-15
c31404 1321 1322 1.487e-15
c31405 1331 1324 1.58e-16
c31406 3456 0 6.62e-16
c31407 2557 2871 3.92e-16
c31408 4474 3639 1.96e-16
c31409 4479 3633 1.96e-16
c31410 4767 0 8e-16
c31411 2929 858 1.58e-16
c31412 0 178 1.26072e-13
c31413 5188 1 1.88e-16
c31414 5032 5045 1.96e-16
c31415 2196 1681 1.58e-16
c31416 2182 2218 1.58e-16
c31417 1426 662 1.84e-16
c31418 74 71 2.142e-15
c31419 4634 5514 1.58e-16
c31420 2541 2853 1.58e-16
c31421 1161 1162 8.58e-16
c31422 3900 4387 1.58e-16
c31423 3245 762 1.58e-16
c31424 3879 0 8.28e-14
c31425 3133 2611 1.96e-16
c31426 3128 2617 1.96e-16
c31427 1328 1 3.358e-15
c31428 1937 1550 1.532e-15
c31429 1943 1942 5.65e-16
c31430 1706 1781 1.58e-16
c31431 1690 1769 1.58e-16
c31432 3030 767 3.15e-16
c31433 595 2209 1.58e-16
c31434 602 2206 1.832e-15
c31435 295 1 4.92e-16
c31436 5393 5277 1.52e-16
c31437 4844 5081 6.9e-16
c31438 3397 3174 1.58e-16
c31439 3676 3688 2.32e-16
c31440 657 3498 2.65e-16
c31441 3728 3743 3.25e-16
c31442 3866 858 1.58e-16
c31443 5422 1 9.04e-16
c31444 3370 852 1.58e-16
c31445 1397 647 3.15e-16
c31446 1415 1406 3.92e-16
c31447 981 1409 5.66e-16
c31448 3656 812 2.33e-16
c31449 4838 149 1.88e-16
c31450 3064 1 6.15e-16
c31451 2812 2809 3.01e-16
c31452 2808 2805 6.44e-16
c31453 1281 1251 5.69e-16
c31454 3548 4365 1.58e-16
c31455 1811 717 1.58e-16
c31456 2545 2458 1.58e-16
c31457 1345 1487 3.92e-16
c31458 762 769 1.6e-16
c31459 1708 1363 5.5e-16
c31460 3617 762 2.65e-16
c31461 4209 1 4.7375e-14
c31462 4674 4299 4.9e-16
c31463 4571 858 1.33e-16
c31464 4919 4920 3.92e-16
c31465 2798 837 1.58e-16
c31466 1835 0 1.6491e-14
c31467 1755 1752 5.5e-16
c31468 3409 3535 1.58e-16
c31469 747 1888 1.58e-16
c31470 421 291 1.88e-16
c31471 902 901 1.159e-15
c31472 4571 4673 3.92e-16
c31473 595 2166 1.655e-15
c31474 602 2578 3.64e-16
c31475 2257 1 5.808e-15
c31476 2254 2255 1.35e-16
c31477 161 1 1.65e-15
c31478 1508 732 1.58e-16
c31479 3047 0 1.4914e-14
c31480 146 37 1.88e-16
c31481 4284 4285 2.48e-16
c31482 4389 737 5.03e-16
c31483 2535 2452 5.5e-16
c31484 2722 2731 3.92e-16
c31485 1690 677 3.15e-16
c31486 1694 662 3.15e-16
c31487 1321 1469 1.58e-16
c31488 1343 1457 1.58e-16
c31489 536 552 3.84e-16
c31490 3610 762 2.72e-16
c31491 3048 2634 1.58e-16
c31492 1496 1493 3.01e-16
c31493 1492 1489 6.44e-16
c31494 4550 3882 1.96e-16
c31495 3886 3900 4.274e-15
c31496 1448 1803 1.58e-16
c31497 3034 792 7.99e-16
c31498 2942 2918 6.73e-16
c31499 944 1 1.816e-15
c31500 3299 2781 2.38e-15
c31501 3222 3220 1.6e-16
c31502 2017 2016 1.6e-16
c31503 2009 2007 2.15e-16
c31504 1694 1918 4.63e-16
c31505 1644 0 3.372e-14
c31506 762 1345 3.58e-16
c31507 4580 4643 1.58e-16
c31508 4571 4655 1.58e-16
c31509 5155 5159 5.6e-16
c31510 5179 5157 9.18e-16
c31511 824 823 1.6e-16
c31512 333 332 5.8e-16
c31513 3208 737 2.33e-16
c31514 5152 236 3.54e-16
c31515 3463 3072 1.136e-15
c31516 1404 647 1.339e-15
c31517 890 767 3.15e-16
c31518 907 1127 3.92e-16
c31519 407 9 5.8e-16
c31520 223 222 3.84e-16
c31521 4685 1 1.4735e-14
c31522 2632 2265 1.58e-16
c31523 920 931 1.58e-16
c31524 3220 1 1.868e-15
c31525 2393 767 1.58e-16
c31526 1737 1319 4.11e-16
c31527 914 0 2.94e-16
c31528 2308 692 1.58e-16
c31529 601 1319 3.15e-16
c31530 627 1352 5.73e-16
c31531 1474 1 5.808e-15
c31532 1706 1522 1.58e-16
c31533 1476 0 3.466e-15
c31534 747 1071 5.73e-16
c31535 187 195 2.218e-15
c31536 4915 4918 1.881e-15
c31537 5010 4919 1.58e-16
c31538 2352 2351 1.6e-16
c31539 4893 4894 8.22e-16
c31540 3296 812 1.58e-16
c31541 3034 737 3.15e-16
c31542 1 12 9.8e-16
c31543 2624 2622 1.6e-16
c31544 2619 2618 2.03e-16
c31545 3270 3259 1.58e-16
c31546 5200 5240 4.39e-16
c31547 4821 526 1.88e-16
c31548 2194 2507 1.58e-16
c31549 2178 2495 1.58e-16
c31550 2545 1 4.57e-15
c31551 2541 2616 1.96e-16
c31552 705 1 1.65e-16
c31553 4351 4362 1.96e-16
c31554 3572 1 1.716e-15
c31555 4608 4607 2.03e-16
c31556 3485 3117 1.96e-16
c31557 537 378 1.88e-16
c31558 3364 2849 1.885e-15
c31559 911 2186 1.829e-15
c31560 2172 797 4.48e-16
c31561 1814 1 1.056e-15
c31562 3288 2770 1.96e-16
c31563 3253 3644 4.11e-16
c31564 4868 0 6.72e-16
c31565 1012 647 1.58e-16
c31566 1013 672 1.58e-16
c31567 5200 5254 9.34e-16
c31568 5240 5251 3.92e-16
c31569 5151 5224 1.03e-16
c31570 2182 2495 1.58e-16
c31571 3668 797 3.64e-16
c31572 4911 64 9.55e-16
c31573 42 9 5.8e-16
c31574 5522 5296 1.666e-15
c31575 2996 1 3.36e-16
c31576 617 3094 1.9e-16
c31577 2969 0 2.6642e-14
c31578 919 1083 1.58e-16
c31579 78 27 1.88e-16
c31580 3429 4247 1.96e-16
c31581 1542 1554 2.32e-16
c31582 3002 3004 1.6e-16
c31583 3900 3667 5.5e-16
c31584 2673 677 1.9e-16
c31585 1807 1806 5.65e-16
c31586 3726 468 1.163e-15
c31587 1077 0 6.29e-16
c31588 1608 0 1.6491e-14
c31589 4316 0 3.6274e-14
c31590 37 320 1.88e-16
c31591 601 3088 1.58e-16
c31592 2779 1 6.15e-16
c31593 909 1068 3.54e-16
c31594 3713 868 1.58e-16
c31595 2775 777 2.72e-16
c31596 59 48 3.84e-16
c31597 56 42 3.84e-16
c31598 2873 2986 1.58e-16
c31599 602 4243 3.64e-16
c31600 595 3381 1.655e-15
c31601 4432 4430 1.6e-16
c31602 5588 5577 3.92e-16
c31603 3267 3264 3.01e-16
c31604 3263 3260 6.44e-16
c31605 1634 1625 3.46e-16
c31606 1726 2219 1.96e-16
c31607 3409 3236 5.5e-16
c31608 2541 2581 1.58e-16
c31609 627 969 1.58e-16
c31610 2007 842 1.832e-15
c31611 1321 1106 5.5e-16
c31612 1331 1559 1.58e-16
c31613 3469 1 4.41e-15
c31614 3090 3092 1.862e-15
c31615 2577 2583 1.418e-15
c31616 2758 752 1.9e-16
c31617 1499 1897 4.36e-16
c31618 1895 1888 1.96e-16
c31619 1208 1 4.59e-16
c31620 372 361 2.45e-16
c31621 1205 0 1.0077e-14
c31622 4303 0 6.62e-16
c31623 3048 3326 3.92e-16
c31624 1783 1 4.41e-15
c31625 458 465 3.54e-16
c31626 3236 3621 1.96e-16
c31627 4571 4745 1.58e-16
c31628 4582 4757 1.58e-16
c31629 4742 4747 5.53e-16
c31630 5205 5195 1.462e-15
c31631 3397 3467 1.58e-16
c31632 1981 2478 1.58e-16
c31633 978 984 1.58e-16
c31634 5447 0 3.1318e-14
c31635 1041 1042 8.58e-16
c31636 2559 2356 1.58e-16
c31637 642 3900 3.58e-16
c31638 3667 4509 2.38e-15
c31639 1812 1414 4.36e-16
c31640 3749 0 2.078e-15
c31641 4652 1 1.749e-15
c31642 1694 1624 1.58e-16
c31643 1587 1 1.056e-15
c31644 4644 0 7.67e-16
c31645 2362 0 1.4092e-14
c31646 0 455 1.79664e-13
c31647 3723 3393 1.96e-16
c31648 5098 5108 1.125e-15
c31649 687 3156 2.4e-16
c31650 107 100 7.76e-16
c31651 64 207 1.88e-16
c31652 3891 3885 1.6e-16
c31653 4345 692 7.68e-16
c31654 2752 762 2.4e-16
c31655 2170 2569 1.58e-16
c31656 4792 767 1.23e-16
c31657 1176 842 1.75e-16
c31658 1011 1016 1.58e-16
c31659 2611 2606 1.642e-15
c31660 836 1 5.57e-16
c31661 4690 4689 8.22e-16
c31662 2541 662 3.15e-16
c31663 172 171 6.4e-16
c31664 3605 792 5.73e-16
c31665 3437 3055 2.48e-16
c31666 2290 2292 2.03e-16
c31667 2148 0 1.65e-16
c31668 3696 837 1.58e-16
c31669 4804 4799 1.536e-15
c31670 4922 236 1.88e-16
c31671 2769 2384 1.96e-16
c31672 3886 3486 1.58e-16
c31673 4515 827 3.64e-16
c31674 3673 868 5.73e-16
c31675 3109 1 5.808e-15
c31676 2781 2390 1.136e-15
c31677 3886 4251 1.58e-16
c31678 3876 3385 5.5e-16
c31679 3111 0 3.466e-15
c31680 922 1190 3.92e-16
c31681 798 0 7.86e-15
c31682 1151 1576 1.58e-16
c31683 1867 1866 9.1e-16
c31684 3048 3262 1.58e-16
c31685 1905 0 3.3578e-14
c31686 592 757 1.96e-16
c31687 4589 4597 1.81e-16
c31688 4567 4327 5.5e-16
c31689 4021 4015 7.45e-16
c31690 4674 5296 6.17e-16
c31691 2194 2235 1.58e-16
c31692 2178 2223 1.58e-16
c31693 2169 2168 3.54e-16
c31694 3463 3469 1.418e-15
c31695 4300 4302 1.862e-15
c31696 4430 752 3.64e-16
c31697 3481 1 1.868e-15
c31698 1510 1061 4.11e-16
c31699 1327 1335 8.73e-16
c31700 3471 0 2.93e-15
c31701 797 0 2.80345e-13
c31702 2921 2944 1.96e-16
c31703 4784 0 8e-16
c31704 2719 3228 7.84e-16
c31705 3160 677 1.832e-15
c31706 2662 672 2.22e-16
c31707 1723 0 8e-16
c31708 2196 2393 1.58e-16
c31709 4586 0 1.23e-16
c31710 677 671 1.74e-16
c31711 203 201 7.1e-16
c31712 193 192 2.84e-16
c31713 3705 3409 1.58e-16
c31714 3818 3821 3.92e-16
c31715 5428 0 1.65e-16
c31716 747 2367 3.79e-16
c31717 2182 2223 1.58e-16
c31718 1443 672 1.58e-16
c31719 147 150 6.67e-16
c31720 5205 0 1.4815e-14
c31721 287 245 9.5e-16
c31722 5358 5326 1.58e-16
c31723 2827 2441 5.66e-16
c31724 4117 4111 7.45e-16
c31725 2136 2127 8.15e-16
c31726 1166 1163 1.984e-15
c31727 2557 2870 1.58e-16
c31728 2541 2858 1.58e-16
c31729 1778 1386 1.96e-16
c31730 1779 1772 6.73e-16
c31731 2535 2288 1.58e-16
c31732 3024 3071 3.92e-16
c31733 1086 0 3.7577e-14
c31734 4411 1 8.43e-16
c31735 4661 4659 2.03e-16
c31736 2803 782 1.58e-16
c31737 3532 677 3.64e-16
c31738 4537 4980 4.78e-16
c31739 3316 827 1.84e-16
c31740 3024 782 4.48e-16
c31741 601 2206 1.58e-16
c31742 911 3038 1.829e-15
c31743 9 448 5.8e-16
c31744 3786 3781 1.96e-16
c31745 4582 4847 1.58e-16
c31746 4030 3918 6.32e-16
c31747 5536 5540 1.96e-16
c31748 3244 0 2.93e-15
c31749 3073 1 1.716e-15
c31750 1281 1295 1.58e-16
c31751 760 1 3.79e-16
c31752 3548 4370 1.58e-16
c31753 1845 702 2.22e-16
c31754 1327 1657 1.96e-16
c31755 1574 1121 1.532e-15
c31756 1580 1579 5.65e-16
c31757 753 0 7.86e-15
c31758 538 1 1.65e-15
c31759 4654 4652 1.6e-16
c31760 3219 777 1.58e-16
c31761 792 596 1.96e-16
c31762 3383 3382 4.57e-16
c31763 3313 3325 2.32e-16
c31764 3409 3540 1.58e-16
c31765 3679 3686 6.73e-16
c31766 4361 1 6.275e-15
c31767 3231 752 1.84e-16
c31768 592 712 1.96e-16
c31769 275 291 3.84e-16
c31770 1 100 2.946e-15
c31771 3589 3208 3.92e-16
c31772 4571 4690 3.92e-16
c31773 5044 5057 9.34e-16
c31774 601 2578 7.68e-16
c31775 2449 2446 3.01e-16
c31776 2445 2442 6.44e-16
c31777 2277 1 2.054e-15
c31778 5532 5543 6.38e-16
c31779 4725 381 1.88e-16
c31780 1278 1231 7.26e-16
c31781 1251 1243 1.96e-16
c31782 3838 3725 1.58e-16
c31783 2559 2469 5.5e-16
c31784 1345 1486 5.42e-16
c31785 1321 1474 1.58e-16
c31786 146 134 1.58e-16
c31787 3043 3044 1.736e-15
c31788 2299 707 1.58e-16
c31789 2495 852 1.58e-16
c31790 642 1708 3.58e-16
c31791 3713 0 1.4092e-14
c31792 4175 37 1.88e-16
c31793 4012 1 4.64e-16
c31794 1752 1759 1.96e-16
c31795 777 1127 2.68e-16
c31796 4463 4825 1.58e-16
c31797 1694 1708 4.274e-15
c31798 2159 1690 1.96e-16
c31799 1327 1 2.824e-15
c31800 84 88 1.58e-16
c31801 4558 1 1.96e-16
c31802 25 22 7.06e-16
c31803 3208 3590 2.48e-16
c31804 4580 4660 1.58e-16
c31805 4571 4672 1.58e-16
c31806 642 2178 4.03e-16
c31807 889 891 8.21e-16
c31808 3202 752 1.58e-16
c31809 3775 3809 1.58e-16
c31810 2810 1 2.054e-15
c31811 883 782 6.45e-16
c31812 909 1142 4.35e-16
c31813 907 1141 1.88e-16
c31814 890 1134 1.58e-16
c31815 2720 2731 1.96e-16
c31816 5324 5377 3.18e-16
c31817 2812 0 8e-16
c31818 2248 1 5.97e-15
c31819 1098 1099 1.21e-16
c31820 1857 722 1.84e-16
c31821 1499 717 2.22e-16
c31822 3391 0 6.78e-16
c31823 3886 3531 5.5e-16
c31824 2401 782 3.15e-16
c31825 939 1 4.03e-16
c31826 3303 2781 1.96e-16
c31827 3983 37 1.88e-16
c31828 2702 3210 2.48e-16
c31829 2328 692 1.58e-16
c31830 627 1761 2.65e-16
c31831 617 1319 1.58e-16
c31832 612 1380 2.22e-16
c31833 1654 1653 1.6e-16
c31834 1646 1644 2.15e-16
c31835 1494 1 2.054e-15
c31836 3718 3898 3.92e-16
c31837 4714 4711 5.5e-16
c31838 642 2182 7.99e-16
c31839 822 1610 1.58e-16
c31840 1926 1924 1.6e-16
c31841 1921 1920 2.03e-16
c31842 747 1534 2.65e-16
c31843 1496 0 8e-16
c31844 37 577 3.84e-16
c31845 3316 812 1.58e-16
c31846 4294 647 7.68e-16
c31847 5365 5363 3.92e-16
c31848 890 931 1.58e-16
c31849 909 955 1.58e-16
c31850 3270 3668 4.36e-16
c31851 4164 4166 4.33e-16
c31852 239 0 1.4515e-14
c31853 5136 91 1.58e-16
c31854 2048 2046 1.186e-15
c31855 1345 722 3.15e-16
c31856 1391 966 1.96e-16
c31857 2557 2633 3.92e-16
c31858 715 1 3.79e-16
c31859 3960 25 7.01e-16
c31860 2306 692 1.339e-15
c31861 1327 1622 1.58e-16
c31862 708 0 7.86e-15
c31863 4542 4538 1.96e-16
c31864 570 563 7.76e-16
c31865 583 581 6.67e-16
c31866 3294 812 1.339e-15
c31867 2261 2259 1.6e-16
c31868 2256 2255 2.03e-16
c31869 822 1567 1.58e-16
c31870 4823 4816 6.73e-16
c31871 4822 4435 1.96e-16
c31872 4885 0 6.72e-16
c31873 1 309 9.8e-16
c31874 9 274 5.8e-16
c31875 1998 2196 5.5e-16
c31876 2522 2512 1.65e-16
c31877 1896 1 5.97e-15
c31878 3287 797 3.15e-16
c31879 5532 526 3.54e-16
c31880 5522 0 1.5838e-14
c31881 762 19 1.41e-15
c31882 3900 732 3.58e-16
c31883 2801 2799 1.6e-16
c31884 1056 722 1.75e-16
c31885 1226 1229 5.98e-16
c31886 632 984 1.58e-16
c31887 3002 0 3.26e-15
c31888 674 25 1.13e-15
c31889 678 19 1.58e-16
c31890 4333 4334 1.35e-16
c31891 4523 4535 2.32e-16
c31892 2486 842 3.15e-16
c31893 1730 1731 9.1e-16
c31894 117 218 1.88e-16
c31895 64 296 2.84e-16
c31896 617 3088 7.38e-16
c31897 1164 1171 2.27e-16
c31898 894 1083 3.54e-16
c31899 3429 4246 1.58e-16
c31900 3418 4254 5.66e-16
c31901 4260 4251 3.92e-16
c31902 3371 1 5.01e-16
c31903 1835 707 1.339e-15
c31904 1331 858 3.15e-16
c31905 1455 1026 3.92e-16
c31906 1459 1460 1.6e-16
c31907 1384 957 1.58e-16
c31908 602 3385 1.58e-16
c31909 601 4243 7.68e-16
c31910 612 3418 1.58e-16
c31911 3876 4315 3.92e-16
c31912 2879 2874 1.078e-15
c31913 4801 4798 3.01e-16
c31914 864 0 1.1593e-14
c31915 3177 3189 2.32e-16
c31916 3673 0 3.6368e-14
c31917 482 483 2.84e-16
c31918 3483 3481 1.6e-16
c31919 3570 722 7.38e-16
c31920 1590 1 4.41e-15
c31921 1974 0 6.62e-16
c31922 696 685 7.23e-16
c31923 3387 3654 1.58e-16
c31924 1088 722 3.57e-16
c31925 1068 1081 1.58e-16
c31926 5320 5316 3.54e-16
c31927 4922 4905 1.535e-15
c31928 1568 782 7.68e-16
c31929 3882 4314 1.58e-16
c31930 3898 858 1.58e-16
c31931 3886 852 7.99e-16
c31932 4804 381 1.88e-16
c31933 3309 822 2.4e-16
c31934 2891 2876 3.25e-16
c31935 2874 2877 6.71e-16
c31936 920 921 4.47e-15
c31937 4337 4334 6.44e-16
c31938 4341 4338 3.01e-16
c31939 1345 1121 5.5e-16
c31940 1211 1210 3.94e-16
c31941 84 37 1.88e-16
c31942 2022 178 7.57e-16
c31943 1 335 1.65e-15
c31944 215 218 1.099e-15
c31945 3397 3472 1.58e-16
c31946 3411 807 3.58e-16
c31947 4571 4762 1.58e-16
c31948 4582 4774 1.58e-16
c31949 5225 5224 5.87e-16
c31950 5101 62 9.15e-16
c31951 997 999 7.84e-16
c31952 592 622 1.96e-16
c31953 1476 707 5.03e-16
c31954 1046 1043 1.984e-15
c31955 396 0 1.5723e-14
c31956 375 37 5.71e-16
c31957 5482 5503 6.16e-16
c31958 5484 5483 5.68e-16
c31959 5429 5436 3.18e-16
c31960 5422 5409 1.58e-16
c31961 4742 5391 1.628e-15
c31962 920 1069 1.58e-16
c31963 1091 1086 1.58e-16
c31964 3504 0 1.6491e-14
c31965 4117 0 1.5176e-14
c31966 4669 1 1.749e-15
c31967 3177 717 1.58e-16
c31968 3024 2611 5.5e-16
c31969 3034 3126 1.58e-16
c31970 233 450 1.88e-16
c31971 5217 5195 6.67e-16
c31972 3550 3543 6.73e-16
c31973 3549 3157 1.96e-16
c31974 4661 0 7.67e-16
c31975 2392 1885 2.48e-16
c31976 3321 837 3.79e-16
c31977 3855 3393 3.16e-16
c31978 3397 3387 4.116e-15
c31979 4355 702 2.72e-16
c31980 3514 692 3.15e-16
c31981 612 3058 1.58e-16
c31982 2970 0 2.078e-15
c31983 920 717 3.15e-16
c31984 1466 1016 4.36e-16
c31985 3313 0 3.3874e-14
c31986 4079 19 3.84e-16
c31987 4088 0 2.0707e-14
c31988 4403 3565 4.97e-16
c31989 1667 1211 1.96e-16
c31990 4693 4316 2.48e-16
c31991 320 317 3.54e-16
c31992 4459 0 6.72e-16
c31993 5074 5093 4.78e-16
c31994 3616 777 3.79e-16
c31995 4982 4975 8.96e-16
c31996 3048 837 3.58e-16
c31997 2530 1 1.96e-16
c31998 1678 2209 2.38e-15
c31999 1077 707 4.98e-16
c32000 5262 5209 9.01e-16
c32001 4844 410 1.88e-16
c32002 1106 1102 3.78e-16
c32003 3900 3429 5.5e-16
c32004 919 1204 1.58e-16
c32005 2545 2543 5.93e-16
c32006 625 1 3.79e-16
c32007 1708 1815 5.42e-16
c32008 1684 1803 1.58e-16
c32009 3270 0 6.9481e-14
c32010 4564 4197 2.051e-15
c32011 1873 1869 1.96e-16
c32012 4946 4980 1.58e-16
c32013 3030 2770 1.58e-16
c32014 9 449 6.48e-16
c32015 3236 3591 1.58e-16
c32016 3219 3608 2.386e-15
c32017 3617 3611 1.6e-16
c32018 4567 4344 5.5e-16
c32019 4674 0 3.44156e-13
c32020 5136 5106 1.604e-15
c32021 2485 1964 1.96e-16
c32022 2480 1970 1.96e-16
c32023 2172 2252 1.58e-16
c32024 2194 2240 1.58e-16
c32025 1031 1030 3.94e-16
c32026 3599 752 3.15e-16
c32027 2255 647 1.339e-15
c32028 1708 732 3.58e-16
c32029 628 1 1.65e-16
c32030 3100 1 5.97e-15
c32031 3646 0 6.72e-16
c32032 1687 1324 1.96e-16
c32033 2731 732 2.65e-16
c32034 4491 3650 4.11e-16
c32035 2178 732 4.03e-16
c32036 1164 0 2.7376e-14
c32037 4747 4745 2.15e-16
c32038 4743 4754 1.96e-16
c32039 4801 0 8e-16
c32040 1 476 4.59e-16
c32041 245 252 7.76e-16
c32042 3611 3610 1.6e-16
c32043 2327 0 3.466e-15
c32044 2072 1 1.021e-15
c32045 3911 857 3.1e-16
c32046 5039 5028 7.92e-16
c32047 5087 5066 5.87e-16
c32048 2196 1726 5.5e-16
c32049 1011 662 2.33e-16
c32050 909 837 3.15e-16
c32051 98 1 4.22e-16
c32052 1766 2274 7.84e-16
c32053 105 0 9.795e-15
c32054 4332 662 1.58e-16
c32055 602 2557 4.46e-16
c32056 595 2535 1.511e-15
c32057 2781 2776 1.642e-15
c32058 1327 1317 3.54e-16
c32059 1343 1320 1.58e-16
c32060 2739 747 1.58e-16
c32061 2576 2166 1.96e-16
c32062 3882 3565 5.88e-16
c32063 3876 3571 1.58e-16
c32064 2921 2913 3.54e-16
c32065 2418 807 1.813e-15
c32066 2182 732 7.99e-16
c32067 1397 1386 1.58e-16
c32068 2559 2305 1.58e-16
c32069 2545 2700 1.58e-16
c32070 978 0 4.6723e-14
c32071 4048 0 8.5405e-14
c32072 3048 3088 3.92e-16
c32073 822 1345 3.58e-16
c32074 508 494 1.88e-16
c32075 2125 1 7.49e-16
c32076 248 246 1.58e-16
c32077 3151 677 3.15e-16
c32078 5217 0 1.23e-16
c32079 601 2226 1.58e-16
c32080 2115 0 2.078e-15
c32081 4878 5144 5.5e-16
c32082 890 1022 1.96e-16
c32083 4582 4864 1.58e-16
c32084 2756 2367 2.386e-15
c32085 2739 2384 1.58e-16
c32086 2549 2542 7.37e-16
c32087 70 71 1.482e-15
c32088 3099 1 8.43e-16
c32089 779 1 7.18e-16
c32090 1694 852 7.99e-16
c32091 1706 858 1.58e-16
c32092 632 1386 2.33e-16
c32093 1345 1677 3.54e-16
c32094 1321 1327 4.078e-15
c32095 877 1 5.472e-15
c32096 4226 1 6.66e-16
c32097 3412 3394 1.94e-16
c32098 3386 3406 2.07e-16
c32099 3398 3392 2.267e-15
c32100 601 2204 1.339e-15
c32101 3519 662 1.58e-16
c32102 4378 1 6.275e-15
c32103 3293 3304 1.58e-16
c32104 5579 0 3.23e-15
c32105 612 2170 1.813e-15
c32106 2172 1868 1.58e-16
c32107 2178 1862 5.88e-16
c32108 3801 3804 1.099e-15
c32109 5467 5442 5.87e-16
c32110 5444 5446 6.87e-16
c32111 1345 1491 1.58e-16
c32112 911 918 1.88e-16
c32113 2716 707 4.81e-16
c32114 2333 692 1.58e-16
c32115 1211 1673 3.38e-16
c32116 4199 26 1.96e-16
c32117 2194 692 4.46e-16
c32118 4068 2552 1.96e-16
c32119 4842 4463 1.58e-16
c32120 3316 3323 6.73e-16
c32121 2281 1 8.43e-16
c32122 632 2172 4.48e-16
c32123 2043 2042 1.6e-16
c32124 15 262 5.8e-16
c32125 9 252 5.8e-16
c32126 3732 3796 1.6e-16
c32127 4674 4676 4.93e-16
c32128 4580 4677 1.58e-16
c32129 4571 4689 1.58e-16
c32130 2182 1862 5.5e-16
c32131 5442 439 3.15e-16
c32132 1425 647 1.9e-16
c32133 407 408 7.03e-16
c32134 4685 410 1.88e-16
c32135 2828 0 6.72e-16
c32136 2809 2424 1.96e-16
c32137 2254 2636 2.48e-16
c32138 922 963 1.58e-16
c32139 1056 1491 7.84e-16
c32140 3238 1 9.28e-16
c32141 1759 1750 3.46e-16
c32142 958 0 6.29e-16
c32143 3030 3044 3.92e-16
c32144 3048 3052 1.6e-16
c32145 617 1763 4.81e-16
c32146 627 1380 3.79e-16
c32147 1684 1533 5.5e-16
c32148 1694 1922 1.58e-16
c32149 1550 1918 1.96e-16
c32150 425 424 2.84e-16
c32151 325 354 4.71e-16
c32152 2357 2368 1.96e-16
c32153 2043 0 1.65e-16
c32154 4991 1 3.66e-16
c32155 1749 2256 2.48e-16
c32156 1330 886 1.176e-15
c32157 883 923 3.54e-16
c32158 894 969 1.58e-16
c32159 222 233 3.84e-16
c32160 421 13 1.88e-16
c32161 4589 33 1.88e-16
c32162 4855 0 3.06135e-13
c32163 4070 4075 1.96e-16
c32164 4190 3918 6.32e-16
c32165 734 1 7.18e-16
c32166 3974 37 1.88e-16
c32167 4372 3537 1.96e-16
c32168 4377 3531 1.96e-16
c32169 1343 1639 1.58e-16
c32170 1327 1627 1.58e-16
c32171 1563 1561 1.6e-16
c32172 1558 1557 2.03e-16
c32173 4625 4624 2.03e-16
c32174 1275 1 6.11e-16
c32175 2987 2933 1.791e-15
c32176 1818 1 1.716e-15
c32177 3409 3304 5.5e-16
c32178 4889 4883 1.455e-15
c32179 5197 207 5.5e-16
c32180 2153 2149 1.96e-16
c32181 3393 827 3.15e-16
c32182 2438 1 1.056e-15
c32183 1029 1036 2.27e-16
c32184 45 0 1.051e-14
c32185 3998 3918 6.32e-16
c32186 5514 5505 2.85e-16
c32187 1937 807 1.58e-16
c32188 3574 0 3.3874e-14
c32189 1083 1 1.56e-15
c32190 4172 1 4.64e-16
c32191 3886 3690 1.58e-16
c32192 3030 3189 1.58e-16
c32193 2133 2137 1.202e-15
c32194 3574 3586 2.32e-16
c32195 732 739 1.6e-16
c32196 1 569 9.8e-16
c32197 302 304 2.84e-16
c32198 310 309 3.84e-16
c32199 2408 1902 3.92e-16
c32200 2412 2413 1.6e-16
c32201 3370 3847 5.5e-16
c32202 3531 732 1.58e-16
c32203 4793 5240 3.92e-16
c32204 4776 5200 7.84e-16
c32205 2710 2707 3.01e-16
c32206 2706 2703 6.44e-16
c32207 1158 812 1.58e-16
c32208 642 3409 3.15e-16
c32209 3429 4251 1.58e-16
c32210 919 918 1.88e-16
c32211 3001 3014 1.96e-16
c32212 4143 37 1.88e-16
c32213 3951 1 5.195e-15
c32214 627 3418 5.73e-16
c32215 601 3385 3.15e-16
c32216 3900 4332 3.92e-16
c32217 4440 4441 1.6e-16
c32218 4436 3605 3.92e-16
c32219 722 19 1.676e-15
c32220 3275 2764 1.96e-16
c32221 3943 19 3.45e-16
c32222 3941 0 1.5061e-14
c32223 5144 1 1.672e-15
c32224 1999 1 1.868e-15
c32225 796 794 5.88e-16
c32226 1989 0 2.93e-15
c32227 3387 3659 1.58e-16
c32228 3411 3671 5.42e-16
c32229 3393 3276 1.58e-16
c32230 1088 1089 1.213e-15
c32231 592 850 6.34e-16
c32232 42 48 5.8e-16
c32233 4582 4580 4.506e-15
c32234 1121 782 3.15e-16
c32235 1368 881 1.96e-16
c32236 1131 1134 1.58e-16
c32237 2559 2598 5.42e-16
c32238 2535 2586 1.58e-16
c32239 1448 1420 2.64e-16
c32240 617 983 3.57e-16
c32241 4330 1 1.056e-15
c32242 1915 1914 1.6e-16
c32243 1907 1905 2.15e-16
c32244 632 2270 1.58e-16
c32245 3030 717 4.03e-16
c32246 88 368 1.88e-16
c32247 5314 5318 1.088e-15
c32248 1 552 4.22e-16
c32249 3393 812 3.15e-16
c32250 4571 4779 1.58e-16
c32251 4582 4791 1.58e-16
c32252 4821 207 1.88e-16
c32253 4861 468 1.88e-16
c32254 2588 0 3.466e-15
c32255 2504 1987 1.96e-16
c32256 2505 2498 6.73e-16
c32257 797 790 5.58e-16
c32258 3952 3950 1.76e-16
c32259 3165 0 8e-16
c32260 777 2373 5.73e-16
c32261 1496 707 1.09e-16
c32262 612 3393 4.03e-16
c32263 3684 3673 1.58e-16
c32264 2957 2509 4.06e-16
c32265 858 26 7.12e-16
c32266 3366 3362 1.96e-16
c32267 747 1100 1.85e-16
c32268 4686 1 1.749e-15
c32269 3197 717 1.58e-16
c32270 2541 852 4.03e-16
c32271 2036 2064 4.39e-16
c32272 1397 0 6.9481e-14
c32273 1591 1 1.716e-15
c32274 468 471 4.6e-16
c32275 3168 3157 1.58e-16
c32276 2186 1 8.822e-15
c32277 4678 0 7.67e-16
c32278 1868 0 3.6368e-14
c32279 1989 1991 2.03e-16
c32280 26 201 1.03e-15
c32281 3780 3775 3.54e-16
c32282 4922 178 1.88e-16
c32283 612 3078 1.58e-16
c32284 1147 1148 7.46e-16
c32285 4236 3384 1.96e-16
c32286 4241 3381 1.96e-16
c32287 2595 2203 1.96e-16
c32288 2596 2589 6.73e-16
c32289 1655 842 4.81e-16
c32290 537 494 1.88e-16
c32291 3886 4468 4.63e-16
c32292 3333 0 1.4092e-14
c32293 1052 0 1.0183e-14
c32294 2356 752 1.75e-16
c32295 1690 2020 1.96e-16
c32296 632 0 2.80371e-13
c32297 3167 3160 1.96e-16
c32298 2559 702 3.58e-16
c32299 1971 1973 1.862e-15
c32300 1584 1590 1.418e-15
c32301 1601 1573 2.64e-16
c32302 4563 4578 3.92e-16
c32303 5072 5074 1.721e-15
c32304 3168 717 1.813e-15
c32305 3454 3066 4.97e-16
c32306 3693 3700 1.96e-16
c32307 3893 3899 1.988e-15
c32308 5416 5404 1.74e-16
c32309 890 717 3.35e-16
c32310 592 805 6.34e-16
c32311 2170 2593 1.96e-16
c32312 2203 2588 1.96e-16
c32313 1640 827 1.58e-16
c32314 2178 2440 1.96e-16
c32315 4523 842 1.832e-15
c32316 3311 0 1.6491e-14
c32317 1257 1243 1.609e-15
c32318 1749 647 1.75e-16
c32319 595 965 4.62e-16
c32320 644 1 7.18e-16
c32321 1404 0 1.6491e-14
c32322 3438 3450 2.32e-16
c32323 195 194 6.96e-16
c32324 2302 2300 1.6e-16
c32325 3046 2787 1.58e-16
c32326 3046 677 4.46e-16
c32327 1678 2213 1.96e-16
c32328 1681 2208 1.96e-16
c32329 2097 178 2.51e-16
c32330 2773 2384 2.386e-15
c32331 5189 5188 2.67e-16
c32332 2182 2440 4.63e-16
c32333 2196 792 3.58e-16
c32334 877 1317 4.65e-16
c32335 920 842 3.69e-16
c32336 5501 5486 6.67e-16
c32337 5476 5478 5.48e-16
c32338 3165 3162 3.01e-16
c32339 2663 2657 1.6e-16
c32340 1532 1523 3.46e-16
c32341 1343 1367 1.58e-16
c32342 1327 1355 1.58e-16
c32343 3435 0 3.6368e-14
c32344 3034 2764 5.5e-16
c32345 1352 1 4.41e-15
c32346 1736 0 6.62e-16
c32347 4818 0 8e-16
c32348 3409 3383 1.58e-16
c32349 3393 3406 1.58e-16
c32350 2651 692 1.75e-16
c32351 2545 837 7.99e-16
c32352 2345 1 2.054e-15
c32353 2065 2066 2.67e-16
c32354 2073 2062 6.73e-16
c32355 4571 4724 3.92e-16
c32356 339 335 1.58e-16
c32357 3530 3521 3.46e-16
c32358 2347 0 8e-16
c32359 747 2385 2.65e-16
c32360 5452 5459 3.54e-16
c32361 5450 5490 1.062e-15
c32362 3883 3881 8.67e-16
c32363 2657 2656 1.6e-16
c32364 601 2557 4.46e-16
c32365 911 3872 1.88e-16
c32366 4215 3890 5.8e-16
c32367 1321 877 3.54e-16
c32368 3886 4433 1.58e-16
c32369 3898 3582 5.5e-16
c32370 3900 3588 1.58e-16
c32371 3650 4485 1.96e-16
c32372 2196 737 3.15e-16
c32373 1397 1795 4.36e-16
c32374 1793 1786 1.96e-16
c32375 642 922 3.15e-16
c32376 2545 2705 1.58e-16
c32377 1012 0 1.8851e-14
c32378 1690 1985 1.58e-16
c32379 4590 0 1.6462e-14
c32380 4678 4676 2.03e-16
c32381 210 207 4.6e-16
c32382 197 204 3.54e-16
c32383 201 187 3.84e-16
c32384 565 455 1.88e-16
c32385 33 354 1.88e-16
c32386 1862 2379 2.38e-15
c32387 627 2240 1.58e-16
c32388 617 2226 1.84e-16
c32389 751 749 5.88e-16
c32390 4905 4900 7.46e-16
c32391 2699 1 1.056e-15
c32392 1766 2272 3.92e-16
c32393 2277 2276 1.6e-16
c32394 907 677 4.8e-16
c32395 883 1037 3.92e-16
c32396 890 1036 1.88e-16
c32397 277 283 1.372e-15
c32398 276 275 1.88e-16
c32399 165 175 1.88e-16
c32400 2833 822 2.65e-16
c32401 4567 1 4.476e-15
c32402 4582 4881 1.58e-16
c32403 4668 468 1.88e-16
c32404 3272 1 9.28e-16
c32405 2567 2570 6.44e-16
c32406 5558 5561 7.46e-16
c32407 4215 4208 2.697e-15
c32408 4397 4390 6.73e-16
c32409 4396 3554 1.96e-16
c32410 1834 722 1.75e-16
c32411 3634 1 1.868e-15
c32412 3891 0 6.35e-16
c32413 4671 4669 1.6e-16
c32414 3158 2645 1.532e-15
c32415 2793 797 1.84e-16
c32416 4407 0 1.4092e-14
c32417 2708 722 1.84e-16
c32418 1888 1 5.808e-15
c32419 1853 1855 2.03e-16
c32420 3839 4546 1.96e-16
c32421 5022 3751 6.26e-16
c32422 2821 842 1.75e-16
c32423 4395 1 6.275e-15
c32424 3333 3330 5.5e-16
c32425 2736 752 2.33e-16
c32426 762 1522 1.58e-16
c32427 1890 0 3.466e-15
c32428 4861 4865 1.81e-16
c32429 5262 5157 1.58e-16
c32430 3883 3390 1.939e-15
c32431 627 2170 1.58e-16
c32432 118 122 6.38e-16
c32433 3397 752 3.15e-16
c32434 2457 1947 1.96e-16
c32435 101 9 6.48e-16
c32436 3075 0 3.3874e-14
c32437 4861 64 1.88e-16
c32438 543 15 4.88e-16
c32439 3159 2645 4.97e-16
c32440 534 0 9.795e-15
c32441 3394 3404 5.8e-16
c32442 1835 1837 1.862e-15
c32443 1448 1454 1.418e-15
c32444 1465 1437 2.64e-16
c32445 4033 1 1.4213e-14
c32446 1769 1771 2.15e-16
c32447 792 1134 1.58e-16
c32448 3046 3241 3.92e-16
c32449 1709 1 2.86e-16
c32450 687 2299 3.79e-16
c32451 822 19 1.41e-15
c32452 15 195 4.88e-16
c32453 1 181 5.62e-16
c32454 114 26 1.03e-15
c32455 3409 732 3.15e-16
c32456 4691 4698 1.81e-16
c32457 4580 4694 1.58e-16
c32458 4571 4706 1.58e-16
c32459 1936 2444 7.84e-16
c32460 2178 2175 1.123e-15
c32461 3831 3830 1.6e-16
c32462 3806 3361 6.55e-16
c32463 3006 2486 5.69e-16
c32464 894 1156 1.58e-16
c32465 907 1128 3.54e-16
c32466 64 497 1.88e-16
c32467 4181 4182 3.15e-16
c32468 1488 737 1.75e-16
c32469 1061 1474 1.58e-16
c32470 3018 0 4.7674e-14
c32471 59 107 1.88e-16
c32472 3616 4455 2.386e-15
c32473 4464 4458 1.6e-16
c32474 4606 5536 3.65e-16
c32475 2419 782 7.68e-16
c32476 969 1 2.972e-15
c32477 3315 2798 4.11e-16
c32478 970 0 6.29e-16
c32479 4007 37 1.88e-16
c32480 4008 26 1.075e-15
c32481 1659 1196 1.477e-15
c32482 1071 1 4.044e-15
c32483 4546 3701 9.7e-16
c32484 4731 4728 5.5e-16
c32485 1708 1550 5.5e-16
c32486 1509 0 6.62e-16
c32487 5010 4977 1.58e-16
c32488 2182 2175 1.58e-16
c32489 632 3122 1.58e-16
c32490 1119 752 8.3e-16
c32491 280 0 1.5723e-14
c32492 4086 4085 3.15e-16
c32493 1414 647 3.15e-16
c32494 1136 807 1.813e-15
c32495 2327 707 5.03e-16
c32496 1121 1555 1.96e-16
c32497 3393 747 4.03e-16
c32498 2611 3121 1.58e-16
c32499 1931 1922 3.92e-16
c32500 1539 1925 5.66e-16
c32501 1690 1748 1.96e-16
c32502 3030 3380 2e-16
c32503 1844 1 8.43e-16
c32504 4839 4452 1.96e-16
c32505 233 26 8.41e-16
c32506 3411 3140 1.58e-16
c32507 3671 3672 9.1e-16
c32508 2454 1 9.28e-16
c32509 2424 0 3.6368e-14
c32510 3989 3990 3.15e-16
c32511 3038 1 8.822e-15
c32512 5538 526 5.5e-16
c32513 1519 722 4.81e-16
c32514 3882 752 3.15e-16
c32515 366 0 9.795e-15
c32516 2504 842 3.64e-16
c32517 580 563 1.138e-15
c32518 3046 3206 1.58e-16
c32519 3030 3194 1.58e-16
c32520 1647 1 2.054e-15
c32521 1649 0 8e-16
c32522 911 2170 1.88e-16
c32523 602 2536 5.18e-16
c32524 2012 2009 3.01e-16
c32525 2008 2005 6.44e-16
c32526 737 728 1.078e-15
c32527 0 313 1.4803e-14
c32528 37 316 1.88e-16
c32529 3387 702 3.15e-16
c32530 3980 3974 1.96e-16
c32531 5152 5155 1.075e-15
c32532 4776 439 1.88e-16
c32533 5326 294 1.58e-16
c32534 361 364 2.142e-15
c32535 375 377 7.1e-16
c32536 5436 5426 3.92e-16
c32537 5388 5379 2.85e-16
c32538 3429 4271 2.38e-15
c32539 2620 2632 2.32e-16
c32540 1472 1031 1.532e-15
c32541 1478 1477 5.65e-16
c32542 617 608 1.078e-15
c32543 642 971 1.813e-15
c32544 612 3446 2.22e-16
c32545 617 3385 1.58e-16
c32546 627 4277 2.65e-16
c32547 3958 26 4.48e-16
c32548 4818 4815 3.01e-16
c32549 895 0 1.27e-14
c32550 3197 3194 5.5e-16
c32551 2600 647 1.75e-16
c32552 465 450 1.88e-16
c32553 3491 3492 1.6e-16
c32554 3487 3106 3.92e-16
c32555 2347 2344 3.01e-16
c32556 2343 2340 6.44e-16
c32557 706 704 5.88e-16
c32558 3411 3676 1.58e-16
c32559 3397 3689 4.63e-16
c32560 920 925 3.92e-16
c32561 8 1 1.65e-15
c32562 4589 526 5.8e-16
c32563 2214 0 6.904e-14
c32564 1387 957 1.532e-15
c32565 4242 3384 1.136e-15
c32566 3876 4319 1.58e-16
c32567 3900 4331 5.42e-16
c32568 4349 3514 1.96e-16
c32569 4668 64 1.88e-16
c32570 2559 2603 1.58e-16
c32571 1331 1146 1.58e-16
c32572 900 0 5.86e-16
c32573 4346 1 9.28e-16
c32574 3633 822 1.58e-16
c32575 1708 1707 1.866e-15
c32576 535 580 1.88e-16
c32577 2103 2117 2.102e-15
c32578 15 512 6.58e-16
c32579 4571 4796 1.58e-16
c32580 4582 4808 1.58e-16
c32581 5239 5241 3.92e-16
c32582 1998 1987 1.58e-16
c32583 1012 1013 7.46e-16
c32584 807 805 3.327e-15
c32585 102 88 1.88e-16
c32586 3918 3942 2.48e-16
c32587 2923 1 1.021e-15
c32588 1218 858 1.58e-16
c32589 59 1 4.22e-16
c32590 3503 4336 7.84e-16
c32591 4458 782 1.58e-16
c32592 919 1100 3.92e-16
c32593 922 1099 2.54e-16
c32594 627 3393 4.03e-16
c32595 1941 782 1.9e-16
c32596 1552 1551 1.6e-16
c32597 1544 1542 2.15e-16
c32598 1321 1419 3.92e-16
c32599 4591 4592 2.48e-16
c32600 4596 4595 2.83e-16
c32601 4599 3870 1.96e-16
c32602 4134 1 7.08e-16
c32603 2957 2521 2.107e-15
c32604 2657 662 1.58e-16
c32605 612 1368 2.4e-16
c32606 3030 2838 1.58e-16
c32607 1617 1 8.43e-16
c32608 3387 3485 3.92e-16
c32609 4703 1 1.749e-15
c32610 2072 2070 1.09e-15
c32611 596 640 2.45e-16
c32612 1 321 1.456e-15
c32613 233 187 1.88e-16
c32614 4695 0 7.67e-16
c32615 3564 3557 1.96e-16
c32616 3168 3566 4.36e-16
c32617 717 723 1.097e-15
c32618 4580 4564 1.632e-15
c32619 4563 4581 6.81e-16
c32620 4827 352 1.88e-16
c32621 2196 2303 5.42e-16
c32622 890 1235 1.58e-16
c32623 3862 3855 2.15e-16
c32624 2683 2299 1.58e-16
c32625 922 732 3.15e-16
c32626 687 691 2.19e-16
c32627 1327 1418 1.58e-16
c32628 2214 2203 1.58e-16
c32629 1196 1194 1.931e-15
c32630 2541 2768 1.58e-16
c32631 3003 852 2.8e-16
c32632 2070 2125 3.18e-16
c32633 1626 1628 2.03e-16
c32634 3656 1 4.41e-15
c32635 541 535 5.8e-16
c32636 2393 2405 2.32e-16
c32637 4490 0 6.62e-16
c32638 2183 0 1.157e-14
c32639 3387 3869 3.54e-16
c32640 4952 4941 7.27e-16
c32641 5068 1 2.53e-16
c32642 4954 4969 3.92e-16
c32643 3030 842 3.15e-16
c32644 3034 827 3.15e-16
c32645 2308 1800 7.84e-16
c32646 2232 1715 1.96e-16
c32647 3397 3625 1.58e-16
c32648 2754 0 1.6491e-14
c32649 1327 837 4.03e-16
c32650 2194 2457 3.92e-16
c32651 4640 5473 3.92e-16
c32652 4634 5447 1.152e-15
c32653 4623 5412 5.87e-16
c32654 3327 3355 2.64e-16
c32655 1355 877 2.386e-15
c32656 4407 4404 5.5e-16
c32657 1766 672 5.73e-16
c32658 2012 842 1.09e-16
c32659 1608 1610 1.862e-15
c32660 1151 1161 1.418e-15
c32661 1706 1437 1.58e-16
c32662 4994 4946 9.29e-16
c32663 1556 0 3.6368e-14
c32664 435 433 7.1e-16
c32665 4878 120 1.88e-16
c32666 4753 439 1.88e-16
c32667 2178 2439 1.58e-16
c32668 1345 672 3.58e-16
c32669 1353 880 3.92e-16
c32670 1357 1358 1.6e-16
c32671 3798 3355 9.1e-16
c32672 3925 3919 7.55e-16
c32673 5417 381 7.46e-16
c32674 2541 2538 1.123e-15
c32675 1690 752 3.15e-16
c32676 3677 0 6.62e-16
c32677 4223 4225 2.254e-15
c32678 3075 3087 2.32e-16
c32679 1321 1384 1.58e-16
c32680 4513 4504 3.46e-16
c32681 2457 812 7.38e-16
c32682 2211 2208 3.01e-16
c32683 2207 2204 6.44e-16
c32684 1761 1 1.868e-15
c32685 1751 0 2.93e-15
c32686 534 542 1.58e-16
c32687 4764 4762 2.15e-16
c32688 4760 4771 1.96e-16
c32689 4835 0 8e-16
c32690 3393 3021 1.58e-16
c32691 3411 3433 5.42e-16
c32692 3387 3421 1.58e-16
c32693 3186 692 3.64e-16
c32694 2367 1 5.97e-15
c32695 642 2237 1.58e-16
c32696 632 2612 7.68e-16
c32697 4571 4741 3.92e-16
c32698 4725 4350 4.9e-16
c32699 2196 1919 1.58e-16
c32700 2182 2439 1.58e-16
c32701 5025 5062 5.48e-16
c32702 2363 0 6.72e-16
c32703 1031 662 3.57e-16
c32704 890 842 3.15e-16
c32705 907 1202 3.92e-16
c32706 3877 3881 1.988e-15
c32707 3888 3887 6.97e-16
c32708 2963 294 9.36e-16
c32709 617 2557 4.46e-16
c32710 919 692 3.15e-16
c32711 920 1023 1.58e-16
c32712 957 956 3.94e-16
c32713 64 209 1.88e-16
c32714 2854 2486 1.96e-16
c32715 911 3393 7.6e-16
c32716 3296 1 5.808e-15
c32717 3886 4438 1.58e-16
c32718 3876 3599 5.5e-16
c32719 1936 807 1.58e-16
c32720 3356 2838 1.96e-16
c32721 2770 792 1.58e-16
c32722 1696 1695 6.97e-16
c32723 1697 1693 1.71e-16
c32724 1706 2002 1.58e-16
c32725 1690 1990 1.58e-16
c32726 4607 0 1.6462e-14
c32727 1955 1573 2.48e-16
c32728 30 499 3.84e-16
c32729 2106 1 4.071e-15
c32730 3917 3914 5.5e-16
c32731 2131 0 1.2027e-14
c32732 186 185 6.67e-16
c32733 5389 265 3.54e-16
c32734 3034 812 3.15e-16
c32735 2715 1 9.28e-16
c32736 2755 2373 2.48e-16
c32737 3285 1 6.15e-16
c32738 1812 677 7.68e-16
c32739 1805 662 1.9e-16
c32740 986 1432 4.36e-16
c32741 1430 1423 1.96e-16
c32742 612 3034 7.99e-16
c32743 1328 1330 3.67e-16
c32744 4043 25 4.68e-16
c32745 2368 722 3.64e-16
c32746 657 1397 1.813e-15
c32747 3253 1 5.97e-15
c32748 911 1685 2.09e-16
c32749 1378 1 6.15e-16
c32750 3018 3430 4.36e-16
c32751 3428 3421 1.96e-16
c32752 1908 1 2.054e-15
c32753 262 247 1.88e-16
c32754 258 259 6.4e-16
c32755 244 252 1.58e-16
c32756 4950 4957 1.96e-16
c32757 3356 842 3.64e-16
c32758 2273 1760 4.97e-16
c32759 4412 1 6.275e-15
c32760 1910 0 8e-16
c32761 1067 692 1.58e-16
c32762 5136 5115 2.85e-16
c32763 4827 294 1.88e-16
c32764 4702 352 1.88e-16
c32765 910 3018 1.58e-16
c32766 2833 2827 1.6e-16
c32767 3095 0 1.4092e-14
c32768 2518 2526 4.06e-16
c32769 919 1158 1.58e-16
c32770 397 396 3.84e-16
c32771 389 388 6.67e-16
c32772 3480 3469 1.58e-16
c32773 4301 3463 4.97e-16
c32774 1590 837 5.73e-16
c32775 1136 1572 1.96e-16
c32776 1321 1071 1.58e-16
c32777 1327 1061 5.88e-16
c32778 2533 3043 2.79e-16
c32779 3401 3392 5.71e-16
c32780 4217 19 7.04e-16
c32781 1152 0 6.29e-16
c32782 777 1128 1.58e-16
c32783 542 146 1.88e-16
c32784 3330 3337 1.96e-16
c32785 3700 3691 3.46e-16
c32786 1713 0 2.96e-16
c32787 3370 3372 3.2e-16
c32788 1 362 1.073e-15
c32789 1947 2456 1.58e-16
c32790 129 137 2.218e-15
c32791 4691 5283 6.58e-16
c32792 909 1143 3.54e-16
c32793 2859 0 6.62e-16
c32794 280 281 3.84e-16
c32795 3882 3883 1.239e-15
c32796 4219 4164 1.88e-16
c32797 2663 2265 4.36e-16
c32798 1897 737 3.64e-16
c32799 657 1404 1.58e-16
c32800 1913 782 3.15e-16
c32801 1684 1420 1.58e-16
c32802 1771 1767 1.96e-16
c32803 4845 4463 1.443e-15
c32804 3046 2532 1.58e-16
c32805 1534 1 1.868e-15
c32806 1524 0 2.93e-15
c32807 0 267 5.6293e-14
c32808 5284 352 4.44e-16
c32809 4531 4991 1.112e-15
c32810 400 390 8.86e-16
c32811 59 363 1.88e-16
c32812 4300 662 1.339e-15
c32813 2656 2265 4.11e-16
c32814 5136 5051 8.28e-16
c32815 4120 4068 1.88e-16
c32816 2949 2965 9.55e-16
c32817 1596 812 1.84e-16
c32818 632 3452 2.33e-16
c32819 1297 1294 3.92e-16
c32820 1281 1270 1.96e-16
c32821 146 281 1.88e-16
c32822 2322 717 1.58e-16
c32823 2347 707 1.09e-16
c32824 1196 1660 4.78e-16
c32825 1345 1644 1.58e-16
c32826 1471 1472 1.35e-16
c32827 1342 1 2.94e-16
c32828 4642 4641 2.03e-16
c32829 1550 1922 1.58e-16
c32830 1706 1765 3.92e-16
c32831 204 484 1.88e-16
c32832 1334 0 6.35e-16
c32833 3506 672 1.58e-16
c32834 4980 3718 1.58e-16
c32835 4546 1 4.019e-15
c32836 4919 4918 1.334e-15
c32837 216 224 2.218e-15
c32838 420 0 1.5696e-14
c32839 295 292 6.67e-16
c32840 1 120 3.36e-15
c32841 421 27 1.88e-16
c32842 3387 3151 5.5e-16
c32843 3338 868 3.79e-16
c32844 5136 5274 3.54e-16
c32845 2467 1 6.15e-16
c32846 1042 677 1.58e-16
c32847 1023 1029 1.58e-16
c32848 4090 4088 7.1e-16
c32849 5044 5046 1.062e-15
c32850 1283 1243 3.78e-16
c32851 1280 1231 1.96e-16
c32852 1076 1074 1.931e-15
c32853 5533 5535 1.377e-15
c32854 5514 5484 1.604e-15
c32855 657 1012 1.58e-16
c32856 1567 797 3.15e-16
c32857 1958 807 2.72e-16
c32858 1568 1559 3.92e-16
c32859 1116 1562 5.66e-16
c32860 3718 3327 1.136e-15
c32861 4193 1 3.79e-14
c32862 1998 842 3.15e-16
c32863 1819 1437 2.48e-16
c32864 1231 0 2.9078e-14
c32865 4897 4907 1.008e-15
c32866 4175 0 1.8008e-14
c32867 3308 3309 9.1e-16
c32868 3024 3223 1.58e-16
c32869 3046 3211 1.58e-16
c32870 1820 0 3.3874e-14
c32871 1664 1 1.871e-15
c32872 3409 3519 3.92e-16
c32873 17 5 8.86e-16
c32874 426 508 1.88e-16
c32875 5230 5232 1.96e-16
c32876 1663 0 3.792e-15
c32877 2425 1913 1.532e-15
c32878 2431 2430 5.65e-16
c32879 59 131 1.88e-16
c32880 3035 0 1.157e-14
c32881 2718 2333 1.96e-16
c32882 542 320 1.88e-16
c32883 3882 4536 1.96e-16
c32884 2920 2925 3.07e-16
c32885 2535 2803 3.92e-16
c32886 918 1 3.955e-15
c32887 4001 1 9.475e-15
c32888 4167 37 1.88e-16
c32889 4168 26 1.075e-15
c32890 627 3446 3.79e-16
c32891 617 4279 4.81e-16
c32892 1550 1101 1.136e-15
c32893 3983 0 2.1578e-14
c32894 1649 1646 3.01e-16
c32895 1645 1642 6.44e-16
c32896 4713 4714 1.6e-16
c32897 4709 4327 1.443e-15
c32898 297 296 3.84e-16
c32899 117 334 1.88e-16
c32900 889 886 7.84e-16
c32901 2255 0 1.6491e-14
c32902 2017 1 9.28e-16
c32903 3338 3868 1.23e-16
c32904 4810 5232 1.344e-15
c32905 632 3092 1.58e-16
c32906 1102 1083 1.546e-15
c32907 596 863 3.134e-15
c32908 237 1 4.92e-16
c32909 5326 5347 1.96e-16
c32910 2790 2407 7.84e-16
c32911 2541 2802 1.58e-16
c32912 1574 797 1.339e-15
c32913 3900 4336 1.58e-16
c32914 2541 2237 1.58e-16
c32915 3194 3201 1.96e-16
c32916 3107 2594 1.532e-15
c32917 3113 3112 5.65e-16
c32918 3106 3117 1.58e-16
c32919 3100 3488 4.97e-16
c32920 4359 1 6.15e-16
c32921 4915 4916 3.18e-16
c32922 792 921 3.15e-16
c32923 5010 31 3.84e-16
c32924 3309 797 1.58e-16
c32925 2892 2879 1.58e-16
c32926 1953 1954 1.35e-16
c32927 4571 4813 1.58e-16
c32928 4582 4825 1.58e-16
c32929 2707 2322 1.96e-16
c32930 1998 2525 4.69e-16
c32931 2510 2515 2.029e-15
c32932 1381 1375 1.6e-16
c32933 881 1372 2.386e-15
c32934 3178 0 6.62e-16
c32935 3514 4348 1.58e-16
c32936 2535 762 3.15e-16
c32937 2015 2528 1.58e-16
c32938 3557 1 5.808e-15
c32939 2594 3108 4.97e-16
c32940 3559 0 3.466e-15
c32941 1708 1683 2.38e-16
c32942 1684 1680 3.54e-16
c32943 3208 747 1.58e-16
c32944 4525 4523 2.15e-16
c32945 4533 4532 1.6e-16
c32946 1618 1613 1.642e-15
c32947 3034 2651 1.58e-16
c32948 3411 3502 3.92e-16
c32949 4708 497 1.88e-16
c32950 2196 2308 1.58e-16
c32951 921 737 3.15e-16
c32952 59 310 1.88e-16
c32953 3327 858 1.75e-16
c32954 2535 2401 5.5e-16
c32955 2691 2697 1.6e-16
c32956 2688 2299 2.386e-15
c32957 2316 2671 1.58e-16
c32958 4253 3385 4.11e-16
c32959 2214 2612 4.36e-16
c32960 1850 692 1.58e-16
c32961 1461 1459 1.6e-16
c32962 1456 1455 2.03e-16
c32963 1206 1208 7.72e-16
c32964 595 603 1.097e-15
c32965 3882 4501 1.58e-16
c32966 2041 2998 1.33e-16
c32967 3034 747 7.99e-16
c32968 1718 1716 1.862e-15
c32969 4515 1 1.868e-15
c32970 3187 3186 1.6e-16
c32971 2001 1999 1.6e-16
c32972 1694 1867 4.63e-16
c32973 1593 0 3.3592e-14
c32974 479 477 1.88e-16
c32975 316 317 6.4e-16
c32976 567 568 6.67e-16
c32977 3555 732 1.58e-16
c32978 3024 858 4.48e-16
c32979 2320 1811 1.58e-16
c32980 1726 1715 1.58e-16
c32981 5286 5300 1.455e-15
c32982 5262 5240 1.58e-16
c32983 2771 2390 3.92e-16
c32984 2172 2474 3.92e-16
c32985 2890 2874 9.43e-16
c32986 871 1 1.65e-16
c32987 3920 0 3.3562e-14
c32988 3172 3173 9.1e-16
c32989 1684 1454 1.58e-16
c32990 1690 1448 5.88e-16
c32991 1423 1 5.808e-15
c32992 1425 0 3.466e-15
c32993 3458 3455 5.5e-16
c32994 642 2260 1.58e-16
c32995 362 363 1.88e-16
c32996 484 175 1.88e-16
c32997 4905 4946 2.45e-16
c32998 2306 1800 3.92e-16
c32999 3034 3342 1.58e-16
c33000 1682 2225 4.11e-16
c33001 3253 3225 2.64e-16
c33002 2194 2456 1.58e-16
c33003 2178 2444 1.58e-16
c33004 2172 1749 1.58e-16
c33005 361 19 3.84e-16
c33006 2541 2540 3.15e-16
c33007 652 1 5.62e-16
c33008 4323 4322 5.65e-16
c33009 3513 1 8.43e-16
c33010 3692 0 2.93e-15
c33011 4125 1 6.78e-16
c33012 2951 2952 3.54e-16
c33013 2764 767 3.15e-16
c33014 1380 1 5.97e-15
c33015 85 42 1.88e-16
c33016 2730 2736 1.418e-15
c33017 4852 0 8e-16
c33018 3397 3451 4.63e-16
c33019 3411 3438 1.58e-16
c33020 2679 692 3.15e-16
c33021 632 2231 3.15e-16
c33022 5192 5190 8.35e-16
c33023 2182 2444 1.58e-16
c33024 557 553 1.059e-15
c33025 3542 3538 1.96e-16
c33026 3242 782 1.75e-16
c33027 3951 857 1.88e-16
c33028 2165 1 9.43e-16
c33029 5450 5491 1.817e-15
c33030 4804 5265 5.5e-16
c33031 1460 692 1.84e-16
c33032 883 858 6.45e-16
c33033 909 1217 4.35e-16
c33034 907 1216 1.88e-16
c33035 890 1209 1.58e-16
c33036 2739 1 5.808e-15
c33037 59 339 1.88e-16
c33038 3316 1 2.054e-15
c33039 612 596 1.96e-16
c33040 2265 662 3.15e-16
c33041 3829 1 3.36e-16
c33042 4068 19 3.84e-16
c33043 3245 3244 2.48e-16
c33044 1707 1701 1.988e-15
c33045 2062 2067 3.54e-16
c33046 4624 0 1.6462e-14
c33047 4695 4693 2.03e-16
c33048 1557 0 1.6491e-14
c33049 777 1562 1.58e-16
c33050 333 331 2.84e-16
c33051 5072 5069 7.81e-16
c33052 1879 1868 1.58e-16
c33053 3883 3890 7.37e-16
c33054 5004 4977 9.02e-16
c33055 2728 1 6.15e-16
c33056 2294 2295 5.65e-16
c33057 894 692 3.15e-16
c33058 890 1023 3.54e-16
c33059 909 1044 1.58e-16
c33060 2853 2486 1.58e-16
c33061 4567 4531 3.92e-16
c33062 5170 5173 1.817e-15
c33063 687 3504 1.58e-16
c33064 3294 1 1.716e-15
c33065 1345 797 3.15e-16
c33066 627 3034 7.99e-16
c33067 3867 1 7.21e-16
c33068 3882 4264 1.96e-16
c33069 825 1 1.65e-16
c33070 672 19 1.41e-15
c33071 3670 1 1.056e-15
c33072 3338 0 7.0008e-14
c33073 1592 1146 2.48e-16
c33074 1387 1 1.716e-15
c33075 792 794 5.59e-16
c33076 4688 4686 1.6e-16
c33077 3022 3018 1.58e-16
c33078 5291 354 3.19e-16
c33079 4903 4957 1.137e-15
c33080 4979 4980 1.624e-15
c33081 2300 1777 4.36e-16
c33082 4429 1 6.275e-15
c33083 4691 1 1.3956e-14
c33084 3715 3712 3.01e-16
c33085 3710 3397 1.58e-16
c33086 3722 3387 1.58e-16
c33087 4821 497 1.88e-16
c33088 2015 2051 2.31e-16
c33089 1545 752 1.58e-16
c33090 3900 807 3.58e-16
c33091 2756 2763 1.96e-16
c33092 607 1 5.62e-16
c33093 537 426 1.88e-16
c33094 1999 837 2.65e-16
c33095 1345 1086 1.58e-16
c33096 1343 1076 5.5e-16
c33097 1331 1537 1.58e-16
c33098 3418 1 4.41e-15
c33099 2529 3067 4.36e-16
c33100 3065 3058 1.96e-16
c33101 1865 1863 1.6e-16
c33102 4252 0 6.62e-16
c33103 5281 5285 5.6e-16
c33104 3606 3607 2.03e-16
c33105 3887 3401 1.018e-15
c33106 2031 2046 1.96e-16
c33107 923 962 1.96e-16
c33108 465 26 8.41e-16
c33109 459 0 6.224e-15
c33110 268 265 4.6e-16
c33111 2470 2464 1.6e-16
c33112 1947 2461 2.386e-15
c33113 1953 2469 1.136e-15
c33114 1964 2444 1.58e-16
c33115 2194 2219 3.92e-16
c33116 392 204 1.88e-16
c33117 1438 677 1.339e-15
c33118 894 1158 3.54e-16
c33119 4209 4207 1.76e-16
c33120 1516 737 3.15e-16
c33121 1327 1330 1.96e-16
c33122 998 1 4.59e-16
c33123 4052 1 6.78e-16
c33124 3337 3328 3.46e-16
c33125 1414 1386 2.64e-16
c33126 995 0 1.0077e-14
c33127 3024 2566 1.58e-16
c33128 3030 2533 5.5e-16
c33129 1694 1573 1.58e-16
c33130 0 163 9.795e-15
c33131 5032 5028 7.1e-16
c33132 5034 5049 1.96e-16
c33133 2538 2175 1.96e-16
c33134 3830 3775 3.18e-16
c33135 2078 0 6.0252e-14
c33136 1118 767 1.58e-16
c33137 159 165 3.84e-16
c33138 4514 4876 1.58e-16
c33139 74 88 1.58e-16
c33140 1419 1418 9.1e-16
c33141 3872 1 2.346e-15
c33142 1206 1327 1.58e-16
c33143 780 1 1.65e-16
c33144 1550 1942 2.38e-15
c33145 1684 1782 3.92e-16
c33146 1349 0 1.23e-16
c33147 612 2219 2.4e-16
c33148 5383 5385 1.609e-15
c33149 5291 5387 9.36e-16
c33150 3411 3168 5.5e-16
c33151 2866 3360 1.96e-16
c33152 2476 1 1.716e-15
c33153 5561 0 2.3865e-14
c33154 3058 1 5.808e-15
c33155 911 3034 3.45e-16
c33156 1270 1243 1.58e-16
c33157 1086 1088 7.72e-16
c33158 2806 2807 2.48e-16
c33159 3060 0 3.466e-15
c33160 920 1144 1.58e-16
c33161 3129 3130 5.65e-16
c33162 1121 1559 1.58e-16
c33163 2514 852 2.42e-16
c33164 1840 0 1.4092e-14
c33165 5025 180 6.66e-16
c33166 2024 2023 5.87e-16
c33167 1 264 4.92e-16
c33168 166 15 4.88e-16
c33169 1749 0 3.6368e-14
c33170 143 37 5.71e-16
c33171 3554 737 1.75e-16
c33172 5412 5411 5.25e-16
c33173 4295 4288 6.73e-16
c33174 4294 3452 1.96e-16
c33175 922 980 3.92e-16
c33176 3386 1 2.259e-15
c33177 1867 732 2.4e-16
c33178 1490 1491 2.48e-16
c33179 538 535 2.142e-15
c33180 3876 3882 4.078e-15
c33181 3900 4556 3.54e-16
c33182 2918 2931 8.07e-16
c33183 2880 2882 1.96e-16
c33184 2559 2820 3.92e-16
c33185 1751 1753 2.03e-16
c33186 4835 4832 3.01e-16
c33187 2611 672 1.58e-16
c33188 3137 647 4.81e-16
c33189 1624 2007 7.84e-16
c33190 49 305 1.88e-16
c33191 430 436 1.58e-16
c33192 5530 584 9.1e-16
c33193 642 3112 1.58e-16
c33194 2355 1845 1.96e-16
c33195 1409 647 1.84e-16
c33196 379 382 6.67e-16
c33197 407 1 4.22e-16
c33198 4838 1 3.4874e-14
c33199 2866 868 2.22e-16
c33200 4617 0 4.5538e-13
c33201 3633 3242 1.136e-15
c33202 4071 4070 1.58e-16
c33203 3882 3520 1.58e-16
c33204 1319 1352 1.418e-15
c33205 898 0 8.1372e-14
c33206 1331 1166 5.5e-16
c33207 735 1 1.65e-16
c33208 1041 0 3.7577e-14
c33209 2189 1687 1.159e-15
c33210 4368 1 1.716e-15
c33211 4446 4441 1.642e-15
c33212 4541 0 6.78e-16
c33213 1708 1730 5.42e-16
c33214 1684 1718 1.58e-16
c33215 436 484 1.88e-16
c33216 2407 1 4.41e-15
c33217 2621 0 6.62e-16
c33218 1 41 4.59e-16
c33219 642 3083 1.813e-15
c33220 4571 4830 1.58e-16
c33221 4582 4842 1.58e-16
c33222 2717 2350 1.58e-16
c33223 64 412 1.88e-16
c33224 4464 797 7.68e-16
c33225 4702 5347 1.96e-16
c33226 3193 0 2.93e-15
c33227 3017 1 9.43e-16
c33228 1254 1262 3.92e-16
c33229 3531 4336 1.58e-16
c33230 3514 4353 2.386e-15
c33231 4362 4356 1.6e-16
c33232 1811 662 1.58e-16
c33233 1708 807 3.58e-16
c33234 1327 1606 1.96e-16
c33235 2559 777 3.58e-16
c33236 691 19 1.96e-16
c33237 3577 1 2.054e-15
c33238 4608 4609 2.48e-16
c33239 4613 4612 2.83e-16
c33240 4616 3874 1.96e-16
c33241 2545 2557 4.369e-15
c33242 3013 2541 6.89e-16
c33243 2178 807 4.03e-16
c33244 747 596 1.96e-16
c33245 3117 647 3.15e-16
c33246 3134 672 3.79e-16
c33247 3048 2855 1.58e-16
c33248 3046 2849 5.5e-16
c33249 2781 807 1.813e-15
c33250 3642 3640 1.862e-15
c33251 2696 732 1.813e-15
c33252 2131 2022 6.31e-16
c33253 2138 2133 9.94e-16
c33254 1658 2106 4.06e-16
c33255 1 525 4.92e-16
c33256 276 204 1.88e-16
c33257 5232 5241 1.96e-16
c33258 0 531 2.87e-16
c33259 3584 3583 1.6e-16
c33260 2414 2412 1.6e-16
c33261 2409 2408 2.03e-16
c33262 2194 1800 1.58e-16
c33263 2240 1 5.808e-15
c33264 42 1 2.946e-15
c33265 592 852 5.8e-16
c33266 617 2583 2.33e-16
c33267 2982 0 1.2027e-14
c33268 1175 812 5.74e-16
c33269 53 0 6.224e-15
c33270 392 175 1.88e-16
c33271 146 565 1.88e-16
c33272 4372 722 5.03e-16
c33273 1345 1435 5.42e-16
c33274 1321 1423 1.58e-16
c33275 4159 4150 1.96e-16
c33276 3002 3001 1.6e-16
c33277 1031 1453 1.96e-16
c33278 612 1372 1.58e-16
c33279 3882 4506 1.58e-16
c33280 3898 4518 1.58e-16
c33281 2461 827 1.58e-16
c33282 2182 807 7.99e-16
c33283 2559 2785 5.42e-16
c33284 1053 0 4.6723e-14
c33285 4132 37 1.88e-16
c33286 3937 1 2.207e-15
c33287 4143 0 1.8062e-14
c33288 4437 4436 2.03e-16
c33289 4442 4440 1.6e-16
c33290 687 1816 2.4e-16
c33291 2106 2070 1.58e-16
c33292 2535 722 4.48e-16
c33293 595 1721 1.58e-16
c33294 602 1718 1.832e-15
c33295 1613 0 1.4092e-14
c33296 507 505 2.84e-16
c33297 513 508 1.88e-16
c33298 3569 3570 9.1e-16
c33299 4563 3870 1.58e-16
c33300 4571 3873 1.58e-16
c33301 2229 1 6.15e-16
c33302 801 790 7.23e-16
c33303 793 794 1.6e-16
c33304 3191 722 2.33e-16
c33305 2773 1 5.808e-15
c33306 2328 2334 1.6e-16
c33307 2325 1811 2.386e-15
c33308 1828 2308 1.58e-16
c33309 890 1097 1.96e-16
c33310 4838 5081 7.87e-16
c33311 2686 2299 1.532e-15
c33312 1726 2249 4.36e-16
c33313 5321 5331 1.462e-15
c33314 2775 0 3.466e-15
c33315 2170 1 5.277e-15
c33316 73 72 1.88e-16
c33317 1448 702 1.813e-15
c33318 617 3436 1.339e-15
c33319 3171 1 1.056e-15
c33320 1368 957 1.96e-16
c33321 4520 4571 1.58e-16
c33322 4514 4563 5.88e-16
c33323 717 25 1.58e-16
c33324 3175 3179 1.96e-16
c33325 2291 677 1.58e-16
c33326 612 1315 1.58e-16
c33327 1638 1636 1.6e-16
c33328 1708 1471 1.58e-16
c33329 1706 1465 5.5e-16
c33330 1694 1866 1.58e-16
c33331 1910 1907 3.01e-16
c33332 1906 1903 6.44e-16
c33333 484 349 1.88e-16
c33334 455 262 1.88e-16
c33335 5034 0 3.8148e-14
c33336 3387 3638 3.92e-16
c33337 5319 5318 8.03e-16
c33338 1074 732 1.58e-16
c33339 592 832 1.96e-16
c33340 3636 3634 1.6e-16
c33341 993 994 1.21e-16
c33342 4047 4040 1.88e-16
c33343 2475 2503 2.64e-16
c33344 2497 2493 1.96e-16
c33345 2172 2473 1.58e-16
c33346 2194 2461 1.58e-16
c33347 2557 2582 3.92e-16
c33348 1327 1571 1.58e-16
c33349 642 1343 3.15e-16
c33350 602 3397 3.15e-16
c33351 397 146 1.88e-16
c33352 3095 3092 5.5e-16
c33353 2955 2951 6.22e-16
c33354 657 2255 1.58e-16
c33355 2194 767 4.46e-16
c33356 1797 1 1.056e-15
c33357 1414 0 6.915e-14
c33358 3393 3066 5.88e-16
c33359 4777 4788 1.96e-16
c33360 2385 1 1.868e-15
c33361 782 798 1.621e-15
c33362 1 214 4.22e-16
c33363 2196 1947 5.5e-16
c33364 3651 782 3.64e-16
c33365 5457 0 1.4815e-14
c33366 5141 5025 1.52e-16
c33367 2375 0 2.93e-15
c33368 3770 3769 3.54e-16
c33369 3765 3772 8.94e-16
c33370 3027 2538 1.96e-16
c33371 2780 2773 1.96e-16
c33372 4564 3890 2.035e-15
c33373 2671 2670 2.48e-16
c33374 1331 966 1.58e-16
c33375 692 1 3.1284e-14
c33376 627 596 1.96e-16
c33377 4104 1 5.1e-16
c33378 4316 4317 1.35e-16
c33379 2461 812 1.832e-15
c33380 1964 807 2.22e-16
c33381 1760 1369 1.136e-15
c33382 822 1163 1.58e-16
c33383 1708 2007 1.58e-16
c33384 1834 1835 1.35e-16
c33385 3624 3623 2.03e-16
c33386 3629 3627 1.6e-16
c33387 4641 0 1.6462e-14
c33388 1972 1584 4.97e-16
c33389 0 424 9.795e-15
c33390 565 320 1.88e-16
c33391 33 439 1.88e-16
c33392 4563 4559 4.38e-16
c33393 5025 5097 4.16e-16
c33394 3559 707 1.9e-16
c33395 3893 3881 3.225e-15
c33396 4954 4944 5.37e-16
c33397 2737 1 1.716e-15
c33398 883 1038 3.54e-16
c33399 894 1059 1.58e-16
c33400 952 953 8.96e-16
c33401 106 100 5.8e-16
c33402 88 136 1.88e-16
c33403 2858 2486 1.58e-16
c33404 3320 1 8.43e-16
c33405 3898 4281 3.92e-16
c33406 4528 842 1.09e-16
c33407 835 1 3.79e-16
c33408 828 0 7.86e-15
c33409 1413 1 8.43e-16
c33410 595 1331 9.84e-16
c33411 1956 1968 2.32e-16
c33412 175 168 3.54e-16
c33413 3448 3447 1.6e-16
c33414 3440 3438 2.15e-16
c33415 1539 1 4.41e-15
c33416 1923 0 6.62e-16
c33417 4446 1 6.275e-15
c33418 4878 4889 1.88e-16
c33419 4922 4919 1.58e-16
c33420 5283 5280 3.54e-16
c33421 5300 5301 3.92e-16
c33422 4134 857 1.88e-16
c33423 4022 4015 2.45e-16
c33424 3882 4263 1.58e-16
c33425 2600 0 3.5142e-14
c33426 602 936 5.16e-16
c33427 794 25 1.13e-15
c33428 798 19 1.58e-16
c33429 1524 1526 2.03e-16
c33430 602 3882 3.15e-16
c33431 595 3898 3.15e-16
c33432 4277 1 1.868e-15
c33433 2533 2529 1.58e-16
c33434 2787 2788 1.35e-16
c33435 1158 1 1.56e-15
c33436 255 256 1.58e-16
c33437 3433 3434 9.1e-16
c33438 4267 0 2.93e-15
c33439 4847 4854 1.96e-16
c33440 1913 1522 1.136e-15
c33441 276 175 1.88e-16
c33442 3893 3390 1.159e-15
c33443 4589 3870 5.2e-16
c33444 4580 4333 1.58e-16
c33445 5136 5074 6.96e-16
c33446 2172 2236 3.92e-16
c33447 397 320 1.88e-16
c33448 5452 5442 1.021e-15
c33449 5450 5471 1.96e-16
c33450 1026 1027 8.58e-16
c33451 4305 4302 5.5e-16
c33452 1506 1508 1.862e-15
c33453 1061 1071 1.418e-15
c33454 657 1425 2.72e-16
c33455 1020 1 3.06e-16
c33456 797 19 1.676e-15
c33457 4054 1 7.08e-16
c33458 4675 4299 3.92e-16
c33459 2425 797 1.339e-15
c33460 2866 0 6.0538e-14
c33461 4598 1 6.42e-16
c33462 2730 3224 1.96e-16
c33463 3048 2583 1.58e-16
c33464 3046 2577 5.5e-16
c33465 3034 3104 1.58e-16
c33466 1552 1 9.28e-16
c33467 3504 3506 1.862e-15
c33468 4588 0 3.22e-16
c33469 677 670 5.58e-16
c33470 0 368 1.45066e-13
c33471 193 204 3.84e-16
c33472 208 205 6.67e-16
c33473 209 210 3.84e-16
c33474 2540 2175 7.67e-16
c33475 2383 2374 3.46e-16
c33476 5238 0 1.65e-16
c33477 756 745 7.23e-16
c33478 4321 662 1.9e-16
c33479 4328 677 7.68e-16
c33480 2848 2452 1.96e-16
c33481 1140 767 6.48e-16
c33482 3882 3896 3.92e-16
c33483 4514 4893 1.58e-16
c33484 2671 0 3.3717e-14
c33485 3248 0 1.4092e-14
c33486 3393 1 2.824e-15
c33487 4389 4385 1.96e-16
c33488 2545 2684 4.63e-16
c33489 3387 777 3.15e-16
c33490 4659 4658 2.03e-16
c33491 305 194 1.88e-16
c33492 4408 0 6.72e-16
c33493 3582 762 1.813e-15
c33494 745 746 6.67e-16
c33495 422 426 1.58e-16
c33496 1 448 2.946e-15
c33497 4108 4116 6.67e-16
c33498 4114 4104 7.1e-16
c33499 4844 4847 6.02e-16
c33500 2748 2356 1.96e-16
c33501 2542 2544 3.67e-16
c33502 3571 3572 1.35e-16
c33503 3078 1 2.054e-15
c33504 1311 1299 1.18e-15
c33505 3656 837 5.73e-16
c33506 3080 0 8e-16
c33507 2751 2752 9.1e-16
c33508 749 25 1.13e-15
c33509 753 19 1.58e-16
c33510 1121 1579 2.38e-15
c33511 3219 0 6.9481e-14
c33512 1836 1448 4.97e-16
c33513 3030 2719 1.58e-16
c33514 1685 1 2.606e-15
c33515 4915 352 1.88e-16
c33516 827 818 1.078e-15
c33517 1 186 4.59e-16
c33518 15 158 5.8e-16
c33519 223 247 1.88e-16
c33520 3219 3586 1.58e-16
c33521 3208 3594 5.66e-16
c33522 3600 3591 3.92e-16
c33523 5044 5048 2.95e-16
c33524 4810 323 1.88e-16
c33525 2443 2444 2.48e-16
c33526 944 889 3.84e-16
c33527 1231 1226 1.56e-15
c33528 3804 3806 1.133e-15
c33529 64 468 1.88e-16
c33530 2535 822 3.15e-16
c33531 919 994 1.58e-16
c33532 537 513 1.88e-16
c33533 3613 0 8e-16
c33534 3432 1 1.056e-15
c33535 2196 827 3.15e-16
c33536 1820 1832 2.32e-16
c33537 632 1402 7.38e-16
c33538 1127 0 1.0183e-14
c33539 4014 1 6.76e-16
c33540 4184 37 5.71e-16
c33541 3886 4383 4.63e-16
c33542 1684 1690 4.078e-15
c33543 4568 1 3.009e-15
c33544 4730 4731 1.6e-16
c33545 4726 4344 1.443e-15
c33546 4746 0 7.67e-16
c33547 2713 3206 1.58e-16
c33548 1690 1935 1.96e-16
c33549 3591 3593 2.15e-16
c33550 4573 0 6.35e-16
c33551 5036 5033 2.05e-15
c33552 5324 5366 3.15e-16
c33553 4787 236 1.88e-16
c33554 3728 3726 8.88e-16
c33555 3403 0 5.86e-16
c33556 2048 2045 1.84e-16
c33557 2136 2044 1.772e-15
c33558 1769 647 1.58e-16
c33559 1595 797 1.9e-16
c33560 3898 3537 1.58e-16
c33561 2929 2937 1.96e-16
c33562 2559 2819 5.42e-16
c33563 2535 2807 1.58e-16
c33564 2559 2254 1.58e-16
c33565 2557 2248 5.5e-16
c33566 2545 2649 1.58e-16
c33567 3992 37 5.71e-16
c33568 1191 1644 7.84e-16
c33569 3211 3213 2.15e-16
c33570 2786 767 1.58e-16
c33571 1924 1533 4.11e-16
c33572 1708 1735 1.58e-16
c33573 4889 1 9.38e-16
c33574 3364 3048 3.25e-16
c33575 3046 752 4.46e-16
c33576 3202 2685 1.136e-15
c33577 233 15 5.8e-16
c33578 4827 5047 8.41e-16
c33579 2636 0 2.93e-15
c33580 230 25 7.06e-16
c33581 238 33 1.88e-16
c33582 2722 2350 1.58e-16
c33583 2194 2196 4.506e-15
c33584 1343 732 3.15e-16
c33585 4474 807 2.72e-16
c33586 3633 797 3.15e-16
c33587 3226 762 1.58e-16
c33588 1343 1623 3.92e-16
c33589 704 25 1.13e-15
c33590 708 19 1.58e-16
c33591 367 0 1.5723e-14
c33592 4538 3701 1.477e-15
c33593 576 580 1.58e-16
c33594 569 563 5.8e-16
c33595 2259 1743 4.11e-16
c33596 595 1706 3.15e-16
c33597 602 1690 3.15e-16
c33598 3034 2679 5.5e-16
c33599 4709 1 1.806e-15
c33600 3214 737 1.84e-16
c33601 1694 1652 3.92e-16
c33602 1670 2144 5.5e-16
c33603 1 274 2.946e-15
c33604 2524 2196 6.7e-16
c33605 5168 5152 7.48e-16
c33606 2408 0 1.6491e-14
c33607 777 2413 1.58e-16
c33608 1913 2406 1.96e-16
c33609 2172 1817 1.58e-16
c33610 2178 1811 5.88e-16
c33611 3310 3304 1.418e-15
c33612 375 332 1.88e-16
c33613 392 349 1.88e-16
c33614 4275 4266 3.46e-16
c33615 2630 2629 1.6e-16
c33616 151 64 1.88e-16
c33617 3013 3003 3.13e-16
c33618 627 1372 1.58e-16
c33619 2481 827 1.58e-16
c33620 2478 868 1.58e-16
c33621 2196 812 3.15e-16
c33622 762 1112 2.68e-16
c33623 1087 0 1.8851e-14
c33624 3279 3277 1.862e-15
c33625 2770 2764 1.418e-15
c33626 3030 3173 1.96e-16
c33627 2781 2753 2.64e-16
c33628 3192 3203 1.96e-16
c33629 601 1718 1.58e-16
c33630 4533 1 9.28e-16
c33631 3572 3576 1.96e-16
c33632 3661 807 2.72e-16
c33633 4563 3874 5.5e-16
c33634 4571 4231 1.58e-16
c33635 2182 1811 5.5e-16
c33636 2238 1 1.716e-15
c33637 612 2196 3.58e-16
c33638 3493 3491 1.6e-16
c33639 3270 3265 1.642e-15
c33640 3185 737 1.58e-16
c33641 907 752 4.8e-16
c33642 883 1112 3.92e-16
c33643 890 1111 1.88e-16
c33644 2614 1 1.056e-15
c33645 2615 2616 9.1e-16
c33646 612 618 1.097e-15
c33647 3367 1 1.871e-15
c33648 1840 707 1.84e-16
c33649 1677 858 3.15e-16
c33650 1466 1457 3.92e-16
c33651 1026 1460 5.66e-16
c33652 1031 1452 1.58e-16
c33653 4156 3918 2.87e-16
c33654 3366 0 3.792e-15
c33655 3187 1 9.28e-16
c33656 2384 767 3.15e-16
c33657 2396 752 1.58e-16
c33658 870 26 2.65e-15
c33659 3932 26 4.58e-16
c33660 2311 677 1.58e-16
c33661 1684 1482 5.5e-16
c33662 1694 1871 1.58e-16
c33663 4604 4605 8.22e-16
c33664 494 477 1.325e-15
c33665 657 1749 5.73e-16
c33666 3579 722 1.09e-16
c33667 2323 1811 1.532e-15
c33668 4915 294 1.88e-16
c33669 3411 3655 3.92e-16
c33670 4719 323 1.88e-16
c33671 2172 2478 1.58e-16
c33672 1321 692 4.48e-16
c33673 383 412 3.75e-16
c33674 2884 2876 3.54e-16
c33675 3914 25 4.68e-16
c33676 4335 4336 2.48e-16
c33677 2289 677 1.339e-15
c33678 2007 852 1.58e-16
c33679 1343 1588 1.58e-16
c33680 1327 1576 1.58e-16
c33681 632 1345 3.15e-16
c33682 1211 1208 1.984e-15
c33683 601 3397 3.15e-16
c33684 1547 1544 3.01e-16
c33685 1543 1540 6.44e-16
c33686 15 340 4.88e-16
c33687 1006 1007 1.238e-15
c33688 3409 807 3.15e-16
c33689 3729 3732 1.96e-16
c33690 4040 4038 3.54e-16
c33691 4759 4384 4.9e-16
c33692 3270 782 3.15e-16
c33693 3029 2538 7.67e-16
c33694 3876 702 3.15e-16
c33695 4451 782 7.38e-16
c33696 5511 5516 9.94e-16
c33697 4742 5396 5.5e-16
c33698 4776 5262 1.596e-15
c33699 1041 707 1.75e-16
c33700 1203 883 4.5e-16
c33701 1232 1224 9.24e-16
c33702 4366 707 7.38e-16
c33703 1925 767 1.58e-16
c33704 2804 2805 1.35e-16
c33705 55 56 6.4e-16
c33706 78 59 1.88e-16
c33707 3509 0 1.4092e-14
c33708 2954 2968 2.102e-15
c33709 602 1357 1.9e-16
c33710 1059 1 2.972e-15
c33711 3886 3639 1.58e-16
c33712 2650 662 7.38e-16
c33713 4117 19 9.67e-16
c33714 1060 0 6.29e-16
c33715 3030 3138 1.58e-16
c33716 3014 858 1.58e-16
c33717 2116 2070 1.062e-15
c33718 4658 0 1.6462e-14
c33719 2181 1 2.56e-15
c33720 552 535 1.325e-15
c33721 5106 5108 1.001e-15
c33722 5104 5100 5.7e-16
c33723 4810 265 1.88e-16
c33724 2403 2402 1.6e-16
c33725 2395 2393 2.15e-16
c33726 4938 4940 8.11e-16
c33727 2308 2307 2.48e-16
c33728 2763 1 8.43e-16
c33729 3520 702 1.58e-16
c33730 2675 2673 1.6e-16
c33731 2670 2669 2.03e-16
c33732 3760 3759 1.6e-16
c33733 4135 4143 9.33e-16
c33734 4136 4134 3.54e-16
c33735 4088 19 7.35e-16
c33736 4402 4413 1.96e-16
c33737 1516 1511 1.642e-15
c33738 3822 0 2.078e-15
c33739 1609 1151 4.97e-16
c33740 4705 4703 1.6e-16
c33741 2835 812 4.81e-16
c33742 3616 0 6.9118e-14
c33743 3553 707 7.38e-16
c33744 1948 1 1.868e-15
c33745 1938 0 2.93e-15
c33746 3387 3608 1.58e-16
c33747 3411 3620 5.42e-16
c33748 3393 3225 1.58e-16
c33749 1053 707 1.58e-16
c33750 4691 410 1.88e-16
c33751 165 88 1.88e-16
c33752 4640 439 5.88e-16
c33753 2537 0 5.96e-16
c33754 1551 767 7.68e-16
c33755 1359 1357 1.6e-16
c33756 1354 1353 2.03e-16
c33757 3882 4268 1.58e-16
c33758 3898 4280 1.58e-16
c33759 602 953 1.58e-16
c33760 1593 1605 2.32e-16
c33761 1691 1335 2.035e-15
c33762 601 3882 3.15e-16
c33763 3446 1 5.97e-15
c33764 4395 4390 1.642e-15
c33765 3085 3084 1.6e-16
c33766 3077 3075 2.15e-16
c33767 1869 1488 3.92e-16
c33768 1873 1874 1.6e-16
c33769 1389 0 3.3846e-14
c33770 1798 1414 1.58e-16
c33771 3514 3123 1.136e-15
c33772 1 449 1.073e-15
c33773 4606 4231 4.9e-16
c33774 4580 4350 1.58e-16
c33775 4725 4729 1.81e-16
c33776 4793 33 1.88e-16
c33777 1031 1028 1.984e-15
c33778 2900 0 1.6161e-14
c33779 920 1040 3.92e-16
c33780 921 1039 2.54e-16
c33781 3070 3071 9.1e-16
c33782 3487 0 1.6491e-14
c33783 1034 1 3.06e-16
c33784 3667 3639 2.64e-16
c33785 3650 3656 1.418e-15
c33786 4487 4489 1.862e-15
c33787 3349 3345 1.96e-16
c33788 1686 1685 6.67e-16
c33789 4615 1 6.42e-16
c33790 4367 4748 5.66e-16
c33791 4754 4745 3.92e-16
c33792 1694 1601 5.5e-16
c33793 3393 3405 6.67e-16
c33794 1817 0 3.6368e-14
c33795 856 854 5.88e-16
c33796 595 26 1.58e-16
c33797 19 491 8.4e-16
c33798 5064 5068 3.54e-16
c33799 102 0 3.0454e-14
c33800 3708 852 1.58e-16
c33801 3497 677 3.15e-16
c33802 920 662 3.69e-16
c33803 3882 3893 1.96e-16
c33804 2691 0 1.4092e-14
c33805 3886 4417 4.63e-16
c33806 657 1414 3.79e-16
c33807 3411 792 3.58e-16
c33808 3141 3143 1.862e-15
c33809 1567 1556 1.58e-16
c33810 258 262 1.58e-16
c33811 4950 4889 1.119e-15
c33812 2987 2957 6.53e-16
c33813 1998 1993 1.642e-15
c33814 2669 0 1.6491e-14
c33815 4770 4384 1.179e-15
c33816 70 88 1.58e-16
c33817 2178 2389 1.96e-16
c33818 4515 837 2.65e-16
c33819 4736 5177 1.96e-16
c33820 1091 1087 3.78e-16
c33821 3096 0 6.72e-16
c33822 919 1175 3.92e-16
c33823 922 1174 2.54e-16
c33824 2535 2475 1.58e-16
c33825 378 379 7.03e-16
c33826 1684 1786 1.58e-16
c33827 4575 4566 7.06e-16
c33828 1353 0 1.6491e-14
c33829 1691 1 3.358e-15
c33830 3692 3694 2.03e-16
c33831 1 350 1.456e-15
c33832 3411 737 3.15e-16
c33833 2478 0 3.3692e-14
c33834 2182 2389 4.63e-16
c33835 2196 747 3.58e-16
c33836 4321 3486 1.96e-16
c33837 5400 0 1.376e-15
c33838 2194 2192 1.96e-16
c33839 2178 2191 1.58e-16
c33840 922 807 3.15e-16
c33841 134 136 1.257e-15
c33842 3582 722 1.58e-16
c33843 4415 737 4.81e-16
c33844 5446 5447 3.54e-16
c33845 1684 702 3.15e-16
c33846 2646 2637 3.92e-16
c33847 2254 2640 5.66e-16
c33848 3448 1 9.28e-16
c33849 2714 717 2.65e-16
c33850 1211 1327 4.3e-16
c33851 4201 25 7.01e-16
c33852 2957 2015 1.12e-15
c33853 4852 4849 3.01e-16
c33854 2713 3211 1.58e-16
c33855 1 252 1.5625e-14
c33856 2278 0 6.72e-16
c33857 19 258 3.45e-16
c33858 657 2600 5.73e-16
c33859 2182 2191 1.58e-16
c33860 996 647 2.33e-16
c33861 395 390 1.482e-15
c33862 4838 410 1.88e-16
c33863 2820 2435 1.96e-16
c33864 2646 2647 1.6e-16
c33865 2637 2639 2.15e-16
c33866 642 646 2.19e-16
c33867 1871 732 1.58e-16
c33868 3410 0 1.4914e-14
c33869 1151 1155 2.03e-16
c33870 3633 4451 1.96e-16
c33871 2559 2824 1.58e-16
c33872 1763 1761 1.6e-16
c33873 1196 1656 1.58e-16
c33874 1690 1934 1.58e-16
c33875 439 442 4.6e-16
c33876 433 432 6.4e-16
c33877 5529 584 3.54e-16
c33878 2368 2362 1.6e-16
c33879 1845 2359 2.386e-15
c33880 1851 2367 1.136e-15
c33881 2266 2267 1.6e-16
c33882 2257 2259 2.15e-16
c33883 2644 2635 3.46e-16
c33884 400 0 1.4803e-14
c33885 4872 31 7.84e-16
c33886 4736 33 1.88e-16
c33887 2742 2350 2.38e-15
c33888 1767 647 1.339e-15
c33889 744 1 5.57e-16
c33890 3213 3209 1.96e-16
c33891 1321 1640 3.92e-16
c33892 3208 1 4.41e-15
c33893 1561 1106 4.11e-16
c33894 4625 4626 2.48e-16
c33895 4630 4629 2.83e-16
c33896 4633 4242 1.96e-16
c33897 4181 1 7.71e-16
c33898 4370 0 3.3724e-14
c33899 2475 858 1.75e-16
c33900 1823 1 2.054e-15
c33901 601 1690 3.15e-16
c33902 3502 662 7.38e-16
c33903 4726 1 1.806e-15
c33904 2149 1635 1.477e-15
c33905 747 1488 5.73e-16
c33906 1825 0 8e-16
c33907 3393 3518 1.58e-16
c33908 1029 662 8.3e-16
c33909 9 43 6.48e-16
c33910 13 5 7.76e-16
c33911 4844 4848 1.81e-16
c33912 0 31 1.16477e-13
c33913 5379 1 7.87e-16
c33914 792 2418 3.79e-16
c33915 2194 1828 5.5e-16
c33916 4468 807 2.4e-16
c33917 5540 5539 5.87e-16
c33918 3033 1 2.56e-15
c33919 1251 1262 7.65e-16
c33920 1243 1245 5.5e-16
c33921 919 767 3.15e-16
c33922 920 1098 1.58e-16
c33923 64 122 1.88e-16
c33924 4281 4280 9.1e-16
c33925 4383 732 2.4e-16
c33926 1343 1011 1.58e-16
c33927 3034 1 4.57e-15
c33928 627 1392 1.58e-16
c33929 3900 4523 1.58e-16
c33930 3701 4539 4.78e-16
c33931 2486 852 1.13e-15
c33932 2316 677 1.58e-16
c33933 3989 1 7.71e-16
c33934 4150 25 3.84e-16
c33935 1738 1737 1.6e-16
c33936 4813 4819 7.25e-16
c33937 3046 3190 3.92e-16
c33938 2133 1667 1.383e-15
c33939 2139 1249 2.12e-16
c33940 601 1738 1.58e-16
c33941 4538 1 1.886e-15
c33942 4716 4713 3.01e-16
c33943 2264 1 8.43e-16
c33944 627 2196 3.58e-16
c33945 722 738 1.621e-15
c33946 732 736 2.19e-16
c33947 4563 4242 5.88e-16
c33948 4571 4248 1.58e-16
c33949 2419 2410 3.92e-16
c33950 1902 2413 5.66e-16
c33951 811 809 5.88e-16
c33952 5368 0 1.65e-16
c33953 2630 1 9.28e-16
c33954 1031 1457 1.58e-16
c33955 3200 1 6.15e-16
c33956 3960 1 5.1e-16
c33957 3605 4441 5.66e-16
c33958 4447 4438 3.92e-16
c33959 687 1820 1.58e-16
c33960 3941 19 9.67e-16
c33961 1026 1 4.044e-15
c33962 2841 842 1.58e-16
c33963 1708 1499 5.5e-16
c33964 2756 767 1.58e-16
c33965 1458 0 6.62e-16
c33966 3409 3671 1.58e-16
c33967 2252 2253 9.1e-16
c33968 737 1097 1.58e-16
c33969 890 908 5.51e-16
c33970 907 891 1.486e-15
c33971 64 585 4.6e-16
c33972 3723 842 1.58e-16
c33973 5523 1 3.36e-16
c33974 2511 1998 4.78e-16
c33975 957 1372 1.58e-16
c33976 1221 1223 1.92e-16
c33977 674 1 7.18e-16
c33978 617 3397 3.15e-16
c33979 1522 1905 7.84e-16
c33980 1225 0 8.78e-16
c33981 4528 4525 3.01e-16
c33982 4794 4805 1.96e-16
c33983 2164 2078 1.6e-16
c33984 3387 3106 1.58e-16
c33985 5200 5158 3.41e-16
c33986 4708 468 1.88e-16
c33987 4915 62 1.88e-16
c33988 2403 1 9.28e-16
c33989 2373 0 3.6012e-14
c33990 0 566 1.051e-14
c33991 3531 3140 1.136e-15
c33992 5311 1 3.36e-16
c33993 1500 707 3.64e-16
c33994 601 1357 5.03e-16
c33995 3362 2849 1.477e-15
c33996 3801 410 1.108e-15
c33997 2753 3261 2.48e-16
c33998 3046 3155 1.58e-16
c33999 3030 3143 1.58e-16
c34000 1596 1 2.054e-15
c34001 5198 5219 1.96e-16
c34002 1598 0 8e-16
c34003 4675 0 1.6462e-14
c34004 304 303 5.8e-16
c34005 3796 3773 1.96e-16
c34006 2196 2287 3.92e-16
c34007 566 564 1.58e-16
c34008 3514 717 1.58e-16
c34009 2299 2667 1.96e-16
c34010 5051 149 1.96e-16
c34011 1653 868 2.65e-16
c34012 1181 827 3.15e-16
c34013 1442 1011 1.96e-16
c34014 101 107 3.84e-16
c34015 3924 1 6.78e-16
c34016 911 2196 3.45e-16
c34017 1976 1973 5.5e-16
c34018 632 19 1.676e-15
c34019 77 15 6.58e-16
c34020 49 450 1.88e-16
c34021 369 373 1.372e-15
c34022 204 570 1.88e-16
c34023 3453 3464 1.96e-16
c34024 2312 2310 1.6e-16
c34025 2307 2306 2.03e-16
c34026 3893 3890 2.109e-15
c34027 3693 827 1.832e-15
c34028 384 1 5.62e-16
c34029 4124 3918 2.87e-16
c34030 5588 5575 1.96e-16
c34031 595 3424 1.58e-16
c34032 602 3421 1.832e-15
c34033 2856 2858 1.862e-15
c34034 3898 4285 1.58e-16
c34035 3876 4297 1.58e-16
c34036 2557 2555 1.96e-16
c34037 2541 2554 1.58e-16
c34038 2559 2562 1.6e-16
c34039 612 967 1.58e-16
c34040 601 953 1.822e-15
c34041 654 1 5.57e-16
c34042 617 3882 3.15e-16
c34043 1667 1659 5.95e-16
c34044 1409 0 1.4092e-14
c34045 363 252 1.88e-16
c34046 632 2253 7.38e-16
c34047 3030 662 3.15e-16
c34048 76 75 6.67e-16
c34049 5201 5190 6.73e-16
c34050 5193 5194 2.67e-16
c34051 1981 1953 2.64e-16
c34052 3937 857 1.88e-16
c34053 5538 497 1.58e-16
c34054 3130 0 6.72e-16
c34055 921 827 3.15e-16
c34056 4421 767 1.58e-16
c34057 5476 5481 1.493e-15
c34058 5493 5492 3.92e-16
c34059 383 64 1.88e-16
c34060 4860 827 1.23e-16
c34061 1536 1534 1.6e-16
c34062 1321 1368 3.92e-16
c34063 2446 812 5.03e-16
c34064 4632 1 6.42e-16
c34065 4378 4757 1.58e-16
c34066 2060 2064 1.845e-15
c34067 1566 1 8.43e-16
c34068 3534 3532 1.6e-16
c34069 2149 1 1.886e-15
c34070 5239 0 3.4847e-14
c34071 1670 0 2.7593e-14
c34072 766 764 5.88e-16
c34073 2860 2469 4.11e-16
c34074 2541 2350 5.88e-16
c34075 3117 0 6.916e-14
c34076 1181 812 3.57e-16
c34077 2969 2966 3.92e-16
c34078 2923 2971 1.062e-15
c34079 2541 2717 1.58e-16
c34080 3862 1 1.106e-15
c34081 4060 25 1.88e-16
c34082 2339 737 1.75e-16
c34083 1706 1986 3.92e-16
c34084 3605 1 4.41e-15
c34085 4592 0 3.485e-14
c34086 4676 4675 2.03e-16
c34087 2535 672 3.15e-16
c34088 2559 647 3.15e-16
c34089 219 225 1.372e-15
c34090 205 204 7.03e-16
c34091 4439 0 6.62e-16
c34092 3523 692 1.58e-16
c34093 4944 4980 1.58e-16
c34094 2274 2283 3.92e-16
c34095 890 662 3.15e-16
c34096 3397 3603 1.58e-16
c34097 3714 3712 1.6e-16
c34098 4127 4118 1.96e-16
c34099 4821 468 1.88e-16
c34100 2569 2568 2.48e-16
c34101 2136 1249 4.35e-16
c34102 1806 672 1.58e-16
c34103 3321 3397 5.5e-16
c34104 2535 2299 5.5e-16
c34105 3886 3384 1.58e-16
c34106 2350 732 3.79e-16
c34107 2559 2492 1.58e-16
c34108 1136 1131 1.58e-16
c34109 595 904 2.61e-16
c34110 609 1 5.57e-16
c34111 3163 2645 2.38e-15
c34112 3625 777 1.58e-16
c34113 5018 3744 1.667e-15
c34114 3048 2736 1.58e-16
c34115 3046 2730 5.5e-16
c34116 3034 3257 1.58e-16
c34117 1505 0 3.6368e-14
c34118 3393 3587 1.96e-16
c34119 2184 2183 6.97e-16
c34120 2185 2181 1.71e-16
c34121 15 465 5.8e-16
c34122 1 469 4.92e-16
c34123 4563 4486 1.58e-16
c34124 4861 4862 9.93e-16
c34125 5278 5281 1.075e-15
c34126 461 37 1.88e-16
c34127 4104 857 3.1e-16
c34128 4787 178 7.67e-16
c34129 4793 526 1.88e-16
c34130 911 3401 1.829e-15
c34131 2178 1681 1.58e-16
c34132 921 812 3.15e-16
c34133 101 1 1.073e-15
c34134 4708 64 1.88e-16
c34135 3461 1 6.15e-16
c34136 3626 0 6.62e-16
c34137 2333 717 3.79e-16
c34138 1840 1837 5.5e-16
c34139 4471 3639 2.48e-16
c34140 2679 2674 1.642e-15
c34141 2194 717 3.15e-16
c34142 1769 1386 7.84e-16
c34143 612 921 3.15e-16
c34144 4571 722 1.33e-16
c34145 3329 3331 2.03e-16
c34146 1708 1952 3.92e-16
c34147 1 169 2.87e-16
c34148 117 25 5.71e-16
c34149 233 247 1.88e-16
c34150 4582 4707 3.92e-16
c34151 0 184 2.87e-16
c34152 2082 1 2.224e-15
c34153 3608 752 1.832e-15
c34154 3822 3775 3.18e-16
c34155 3806 3820 2.102e-15
c34156 5209 1 1.257e-15
c34157 632 2611 3.15e-16
c34158 2182 1681 1.58e-16
c34159 986 662 1.58e-16
c34160 5173 0 3.5057e-14
c34161 2654 1 5.808e-15
c34162 3722 3710 2.32e-16
c34163 632 1406 1.832e-15
c34164 1161 1168 7.95e-16
c34165 3886 4387 1.58e-16
c34166 3876 3548 5.5e-16
c34167 4606 5514 1.96e-16
c34168 2798 2804 1.418e-15
c34169 3254 762 2.65e-16
c34170 968 0 1.4198e-14
c34171 3021 3019 3.54e-16
c34172 1206 1664 8.31e-16
c34173 1706 1951 1.58e-16
c34174 1690 1939 1.58e-16
c34175 1946 1937 3.46e-16
c34176 565 368 1.88e-16
c34177 3530 3134 1.96e-16
c34178 5031 5047 2.109e-15
c34179 3304 3299 1.642e-15
c34180 595 1678 1.655e-15
c34181 602 2215 3.64e-16
c34182 175 570 1.88e-16
c34183 5200 207 7.37e-16
c34184 2664 1 9.28e-16
c34185 907 992 3.92e-16
c34186 273 1 4.59e-16
c34187 2819 2435 1.58e-16
c34188 3293 3676 7.84e-16
c34189 1784 672 1.58e-16
c34190 1404 1406 1.862e-15
c34191 2194 2371 1.58e-16
c34192 3247 762 2.72e-16
c34193 3548 3520 2.64e-16
c34194 1817 707 1.75e-16
c34195 642 1363 1.58e-16
c34196 1331 1487 4.63e-16
c34197 1694 1363 5.5e-16
c34198 596 1 1.2643e-14
c34199 3787 1 3.36e-16
c34200 2691 707 1.84e-16
c34201 617 1690 3.15e-16
c34202 4919 4916 3.92e-16
c34203 2719 737 2.33e-16
c34204 747 1897 2.65e-16
c34205 1841 0 6.72e-16
c34206 229 37 1.88e-16
c34207 236 30 3.84e-16
c34208 3393 3523 1.58e-16
c34209 3409 3140 1.58e-16
c34210 2746 2350 1.96e-16
c34211 837 835 3.327e-15
c34212 2266 1 1.868e-15
c34213 3781 3785 1.583e-15
c34214 4054 857 1.88e-16
c34215 2424 2425 1.35e-16
c34216 2172 1845 5.5e-16
c34217 1517 732 2.65e-16
c34218 129 15 5.8e-16
c34219 1173 1174 1.21e-16
c34220 146 19 3.84e-16
c34221 4287 4283 1.96e-16
c34222 2722 2720 1.862e-15
c34223 1321 1026 1.58e-16
c34224 3398 1 3.009e-15
c34225 3034 2634 1.58e-16
c34226 3707 3882 1.58e-16
c34227 2172 677 4.48e-16
c34228 3024 3207 3.92e-16
c34229 629 628 1.6e-16
c34230 627 1752 1.58e-16
c34231 617 1738 1.84e-16
c34232 2006 2007 2.48e-16
c34233 762 1331 7.99e-16
c34234 898 901 7.46e-16
c34235 19 313 8.82e-16
c34236 37 291 1.88e-16
c34237 4563 4259 5.88e-16
c34238 4571 4265 1.58e-16
c34239 5162 5154 3.54e-16
c34240 1913 2410 1.58e-16
c34241 894 767 3.15e-16
c34242 890 1098 3.54e-16
c34243 909 1119 1.58e-16
c34244 919 931 1.58e-16
c34245 4600 1 9.556e-15
c34246 2237 2265 2.64e-16
c34247 1031 1477 2.38e-15
c34248 2402 767 7.68e-16
c34249 1684 1369 1.58e-16
c34250 1734 1319 4.97e-16
c34251 4820 4811 3.46e-16
c34252 1483 1 1.868e-15
c34253 4539 1 4.03e-16
c34254 2861 842 1.58e-16
c34255 2300 1783 1.96e-16
c34256 822 1146 5.73e-16
c34257 1473 0 2.93e-15
c34258 187 190 2.142e-15
c34259 3106 3492 5.66e-16
c34260 3498 3489 3.92e-16
c34261 3898 762 3.15e-16
c34262 5010 4902 1.58e-16
c34263 642 3105 2.4e-16
c34264 3409 3676 1.58e-16
c34265 14 15 4.88e-16
c34266 5253 5239 1.96e-16
c34267 5229 5200 1.58e-16
c34268 4736 526 1.88e-16
c34269 2194 1987 1.58e-16
c34270 1392 957 2.38e-15
c34271 4821 64 1.88e-16
c34272 3193 3195 2.03e-16
c34273 1345 1593 1.58e-16
c34274 1533 1888 1.58e-16
c34275 450 194 1.88e-16
c34276 3472 647 1.58e-16
c34277 4874 1 8.85e-16
c34278 3298 797 1.9e-16
c34279 88 484 1.88e-16
c34280 3253 3641 4.97e-16
c34281 3393 837 4.03e-16
c34282 5320 1 2.53e-16
c34283 1061 692 3.57e-16
c34284 1260 1246 6.67e-16
c34285 72 9 6.48e-16
c34286 5422 5412 1.58e-16
c34287 74 0 1.051e-14
c34288 1556 782 2.33e-16
c34289 1101 1542 7.84e-16
c34290 1073 1 4.59e-16
c34291 4149 1 7.71e-16
c34292 3886 3667 5.5e-16
c34293 1810 1801 3.46e-16
c34294 4140 26 4.58e-16
c34295 4132 0 2.0391e-14
c34296 4862 4486 3.92e-16
c34297 4874 4873 1.6e-16
c34298 1070 0 1.0077e-14
c34299 3100 2583 1.136e-15
c34300 2036 2100 2.249e-15
c34301 2104 2115 1.96e-16
c34302 1614 0 6.72e-16
c34303 4692 0 1.6462e-14
c34304 911 2531 1.88e-16
c34305 792 1136 3.79e-16
c34306 0 326 1.4515e-14
c34307 19 320 3.84e-16
c34308 3387 647 4.48e-16
c34309 3344 3397 1.58e-16
c34310 4370 707 1.832e-15
c34311 5414 5404 9.99e-16
c34312 5303 5299 1.866e-15
c34313 1163 797 3.57e-16
c34314 1143 1156 1.58e-16
c34315 3873 3871 3.54e-16
c34316 3719 3708 1.96e-16
c34317 4152 4143 3.84e-16
c34318 4156 4157 6.67e-16
c34319 5323 5325 9.16e-16
c34320 1839 692 1.9e-16
c34321 1644 858 1.58e-16
c34322 1196 868 3.79e-16
c34323 3882 4485 1.96e-16
c34324 2982 2873 6.31e-16
c34325 4514 5580 5.69e-16
c34326 2557 2769 3.92e-16
c34327 3839 3806 1.58e-16
c34328 4118 25 3.84e-16
c34329 4423 3588 1.96e-16
c34330 4428 3582 1.96e-16
c34331 535 549 3.84e-16
c34332 4905 4969 1.6e-16
c34333 1811 2304 1.96e-16
c34334 1966 1 9.28e-16
c34335 2759 0 1.4092e-14
c34336 1072 1074 7.84e-16
c34337 4523 852 1.58e-16
c34338 4634 5457 5.91e-16
c34339 601 3421 1.58e-16
c34340 920 1219 1.58e-16
c34341 2541 2169 1.58e-16
c34342 2016 842 3.64e-16
c34343 1613 1610 5.5e-16
c34344 627 967 1.58e-16
c34345 3090 3101 1.96e-16
c34346 4308 1 6.15e-16
c34347 1886 1499 1.532e-15
c34348 1892 1891 5.65e-16
c34349 5000 4999 1.6e-16
c34350 3034 3326 4.63e-16
c34351 747 921 3.15e-16
c34352 5010 323 1.88e-16
c34353 1769 0 3.3691e-14
c34354 448 462 3.84e-16
c34355 4567 4757 1.58e-16
c34356 4580 4361 5.5e-16
c34357 4582 4367 1.58e-16
c34358 3397 3072 1.58e-16
c34359 880 1358 5.66e-16
c34360 1470 702 2.4e-16
c34361 920 852 3.15e-16
c34362 1041 1048 7.95e-16
c34363 3497 4314 1.58e-16
c34364 4441 767 1.58e-16
c34365 5515 381 3.54e-16
c34366 2545 2356 1.58e-16
c34367 1345 1385 3.92e-16
c34368 642 3886 7.99e-16
c34369 4517 4515 1.6e-16
c34370 2640 647 1.58e-16
c34371 2637 672 1.58e-16
c34372 2466 812 1.09e-16
c34373 1801 1414 1.532e-15
c34374 3030 2781 5.88e-16
c34375 4649 1 6.42e-16
c34376 4395 4757 1.58e-16
c34377 4384 4765 5.66e-16
c34378 4771 4762 3.92e-16
c34379 3409 3433 1.58e-16
c34380 2078 2029 2.634e-15
c34381 2036 2033 1.96e-16
c34382 1635 2019 1.58e-16
c34383 1845 0 6.9481e-14
c34384 3723 3411 3.92e-16
c34385 4571 4561 1.152e-15
c34386 4567 4197 1.58e-16
c34387 5165 236 3.94e-16
c34388 5111 5072 3.18e-16
c34389 4334 692 1.339e-15
c34390 5262 5177 8.28e-16
c34391 2557 2367 5.5e-16
c34392 1152 782 4.98e-16
c34393 957 931 6.54e-16
c34394 1181 1179 1.931e-15
c34395 3882 4450 1.58e-16
c34396 3014 2929 3.96e-16
c34397 677 0 2.80577e-13
c34398 2787 0 3.5142e-14
c34399 2557 2734 1.58e-16
c34400 2541 2722 1.58e-16
c34401 687 1414 1.58e-16
c34402 1249 1254 3.01e-16
c34403 1684 2003 3.92e-16
c34404 4609 0 3.4781e-14
c34405 1966 1965 1.6e-16
c34406 1958 1956 2.15e-16
c34407 1743 1738 1.642e-15
c34408 3140 3522 2.48e-16
c34409 5034 5095 1.6e-16
c34410 3443 3440 3.01e-16
c34411 3439 3436 6.44e-16
c34412 436 570 1.88e-16
c34413 3543 692 1.58e-16
c34414 5170 265 1.96e-16
c34415 762 1706 3.15e-16
c34416 3384 3383 3.54e-16
c34417 3281 0 3.466e-15
c34418 3118 1 1.868e-15
c34419 602 3046 4.46e-16
c34420 595 3024 1.511e-15
c34421 2559 2316 5.5e-16
c34422 1372 1 5.808e-15
c34423 1374 0 3.466e-15
c34424 2722 732 1.58e-16
c34425 2272 2283 1.96e-16
c34426 3024 2747 5.5e-16
c34427 3034 3262 1.58e-16
c34428 4563 4503 1.58e-16
c34429 2573 2571 1.6e-16
c34430 596 770 5.28e-16
c34431 4855 352 1.88e-16
c34432 2194 2405 1.58e-16
c34433 2178 2393 1.58e-16
c34434 4674 5484 1.344e-15
c34435 2194 1715 1.58e-16
c34436 4300 4311 1.96e-16
c34437 3470 1 1.716e-15
c34438 1507 1061 4.97e-16
c34439 1345 1349 1.6e-16
c34440 4055 1 4.45e-16
c34441 1781 1397 1.58e-16
c34442 1128 0 4.6547e-14
c34443 627 921 3.15e-16
c34444 1315 1 5.329e-15
c34445 653 652 1.96e-16
c34446 3237 2719 1.96e-16
c34447 3238 3231 6.73e-16
c34448 3169 677 3.64e-16
c34449 2535 797 4.48e-16
c34450 1800 1 4.41e-15
c34451 2044 2056 1.96e-16
c34452 822 2452 3.79e-16
c34453 2182 2393 1.58e-16
c34454 2375 2377 2.03e-16
c34455 2309 0 6.62e-16
c34456 1202 868 2.68e-16
c34457 890 1172 1.96e-16
c34458 2674 1 2.054e-15
c34459 921 993 1.58e-16
c34460 287 288 6.4e-16
c34461 1331 1329 5.93e-16
c34462 1767 1386 3.92e-16
c34463 1771 1772 1.6e-16
c34464 602 907 5.2e-16
c34465 595 883 5.02e-16
VsrcMul2 15 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
VldMulA 3918 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
VldMulB 596 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
VPhi1H 26 0 pwl (0 0 4e-09 0 6e-09 3 2.2e-08 3 
+ 2.4e-08 0 4e-08 0 4.4e-08 0 4.6e-08 3 
+ 6.2e-08 3 6.4e-08 0 8e-08 0 8.4e-08 0 
+ 8.6e-08 3 1.02e-07 3 1.04e-07 0 1.2e-07 0 
+ 1.24e-07 0 1.26e-07 3 1.42e-07 3 1.44e-07 0 
+ 1.6e-07 0 1.64e-07 0 1.66e-07 3 1.82e-07 3 
+ 1.84e-07 0 2e-07 0 2.04e-07 0 2.06e-07 3 
+ 2.22e-07 3 2.24e-07 0 2.4e-07 0 2.44e-07 0 
+ 2.46e-07 3 2.62e-07 3 2.64e-07 0 2.8e-07 0 
+ 2.84e-07 0 2.86e-07 3 3.02e-07 3 3.04e-07 0 
+ 3.2e-07 0 3.24e-07 0 3.26e-07 3 3.42e-07 3 
+ 3.44e-07 0 3.6e-07 0 3.64e-07 0 3.66e-07 3 
+ 3.82e-07 3 3.84e-07 0 4e-07 0 4.04e-07 0 
+ )
VPhi2H 19 0 pwl (0 0 2.6e-08 0 2.8e-08 3 4e-08 3 
+ 4.2e-08 0 6.6e-08 0 6.8e-08 3 8e-08 3 
+ 8.2e-08 0 1.06e-07 0 1.08e-07 3 1.2e-07 3 
+ 1.22e-07 0 1.46e-07 0 1.48e-07 3 1.6e-07 3 
+ 1.62e-07 0 1.86e-07 0 1.88e-07 3 2e-07 3 
+ 2.02e-07 0 2.26e-07 0 2.28e-07 3 2.4e-07 3 
+ 2.42e-07 0 2.66e-07 0 2.68e-07 3 2.8e-07 3 
+ 2.82e-07 0 3.06e-07 0 3.08e-07 3 3.2e-07 3 
+ 3.22e-07 0 3.46e-07 0 3.48e-07 3 3.6e-07 3 
+ 3.62e-07 0 3.86e-07 0 3.88e-07 3 4e-07 3 
+ 4.02e-07 0 4.26e-07 0 )
Vnbus.1 3969 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.2 3952 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.3 3938 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.4 3920 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.5 4001 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.6 3984 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.7 4033 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.8 4016 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.9 4065 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.10 4048 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.11 4097 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.12 4080 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.13 4129 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.14 4112 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.15 4161 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.16 4144 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.17 4193 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.18 4176 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.19 4228 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vnbus.20 4209 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.1 848 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.2 864 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.3 833 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.4 818 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.5 803 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.6 788 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.7 773 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.8 758 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.9 743 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.10 728 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.11 713 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.12 698 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.13 683 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.14 668 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.15 653 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.16 638 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.17 623 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.18 608 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 1.6e-07 0 
+ 1.62e-07 3 2e-07 3 2.02e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.19 590 0 pwl (0 3 4e-08 3 4.2e-08 0 8e-08 0 
+ 8.2e-08 3 1.2e-07 3 1.22e-07 0 2.4e-07 0 
+ 2.42e-07 3 2.8e-07 3 2.82e-07 0 3.2e-07 0 
+ 3.22e-07 3 3.6e-07 3 3.62e-07 0 4e-07 0 
+ 4.02e-07 3 4.4e-07 3 )
Vrbus.20 934 0 pwl (0 0 8e-08 0 8.2e-08 3 1.2e-07 3 
+ 1.22e-07 0 1.6e-07 0 1.62e-07 3 2e-07 3 
+ 2.02e-07 0 3.2e-07 0 4e-07 0 4.02e-07 3 
+ )
VPhi1#test 25 0 pwl (0 0 4e-06 0 )
VsrcMul1 9 0 pwl (0 0 4e-06 0 )
Vreset 37 0 pwl (0 0 4e-06 0 )
VShfAmt 30 0 pwl (0 3 4e-06 3 )
VVdd 1 0 3 
.options device temp=55 
.print TRAN v(26) v(19) v(596) v(584) v(556) v(528) 
+v(499) v(470) v(441) v(412) v(383) v(354) 
+v(325) v(296) v(267) v(238) v(209) v(180) 
+v(151) v(122) v(93) v(64) v(33) v(526) 
+v(497) v(468) v(439) v(410) v(381) v(352) 
+v(323) v(294) v(265) v(236) v(207) v(178) 
+v(149) v(120) v(91) v(62) v(31) 
*.options limpts=50000 itl5=50000
.TRAN 1e-09 4e-07
.end
