vdmos test circuit
vd 3 0 0
vs 2 0 0
vg 4 0 dc 5
vid 3 5 dc 0

.param dtempParam=10
m1 5 4 2 0 irf130 w=0.386 l=2.5u dtemp={dtempParam}
.model irf130 nmos level=18
+ cv=1
+ cve=1
+ vto=3.5
+ rd= 0
+ rs= 0.005
+ lambda=0
+ m=3
+ sigma0=0
+ uo=230
+ vmax=4e4
+ delta=5
+ tox=50nm

.options device temp=15
*
.dc vd 0 50 5 vg 5 15 5
.print dc v(3) v(4) v(2) i(vid)

.step dtempParam list 0 10 20

.end

