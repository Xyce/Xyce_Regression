level=1 diode circuit with .rol statement 
*
R 1 2 0.0001
V2 2 0 0.21
V1 3 0 0.0
D2 1 3 DA lambertw=1

.MODEL DA D (IS=1.0e-09 RS=6.5e-05 N=1.0)

.SENS objfunc={I(V1)} param=DA:IS,DA:RS
.options SENSITIVITY DAKOTAFILE=0  adjoint=0 direct=1  STDOUTPUT=0
.options topology OUTPUTNAMESFILE=true
.DC V2 0.005 0.5 0.005
.print DC v(2) I(V1)  

.rol

.END

