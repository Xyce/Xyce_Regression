*****************************************************
* Test FORMAT=SPLOT without .STEP.  This should
* produce the same .prn file as FORMAT=STD.
*
* This test also ensures that FORMAT=SPLOT produces
* a file with a .prn extension.  It is sufficient to
* just test this for .PRINT TRAN
*****************************************************

V1 1 0 SIN(0 1 1)
R1 1 2 1
R2 2 0 1

.OPTIONS OUTPUT INITIAL_INTERVAL=0.01
.PRINT TRAN FORMAT=SPLOT R1:R R2:R V(1) V(2)
.TRAN 0 1

.END
