Netlist to Test Xygra
YXYGRA R1 1 0  6 0 7 0
+ COIL = { NAME       = FOO  ,BAR,BAZ
+          NUMWINDINGS=1 ,1 ,1   }
v1 1a 0 0
v2 6a 0 0
v3 7a 0 0
r1 1 1a 1
r2 6 6a 1
r3 7 7a 1
*.DC V1 0 5V 1V
.tran 1us 1s
*.PRINT DC V(1) I(V1)
.PRINT tran I(V1)  I(V2)  I(V3)
*comp I(V1) RELTOL=0.02 ABSTOL=1e-6
*comp I(V2) RELTOL=0.02 ABSTOL=1e-6
*comp I(V3) RELTOL=0.02 ABSTOL=1e-6
.model foobar xygra ()
.END
