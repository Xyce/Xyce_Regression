* A test of the measure TRIG and TARG functionality, using the legacy
* TRIG-TARG mode.  So, it tests the RiseFallDelay class.
* See gitlab-ex issue 303 for more details.
*
* These tests cover the following "special" syntaxes, per SON Bug 679.
* These syntaxes are difficult to auto-parse with the tools in MeasureCommon.pm
*
*   TRIG AT=<time>
*   TRIG v(a)=v(b)
*   TARG v(c)=v(d)
*******************************************************************************
*
* a few sources of different types
VS  1  0  SIN(0 1.0 1KHZ 0 0)
VP  2  0  PULSE(-2 3 0.2ms 0.5ms 0.5ms 1ms 2ms )
VDC 3  0  0.7

R1  1  0  100
R2  2  0  100
R3  3  0  100

* use legacy trig-targ mode
.OPTIONS MEASURE USE_LTTM=1

.TRAN 0 3ms 0 0.01ms

.PRINT TRAN FORMAT=NOINDEX V(1) V(2) V(3)

.measure tran m1 TRIG V(1)=0.5  TARG V(2)=0.5
.measure tran m2 TRIG V(1)=v(3) TARG V(2)=0.5
.measure tran m3 TRIG V(1)=0.5  TARG V(2)=V(3)
.measure tran m4 TRIG V(1)=V(3) TARG V(2)=V(3)
.measure tran m5 TRIG AT=1e-3   TARG V(2)=0.5
.measure tran m6 TRIG AT=1e-3   TARG V(2)=V(3)

.END

