Test of .IC with .STEP.  

.ic v(1)=1.0

c1 1 0 1.0e-6
R1 1 2 1K
v1 2 0 0V

.print tran v(1)
.tran 0 5ms
.options timeint reltol=1e-6 abstol=1e-6
.end

