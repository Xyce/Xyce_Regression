Netlist to Test the bsrc with multipliers, subcircuit implicit multiplier, nested subckt baseline
******************************************************************************
VIN 1 0 DC 12V
G 3 0 2 0 0.2
R1 1 2 300
R2 2 0 900
R3 3 0 200
R4 3 0 200
.DC VIN 1 12 1
.PRINT DC V(1) V(2) V(3) 
.END
