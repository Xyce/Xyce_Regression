Resistor sensitivity test.
*
R1 VA B 10.0
R2 B 0 10.0
VA VA 0 5

.dc VA 5 5 1
.print dc v(VA) v(B) I(VA) {2*I(VA)}

.SENS objfunc={I(VA)} param=R1:R,R2:R
.options SENSITIVITY direct=1 adjoint=0  diagnosticfile=1 
.print sens 

.END

