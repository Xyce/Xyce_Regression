R1 1 0 1
R2 1 0 1
R3 1 0 1
R4 1 0 1
R5 1 0 1
R6 1 0 1
v1 1 0 PWL (0 0 1 1)

*.PRINT TRAN V(1) 
.tran 1u 

.end
