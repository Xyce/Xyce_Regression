Netlist to Test the KLU solver
*COMP V(2) OFFSET=-1
I1 1 0 PULSE(0 5V 0 1MS 1MS 10MS 25MS)
L1 2 0 10mH
R1 1 2 0.001
.TRAN 0.1MS 2MS 0MS
.PRINT TRAN V(1) V(2)
.OPTIONS LINSOL TYPE=klu
.END
