Lead current test for switches
*
v1  1  0        PWL(0 0 1U 0 1.01U 5 2U 5 2.01U 0 3U 0 3.01U 5)
S1  2  1  3  0  VSW
S2  0  2  3  0  ISW
v3  0  3        PWL (0 0 2U 0 2.01U 5)
r3  0  3        200
.MODEL VSW VSWITCH(RON=1 ROFF=1MEG VON=1 VOFF=0)
.MODEL ISW ISWITCH (ION=10mA IOFF=0mA RON=1 ROFF=1E6)
.options timeint method=gear
.options nonlin-tran rhstol=1.0e-7
.TRAN 0.02U 4U
*COMP {I(S1)-I(V1)} abstol=1.0e-6 zerotol=1.0e-7
*COMP {I(S2)-I(V1)} abstol=1.0e-6 zerotol=1.0e-7
.PRINT TRAN V(1) V(3) {I(S1)-I(V1)} {I(S2)-I(V1)}

.measure tran maxmag1   max {abs(I(S1)-I(V1))} failvalue=1e-6
.measure tran totalrms1 rms {I(S1)-I(V1)} failvalue=1e-6 
.measure tran maxmag2   max {abs(I(S2)-I(V1))} failvalue=1e-6
.measure tran totalrms2 rms {I(S2)-I(V1)} failvalue=1e-6 

.END
