*Test of dependent parameter handling in mutual inductors

* Because the mutual inductor device was not properly updating its internal
* copies of the coupled inductance list in processParams, using .step on
* any global param that was used in L value expressions would not actually
* cause the simulation to change behavior, even after bug 28's fix of
* global parameter handling during context resolution for MIs.

* This test case .steps a scale factor that is being applied to the inductors
* coupled by the K device, which in this test is a nonlinear-core MI.

* This netlist is one of 3 individual, non-stepped runs that will be
* performed by the test script, and compared to the main .stepped netlist.


.subckt transformer node1 node6
Llead4 node1 0 10
Llead5 node5 node6 50
Llead6 node6 node7 50
Ktrans2 Llead4 Llead5 Llead6 1.0 nlcore

.model nlcore CORE c=0.001

rload3  node5 0 100
rpathtg2 node7 0 1
.ends

Vinput node1 0 sin(0 14 120 0 0)
X1 node1 node6 transformer
rload4  node6 0 100

.tran 0 10m
.print tran v(node1) v(node6)
.options output PRINTFOOTER=false
.end

