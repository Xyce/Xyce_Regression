
.param foobar=1000

R1 1 0 {foobar}
V1 1 0 1

.dc v1 1 1 1
.print DC V(1) I(V1) R1:R
.end
