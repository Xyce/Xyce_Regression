*******************************************************************************
* This netlist is equivalent to Step 1 for the RMSTest.cir netlist.
* It has VS1:VA=2 and VS3:V0=-0.25
*
*******************************************************************************
*
* a few sources of different types
VS1  1  0  SIN(0 2 100Hz 0 0)
VP  2  0  PULSE( 0 100 0.2ms 0.2ms 0.2ms 1ms 2ms )
VS3  3  0  SIN(-0.25 1.0 100HZ 0 0.5)
VS4  4  0  SIN(0.5 -1.0 100HZ 0 0.5)

R1  1  0  100
R2  2  0  100
R3  3  0  100
R4  4  0  100

.TRAN 0  30ms
.PRINT TRAN FORMAT=NOINDEX V(1) V(2) V(3) V(4)

.measure tran rmsAll RMS v(1)
.measure tran rmsTop rms v(2)

* add TO-FROM modifiers
.measure tran sineHalfInterval Rms V(1) from=0 to=0.015

* mix in TDs before and after FROM value.
.measure tran sineTDbetween rms V(1) FROM=0 TO=0.05 TD=0.01
.measure tran sineTDbefore rms V(1) FROM=0.02 TO=0.05 TD=0.01

* these tests should return -1 and -100
.measure tran returnNegOne rms V(1) FROM=0.2e-3 TO=0.25e-3 TD=0.5e-3

.measure tran returnNeg100 rms V(1) FROM=0.2e-3 TO=0.25e-3 TD=0.5e-3 default_val=-100

* add tests for rise/fall/cross.  VS3 and VS4 have a DC offset
* and are damped sinusoids
.measure tran rmsv3fall2 rms v(3) fall=2
.measure tran rmsv4rise1 rms v(4) rise=1
.measure tran rmsv3cross2 rms v(3) cross=2

* test LAST for rise/fall/cross
.measure tran rmsv3falllast rms v(3) fall=last
.measure tran rmsv4riselast rms v(4) rise=last
.measure tran rmsv3crosslast rms v(3) cross=last
.measure tran rmsv4crosslast rms v(4) cross=last

* test RFC_LEVEL keyword
.measure tran rmsv1Rise1RFClevel50 rms V(1) RFC_LEVEL=0.5 RISE=1
.measure tran rmsv1Fall1RFClevel50 rms V(1) RFC_LEVEL=0.5 FALL=1
.measure tran rmsv1Cross1RFClevel50 rms V(1) RFC_LEVEL=0.5 CROSS=1 

*test Failed measures for rise/fall/cross
.measure tran rmsv3fallfail rms v(3) fall=100
.measure tran rmsv4risefail rms v(4) rise=100
.measure tran rmsv3crossfail rms v(3) cross=100

.END

