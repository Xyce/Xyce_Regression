* PMOS Id-Vg with Vb

.include modelcard.pmos

vg 1 0 -1.2
vd 2 0 -0.1
vb 3 0  0.0

m1 2 1 0 3 p1 W=10.0u L=0.09u

.dc vg 0.6 -1.18 -0.02 vb 0 1.2 0.3
.print dc v(1) v(3) i(vd)

.end

