Netlist to test homtopy output and .op
*********************************************************************** 
R1 1 0 1K 
V1 1 0 5V

.options nonlin continuation=1
.options loca conparam=R1
+ initialvalue=500.0 minvalue=-1.0 maxvalue=1500.0
+ initialstepsize=500.0 minstepsize=1.0e-4 maxstepsize=500.0
+ aggressiveness=1.0

.op
.print homotopy V(1) I(V1)
.print dc V(1) I(V1)

.END
