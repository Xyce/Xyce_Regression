*Id-Vd Characteristics for NMOS 

.include "pmos_b3soi.mod"

* --- Voltage Sources ---
vd drain  0 dc 0
vg gate  0 dc 1
vs source 0 dc 0
ve substrate 0 0
 
* --- Transistor ---
.param dtempParam=10
m1 drain gate source substrate  pmos1 W=1e-5 L=1e-6 

* --- DC Analysis ---
.dc vd 0 -1.2 -0.02
.step lin vg -0.4 -1.2 -0.1
.options device temp=25

.step TEMP list 15 25 35

.print dc v(drain) v(gate) i(vd)
.end
