Analog digitizer to test lookup tables in CHILESPICE
* digcs04.cir:  Analog digitizer to test lookup tables in CHILESPICE.  (KDM)  12/15/00
*****************************************************************************
* Tier No.:     1
* Description:  Test of Chilespice code enhancements:
*
*               Lookup Tables
*
* Input/Output: Measure V(3) a common simulation data output (.csd) file can
*               be generated for viewing the signal using PROBE
*****************************************************************************
*.tran 50ns 1ms 0 50ns 
.tran 50ns 10us 
*COMP V(3) reltol=0.02 abstol=1e-6
.print tran PRECISION=10 WIDTH=19 v(3)
*.options acct
*.options nonlin searchmethod=0 strategy=0 in_forcing=0 abstol=1.0e-3 reltol=1.0e-2 rhstol=1.0e-2

Vi    1 0 DC 0  SIN(0 20 1k 0 0 0)
R1    1 0  1k  
Vdig  2 0  PULSE(0 1 0 0.5us 0.5us 2us 10us)
Rdig  2 0  1Meg  
*X_DM1 1 0 3 0 2 Dig_01
RL    3 0  1Meg  


*************************************************************************
*
* Behavioral digitizer (from Temp_sensor_02).  12/15/00
*
*************************************************************************

*.subckt Dig_01 1 2 3 4 Dig

* Input in volts, output digitized.

Rin  1 0  1Meg

BE_Dig 3 0 V = {TABLE { V(2) * (V(1) + 30) / 60 }
*E_Dig 3 0 TABLE V(2)*(V(1)+30)/60 =
+ (0.0000000, 0)
+ (0.0312500, 0)
+ (0.0312813, 1)
+ (0.0625000, 1)
+ (0.0625313, 2)
+ (0.0937500, 2)
+ (0.0937813, 3)
+ (0.1250000, 3)
+ (0.1250313, 4)
+ (0.1562500, 4)
+ (0.1562813, 5)
+ (0.1875000, 5)
+ (0.1875313, 6)
+ (0.2187500, 6)
+ (0.2187813, 7)
+ (0.2500000, 7)
+ (0.2500313, 8)
+ (0.2812500, 8)
+ (0.2812813, 9)
+ (0.3125000, 9)
+ (0.3125313, 10)
+ (0.3437500, 10)
+ (0.3437813, 11)
+ (0.3750000, 11)
+ (0.3750313, 12)
+ (0.4062500, 12)
+ (0.4062813, 13)
+ (0.4375000, 13)
+ (0.4375313, 14)
+ (0.4687500, 14)
+ (0.4687813, 15)
+ (0.5000000, 15)
+ (0.5000313, 16)
+ (0.5312500, 16)
+ (0.5312813, 17)
+ (0.5625000, 17)
+ (0.5625313, 18)
+ (0.5937500, 18)
+ (0.5937813, 19)
+ (0.6250000, 19)
+ (0.6250313, 20)
+ (0.6562500, 20)
+ (0.6562813, 21)
+ (0.6875000, 21)
+ (0.6875313, 22)
+ (0.7187500, 22)
+ (0.7187813, 23)
+ (0.7500000, 23)
+ (0.7500313, 24)
+ (0.7812500, 24)
+ (0.7812813, 25)
+ (0.8125000, 25)
+ (0.8125313, 26)
+ (0.8437500, 26)
+ (0.8437813, 27)
+ (0.8750000, 27)
+ (0.8750313, 28)
+ (0.9062500, 28)
+ (0.9062813, 29)
+ (0.9375000, 29)
+ (0.9375313, 30)
+ (0.9687500, 30)
+ (0.9687813, 31)
+ (1.0000000, 31) }
*+ (1.0000000, 31)

*.ends


.END
