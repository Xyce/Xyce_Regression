branched cable simulation - rallpack 2 - level1 neuron


.tran 0 0.25  
.options output initial_interval=5.0e-5
.options linsol type=klu

* rallpack 2 calls for a steady current input.  But we need to use PULSE so
* that the current will be off during dcop calculation
Iin 0 n0 PULSE( 0 1.0e-10 1.0e-12 0.0 0.0 1.0e10 1.0e10)

* membrane properties (from rallpack2 README file)
* Ra = 1.0 ohms meter
* Rm = 4.0 ohms meter^2
* Cm = 0.01 F/m^2
* Em = -0.065 Volts
* confirmed that these are the same parameter values as for rallpack1

* axial resistance 1 ohms m
.param Ra = 1.0	; [ohm m]

* specific membrane capacitance 0.01 F/m^2 
.param memC = { 0.01 } ; [F/m^2]

* leak current has membrane resistivity of 4 ohms m^2, with reversal potential of -65mV
.param rm = { 4.0 }    ; [ohm m^2]
.param memG = { 1 / rm }                  ; [1/(ohm m^2)]
.param revE = -0.065                      ; [V]

* neuron model - for level 1 neuron, have to specify actual capacitance and resistances, 
* which depend on surface area - and surface area is different at each level
  
.param SA0 = 1.6085e-09
.model level0Params neuron level=1 cMem={memC*SA0}  gMem={memG*SA0} eLeak={revE} gNa=0.0 gK=0.0 vRest={revE}
.param SA1 = 8.04348e-10
.model level1Params neuron level=1 cMem={memC*SA1}  gMem={memG*SA1} eLeak={revE} gNa=0.0 gK=0.0 vRest={revE}
.param SA2 = 4.02174e-10
.model level2Params neuron level=1 cMem={memC*SA2}  gMem={memG*SA2} eLeak={revE} gNa=0.0 gK=0.0 vRest={revE}
.param SA3 = 2.01062e-10
.model level3Params neuron level=1 cMem={memC*SA3}  gMem={memG*SA3} eLeak={revE} gNa=0.0 gK=0.0 vRest={revE}
.param SA4 = 1.00544e-10
.model level4Params neuron level=1 cMem={memC*SA4}  gMem={memG*SA4} eLeak={revE} gNa=0.0 gK=0.0 vRest={revE}
.param SA5 = 5.02559e-11
.model level5Params neuron level=1 cMem={memC*SA5}  gMem={memG*SA5} eLeak={revE} gNa=0.0 gK=0.0 vRest={revE}
.param SA6 = 2.51327e-11
.model level6Params neuron level=1 cMem={memC*SA6}  gMem={memG*SA6} eLeak={revE} gNa=0.0 gK=0.0 vRest={revE}
.param SA7 = 1.25679e-11
.model level7Params neuron level=1 cMem={memC*SA7}  gMem={memG*SA7} eLeak={revE} gNa=0.0 gK=0.0 vRest={revE}
.param SA8 = 6.28595e-12
.model level8Params neuron level=1 cMem={memC*SA8}  gMem={memG*SA8} eLeak={revE} gNa=0.0 gK=0.0 vRest={revE}
.param SA9 = 3.14159e-12
.model level9Params neuron level=1 cMem={memC*SA9}  gMem={memG*SA9} eLeak={revE} gNa=0.0 gK=0.0 vRest={revE}

.param level0R = {Ra*3.2e-05/(2*3.14159*6.4e-11)}
.param level1R = {Ra*2.54e-05/(2*3.14159*2.54016e-11)}
.param level2R = {Ra*2.016e-05/(2*3.14159*1.00806e-11)}
.param level3R = {Ra*1.6e-05/(2*3.14159*4e-12)}
.param level4R = {Ra*1.27e-05/(2*3.14159*1.5876e-12)}
.param level5R = {Ra*1.008e-05/(2*3.14159*6.29642e-13)}
.param level6R = {Ra*8e-06/(2*3.14159*2.5e-13)}
.param level7R = {Ra*6.35e-06/(2*3.14159*9.9225e-14)}
.param level8R = {Ra*5.04e-06/(2*3.14159*3.94023e-14)}
.param level9R = {Ra*4e-06/(2*3.14159*1.5625e-14)}

R001 n0 n00mid {level0R}
yneuron neuron00 n00mid 0 level0Params 
R002 n00mid n00 {level0R}
R0001 n00 n000mid {level1R}
yneuron neuron000 n000mid 0 level1Params 
R0002 n000mid n000 {level1R}
R00001 n000 n0000mid {level2R}
yneuron neuron0000 n0000mid 0 level2Params 
R00002 n0000mid n0000 {level2R}
R000001 n0000 n00000mid {level3R}
yneuron neuron00000 n00000mid 0 level3Params 
R000002 n00000mid n00000 {level3R}
R0000001 n00000 n000000mid {level4R}
yneuron neuron000000 n000000mid 0 level4Params 
R0000002 n000000mid n000000 {level4R}
R00000001 n000000 n0000000mid {level5R}
yneuron neuron0000000 n0000000mid 0 level5Params 
R00000002 n0000000mid n0000000 {level5R}
R000000001 n0000000 n00000000mid {level6R}
yneuron neuron00000000 n00000000mid 0 level6Params 
R000000002 n00000000mid n00000000 {level6R}
R0000000001 n00000000 n000000000mid {level7R}
yneuron neuron000000000 n000000000mid 0 level7Params 
R0000000002 n000000000mid n000000000 {level7R}
R00000000001 n000000000 n0000000000mid {level8R}
yneuron neuron0000000000 n0000000000mid 0 level8Params 
R00000000002 n0000000000mid n0000000000 {level8R}
R000000000001 n0000000000 n00000000000mid {level9R}
yneuron neuron00000000000 n00000000000mid 0 level9Params 
R000000000002 n00000000000mid n00000000000 {level9R}
R000000000011 n0000000000 n00000000001mid {level9R}
yneuron neuron00000000001 n00000000001mid 0 level9Params 
R000000000012 n00000000001mid n00000000001 {level9R}
R00000000011 n000000000 n0000000001mid {level8R}
yneuron neuron0000000001 n0000000001mid 0 level8Params 
R00000000012 n0000000001mid n0000000001 {level8R}
R000000000101 n0000000001 n00000000010mid {level9R}
yneuron neuron00000000010 n00000000010mid 0 level9Params 
R000000000102 n00000000010mid n00000000010 {level9R}
R000000000111 n0000000001 n00000000011mid {level9R}
yneuron neuron00000000011 n00000000011mid 0 level9Params 
R000000000112 n00000000011mid n00000000011 {level9R}
R0000000011 n00000000 n000000001mid {level7R}
yneuron neuron000000001 n000000001mid 0 level7Params 
R0000000012 n000000001mid n000000001 {level7R}
R00000000101 n000000001 n0000000010mid {level8R}
yneuron neuron0000000010 n0000000010mid 0 level8Params 
R00000000102 n0000000010mid n0000000010 {level8R}
R000000001001 n0000000010 n00000000100mid {level9R}
yneuron neuron00000000100 n00000000100mid 0 level9Params 
R000000001002 n00000000100mid n00000000100 {level9R}
R000000001011 n0000000010 n00000000101mid {level9R}
yneuron neuron00000000101 n00000000101mid 0 level9Params 
R000000001012 n00000000101mid n00000000101 {level9R}
R00000000111 n000000001 n0000000011mid {level8R}
yneuron neuron0000000011 n0000000011mid 0 level8Params 
R00000000112 n0000000011mid n0000000011 {level8R}
R000000001101 n0000000011 n00000000110mid {level9R}
yneuron neuron00000000110 n00000000110mid 0 level9Params 
R000000001102 n00000000110mid n00000000110 {level9R}
R000000001111 n0000000011 n00000000111mid {level9R}
yneuron neuron00000000111 n00000000111mid 0 level9Params 
R000000001112 n00000000111mid n00000000111 {level9R}
R000000011 n0000000 n00000001mid {level6R}
yneuron neuron00000001 n00000001mid 0 level6Params 
R000000012 n00000001mid n00000001 {level6R}
R0000000101 n00000001 n000000010mid {level7R}
yneuron neuron000000010 n000000010mid 0 level7Params 
R0000000102 n000000010mid n000000010 {level7R}
R00000001001 n000000010 n0000000100mid {level8R}
yneuron neuron0000000100 n0000000100mid 0 level8Params 
R00000001002 n0000000100mid n0000000100 {level8R}
R000000010001 n0000000100 n00000001000mid {level9R}
yneuron neuron00000001000 n00000001000mid 0 level9Params 
R000000010002 n00000001000mid n00000001000 {level9R}
R000000010011 n0000000100 n00000001001mid {level9R}
yneuron neuron00000001001 n00000001001mid 0 level9Params 
R000000010012 n00000001001mid n00000001001 {level9R}
R00000001011 n000000010 n0000000101mid {level8R}
yneuron neuron0000000101 n0000000101mid 0 level8Params 
R00000001012 n0000000101mid n0000000101 {level8R}
R000000010101 n0000000101 n00000001010mid {level9R}
yneuron neuron00000001010 n00000001010mid 0 level9Params 
R000000010102 n00000001010mid n00000001010 {level9R}
R000000010111 n0000000101 n00000001011mid {level9R}
yneuron neuron00000001011 n00000001011mid 0 level9Params 
R000000010112 n00000001011mid n00000001011 {level9R}
R0000000111 n00000001 n000000011mid {level7R}
yneuron neuron000000011 n000000011mid 0 level7Params 
R0000000112 n000000011mid n000000011 {level7R}
R00000001101 n000000011 n0000000110mid {level8R}
yneuron neuron0000000110 n0000000110mid 0 level8Params 
R00000001102 n0000000110mid n0000000110 {level8R}
R000000011001 n0000000110 n00000001100mid {level9R}
yneuron neuron00000001100 n00000001100mid 0 level9Params 
R000000011002 n00000001100mid n00000001100 {level9R}
R000000011011 n0000000110 n00000001101mid {level9R}
yneuron neuron00000001101 n00000001101mid 0 level9Params 
R000000011012 n00000001101mid n00000001101 {level9R}
R00000001111 n000000011 n0000000111mid {level8R}
yneuron neuron0000000111 n0000000111mid 0 level8Params 
R00000001112 n0000000111mid n0000000111 {level8R}
R000000011101 n0000000111 n00000001110mid {level9R}
yneuron neuron00000001110 n00000001110mid 0 level9Params 
R000000011102 n00000001110mid n00000001110 {level9R}
R000000011111 n0000000111 n00000001111mid {level9R}
yneuron neuron00000001111 n00000001111mid 0 level9Params 
R000000011112 n00000001111mid n00000001111 {level9R}
R00000011 n000000 n0000001mid {level5R}
yneuron neuron0000001 n0000001mid 0 level5Params 
R00000012 n0000001mid n0000001 {level5R}
R000000101 n0000001 n00000010mid {level6R}
yneuron neuron00000010 n00000010mid 0 level6Params 
R000000102 n00000010mid n00000010 {level6R}
R0000001001 n00000010 n000000100mid {level7R}
yneuron neuron000000100 n000000100mid 0 level7Params 
R0000001002 n000000100mid n000000100 {level7R}
R00000010001 n000000100 n0000001000mid {level8R}
yneuron neuron0000001000 n0000001000mid 0 level8Params 
R00000010002 n0000001000mid n0000001000 {level8R}
R000000100001 n0000001000 n00000010000mid {level9R}
yneuron neuron00000010000 n00000010000mid 0 level9Params 
R000000100002 n00000010000mid n00000010000 {level9R}
R000000100011 n0000001000 n00000010001mid {level9R}
yneuron neuron00000010001 n00000010001mid 0 level9Params 
R000000100012 n00000010001mid n00000010001 {level9R}
R00000010011 n000000100 n0000001001mid {level8R}
yneuron neuron0000001001 n0000001001mid 0 level8Params 
R00000010012 n0000001001mid n0000001001 {level8R}
R000000100101 n0000001001 n00000010010mid {level9R}
yneuron neuron00000010010 n00000010010mid 0 level9Params 
R000000100102 n00000010010mid n00000010010 {level9R}
R000000100111 n0000001001 n00000010011mid {level9R}
yneuron neuron00000010011 n00000010011mid 0 level9Params 
R000000100112 n00000010011mid n00000010011 {level9R}
R0000001011 n00000010 n000000101mid {level7R}
yneuron neuron000000101 n000000101mid 0 level7Params 
R0000001012 n000000101mid n000000101 {level7R}
R00000010101 n000000101 n0000001010mid {level8R}
yneuron neuron0000001010 n0000001010mid 0 level8Params 
R00000010102 n0000001010mid n0000001010 {level8R}
R000000101001 n0000001010 n00000010100mid {level9R}
yneuron neuron00000010100 n00000010100mid 0 level9Params 
R000000101002 n00000010100mid n00000010100 {level9R}
R000000101011 n0000001010 n00000010101mid {level9R}
yneuron neuron00000010101 n00000010101mid 0 level9Params 
R000000101012 n00000010101mid n00000010101 {level9R}
R00000010111 n000000101 n0000001011mid {level8R}
yneuron neuron0000001011 n0000001011mid 0 level8Params 
R00000010112 n0000001011mid n0000001011 {level8R}
R000000101101 n0000001011 n00000010110mid {level9R}
yneuron neuron00000010110 n00000010110mid 0 level9Params 
R000000101102 n00000010110mid n00000010110 {level9R}
R000000101111 n0000001011 n00000010111mid {level9R}
yneuron neuron00000010111 n00000010111mid 0 level9Params 
R000000101112 n00000010111mid n00000010111 {level9R}
R000000111 n0000001 n00000011mid {level6R}
yneuron neuron00000011 n00000011mid 0 level6Params 
R000000112 n00000011mid n00000011 {level6R}
R0000001101 n00000011 n000000110mid {level7R}
yneuron neuron000000110 n000000110mid 0 level7Params 
R0000001102 n000000110mid n000000110 {level7R}
R00000011001 n000000110 n0000001100mid {level8R}
yneuron neuron0000001100 n0000001100mid 0 level8Params 
R00000011002 n0000001100mid n0000001100 {level8R}
R000000110001 n0000001100 n00000011000mid {level9R}
yneuron neuron00000011000 n00000011000mid 0 level9Params 
R000000110002 n00000011000mid n00000011000 {level9R}
R000000110011 n0000001100 n00000011001mid {level9R}
yneuron neuron00000011001 n00000011001mid 0 level9Params 
R000000110012 n00000011001mid n00000011001 {level9R}
R00000011011 n000000110 n0000001101mid {level8R}
yneuron neuron0000001101 n0000001101mid 0 level8Params 
R00000011012 n0000001101mid n0000001101 {level8R}
R000000110101 n0000001101 n00000011010mid {level9R}
yneuron neuron00000011010 n00000011010mid 0 level9Params 
R000000110102 n00000011010mid n00000011010 {level9R}
R000000110111 n0000001101 n00000011011mid {level9R}
yneuron neuron00000011011 n00000011011mid 0 level9Params 
R000000110112 n00000011011mid n00000011011 {level9R}
R0000001111 n00000011 n000000111mid {level7R}
yneuron neuron000000111 n000000111mid 0 level7Params 
R0000001112 n000000111mid n000000111 {level7R}
R00000011101 n000000111 n0000001110mid {level8R}
yneuron neuron0000001110 n0000001110mid 0 level8Params 
R00000011102 n0000001110mid n0000001110 {level8R}
R000000111001 n0000001110 n00000011100mid {level9R}
yneuron neuron00000011100 n00000011100mid 0 level9Params 
R000000111002 n00000011100mid n00000011100 {level9R}
R000000111011 n0000001110 n00000011101mid {level9R}
yneuron neuron00000011101 n00000011101mid 0 level9Params 
R000000111012 n00000011101mid n00000011101 {level9R}
R00000011111 n000000111 n0000001111mid {level8R}
yneuron neuron0000001111 n0000001111mid 0 level8Params 
R00000011112 n0000001111mid n0000001111 {level8R}
R000000111101 n0000001111 n00000011110mid {level9R}
yneuron neuron00000011110 n00000011110mid 0 level9Params 
R000000111102 n00000011110mid n00000011110 {level9R}
R000000111111 n0000001111 n00000011111mid {level9R}
yneuron neuron00000011111 n00000011111mid 0 level9Params 
R000000111112 n00000011111mid n00000011111 {level9R}
R0000011 n00000 n000001mid {level4R}
yneuron neuron000001 n000001mid 0 level4Params 
R0000012 n000001mid n000001 {level4R}
R00000101 n000001 n0000010mid {level5R}
yneuron neuron0000010 n0000010mid 0 level5Params 
R00000102 n0000010mid n0000010 {level5R}
R000001001 n0000010 n00000100mid {level6R}
yneuron neuron00000100 n00000100mid 0 level6Params 
R000001002 n00000100mid n00000100 {level6R}
R0000010001 n00000100 n000001000mid {level7R}
yneuron neuron000001000 n000001000mid 0 level7Params 
R0000010002 n000001000mid n000001000 {level7R}
R00000100001 n000001000 n0000010000mid {level8R}
yneuron neuron0000010000 n0000010000mid 0 level8Params 
R00000100002 n0000010000mid n0000010000 {level8R}
R000001000001 n0000010000 n00000100000mid {level9R}
yneuron neuron00000100000 n00000100000mid 0 level9Params 
R000001000002 n00000100000mid n00000100000 {level9R}
R000001000011 n0000010000 n00000100001mid {level9R}
yneuron neuron00000100001 n00000100001mid 0 level9Params 
R000001000012 n00000100001mid n00000100001 {level9R}
R00000100011 n000001000 n0000010001mid {level8R}
yneuron neuron0000010001 n0000010001mid 0 level8Params 
R00000100012 n0000010001mid n0000010001 {level8R}
R000001000101 n0000010001 n00000100010mid {level9R}
yneuron neuron00000100010 n00000100010mid 0 level9Params 
R000001000102 n00000100010mid n00000100010 {level9R}
R000001000111 n0000010001 n00000100011mid {level9R}
yneuron neuron00000100011 n00000100011mid 0 level9Params 
R000001000112 n00000100011mid n00000100011 {level9R}
R0000010011 n00000100 n000001001mid {level7R}
yneuron neuron000001001 n000001001mid 0 level7Params 
R0000010012 n000001001mid n000001001 {level7R}
R00000100101 n000001001 n0000010010mid {level8R}
yneuron neuron0000010010 n0000010010mid 0 level8Params 
R00000100102 n0000010010mid n0000010010 {level8R}
R000001001001 n0000010010 n00000100100mid {level9R}
yneuron neuron00000100100 n00000100100mid 0 level9Params 
R000001001002 n00000100100mid n00000100100 {level9R}
R000001001011 n0000010010 n00000100101mid {level9R}
yneuron neuron00000100101 n00000100101mid 0 level9Params 
R000001001012 n00000100101mid n00000100101 {level9R}
R00000100111 n000001001 n0000010011mid {level8R}
yneuron neuron0000010011 n0000010011mid 0 level8Params 
R00000100112 n0000010011mid n0000010011 {level8R}
R000001001101 n0000010011 n00000100110mid {level9R}
yneuron neuron00000100110 n00000100110mid 0 level9Params 
R000001001102 n00000100110mid n00000100110 {level9R}
R000001001111 n0000010011 n00000100111mid {level9R}
yneuron neuron00000100111 n00000100111mid 0 level9Params 
R000001001112 n00000100111mid n00000100111 {level9R}
R000001011 n0000010 n00000101mid {level6R}
yneuron neuron00000101 n00000101mid 0 level6Params 
R000001012 n00000101mid n00000101 {level6R}
R0000010101 n00000101 n000001010mid {level7R}
yneuron neuron000001010 n000001010mid 0 level7Params 
R0000010102 n000001010mid n000001010 {level7R}
R00000101001 n000001010 n0000010100mid {level8R}
yneuron neuron0000010100 n0000010100mid 0 level8Params 
R00000101002 n0000010100mid n0000010100 {level8R}
R000001010001 n0000010100 n00000101000mid {level9R}
yneuron neuron00000101000 n00000101000mid 0 level9Params 
R000001010002 n00000101000mid n00000101000 {level9R}
R000001010011 n0000010100 n00000101001mid {level9R}
yneuron neuron00000101001 n00000101001mid 0 level9Params 
R000001010012 n00000101001mid n00000101001 {level9R}
R00000101011 n000001010 n0000010101mid {level8R}
yneuron neuron0000010101 n0000010101mid 0 level8Params 
R00000101012 n0000010101mid n0000010101 {level8R}
R000001010101 n0000010101 n00000101010mid {level9R}
yneuron neuron00000101010 n00000101010mid 0 level9Params 
R000001010102 n00000101010mid n00000101010 {level9R}
R000001010111 n0000010101 n00000101011mid {level9R}
yneuron neuron00000101011 n00000101011mid 0 level9Params 
R000001010112 n00000101011mid n00000101011 {level9R}
R0000010111 n00000101 n000001011mid {level7R}
yneuron neuron000001011 n000001011mid 0 level7Params 
R0000010112 n000001011mid n000001011 {level7R}
R00000101101 n000001011 n0000010110mid {level8R}
yneuron neuron0000010110 n0000010110mid 0 level8Params 
R00000101102 n0000010110mid n0000010110 {level8R}
R000001011001 n0000010110 n00000101100mid {level9R}
yneuron neuron00000101100 n00000101100mid 0 level9Params 
R000001011002 n00000101100mid n00000101100 {level9R}
R000001011011 n0000010110 n00000101101mid {level9R}
yneuron neuron00000101101 n00000101101mid 0 level9Params 
R000001011012 n00000101101mid n00000101101 {level9R}
R00000101111 n000001011 n0000010111mid {level8R}
yneuron neuron0000010111 n0000010111mid 0 level8Params 
R00000101112 n0000010111mid n0000010111 {level8R}
R000001011101 n0000010111 n00000101110mid {level9R}
yneuron neuron00000101110 n00000101110mid 0 level9Params 
R000001011102 n00000101110mid n00000101110 {level9R}
R000001011111 n0000010111 n00000101111mid {level9R}
yneuron neuron00000101111 n00000101111mid 0 level9Params 
R000001011112 n00000101111mid n00000101111 {level9R}
R00000111 n000001 n0000011mid {level5R}
yneuron neuron0000011 n0000011mid 0 level5Params 
R00000112 n0000011mid n0000011 {level5R}
R000001101 n0000011 n00000110mid {level6R}
yneuron neuron00000110 n00000110mid 0 level6Params 
R000001102 n00000110mid n00000110 {level6R}
R0000011001 n00000110 n000001100mid {level7R}
yneuron neuron000001100 n000001100mid 0 level7Params 
R0000011002 n000001100mid n000001100 {level7R}
R00000110001 n000001100 n0000011000mid {level8R}
yneuron neuron0000011000 n0000011000mid 0 level8Params 
R00000110002 n0000011000mid n0000011000 {level8R}
R000001100001 n0000011000 n00000110000mid {level9R}
yneuron neuron00000110000 n00000110000mid 0 level9Params 
R000001100002 n00000110000mid n00000110000 {level9R}
R000001100011 n0000011000 n00000110001mid {level9R}
yneuron neuron00000110001 n00000110001mid 0 level9Params 
R000001100012 n00000110001mid n00000110001 {level9R}
R00000110011 n000001100 n0000011001mid {level8R}
yneuron neuron0000011001 n0000011001mid 0 level8Params 
R00000110012 n0000011001mid n0000011001 {level8R}
R000001100101 n0000011001 n00000110010mid {level9R}
yneuron neuron00000110010 n00000110010mid 0 level9Params 
R000001100102 n00000110010mid n00000110010 {level9R}
R000001100111 n0000011001 n00000110011mid {level9R}
yneuron neuron00000110011 n00000110011mid 0 level9Params 
R000001100112 n00000110011mid n00000110011 {level9R}
R0000011011 n00000110 n000001101mid {level7R}
yneuron neuron000001101 n000001101mid 0 level7Params 
R0000011012 n000001101mid n000001101 {level7R}
R00000110101 n000001101 n0000011010mid {level8R}
yneuron neuron0000011010 n0000011010mid 0 level8Params 
R00000110102 n0000011010mid n0000011010 {level8R}
R000001101001 n0000011010 n00000110100mid {level9R}
yneuron neuron00000110100 n00000110100mid 0 level9Params 
R000001101002 n00000110100mid n00000110100 {level9R}
R000001101011 n0000011010 n00000110101mid {level9R}
yneuron neuron00000110101 n00000110101mid 0 level9Params 
R000001101012 n00000110101mid n00000110101 {level9R}
R00000110111 n000001101 n0000011011mid {level8R}
yneuron neuron0000011011 n0000011011mid 0 level8Params 
R00000110112 n0000011011mid n0000011011 {level8R}
R000001101101 n0000011011 n00000110110mid {level9R}
yneuron neuron00000110110 n00000110110mid 0 level9Params 
R000001101102 n00000110110mid n00000110110 {level9R}
R000001101111 n0000011011 n00000110111mid {level9R}
yneuron neuron00000110111 n00000110111mid 0 level9Params 
R000001101112 n00000110111mid n00000110111 {level9R}
R000001111 n0000011 n00000111mid {level6R}
yneuron neuron00000111 n00000111mid 0 level6Params 
R000001112 n00000111mid n00000111 {level6R}
R0000011101 n00000111 n000001110mid {level7R}
yneuron neuron000001110 n000001110mid 0 level7Params 
R0000011102 n000001110mid n000001110 {level7R}
R00000111001 n000001110 n0000011100mid {level8R}
yneuron neuron0000011100 n0000011100mid 0 level8Params 
R00000111002 n0000011100mid n0000011100 {level8R}
R000001110001 n0000011100 n00000111000mid {level9R}
yneuron neuron00000111000 n00000111000mid 0 level9Params 
R000001110002 n00000111000mid n00000111000 {level9R}
R000001110011 n0000011100 n00000111001mid {level9R}
yneuron neuron00000111001 n00000111001mid 0 level9Params 
R000001110012 n00000111001mid n00000111001 {level9R}
R00000111011 n000001110 n0000011101mid {level8R}
yneuron neuron0000011101 n0000011101mid 0 level8Params 
R00000111012 n0000011101mid n0000011101 {level8R}
R000001110101 n0000011101 n00000111010mid {level9R}
yneuron neuron00000111010 n00000111010mid 0 level9Params 
R000001110102 n00000111010mid n00000111010 {level9R}
R000001110111 n0000011101 n00000111011mid {level9R}
yneuron neuron00000111011 n00000111011mid 0 level9Params 
R000001110112 n00000111011mid n00000111011 {level9R}
R0000011111 n00000111 n000001111mid {level7R}
yneuron neuron000001111 n000001111mid 0 level7Params 
R0000011112 n000001111mid n000001111 {level7R}
R00000111101 n000001111 n0000011110mid {level8R}
yneuron neuron0000011110 n0000011110mid 0 level8Params 
R00000111102 n0000011110mid n0000011110 {level8R}
R000001111001 n0000011110 n00000111100mid {level9R}
yneuron neuron00000111100 n00000111100mid 0 level9Params 
R000001111002 n00000111100mid n00000111100 {level9R}
R000001111011 n0000011110 n00000111101mid {level9R}
yneuron neuron00000111101 n00000111101mid 0 level9Params 
R000001111012 n00000111101mid n00000111101 {level9R}
R00000111111 n000001111 n0000011111mid {level8R}
yneuron neuron0000011111 n0000011111mid 0 level8Params 
R00000111112 n0000011111mid n0000011111 {level8R}
R000001111101 n0000011111 n00000111110mid {level9R}
yneuron neuron00000111110 n00000111110mid 0 level9Params 
R000001111102 n00000111110mid n00000111110 {level9R}
R000001111111 n0000011111 n00000111111mid {level9R}
yneuron neuron00000111111 n00000111111mid 0 level9Params 
R000001111112 n00000111111mid n00000111111 {level9R}
R000011 n0000 n00001mid {level3R}
yneuron neuron00001 n00001mid 0 level3Params 
R000012 n00001mid n00001 {level3R}
R0000101 n00001 n000010mid {level4R}
yneuron neuron000010 n000010mid 0 level4Params 
R0000102 n000010mid n000010 {level4R}
R00001001 n000010 n0000100mid {level5R}
yneuron neuron0000100 n0000100mid 0 level5Params 
R00001002 n0000100mid n0000100 {level5R}
R000010001 n0000100 n00001000mid {level6R}
yneuron neuron00001000 n00001000mid 0 level6Params 
R000010002 n00001000mid n00001000 {level6R}
R0000100001 n00001000 n000010000mid {level7R}
yneuron neuron000010000 n000010000mid 0 level7Params 
R0000100002 n000010000mid n000010000 {level7R}
R00001000001 n000010000 n0000100000mid {level8R}
yneuron neuron0000100000 n0000100000mid 0 level8Params 
R00001000002 n0000100000mid n0000100000 {level8R}
R000010000001 n0000100000 n00001000000mid {level9R}
yneuron neuron00001000000 n00001000000mid 0 level9Params 
R000010000002 n00001000000mid n00001000000 {level9R}
R000010000011 n0000100000 n00001000001mid {level9R}
yneuron neuron00001000001 n00001000001mid 0 level9Params 
R000010000012 n00001000001mid n00001000001 {level9R}
R00001000011 n000010000 n0000100001mid {level8R}
yneuron neuron0000100001 n0000100001mid 0 level8Params 
R00001000012 n0000100001mid n0000100001 {level8R}
R000010000101 n0000100001 n00001000010mid {level9R}
yneuron neuron00001000010 n00001000010mid 0 level9Params 
R000010000102 n00001000010mid n00001000010 {level9R}
R000010000111 n0000100001 n00001000011mid {level9R}
yneuron neuron00001000011 n00001000011mid 0 level9Params 
R000010000112 n00001000011mid n00001000011 {level9R}
R0000100011 n00001000 n000010001mid {level7R}
yneuron neuron000010001 n000010001mid 0 level7Params 
R0000100012 n000010001mid n000010001 {level7R}
R00001000101 n000010001 n0000100010mid {level8R}
yneuron neuron0000100010 n0000100010mid 0 level8Params 
R00001000102 n0000100010mid n0000100010 {level8R}
R000010001001 n0000100010 n00001000100mid {level9R}
yneuron neuron00001000100 n00001000100mid 0 level9Params 
R000010001002 n00001000100mid n00001000100 {level9R}
R000010001011 n0000100010 n00001000101mid {level9R}
yneuron neuron00001000101 n00001000101mid 0 level9Params 
R000010001012 n00001000101mid n00001000101 {level9R}
R00001000111 n000010001 n0000100011mid {level8R}
yneuron neuron0000100011 n0000100011mid 0 level8Params 
R00001000112 n0000100011mid n0000100011 {level8R}
R000010001101 n0000100011 n00001000110mid {level9R}
yneuron neuron00001000110 n00001000110mid 0 level9Params 
R000010001102 n00001000110mid n00001000110 {level9R}
R000010001111 n0000100011 n00001000111mid {level9R}
yneuron neuron00001000111 n00001000111mid 0 level9Params 
R000010001112 n00001000111mid n00001000111 {level9R}
R000010011 n0000100 n00001001mid {level6R}
yneuron neuron00001001 n00001001mid 0 level6Params 
R000010012 n00001001mid n00001001 {level6R}
R0000100101 n00001001 n000010010mid {level7R}
yneuron neuron000010010 n000010010mid 0 level7Params 
R0000100102 n000010010mid n000010010 {level7R}
R00001001001 n000010010 n0000100100mid {level8R}
yneuron neuron0000100100 n0000100100mid 0 level8Params 
R00001001002 n0000100100mid n0000100100 {level8R}
R000010010001 n0000100100 n00001001000mid {level9R}
yneuron neuron00001001000 n00001001000mid 0 level9Params 
R000010010002 n00001001000mid n00001001000 {level9R}
R000010010011 n0000100100 n00001001001mid {level9R}
yneuron neuron00001001001 n00001001001mid 0 level9Params 
R000010010012 n00001001001mid n00001001001 {level9R}
R00001001011 n000010010 n0000100101mid {level8R}
yneuron neuron0000100101 n0000100101mid 0 level8Params 
R00001001012 n0000100101mid n0000100101 {level8R}
R000010010101 n0000100101 n00001001010mid {level9R}
yneuron neuron00001001010 n00001001010mid 0 level9Params 
R000010010102 n00001001010mid n00001001010 {level9R}
R000010010111 n0000100101 n00001001011mid {level9R}
yneuron neuron00001001011 n00001001011mid 0 level9Params 
R000010010112 n00001001011mid n00001001011 {level9R}
R0000100111 n00001001 n000010011mid {level7R}
yneuron neuron000010011 n000010011mid 0 level7Params 
R0000100112 n000010011mid n000010011 {level7R}
R00001001101 n000010011 n0000100110mid {level8R}
yneuron neuron0000100110 n0000100110mid 0 level8Params 
R00001001102 n0000100110mid n0000100110 {level8R}
R000010011001 n0000100110 n00001001100mid {level9R}
yneuron neuron00001001100 n00001001100mid 0 level9Params 
R000010011002 n00001001100mid n00001001100 {level9R}
R000010011011 n0000100110 n00001001101mid {level9R}
yneuron neuron00001001101 n00001001101mid 0 level9Params 
R000010011012 n00001001101mid n00001001101 {level9R}
R00001001111 n000010011 n0000100111mid {level8R}
yneuron neuron0000100111 n0000100111mid 0 level8Params 
R00001001112 n0000100111mid n0000100111 {level8R}
R000010011101 n0000100111 n00001001110mid {level9R}
yneuron neuron00001001110 n00001001110mid 0 level9Params 
R000010011102 n00001001110mid n00001001110 {level9R}
R000010011111 n0000100111 n00001001111mid {level9R}
yneuron neuron00001001111 n00001001111mid 0 level9Params 
R000010011112 n00001001111mid n00001001111 {level9R}
R00001011 n000010 n0000101mid {level5R}
yneuron neuron0000101 n0000101mid 0 level5Params 
R00001012 n0000101mid n0000101 {level5R}
R000010101 n0000101 n00001010mid {level6R}
yneuron neuron00001010 n00001010mid 0 level6Params 
R000010102 n00001010mid n00001010 {level6R}
R0000101001 n00001010 n000010100mid {level7R}
yneuron neuron000010100 n000010100mid 0 level7Params 
R0000101002 n000010100mid n000010100 {level7R}
R00001010001 n000010100 n0000101000mid {level8R}
yneuron neuron0000101000 n0000101000mid 0 level8Params 
R00001010002 n0000101000mid n0000101000 {level8R}
R000010100001 n0000101000 n00001010000mid {level9R}
yneuron neuron00001010000 n00001010000mid 0 level9Params 
R000010100002 n00001010000mid n00001010000 {level9R}
R000010100011 n0000101000 n00001010001mid {level9R}
yneuron neuron00001010001 n00001010001mid 0 level9Params 
R000010100012 n00001010001mid n00001010001 {level9R}
R00001010011 n000010100 n0000101001mid {level8R}
yneuron neuron0000101001 n0000101001mid 0 level8Params 
R00001010012 n0000101001mid n0000101001 {level8R}
R000010100101 n0000101001 n00001010010mid {level9R}
yneuron neuron00001010010 n00001010010mid 0 level9Params 
R000010100102 n00001010010mid n00001010010 {level9R}
R000010100111 n0000101001 n00001010011mid {level9R}
yneuron neuron00001010011 n00001010011mid 0 level9Params 
R000010100112 n00001010011mid n00001010011 {level9R}
R0000101011 n00001010 n000010101mid {level7R}
yneuron neuron000010101 n000010101mid 0 level7Params 
R0000101012 n000010101mid n000010101 {level7R}
R00001010101 n000010101 n0000101010mid {level8R}
yneuron neuron0000101010 n0000101010mid 0 level8Params 
R00001010102 n0000101010mid n0000101010 {level8R}
R000010101001 n0000101010 n00001010100mid {level9R}
yneuron neuron00001010100 n00001010100mid 0 level9Params 
R000010101002 n00001010100mid n00001010100 {level9R}
R000010101011 n0000101010 n00001010101mid {level9R}
yneuron neuron00001010101 n00001010101mid 0 level9Params 
R000010101012 n00001010101mid n00001010101 {level9R}
R00001010111 n000010101 n0000101011mid {level8R}
yneuron neuron0000101011 n0000101011mid 0 level8Params 
R00001010112 n0000101011mid n0000101011 {level8R}
R000010101101 n0000101011 n00001010110mid {level9R}
yneuron neuron00001010110 n00001010110mid 0 level9Params 
R000010101102 n00001010110mid n00001010110 {level9R}
R000010101111 n0000101011 n00001010111mid {level9R}
yneuron neuron00001010111 n00001010111mid 0 level9Params 
R000010101112 n00001010111mid n00001010111 {level9R}
R000010111 n0000101 n00001011mid {level6R}
yneuron neuron00001011 n00001011mid 0 level6Params 
R000010112 n00001011mid n00001011 {level6R}
R0000101101 n00001011 n000010110mid {level7R}
yneuron neuron000010110 n000010110mid 0 level7Params 
R0000101102 n000010110mid n000010110 {level7R}
R00001011001 n000010110 n0000101100mid {level8R}
yneuron neuron0000101100 n0000101100mid 0 level8Params 
R00001011002 n0000101100mid n0000101100 {level8R}
R000010110001 n0000101100 n00001011000mid {level9R}
yneuron neuron00001011000 n00001011000mid 0 level9Params 
R000010110002 n00001011000mid n00001011000 {level9R}
R000010110011 n0000101100 n00001011001mid {level9R}
yneuron neuron00001011001 n00001011001mid 0 level9Params 
R000010110012 n00001011001mid n00001011001 {level9R}
R00001011011 n000010110 n0000101101mid {level8R}
yneuron neuron0000101101 n0000101101mid 0 level8Params 
R00001011012 n0000101101mid n0000101101 {level8R}
R000010110101 n0000101101 n00001011010mid {level9R}
yneuron neuron00001011010 n00001011010mid 0 level9Params 
R000010110102 n00001011010mid n00001011010 {level9R}
R000010110111 n0000101101 n00001011011mid {level9R}
yneuron neuron00001011011 n00001011011mid 0 level9Params 
R000010110112 n00001011011mid n00001011011 {level9R}
R0000101111 n00001011 n000010111mid {level7R}
yneuron neuron000010111 n000010111mid 0 level7Params 
R0000101112 n000010111mid n000010111 {level7R}
R00001011101 n000010111 n0000101110mid {level8R}
yneuron neuron0000101110 n0000101110mid 0 level8Params 
R00001011102 n0000101110mid n0000101110 {level8R}
R000010111001 n0000101110 n00001011100mid {level9R}
yneuron neuron00001011100 n00001011100mid 0 level9Params 
R000010111002 n00001011100mid n00001011100 {level9R}
R000010111011 n0000101110 n00001011101mid {level9R}
yneuron neuron00001011101 n00001011101mid 0 level9Params 
R000010111012 n00001011101mid n00001011101 {level9R}
R00001011111 n000010111 n0000101111mid {level8R}
yneuron neuron0000101111 n0000101111mid 0 level8Params 
R00001011112 n0000101111mid n0000101111 {level8R}
R000010111101 n0000101111 n00001011110mid {level9R}
yneuron neuron00001011110 n00001011110mid 0 level9Params 
R000010111102 n00001011110mid n00001011110 {level9R}
R000010111111 n0000101111 n00001011111mid {level9R}
yneuron neuron00001011111 n00001011111mid 0 level9Params 
R000010111112 n00001011111mid n00001011111 {level9R}
R0000111 n00001 n000011mid {level4R}
yneuron neuron000011 n000011mid 0 level4Params 
R0000112 n000011mid n000011 {level4R}
R00001101 n000011 n0000110mid {level5R}
yneuron neuron0000110 n0000110mid 0 level5Params 
R00001102 n0000110mid n0000110 {level5R}
R000011001 n0000110 n00001100mid {level6R}
yneuron neuron00001100 n00001100mid 0 level6Params 
R000011002 n00001100mid n00001100 {level6R}
R0000110001 n00001100 n000011000mid {level7R}
yneuron neuron000011000 n000011000mid 0 level7Params 
R0000110002 n000011000mid n000011000 {level7R}
R00001100001 n000011000 n0000110000mid {level8R}
yneuron neuron0000110000 n0000110000mid 0 level8Params 
R00001100002 n0000110000mid n0000110000 {level8R}
R000011000001 n0000110000 n00001100000mid {level9R}
yneuron neuron00001100000 n00001100000mid 0 level9Params 
R000011000002 n00001100000mid n00001100000 {level9R}
R000011000011 n0000110000 n00001100001mid {level9R}
yneuron neuron00001100001 n00001100001mid 0 level9Params 
R000011000012 n00001100001mid n00001100001 {level9R}
R00001100011 n000011000 n0000110001mid {level8R}
yneuron neuron0000110001 n0000110001mid 0 level8Params 
R00001100012 n0000110001mid n0000110001 {level8R}
R000011000101 n0000110001 n00001100010mid {level9R}
yneuron neuron00001100010 n00001100010mid 0 level9Params 
R000011000102 n00001100010mid n00001100010 {level9R}
R000011000111 n0000110001 n00001100011mid {level9R}
yneuron neuron00001100011 n00001100011mid 0 level9Params 
R000011000112 n00001100011mid n00001100011 {level9R}
R0000110011 n00001100 n000011001mid {level7R}
yneuron neuron000011001 n000011001mid 0 level7Params 
R0000110012 n000011001mid n000011001 {level7R}
R00001100101 n000011001 n0000110010mid {level8R}
yneuron neuron0000110010 n0000110010mid 0 level8Params 
R00001100102 n0000110010mid n0000110010 {level8R}
R000011001001 n0000110010 n00001100100mid {level9R}
yneuron neuron00001100100 n00001100100mid 0 level9Params 
R000011001002 n00001100100mid n00001100100 {level9R}
R000011001011 n0000110010 n00001100101mid {level9R}
yneuron neuron00001100101 n00001100101mid 0 level9Params 
R000011001012 n00001100101mid n00001100101 {level9R}
R00001100111 n000011001 n0000110011mid {level8R}
yneuron neuron0000110011 n0000110011mid 0 level8Params 
R00001100112 n0000110011mid n0000110011 {level8R}
R000011001101 n0000110011 n00001100110mid {level9R}
yneuron neuron00001100110 n00001100110mid 0 level9Params 
R000011001102 n00001100110mid n00001100110 {level9R}
R000011001111 n0000110011 n00001100111mid {level9R}
yneuron neuron00001100111 n00001100111mid 0 level9Params 
R000011001112 n00001100111mid n00001100111 {level9R}
R000011011 n0000110 n00001101mid {level6R}
yneuron neuron00001101 n00001101mid 0 level6Params 
R000011012 n00001101mid n00001101 {level6R}
R0000110101 n00001101 n000011010mid {level7R}
yneuron neuron000011010 n000011010mid 0 level7Params 
R0000110102 n000011010mid n000011010 {level7R}
R00001101001 n000011010 n0000110100mid {level8R}
yneuron neuron0000110100 n0000110100mid 0 level8Params 
R00001101002 n0000110100mid n0000110100 {level8R}
R000011010001 n0000110100 n00001101000mid {level9R}
yneuron neuron00001101000 n00001101000mid 0 level9Params 
R000011010002 n00001101000mid n00001101000 {level9R}
R000011010011 n0000110100 n00001101001mid {level9R}
yneuron neuron00001101001 n00001101001mid 0 level9Params 
R000011010012 n00001101001mid n00001101001 {level9R}
R00001101011 n000011010 n0000110101mid {level8R}
yneuron neuron0000110101 n0000110101mid 0 level8Params 
R00001101012 n0000110101mid n0000110101 {level8R}
R000011010101 n0000110101 n00001101010mid {level9R}
yneuron neuron00001101010 n00001101010mid 0 level9Params 
R000011010102 n00001101010mid n00001101010 {level9R}
R000011010111 n0000110101 n00001101011mid {level9R}
yneuron neuron00001101011 n00001101011mid 0 level9Params 
R000011010112 n00001101011mid n00001101011 {level9R}
R0000110111 n00001101 n000011011mid {level7R}
yneuron neuron000011011 n000011011mid 0 level7Params 
R0000110112 n000011011mid n000011011 {level7R}
R00001101101 n000011011 n0000110110mid {level8R}
yneuron neuron0000110110 n0000110110mid 0 level8Params 
R00001101102 n0000110110mid n0000110110 {level8R}
R000011011001 n0000110110 n00001101100mid {level9R}
yneuron neuron00001101100 n00001101100mid 0 level9Params 
R000011011002 n00001101100mid n00001101100 {level9R}
R000011011011 n0000110110 n00001101101mid {level9R}
yneuron neuron00001101101 n00001101101mid 0 level9Params 
R000011011012 n00001101101mid n00001101101 {level9R}
R00001101111 n000011011 n0000110111mid {level8R}
yneuron neuron0000110111 n0000110111mid 0 level8Params 
R00001101112 n0000110111mid n0000110111 {level8R}
R000011011101 n0000110111 n00001101110mid {level9R}
yneuron neuron00001101110 n00001101110mid 0 level9Params 
R000011011102 n00001101110mid n00001101110 {level9R}
R000011011111 n0000110111 n00001101111mid {level9R}
yneuron neuron00001101111 n00001101111mid 0 level9Params 
R000011011112 n00001101111mid n00001101111 {level9R}
R00001111 n000011 n0000111mid {level5R}
yneuron neuron0000111 n0000111mid 0 level5Params 
R00001112 n0000111mid n0000111 {level5R}
R000011101 n0000111 n00001110mid {level6R}
yneuron neuron00001110 n00001110mid 0 level6Params 
R000011102 n00001110mid n00001110 {level6R}
R0000111001 n00001110 n000011100mid {level7R}
yneuron neuron000011100 n000011100mid 0 level7Params 
R0000111002 n000011100mid n000011100 {level7R}
R00001110001 n000011100 n0000111000mid {level8R}
yneuron neuron0000111000 n0000111000mid 0 level8Params 
R00001110002 n0000111000mid n0000111000 {level8R}
R000011100001 n0000111000 n00001110000mid {level9R}
yneuron neuron00001110000 n00001110000mid 0 level9Params 
R000011100002 n00001110000mid n00001110000 {level9R}
R000011100011 n0000111000 n00001110001mid {level9R}
yneuron neuron00001110001 n00001110001mid 0 level9Params 
R000011100012 n00001110001mid n00001110001 {level9R}
R00001110011 n000011100 n0000111001mid {level8R}
yneuron neuron0000111001 n0000111001mid 0 level8Params 
R00001110012 n0000111001mid n0000111001 {level8R}
R000011100101 n0000111001 n00001110010mid {level9R}
yneuron neuron00001110010 n00001110010mid 0 level9Params 
R000011100102 n00001110010mid n00001110010 {level9R}
R000011100111 n0000111001 n00001110011mid {level9R}
yneuron neuron00001110011 n00001110011mid 0 level9Params 
R000011100112 n00001110011mid n00001110011 {level9R}
R0000111011 n00001110 n000011101mid {level7R}
yneuron neuron000011101 n000011101mid 0 level7Params 
R0000111012 n000011101mid n000011101 {level7R}
R00001110101 n000011101 n0000111010mid {level8R}
yneuron neuron0000111010 n0000111010mid 0 level8Params 
R00001110102 n0000111010mid n0000111010 {level8R}
R000011101001 n0000111010 n00001110100mid {level9R}
yneuron neuron00001110100 n00001110100mid 0 level9Params 
R000011101002 n00001110100mid n00001110100 {level9R}
R000011101011 n0000111010 n00001110101mid {level9R}
yneuron neuron00001110101 n00001110101mid 0 level9Params 
R000011101012 n00001110101mid n00001110101 {level9R}
R00001110111 n000011101 n0000111011mid {level8R}
yneuron neuron0000111011 n0000111011mid 0 level8Params 
R00001110112 n0000111011mid n0000111011 {level8R}
R000011101101 n0000111011 n00001110110mid {level9R}
yneuron neuron00001110110 n00001110110mid 0 level9Params 
R000011101102 n00001110110mid n00001110110 {level9R}
R000011101111 n0000111011 n00001110111mid {level9R}
yneuron neuron00001110111 n00001110111mid 0 level9Params 
R000011101112 n00001110111mid n00001110111 {level9R}
R000011111 n0000111 n00001111mid {level6R}
yneuron neuron00001111 n00001111mid 0 level6Params 
R000011112 n00001111mid n00001111 {level6R}
R0000111101 n00001111 n000011110mid {level7R}
yneuron neuron000011110 n000011110mid 0 level7Params 
R0000111102 n000011110mid n000011110 {level7R}
R00001111001 n000011110 n0000111100mid {level8R}
yneuron neuron0000111100 n0000111100mid 0 level8Params 
R00001111002 n0000111100mid n0000111100 {level8R}
R000011110001 n0000111100 n00001111000mid {level9R}
yneuron neuron00001111000 n00001111000mid 0 level9Params 
R000011110002 n00001111000mid n00001111000 {level9R}
R000011110011 n0000111100 n00001111001mid {level9R}
yneuron neuron00001111001 n00001111001mid 0 level9Params 
R000011110012 n00001111001mid n00001111001 {level9R}
R00001111011 n000011110 n0000111101mid {level8R}
yneuron neuron0000111101 n0000111101mid 0 level8Params 
R00001111012 n0000111101mid n0000111101 {level8R}
R000011110101 n0000111101 n00001111010mid {level9R}
yneuron neuron00001111010 n00001111010mid 0 level9Params 
R000011110102 n00001111010mid n00001111010 {level9R}
R000011110111 n0000111101 n00001111011mid {level9R}
yneuron neuron00001111011 n00001111011mid 0 level9Params 
R000011110112 n00001111011mid n00001111011 {level9R}
R0000111111 n00001111 n000011111mid {level7R}
yneuron neuron000011111 n000011111mid 0 level7Params 
R0000111112 n000011111mid n000011111 {level7R}
R00001111101 n000011111 n0000111110mid {level8R}
yneuron neuron0000111110 n0000111110mid 0 level8Params 
R00001111102 n0000111110mid n0000111110 {level8R}
R000011111001 n0000111110 n00001111100mid {level9R}
yneuron neuron00001111100 n00001111100mid 0 level9Params 
R000011111002 n00001111100mid n00001111100 {level9R}
R000011111011 n0000111110 n00001111101mid {level9R}
yneuron neuron00001111101 n00001111101mid 0 level9Params 
R000011111012 n00001111101mid n00001111101 {level9R}
R00001111111 n000011111 n0000111111mid {level8R}
yneuron neuron0000111111 n0000111111mid 0 level8Params 
R00001111112 n0000111111mid n0000111111 {level8R}
R000011111101 n0000111111 n00001111110mid {level9R}
yneuron neuron00001111110 n00001111110mid 0 level9Params 
R000011111102 n00001111110mid n00001111110 {level9R}
R000011111111 n0000111111 n00001111111mid {level9R}
yneuron neuron00001111111 n00001111111mid 0 level9Params 
R000011111112 n00001111111mid n00001111111 {level9R}
R00011 n000 n0001mid {level2R}
yneuron neuron0001 n0001mid 0 level2Params 
R00012 n0001mid n0001 {level2R}
R000101 n0001 n00010mid {level3R}
yneuron neuron00010 n00010mid 0 level3Params 
R000102 n00010mid n00010 {level3R}
R0001001 n00010 n000100mid {level4R}
yneuron neuron000100 n000100mid 0 level4Params 
R0001002 n000100mid n000100 {level4R}
R00010001 n000100 n0001000mid {level5R}
yneuron neuron0001000 n0001000mid 0 level5Params 
R00010002 n0001000mid n0001000 {level5R}
R000100001 n0001000 n00010000mid {level6R}
yneuron neuron00010000 n00010000mid 0 level6Params 
R000100002 n00010000mid n00010000 {level6R}
R0001000001 n00010000 n000100000mid {level7R}
yneuron neuron000100000 n000100000mid 0 level7Params 
R0001000002 n000100000mid n000100000 {level7R}
R00010000001 n000100000 n0001000000mid {level8R}
yneuron neuron0001000000 n0001000000mid 0 level8Params 
R00010000002 n0001000000mid n0001000000 {level8R}
R000100000001 n0001000000 n00010000000mid {level9R}
yneuron neuron00010000000 n00010000000mid 0 level9Params 
R000100000002 n00010000000mid n00010000000 {level9R}
R000100000011 n0001000000 n00010000001mid {level9R}
yneuron neuron00010000001 n00010000001mid 0 level9Params 
R000100000012 n00010000001mid n00010000001 {level9R}
R00010000011 n000100000 n0001000001mid {level8R}
yneuron neuron0001000001 n0001000001mid 0 level8Params 
R00010000012 n0001000001mid n0001000001 {level8R}
R000100000101 n0001000001 n00010000010mid {level9R}
yneuron neuron00010000010 n00010000010mid 0 level9Params 
R000100000102 n00010000010mid n00010000010 {level9R}
R000100000111 n0001000001 n00010000011mid {level9R}
yneuron neuron00010000011 n00010000011mid 0 level9Params 
R000100000112 n00010000011mid n00010000011 {level9R}
R0001000011 n00010000 n000100001mid {level7R}
yneuron neuron000100001 n000100001mid 0 level7Params 
R0001000012 n000100001mid n000100001 {level7R}
R00010000101 n000100001 n0001000010mid {level8R}
yneuron neuron0001000010 n0001000010mid 0 level8Params 
R00010000102 n0001000010mid n0001000010 {level8R}
R000100001001 n0001000010 n00010000100mid {level9R}
yneuron neuron00010000100 n00010000100mid 0 level9Params 
R000100001002 n00010000100mid n00010000100 {level9R}
R000100001011 n0001000010 n00010000101mid {level9R}
yneuron neuron00010000101 n00010000101mid 0 level9Params 
R000100001012 n00010000101mid n00010000101 {level9R}
R00010000111 n000100001 n0001000011mid {level8R}
yneuron neuron0001000011 n0001000011mid 0 level8Params 
R00010000112 n0001000011mid n0001000011 {level8R}
R000100001101 n0001000011 n00010000110mid {level9R}
yneuron neuron00010000110 n00010000110mid 0 level9Params 
R000100001102 n00010000110mid n00010000110 {level9R}
R000100001111 n0001000011 n00010000111mid {level9R}
yneuron neuron00010000111 n00010000111mid 0 level9Params 
R000100001112 n00010000111mid n00010000111 {level9R}
R000100011 n0001000 n00010001mid {level6R}
yneuron neuron00010001 n00010001mid 0 level6Params 
R000100012 n00010001mid n00010001 {level6R}
R0001000101 n00010001 n000100010mid {level7R}
yneuron neuron000100010 n000100010mid 0 level7Params 
R0001000102 n000100010mid n000100010 {level7R}
R00010001001 n000100010 n0001000100mid {level8R}
yneuron neuron0001000100 n0001000100mid 0 level8Params 
R00010001002 n0001000100mid n0001000100 {level8R}
R000100010001 n0001000100 n00010001000mid {level9R}
yneuron neuron00010001000 n00010001000mid 0 level9Params 
R000100010002 n00010001000mid n00010001000 {level9R}
R000100010011 n0001000100 n00010001001mid {level9R}
yneuron neuron00010001001 n00010001001mid 0 level9Params 
R000100010012 n00010001001mid n00010001001 {level9R}
R00010001011 n000100010 n0001000101mid {level8R}
yneuron neuron0001000101 n0001000101mid 0 level8Params 
R00010001012 n0001000101mid n0001000101 {level8R}
R000100010101 n0001000101 n00010001010mid {level9R}
yneuron neuron00010001010 n00010001010mid 0 level9Params 
R000100010102 n00010001010mid n00010001010 {level9R}
R000100010111 n0001000101 n00010001011mid {level9R}
yneuron neuron00010001011 n00010001011mid 0 level9Params 
R000100010112 n00010001011mid n00010001011 {level9R}
R0001000111 n00010001 n000100011mid {level7R}
yneuron neuron000100011 n000100011mid 0 level7Params 
R0001000112 n000100011mid n000100011 {level7R}
R00010001101 n000100011 n0001000110mid {level8R}
yneuron neuron0001000110 n0001000110mid 0 level8Params 
R00010001102 n0001000110mid n0001000110 {level8R}
R000100011001 n0001000110 n00010001100mid {level9R}
yneuron neuron00010001100 n00010001100mid 0 level9Params 
R000100011002 n00010001100mid n00010001100 {level9R}
R000100011011 n0001000110 n00010001101mid {level9R}
yneuron neuron00010001101 n00010001101mid 0 level9Params 
R000100011012 n00010001101mid n00010001101 {level9R}
R00010001111 n000100011 n0001000111mid {level8R}
yneuron neuron0001000111 n0001000111mid 0 level8Params 
R00010001112 n0001000111mid n0001000111 {level8R}
R000100011101 n0001000111 n00010001110mid {level9R}
yneuron neuron00010001110 n00010001110mid 0 level9Params 
R000100011102 n00010001110mid n00010001110 {level9R}
R000100011111 n0001000111 n00010001111mid {level9R}
yneuron neuron00010001111 n00010001111mid 0 level9Params 
R000100011112 n00010001111mid n00010001111 {level9R}
R00010011 n000100 n0001001mid {level5R}
yneuron neuron0001001 n0001001mid 0 level5Params 
R00010012 n0001001mid n0001001 {level5R}
R000100101 n0001001 n00010010mid {level6R}
yneuron neuron00010010 n00010010mid 0 level6Params 
R000100102 n00010010mid n00010010 {level6R}
R0001001001 n00010010 n000100100mid {level7R}
yneuron neuron000100100 n000100100mid 0 level7Params 
R0001001002 n000100100mid n000100100 {level7R}
R00010010001 n000100100 n0001001000mid {level8R}
yneuron neuron0001001000 n0001001000mid 0 level8Params 
R00010010002 n0001001000mid n0001001000 {level8R}
R000100100001 n0001001000 n00010010000mid {level9R}
yneuron neuron00010010000 n00010010000mid 0 level9Params 
R000100100002 n00010010000mid n00010010000 {level9R}
R000100100011 n0001001000 n00010010001mid {level9R}
yneuron neuron00010010001 n00010010001mid 0 level9Params 
R000100100012 n00010010001mid n00010010001 {level9R}
R00010010011 n000100100 n0001001001mid {level8R}
yneuron neuron0001001001 n0001001001mid 0 level8Params 
R00010010012 n0001001001mid n0001001001 {level8R}
R000100100101 n0001001001 n00010010010mid {level9R}
yneuron neuron00010010010 n00010010010mid 0 level9Params 
R000100100102 n00010010010mid n00010010010 {level9R}
R000100100111 n0001001001 n00010010011mid {level9R}
yneuron neuron00010010011 n00010010011mid 0 level9Params 
R000100100112 n00010010011mid n00010010011 {level9R}
R0001001011 n00010010 n000100101mid {level7R}
yneuron neuron000100101 n000100101mid 0 level7Params 
R0001001012 n000100101mid n000100101 {level7R}
R00010010101 n000100101 n0001001010mid {level8R}
yneuron neuron0001001010 n0001001010mid 0 level8Params 
R00010010102 n0001001010mid n0001001010 {level8R}
R000100101001 n0001001010 n00010010100mid {level9R}
yneuron neuron00010010100 n00010010100mid 0 level9Params 
R000100101002 n00010010100mid n00010010100 {level9R}
R000100101011 n0001001010 n00010010101mid {level9R}
yneuron neuron00010010101 n00010010101mid 0 level9Params 
R000100101012 n00010010101mid n00010010101 {level9R}
R00010010111 n000100101 n0001001011mid {level8R}
yneuron neuron0001001011 n0001001011mid 0 level8Params 
R00010010112 n0001001011mid n0001001011 {level8R}
R000100101101 n0001001011 n00010010110mid {level9R}
yneuron neuron00010010110 n00010010110mid 0 level9Params 
R000100101102 n00010010110mid n00010010110 {level9R}
R000100101111 n0001001011 n00010010111mid {level9R}
yneuron neuron00010010111 n00010010111mid 0 level9Params 
R000100101112 n00010010111mid n00010010111 {level9R}
R000100111 n0001001 n00010011mid {level6R}
yneuron neuron00010011 n00010011mid 0 level6Params 
R000100112 n00010011mid n00010011 {level6R}
R0001001101 n00010011 n000100110mid {level7R}
yneuron neuron000100110 n000100110mid 0 level7Params 
R0001001102 n000100110mid n000100110 {level7R}
R00010011001 n000100110 n0001001100mid {level8R}
yneuron neuron0001001100 n0001001100mid 0 level8Params 
R00010011002 n0001001100mid n0001001100 {level8R}
R000100110001 n0001001100 n00010011000mid {level9R}
yneuron neuron00010011000 n00010011000mid 0 level9Params 
R000100110002 n00010011000mid n00010011000 {level9R}
R000100110011 n0001001100 n00010011001mid {level9R}
yneuron neuron00010011001 n00010011001mid 0 level9Params 
R000100110012 n00010011001mid n00010011001 {level9R}
R00010011011 n000100110 n0001001101mid {level8R}
yneuron neuron0001001101 n0001001101mid 0 level8Params 
R00010011012 n0001001101mid n0001001101 {level8R}
R000100110101 n0001001101 n00010011010mid {level9R}
yneuron neuron00010011010 n00010011010mid 0 level9Params 
R000100110102 n00010011010mid n00010011010 {level9R}
R000100110111 n0001001101 n00010011011mid {level9R}
yneuron neuron00010011011 n00010011011mid 0 level9Params 
R000100110112 n00010011011mid n00010011011 {level9R}
R0001001111 n00010011 n000100111mid {level7R}
yneuron neuron000100111 n000100111mid 0 level7Params 
R0001001112 n000100111mid n000100111 {level7R}
R00010011101 n000100111 n0001001110mid {level8R}
yneuron neuron0001001110 n0001001110mid 0 level8Params 
R00010011102 n0001001110mid n0001001110 {level8R}
R000100111001 n0001001110 n00010011100mid {level9R}
yneuron neuron00010011100 n00010011100mid 0 level9Params 
R000100111002 n00010011100mid n00010011100 {level9R}
R000100111011 n0001001110 n00010011101mid {level9R}
yneuron neuron00010011101 n00010011101mid 0 level9Params 
R000100111012 n00010011101mid n00010011101 {level9R}
R00010011111 n000100111 n0001001111mid {level8R}
yneuron neuron0001001111 n0001001111mid 0 level8Params 
R00010011112 n0001001111mid n0001001111 {level8R}
R000100111101 n0001001111 n00010011110mid {level9R}
yneuron neuron00010011110 n00010011110mid 0 level9Params 
R000100111102 n00010011110mid n00010011110 {level9R}
R000100111111 n0001001111 n00010011111mid {level9R}
yneuron neuron00010011111 n00010011111mid 0 level9Params 
R000100111112 n00010011111mid n00010011111 {level9R}
R0001011 n00010 n000101mid {level4R}
yneuron neuron000101 n000101mid 0 level4Params 
R0001012 n000101mid n000101 {level4R}
R00010101 n000101 n0001010mid {level5R}
yneuron neuron0001010 n0001010mid 0 level5Params 
R00010102 n0001010mid n0001010 {level5R}
R000101001 n0001010 n00010100mid {level6R}
yneuron neuron00010100 n00010100mid 0 level6Params 
R000101002 n00010100mid n00010100 {level6R}
R0001010001 n00010100 n000101000mid {level7R}
yneuron neuron000101000 n000101000mid 0 level7Params 
R0001010002 n000101000mid n000101000 {level7R}
R00010100001 n000101000 n0001010000mid {level8R}
yneuron neuron0001010000 n0001010000mid 0 level8Params 
R00010100002 n0001010000mid n0001010000 {level8R}
R000101000001 n0001010000 n00010100000mid {level9R}
yneuron neuron00010100000 n00010100000mid 0 level9Params 
R000101000002 n00010100000mid n00010100000 {level9R}
R000101000011 n0001010000 n00010100001mid {level9R}
yneuron neuron00010100001 n00010100001mid 0 level9Params 
R000101000012 n00010100001mid n00010100001 {level9R}
R00010100011 n000101000 n0001010001mid {level8R}
yneuron neuron0001010001 n0001010001mid 0 level8Params 
R00010100012 n0001010001mid n0001010001 {level8R}
R000101000101 n0001010001 n00010100010mid {level9R}
yneuron neuron00010100010 n00010100010mid 0 level9Params 
R000101000102 n00010100010mid n00010100010 {level9R}
R000101000111 n0001010001 n00010100011mid {level9R}
yneuron neuron00010100011 n00010100011mid 0 level9Params 
R000101000112 n00010100011mid n00010100011 {level9R}
R0001010011 n00010100 n000101001mid {level7R}
yneuron neuron000101001 n000101001mid 0 level7Params 
R0001010012 n000101001mid n000101001 {level7R}
R00010100101 n000101001 n0001010010mid {level8R}
yneuron neuron0001010010 n0001010010mid 0 level8Params 
R00010100102 n0001010010mid n0001010010 {level8R}
R000101001001 n0001010010 n00010100100mid {level9R}
yneuron neuron00010100100 n00010100100mid 0 level9Params 
R000101001002 n00010100100mid n00010100100 {level9R}
R000101001011 n0001010010 n00010100101mid {level9R}
yneuron neuron00010100101 n00010100101mid 0 level9Params 
R000101001012 n00010100101mid n00010100101 {level9R}
R00010100111 n000101001 n0001010011mid {level8R}
yneuron neuron0001010011 n0001010011mid 0 level8Params 
R00010100112 n0001010011mid n0001010011 {level8R}
R000101001101 n0001010011 n00010100110mid {level9R}
yneuron neuron00010100110 n00010100110mid 0 level9Params 
R000101001102 n00010100110mid n00010100110 {level9R}
R000101001111 n0001010011 n00010100111mid {level9R}
yneuron neuron00010100111 n00010100111mid 0 level9Params 
R000101001112 n00010100111mid n00010100111 {level9R}
R000101011 n0001010 n00010101mid {level6R}
yneuron neuron00010101 n00010101mid 0 level6Params 
R000101012 n00010101mid n00010101 {level6R}
R0001010101 n00010101 n000101010mid {level7R}
yneuron neuron000101010 n000101010mid 0 level7Params 
R0001010102 n000101010mid n000101010 {level7R}
R00010101001 n000101010 n0001010100mid {level8R}
yneuron neuron0001010100 n0001010100mid 0 level8Params 
R00010101002 n0001010100mid n0001010100 {level8R}
R000101010001 n0001010100 n00010101000mid {level9R}
yneuron neuron00010101000 n00010101000mid 0 level9Params 
R000101010002 n00010101000mid n00010101000 {level9R}
R000101010011 n0001010100 n00010101001mid {level9R}
yneuron neuron00010101001 n00010101001mid 0 level9Params 
R000101010012 n00010101001mid n00010101001 {level9R}
R00010101011 n000101010 n0001010101mid {level8R}
yneuron neuron0001010101 n0001010101mid 0 level8Params 
R00010101012 n0001010101mid n0001010101 {level8R}
R000101010101 n0001010101 n00010101010mid {level9R}
yneuron neuron00010101010 n00010101010mid 0 level9Params 
R000101010102 n00010101010mid n00010101010 {level9R}
R000101010111 n0001010101 n00010101011mid {level9R}
yneuron neuron00010101011 n00010101011mid 0 level9Params 
R000101010112 n00010101011mid n00010101011 {level9R}
R0001010111 n00010101 n000101011mid {level7R}
yneuron neuron000101011 n000101011mid 0 level7Params 
R0001010112 n000101011mid n000101011 {level7R}
R00010101101 n000101011 n0001010110mid {level8R}
yneuron neuron0001010110 n0001010110mid 0 level8Params 
R00010101102 n0001010110mid n0001010110 {level8R}
R000101011001 n0001010110 n00010101100mid {level9R}
yneuron neuron00010101100 n00010101100mid 0 level9Params 
R000101011002 n00010101100mid n00010101100 {level9R}
R000101011011 n0001010110 n00010101101mid {level9R}
yneuron neuron00010101101 n00010101101mid 0 level9Params 
R000101011012 n00010101101mid n00010101101 {level9R}
R00010101111 n000101011 n0001010111mid {level8R}
yneuron neuron0001010111 n0001010111mid 0 level8Params 
R00010101112 n0001010111mid n0001010111 {level8R}
R000101011101 n0001010111 n00010101110mid {level9R}
yneuron neuron00010101110 n00010101110mid 0 level9Params 
R000101011102 n00010101110mid n00010101110 {level9R}
R000101011111 n0001010111 n00010101111mid {level9R}
yneuron neuron00010101111 n00010101111mid 0 level9Params 
R000101011112 n00010101111mid n00010101111 {level9R}
R00010111 n000101 n0001011mid {level5R}
yneuron neuron0001011 n0001011mid 0 level5Params 
R00010112 n0001011mid n0001011 {level5R}
R000101101 n0001011 n00010110mid {level6R}
yneuron neuron00010110 n00010110mid 0 level6Params 
R000101102 n00010110mid n00010110 {level6R}
R0001011001 n00010110 n000101100mid {level7R}
yneuron neuron000101100 n000101100mid 0 level7Params 
R0001011002 n000101100mid n000101100 {level7R}
R00010110001 n000101100 n0001011000mid {level8R}
yneuron neuron0001011000 n0001011000mid 0 level8Params 
R00010110002 n0001011000mid n0001011000 {level8R}
R000101100001 n0001011000 n00010110000mid {level9R}
yneuron neuron00010110000 n00010110000mid 0 level9Params 
R000101100002 n00010110000mid n00010110000 {level9R}
R000101100011 n0001011000 n00010110001mid {level9R}
yneuron neuron00010110001 n00010110001mid 0 level9Params 
R000101100012 n00010110001mid n00010110001 {level9R}
R00010110011 n000101100 n0001011001mid {level8R}
yneuron neuron0001011001 n0001011001mid 0 level8Params 
R00010110012 n0001011001mid n0001011001 {level8R}
R000101100101 n0001011001 n00010110010mid {level9R}
yneuron neuron00010110010 n00010110010mid 0 level9Params 
R000101100102 n00010110010mid n00010110010 {level9R}
R000101100111 n0001011001 n00010110011mid {level9R}
yneuron neuron00010110011 n00010110011mid 0 level9Params 
R000101100112 n00010110011mid n00010110011 {level9R}
R0001011011 n00010110 n000101101mid {level7R}
yneuron neuron000101101 n000101101mid 0 level7Params 
R0001011012 n000101101mid n000101101 {level7R}
R00010110101 n000101101 n0001011010mid {level8R}
yneuron neuron0001011010 n0001011010mid 0 level8Params 
R00010110102 n0001011010mid n0001011010 {level8R}
R000101101001 n0001011010 n00010110100mid {level9R}
yneuron neuron00010110100 n00010110100mid 0 level9Params 
R000101101002 n00010110100mid n00010110100 {level9R}
R000101101011 n0001011010 n00010110101mid {level9R}
yneuron neuron00010110101 n00010110101mid 0 level9Params 
R000101101012 n00010110101mid n00010110101 {level9R}
R00010110111 n000101101 n0001011011mid {level8R}
yneuron neuron0001011011 n0001011011mid 0 level8Params 
R00010110112 n0001011011mid n0001011011 {level8R}
R000101101101 n0001011011 n00010110110mid {level9R}
yneuron neuron00010110110 n00010110110mid 0 level9Params 
R000101101102 n00010110110mid n00010110110 {level9R}
R000101101111 n0001011011 n00010110111mid {level9R}
yneuron neuron00010110111 n00010110111mid 0 level9Params 
R000101101112 n00010110111mid n00010110111 {level9R}
R000101111 n0001011 n00010111mid {level6R}
yneuron neuron00010111 n00010111mid 0 level6Params 
R000101112 n00010111mid n00010111 {level6R}
R0001011101 n00010111 n000101110mid {level7R}
yneuron neuron000101110 n000101110mid 0 level7Params 
R0001011102 n000101110mid n000101110 {level7R}
R00010111001 n000101110 n0001011100mid {level8R}
yneuron neuron0001011100 n0001011100mid 0 level8Params 
R00010111002 n0001011100mid n0001011100 {level8R}
R000101110001 n0001011100 n00010111000mid {level9R}
yneuron neuron00010111000 n00010111000mid 0 level9Params 
R000101110002 n00010111000mid n00010111000 {level9R}
R000101110011 n0001011100 n00010111001mid {level9R}
yneuron neuron00010111001 n00010111001mid 0 level9Params 
R000101110012 n00010111001mid n00010111001 {level9R}
R00010111011 n000101110 n0001011101mid {level8R}
yneuron neuron0001011101 n0001011101mid 0 level8Params 
R00010111012 n0001011101mid n0001011101 {level8R}
R000101110101 n0001011101 n00010111010mid {level9R}
yneuron neuron00010111010 n00010111010mid 0 level9Params 
R000101110102 n00010111010mid n00010111010 {level9R}
R000101110111 n0001011101 n00010111011mid {level9R}
yneuron neuron00010111011 n00010111011mid 0 level9Params 
R000101110112 n00010111011mid n00010111011 {level9R}
R0001011111 n00010111 n000101111mid {level7R}
yneuron neuron000101111 n000101111mid 0 level7Params 
R0001011112 n000101111mid n000101111 {level7R}
R00010111101 n000101111 n0001011110mid {level8R}
yneuron neuron0001011110 n0001011110mid 0 level8Params 
R00010111102 n0001011110mid n0001011110 {level8R}
R000101111001 n0001011110 n00010111100mid {level9R}
yneuron neuron00010111100 n00010111100mid 0 level9Params 
R000101111002 n00010111100mid n00010111100 {level9R}
R000101111011 n0001011110 n00010111101mid {level9R}
yneuron neuron00010111101 n00010111101mid 0 level9Params 
R000101111012 n00010111101mid n00010111101 {level9R}
R00010111111 n000101111 n0001011111mid {level8R}
yneuron neuron0001011111 n0001011111mid 0 level8Params 
R00010111112 n0001011111mid n0001011111 {level8R}
R000101111101 n0001011111 n00010111110mid {level9R}
yneuron neuron00010111110 n00010111110mid 0 level9Params 
R000101111102 n00010111110mid n00010111110 {level9R}
R000101111111 n0001011111 n00010111111mid {level9R}
yneuron neuron00010111111 n00010111111mid 0 level9Params 
R000101111112 n00010111111mid n00010111111 {level9R}
R000111 n0001 n00011mid {level3R}
yneuron neuron00011 n00011mid 0 level3Params 
R000112 n00011mid n00011 {level3R}
R0001101 n00011 n000110mid {level4R}
yneuron neuron000110 n000110mid 0 level4Params 
R0001102 n000110mid n000110 {level4R}
R00011001 n000110 n0001100mid {level5R}
yneuron neuron0001100 n0001100mid 0 level5Params 
R00011002 n0001100mid n0001100 {level5R}
R000110001 n0001100 n00011000mid {level6R}
yneuron neuron00011000 n00011000mid 0 level6Params 
R000110002 n00011000mid n00011000 {level6R}
R0001100001 n00011000 n000110000mid {level7R}
yneuron neuron000110000 n000110000mid 0 level7Params 
R0001100002 n000110000mid n000110000 {level7R}
R00011000001 n000110000 n0001100000mid {level8R}
yneuron neuron0001100000 n0001100000mid 0 level8Params 
R00011000002 n0001100000mid n0001100000 {level8R}
R000110000001 n0001100000 n00011000000mid {level9R}
yneuron neuron00011000000 n00011000000mid 0 level9Params 
R000110000002 n00011000000mid n00011000000 {level9R}
R000110000011 n0001100000 n00011000001mid {level9R}
yneuron neuron00011000001 n00011000001mid 0 level9Params 
R000110000012 n00011000001mid n00011000001 {level9R}
R00011000011 n000110000 n0001100001mid {level8R}
yneuron neuron0001100001 n0001100001mid 0 level8Params 
R00011000012 n0001100001mid n0001100001 {level8R}
R000110000101 n0001100001 n00011000010mid {level9R}
yneuron neuron00011000010 n00011000010mid 0 level9Params 
R000110000102 n00011000010mid n00011000010 {level9R}
R000110000111 n0001100001 n00011000011mid {level9R}
yneuron neuron00011000011 n00011000011mid 0 level9Params 
R000110000112 n00011000011mid n00011000011 {level9R}
R0001100011 n00011000 n000110001mid {level7R}
yneuron neuron000110001 n000110001mid 0 level7Params 
R0001100012 n000110001mid n000110001 {level7R}
R00011000101 n000110001 n0001100010mid {level8R}
yneuron neuron0001100010 n0001100010mid 0 level8Params 
R00011000102 n0001100010mid n0001100010 {level8R}
R000110001001 n0001100010 n00011000100mid {level9R}
yneuron neuron00011000100 n00011000100mid 0 level9Params 
R000110001002 n00011000100mid n00011000100 {level9R}
R000110001011 n0001100010 n00011000101mid {level9R}
yneuron neuron00011000101 n00011000101mid 0 level9Params 
R000110001012 n00011000101mid n00011000101 {level9R}
R00011000111 n000110001 n0001100011mid {level8R}
yneuron neuron0001100011 n0001100011mid 0 level8Params 
R00011000112 n0001100011mid n0001100011 {level8R}
R000110001101 n0001100011 n00011000110mid {level9R}
yneuron neuron00011000110 n00011000110mid 0 level9Params 
R000110001102 n00011000110mid n00011000110 {level9R}
R000110001111 n0001100011 n00011000111mid {level9R}
yneuron neuron00011000111 n00011000111mid 0 level9Params 
R000110001112 n00011000111mid n00011000111 {level9R}
R000110011 n0001100 n00011001mid {level6R}
yneuron neuron00011001 n00011001mid 0 level6Params 
R000110012 n00011001mid n00011001 {level6R}
R0001100101 n00011001 n000110010mid {level7R}
yneuron neuron000110010 n000110010mid 0 level7Params 
R0001100102 n000110010mid n000110010 {level7R}
R00011001001 n000110010 n0001100100mid {level8R}
yneuron neuron0001100100 n0001100100mid 0 level8Params 
R00011001002 n0001100100mid n0001100100 {level8R}
R000110010001 n0001100100 n00011001000mid {level9R}
yneuron neuron00011001000 n00011001000mid 0 level9Params 
R000110010002 n00011001000mid n00011001000 {level9R}
R000110010011 n0001100100 n00011001001mid {level9R}
yneuron neuron00011001001 n00011001001mid 0 level9Params 
R000110010012 n00011001001mid n00011001001 {level9R}
R00011001011 n000110010 n0001100101mid {level8R}
yneuron neuron0001100101 n0001100101mid 0 level8Params 
R00011001012 n0001100101mid n0001100101 {level8R}
R000110010101 n0001100101 n00011001010mid {level9R}
yneuron neuron00011001010 n00011001010mid 0 level9Params 
R000110010102 n00011001010mid n00011001010 {level9R}
R000110010111 n0001100101 n00011001011mid {level9R}
yneuron neuron00011001011 n00011001011mid 0 level9Params 
R000110010112 n00011001011mid n00011001011 {level9R}
R0001100111 n00011001 n000110011mid {level7R}
yneuron neuron000110011 n000110011mid 0 level7Params 
R0001100112 n000110011mid n000110011 {level7R}
R00011001101 n000110011 n0001100110mid {level8R}
yneuron neuron0001100110 n0001100110mid 0 level8Params 
R00011001102 n0001100110mid n0001100110 {level8R}
R000110011001 n0001100110 n00011001100mid {level9R}
yneuron neuron00011001100 n00011001100mid 0 level9Params 
R000110011002 n00011001100mid n00011001100 {level9R}
R000110011011 n0001100110 n00011001101mid {level9R}
yneuron neuron00011001101 n00011001101mid 0 level9Params 
R000110011012 n00011001101mid n00011001101 {level9R}
R00011001111 n000110011 n0001100111mid {level8R}
yneuron neuron0001100111 n0001100111mid 0 level8Params 
R00011001112 n0001100111mid n0001100111 {level8R}
R000110011101 n0001100111 n00011001110mid {level9R}
yneuron neuron00011001110 n00011001110mid 0 level9Params 
R000110011102 n00011001110mid n00011001110 {level9R}
R000110011111 n0001100111 n00011001111mid {level9R}
yneuron neuron00011001111 n00011001111mid 0 level9Params 
R000110011112 n00011001111mid n00011001111 {level9R}
R00011011 n000110 n0001101mid {level5R}
yneuron neuron0001101 n0001101mid 0 level5Params 
R00011012 n0001101mid n0001101 {level5R}
R000110101 n0001101 n00011010mid {level6R}
yneuron neuron00011010 n00011010mid 0 level6Params 
R000110102 n00011010mid n00011010 {level6R}
R0001101001 n00011010 n000110100mid {level7R}
yneuron neuron000110100 n000110100mid 0 level7Params 
R0001101002 n000110100mid n000110100 {level7R}
R00011010001 n000110100 n0001101000mid {level8R}
yneuron neuron0001101000 n0001101000mid 0 level8Params 
R00011010002 n0001101000mid n0001101000 {level8R}
R000110100001 n0001101000 n00011010000mid {level9R}
yneuron neuron00011010000 n00011010000mid 0 level9Params 
R000110100002 n00011010000mid n00011010000 {level9R}
R000110100011 n0001101000 n00011010001mid {level9R}
yneuron neuron00011010001 n00011010001mid 0 level9Params 
R000110100012 n00011010001mid n00011010001 {level9R}
R00011010011 n000110100 n0001101001mid {level8R}
yneuron neuron0001101001 n0001101001mid 0 level8Params 
R00011010012 n0001101001mid n0001101001 {level8R}
R000110100101 n0001101001 n00011010010mid {level9R}
yneuron neuron00011010010 n00011010010mid 0 level9Params 
R000110100102 n00011010010mid n00011010010 {level9R}
R000110100111 n0001101001 n00011010011mid {level9R}
yneuron neuron00011010011 n00011010011mid 0 level9Params 
R000110100112 n00011010011mid n00011010011 {level9R}
R0001101011 n00011010 n000110101mid {level7R}
yneuron neuron000110101 n000110101mid 0 level7Params 
R0001101012 n000110101mid n000110101 {level7R}
R00011010101 n000110101 n0001101010mid {level8R}
yneuron neuron0001101010 n0001101010mid 0 level8Params 
R00011010102 n0001101010mid n0001101010 {level8R}
R000110101001 n0001101010 n00011010100mid {level9R}
yneuron neuron00011010100 n00011010100mid 0 level9Params 
R000110101002 n00011010100mid n00011010100 {level9R}
R000110101011 n0001101010 n00011010101mid {level9R}
yneuron neuron00011010101 n00011010101mid 0 level9Params 
R000110101012 n00011010101mid n00011010101 {level9R}
R00011010111 n000110101 n0001101011mid {level8R}
yneuron neuron0001101011 n0001101011mid 0 level8Params 
R00011010112 n0001101011mid n0001101011 {level8R}
R000110101101 n0001101011 n00011010110mid {level9R}
yneuron neuron00011010110 n00011010110mid 0 level9Params 
R000110101102 n00011010110mid n00011010110 {level9R}
R000110101111 n0001101011 n00011010111mid {level9R}
yneuron neuron00011010111 n00011010111mid 0 level9Params 
R000110101112 n00011010111mid n00011010111 {level9R}
R000110111 n0001101 n00011011mid {level6R}
yneuron neuron00011011 n00011011mid 0 level6Params 
R000110112 n00011011mid n00011011 {level6R}
R0001101101 n00011011 n000110110mid {level7R}
yneuron neuron000110110 n000110110mid 0 level7Params 
R0001101102 n000110110mid n000110110 {level7R}
R00011011001 n000110110 n0001101100mid {level8R}
yneuron neuron0001101100 n0001101100mid 0 level8Params 
R00011011002 n0001101100mid n0001101100 {level8R}
R000110110001 n0001101100 n00011011000mid {level9R}
yneuron neuron00011011000 n00011011000mid 0 level9Params 
R000110110002 n00011011000mid n00011011000 {level9R}
R000110110011 n0001101100 n00011011001mid {level9R}
yneuron neuron00011011001 n00011011001mid 0 level9Params 
R000110110012 n00011011001mid n00011011001 {level9R}
R00011011011 n000110110 n0001101101mid {level8R}
yneuron neuron0001101101 n0001101101mid 0 level8Params 
R00011011012 n0001101101mid n0001101101 {level8R}
R000110110101 n0001101101 n00011011010mid {level9R}
yneuron neuron00011011010 n00011011010mid 0 level9Params 
R000110110102 n00011011010mid n00011011010 {level9R}
R000110110111 n0001101101 n00011011011mid {level9R}
yneuron neuron00011011011 n00011011011mid 0 level9Params 
R000110110112 n00011011011mid n00011011011 {level9R}
R0001101111 n00011011 n000110111mid {level7R}
yneuron neuron000110111 n000110111mid 0 level7Params 
R0001101112 n000110111mid n000110111 {level7R}
R00011011101 n000110111 n0001101110mid {level8R}
yneuron neuron0001101110 n0001101110mid 0 level8Params 
R00011011102 n0001101110mid n0001101110 {level8R}
R000110111001 n0001101110 n00011011100mid {level9R}
yneuron neuron00011011100 n00011011100mid 0 level9Params 
R000110111002 n00011011100mid n00011011100 {level9R}
R000110111011 n0001101110 n00011011101mid {level9R}
yneuron neuron00011011101 n00011011101mid 0 level9Params 
R000110111012 n00011011101mid n00011011101 {level9R}
R00011011111 n000110111 n0001101111mid {level8R}
yneuron neuron0001101111 n0001101111mid 0 level8Params 
R00011011112 n0001101111mid n0001101111 {level8R}
R000110111101 n0001101111 n00011011110mid {level9R}
yneuron neuron00011011110 n00011011110mid 0 level9Params 
R000110111102 n00011011110mid n00011011110 {level9R}
R000110111111 n0001101111 n00011011111mid {level9R}
yneuron neuron00011011111 n00011011111mid 0 level9Params 
R000110111112 n00011011111mid n00011011111 {level9R}
R0001111 n00011 n000111mid {level4R}
yneuron neuron000111 n000111mid 0 level4Params 
R0001112 n000111mid n000111 {level4R}
R00011101 n000111 n0001110mid {level5R}
yneuron neuron0001110 n0001110mid 0 level5Params 
R00011102 n0001110mid n0001110 {level5R}
R000111001 n0001110 n00011100mid {level6R}
yneuron neuron00011100 n00011100mid 0 level6Params 
R000111002 n00011100mid n00011100 {level6R}
R0001110001 n00011100 n000111000mid {level7R}
yneuron neuron000111000 n000111000mid 0 level7Params 
R0001110002 n000111000mid n000111000 {level7R}
R00011100001 n000111000 n0001110000mid {level8R}
yneuron neuron0001110000 n0001110000mid 0 level8Params 
R00011100002 n0001110000mid n0001110000 {level8R}
R000111000001 n0001110000 n00011100000mid {level9R}
yneuron neuron00011100000 n00011100000mid 0 level9Params 
R000111000002 n00011100000mid n00011100000 {level9R}
R000111000011 n0001110000 n00011100001mid {level9R}
yneuron neuron00011100001 n00011100001mid 0 level9Params 
R000111000012 n00011100001mid n00011100001 {level9R}
R00011100011 n000111000 n0001110001mid {level8R}
yneuron neuron0001110001 n0001110001mid 0 level8Params 
R00011100012 n0001110001mid n0001110001 {level8R}
R000111000101 n0001110001 n00011100010mid {level9R}
yneuron neuron00011100010 n00011100010mid 0 level9Params 
R000111000102 n00011100010mid n00011100010 {level9R}
R000111000111 n0001110001 n00011100011mid {level9R}
yneuron neuron00011100011 n00011100011mid 0 level9Params 
R000111000112 n00011100011mid n00011100011 {level9R}
R0001110011 n00011100 n000111001mid {level7R}
yneuron neuron000111001 n000111001mid 0 level7Params 
R0001110012 n000111001mid n000111001 {level7R}
R00011100101 n000111001 n0001110010mid {level8R}
yneuron neuron0001110010 n0001110010mid 0 level8Params 
R00011100102 n0001110010mid n0001110010 {level8R}
R000111001001 n0001110010 n00011100100mid {level9R}
yneuron neuron00011100100 n00011100100mid 0 level9Params 
R000111001002 n00011100100mid n00011100100 {level9R}
R000111001011 n0001110010 n00011100101mid {level9R}
yneuron neuron00011100101 n00011100101mid 0 level9Params 
R000111001012 n00011100101mid n00011100101 {level9R}
R00011100111 n000111001 n0001110011mid {level8R}
yneuron neuron0001110011 n0001110011mid 0 level8Params 
R00011100112 n0001110011mid n0001110011 {level8R}
R000111001101 n0001110011 n00011100110mid {level9R}
yneuron neuron00011100110 n00011100110mid 0 level9Params 
R000111001102 n00011100110mid n00011100110 {level9R}
R000111001111 n0001110011 n00011100111mid {level9R}
yneuron neuron00011100111 n00011100111mid 0 level9Params 
R000111001112 n00011100111mid n00011100111 {level9R}
R000111011 n0001110 n00011101mid {level6R}
yneuron neuron00011101 n00011101mid 0 level6Params 
R000111012 n00011101mid n00011101 {level6R}
R0001110101 n00011101 n000111010mid {level7R}
yneuron neuron000111010 n000111010mid 0 level7Params 
R0001110102 n000111010mid n000111010 {level7R}
R00011101001 n000111010 n0001110100mid {level8R}
yneuron neuron0001110100 n0001110100mid 0 level8Params 
R00011101002 n0001110100mid n0001110100 {level8R}
R000111010001 n0001110100 n00011101000mid {level9R}
yneuron neuron00011101000 n00011101000mid 0 level9Params 
R000111010002 n00011101000mid n00011101000 {level9R}
R000111010011 n0001110100 n00011101001mid {level9R}
yneuron neuron00011101001 n00011101001mid 0 level9Params 
R000111010012 n00011101001mid n00011101001 {level9R}
R00011101011 n000111010 n0001110101mid {level8R}
yneuron neuron0001110101 n0001110101mid 0 level8Params 
R00011101012 n0001110101mid n0001110101 {level8R}
R000111010101 n0001110101 n00011101010mid {level9R}
yneuron neuron00011101010 n00011101010mid 0 level9Params 
R000111010102 n00011101010mid n00011101010 {level9R}
R000111010111 n0001110101 n00011101011mid {level9R}
yneuron neuron00011101011 n00011101011mid 0 level9Params 
R000111010112 n00011101011mid n00011101011 {level9R}
R0001110111 n00011101 n000111011mid {level7R}
yneuron neuron000111011 n000111011mid 0 level7Params 
R0001110112 n000111011mid n000111011 {level7R}
R00011101101 n000111011 n0001110110mid {level8R}
yneuron neuron0001110110 n0001110110mid 0 level8Params 
R00011101102 n0001110110mid n0001110110 {level8R}
R000111011001 n0001110110 n00011101100mid {level9R}
yneuron neuron00011101100 n00011101100mid 0 level9Params 
R000111011002 n00011101100mid n00011101100 {level9R}
R000111011011 n0001110110 n00011101101mid {level9R}
yneuron neuron00011101101 n00011101101mid 0 level9Params 
R000111011012 n00011101101mid n00011101101 {level9R}
R00011101111 n000111011 n0001110111mid {level8R}
yneuron neuron0001110111 n0001110111mid 0 level8Params 
R00011101112 n0001110111mid n0001110111 {level8R}
R000111011101 n0001110111 n00011101110mid {level9R}
yneuron neuron00011101110 n00011101110mid 0 level9Params 
R000111011102 n00011101110mid n00011101110 {level9R}
R000111011111 n0001110111 n00011101111mid {level9R}
yneuron neuron00011101111 n00011101111mid 0 level9Params 
R000111011112 n00011101111mid n00011101111 {level9R}
R00011111 n000111 n0001111mid {level5R}
yneuron neuron0001111 n0001111mid 0 level5Params 
R00011112 n0001111mid n0001111 {level5R}
R000111101 n0001111 n00011110mid {level6R}
yneuron neuron00011110 n00011110mid 0 level6Params 
R000111102 n00011110mid n00011110 {level6R}
R0001111001 n00011110 n000111100mid {level7R}
yneuron neuron000111100 n000111100mid 0 level7Params 
R0001111002 n000111100mid n000111100 {level7R}
R00011110001 n000111100 n0001111000mid {level8R}
yneuron neuron0001111000 n0001111000mid 0 level8Params 
R00011110002 n0001111000mid n0001111000 {level8R}
R000111100001 n0001111000 n00011110000mid {level9R}
yneuron neuron00011110000 n00011110000mid 0 level9Params 
R000111100002 n00011110000mid n00011110000 {level9R}
R000111100011 n0001111000 n00011110001mid {level9R}
yneuron neuron00011110001 n00011110001mid 0 level9Params 
R000111100012 n00011110001mid n00011110001 {level9R}
R00011110011 n000111100 n0001111001mid {level8R}
yneuron neuron0001111001 n0001111001mid 0 level8Params 
R00011110012 n0001111001mid n0001111001 {level8R}
R000111100101 n0001111001 n00011110010mid {level9R}
yneuron neuron00011110010 n00011110010mid 0 level9Params 
R000111100102 n00011110010mid n00011110010 {level9R}
R000111100111 n0001111001 n00011110011mid {level9R}
yneuron neuron00011110011 n00011110011mid 0 level9Params 
R000111100112 n00011110011mid n00011110011 {level9R}
R0001111011 n00011110 n000111101mid {level7R}
yneuron neuron000111101 n000111101mid 0 level7Params 
R0001111012 n000111101mid n000111101 {level7R}
R00011110101 n000111101 n0001111010mid {level8R}
yneuron neuron0001111010 n0001111010mid 0 level8Params 
R00011110102 n0001111010mid n0001111010 {level8R}
R000111101001 n0001111010 n00011110100mid {level9R}
yneuron neuron00011110100 n00011110100mid 0 level9Params 
R000111101002 n00011110100mid n00011110100 {level9R}
R000111101011 n0001111010 n00011110101mid {level9R}
yneuron neuron00011110101 n00011110101mid 0 level9Params 
R000111101012 n00011110101mid n00011110101 {level9R}
R00011110111 n000111101 n0001111011mid {level8R}
yneuron neuron0001111011 n0001111011mid 0 level8Params 
R00011110112 n0001111011mid n0001111011 {level8R}
R000111101101 n0001111011 n00011110110mid {level9R}
yneuron neuron00011110110 n00011110110mid 0 level9Params 
R000111101102 n00011110110mid n00011110110 {level9R}
R000111101111 n0001111011 n00011110111mid {level9R}
yneuron neuron00011110111 n00011110111mid 0 level9Params 
R000111101112 n00011110111mid n00011110111 {level9R}
R000111111 n0001111 n00011111mid {level6R}
yneuron neuron00011111 n00011111mid 0 level6Params 
R000111112 n00011111mid n00011111 {level6R}
R0001111101 n00011111 n000111110mid {level7R}
yneuron neuron000111110 n000111110mid 0 level7Params 
R0001111102 n000111110mid n000111110 {level7R}
R00011111001 n000111110 n0001111100mid {level8R}
yneuron neuron0001111100 n0001111100mid 0 level8Params 
R00011111002 n0001111100mid n0001111100 {level8R}
R000111110001 n0001111100 n00011111000mid {level9R}
yneuron neuron00011111000 n00011111000mid 0 level9Params 
R000111110002 n00011111000mid n00011111000 {level9R}
R000111110011 n0001111100 n00011111001mid {level9R}
yneuron neuron00011111001 n00011111001mid 0 level9Params 
R000111110012 n00011111001mid n00011111001 {level9R}
R00011111011 n000111110 n0001111101mid {level8R}
yneuron neuron0001111101 n0001111101mid 0 level8Params 
R00011111012 n0001111101mid n0001111101 {level8R}
R000111110101 n0001111101 n00011111010mid {level9R}
yneuron neuron00011111010 n00011111010mid 0 level9Params 
R000111110102 n00011111010mid n00011111010 {level9R}
R000111110111 n0001111101 n00011111011mid {level9R}
yneuron neuron00011111011 n00011111011mid 0 level9Params 
R000111110112 n00011111011mid n00011111011 {level9R}
R0001111111 n00011111 n000111111mid {level7R}
yneuron neuron000111111 n000111111mid 0 level7Params 
R0001111112 n000111111mid n000111111 {level7R}
R00011111101 n000111111 n0001111110mid {level8R}
yneuron neuron0001111110 n0001111110mid 0 level8Params 
R00011111102 n0001111110mid n0001111110 {level8R}
R000111111001 n0001111110 n00011111100mid {level9R}
yneuron neuron00011111100 n00011111100mid 0 level9Params 
R000111111002 n00011111100mid n00011111100 {level9R}
R000111111011 n0001111110 n00011111101mid {level9R}
yneuron neuron00011111101 n00011111101mid 0 level9Params 
R000111111012 n00011111101mid n00011111101 {level9R}
R00011111111 n000111111 n0001111111mid {level8R}
yneuron neuron0001111111 n0001111111mid 0 level8Params 
R00011111112 n0001111111mid n0001111111 {level8R}
R000111111101 n0001111111 n00011111110mid {level9R}
yneuron neuron00011111110 n00011111110mid 0 level9Params 
R000111111102 n00011111110mid n00011111110 {level9R}
R000111111111 n0001111111 n00011111111mid {level9R}
yneuron neuron00011111111 n00011111111mid 0 level9Params 
R000111111112 n00011111111mid n00011111111 {level9R}
R0011 n00 n001mid {level1R}
yneuron neuron001 n001mid 0 level1Params 
R0012 n001mid n001 {level1R}
R00101 n001 n0010mid {level2R}
yneuron neuron0010 n0010mid 0 level2Params 
R00102 n0010mid n0010 {level2R}
R001001 n0010 n00100mid {level3R}
yneuron neuron00100 n00100mid 0 level3Params 
R001002 n00100mid n00100 {level3R}
R0010001 n00100 n001000mid {level4R}
yneuron neuron001000 n001000mid 0 level4Params 
R0010002 n001000mid n001000 {level4R}
R00100001 n001000 n0010000mid {level5R}
yneuron neuron0010000 n0010000mid 0 level5Params 
R00100002 n0010000mid n0010000 {level5R}
R001000001 n0010000 n00100000mid {level6R}
yneuron neuron00100000 n00100000mid 0 level6Params 
R001000002 n00100000mid n00100000 {level6R}
R0010000001 n00100000 n001000000mid {level7R}
yneuron neuron001000000 n001000000mid 0 level7Params 
R0010000002 n001000000mid n001000000 {level7R}
R00100000001 n001000000 n0010000000mid {level8R}
yneuron neuron0010000000 n0010000000mid 0 level8Params 
R00100000002 n0010000000mid n0010000000 {level8R}
R001000000001 n0010000000 n00100000000mid {level9R}
yneuron neuron00100000000 n00100000000mid 0 level9Params 
R001000000002 n00100000000mid n00100000000 {level9R}
R001000000011 n0010000000 n00100000001mid {level9R}
yneuron neuron00100000001 n00100000001mid 0 level9Params 
R001000000012 n00100000001mid n00100000001 {level9R}
R00100000011 n001000000 n0010000001mid {level8R}
yneuron neuron0010000001 n0010000001mid 0 level8Params 
R00100000012 n0010000001mid n0010000001 {level8R}
R001000000101 n0010000001 n00100000010mid {level9R}
yneuron neuron00100000010 n00100000010mid 0 level9Params 
R001000000102 n00100000010mid n00100000010 {level9R}
R001000000111 n0010000001 n00100000011mid {level9R}
yneuron neuron00100000011 n00100000011mid 0 level9Params 
R001000000112 n00100000011mid n00100000011 {level9R}
R0010000011 n00100000 n001000001mid {level7R}
yneuron neuron001000001 n001000001mid 0 level7Params 
R0010000012 n001000001mid n001000001 {level7R}
R00100000101 n001000001 n0010000010mid {level8R}
yneuron neuron0010000010 n0010000010mid 0 level8Params 
R00100000102 n0010000010mid n0010000010 {level8R}
R001000001001 n0010000010 n00100000100mid {level9R}
yneuron neuron00100000100 n00100000100mid 0 level9Params 
R001000001002 n00100000100mid n00100000100 {level9R}
R001000001011 n0010000010 n00100000101mid {level9R}
yneuron neuron00100000101 n00100000101mid 0 level9Params 
R001000001012 n00100000101mid n00100000101 {level9R}
R00100000111 n001000001 n0010000011mid {level8R}
yneuron neuron0010000011 n0010000011mid 0 level8Params 
R00100000112 n0010000011mid n0010000011 {level8R}
R001000001101 n0010000011 n00100000110mid {level9R}
yneuron neuron00100000110 n00100000110mid 0 level9Params 
R001000001102 n00100000110mid n00100000110 {level9R}
R001000001111 n0010000011 n00100000111mid {level9R}
yneuron neuron00100000111 n00100000111mid 0 level9Params 
R001000001112 n00100000111mid n00100000111 {level9R}
R001000011 n0010000 n00100001mid {level6R}
yneuron neuron00100001 n00100001mid 0 level6Params 
R001000012 n00100001mid n00100001 {level6R}
R0010000101 n00100001 n001000010mid {level7R}
yneuron neuron001000010 n001000010mid 0 level7Params 
R0010000102 n001000010mid n001000010 {level7R}
R00100001001 n001000010 n0010000100mid {level8R}
yneuron neuron0010000100 n0010000100mid 0 level8Params 
R00100001002 n0010000100mid n0010000100 {level8R}
R001000010001 n0010000100 n00100001000mid {level9R}
yneuron neuron00100001000 n00100001000mid 0 level9Params 
R001000010002 n00100001000mid n00100001000 {level9R}
R001000010011 n0010000100 n00100001001mid {level9R}
yneuron neuron00100001001 n00100001001mid 0 level9Params 
R001000010012 n00100001001mid n00100001001 {level9R}
R00100001011 n001000010 n0010000101mid {level8R}
yneuron neuron0010000101 n0010000101mid 0 level8Params 
R00100001012 n0010000101mid n0010000101 {level8R}
R001000010101 n0010000101 n00100001010mid {level9R}
yneuron neuron00100001010 n00100001010mid 0 level9Params 
R001000010102 n00100001010mid n00100001010 {level9R}
R001000010111 n0010000101 n00100001011mid {level9R}
yneuron neuron00100001011 n00100001011mid 0 level9Params 
R001000010112 n00100001011mid n00100001011 {level9R}
R0010000111 n00100001 n001000011mid {level7R}
yneuron neuron001000011 n001000011mid 0 level7Params 
R0010000112 n001000011mid n001000011 {level7R}
R00100001101 n001000011 n0010000110mid {level8R}
yneuron neuron0010000110 n0010000110mid 0 level8Params 
R00100001102 n0010000110mid n0010000110 {level8R}
R001000011001 n0010000110 n00100001100mid {level9R}
yneuron neuron00100001100 n00100001100mid 0 level9Params 
R001000011002 n00100001100mid n00100001100 {level9R}
R001000011011 n0010000110 n00100001101mid {level9R}
yneuron neuron00100001101 n00100001101mid 0 level9Params 
R001000011012 n00100001101mid n00100001101 {level9R}
R00100001111 n001000011 n0010000111mid {level8R}
yneuron neuron0010000111 n0010000111mid 0 level8Params 
R00100001112 n0010000111mid n0010000111 {level8R}
R001000011101 n0010000111 n00100001110mid {level9R}
yneuron neuron00100001110 n00100001110mid 0 level9Params 
R001000011102 n00100001110mid n00100001110 {level9R}
R001000011111 n0010000111 n00100001111mid {level9R}
yneuron neuron00100001111 n00100001111mid 0 level9Params 
R001000011112 n00100001111mid n00100001111 {level9R}
R00100011 n001000 n0010001mid {level5R}
yneuron neuron0010001 n0010001mid 0 level5Params 
R00100012 n0010001mid n0010001 {level5R}
R001000101 n0010001 n00100010mid {level6R}
yneuron neuron00100010 n00100010mid 0 level6Params 
R001000102 n00100010mid n00100010 {level6R}
R0010001001 n00100010 n001000100mid {level7R}
yneuron neuron001000100 n001000100mid 0 level7Params 
R0010001002 n001000100mid n001000100 {level7R}
R00100010001 n001000100 n0010001000mid {level8R}
yneuron neuron0010001000 n0010001000mid 0 level8Params 
R00100010002 n0010001000mid n0010001000 {level8R}
R001000100001 n0010001000 n00100010000mid {level9R}
yneuron neuron00100010000 n00100010000mid 0 level9Params 
R001000100002 n00100010000mid n00100010000 {level9R}
R001000100011 n0010001000 n00100010001mid {level9R}
yneuron neuron00100010001 n00100010001mid 0 level9Params 
R001000100012 n00100010001mid n00100010001 {level9R}
R00100010011 n001000100 n0010001001mid {level8R}
yneuron neuron0010001001 n0010001001mid 0 level8Params 
R00100010012 n0010001001mid n0010001001 {level8R}
R001000100101 n0010001001 n00100010010mid {level9R}
yneuron neuron00100010010 n00100010010mid 0 level9Params 
R001000100102 n00100010010mid n00100010010 {level9R}
R001000100111 n0010001001 n00100010011mid {level9R}
yneuron neuron00100010011 n00100010011mid 0 level9Params 
R001000100112 n00100010011mid n00100010011 {level9R}
R0010001011 n00100010 n001000101mid {level7R}
yneuron neuron001000101 n001000101mid 0 level7Params 
R0010001012 n001000101mid n001000101 {level7R}
R00100010101 n001000101 n0010001010mid {level8R}
yneuron neuron0010001010 n0010001010mid 0 level8Params 
R00100010102 n0010001010mid n0010001010 {level8R}
R001000101001 n0010001010 n00100010100mid {level9R}
yneuron neuron00100010100 n00100010100mid 0 level9Params 
R001000101002 n00100010100mid n00100010100 {level9R}
R001000101011 n0010001010 n00100010101mid {level9R}
yneuron neuron00100010101 n00100010101mid 0 level9Params 
R001000101012 n00100010101mid n00100010101 {level9R}
R00100010111 n001000101 n0010001011mid {level8R}
yneuron neuron0010001011 n0010001011mid 0 level8Params 
R00100010112 n0010001011mid n0010001011 {level8R}
R001000101101 n0010001011 n00100010110mid {level9R}
yneuron neuron00100010110 n00100010110mid 0 level9Params 
R001000101102 n00100010110mid n00100010110 {level9R}
R001000101111 n0010001011 n00100010111mid {level9R}
yneuron neuron00100010111 n00100010111mid 0 level9Params 
R001000101112 n00100010111mid n00100010111 {level9R}
R001000111 n0010001 n00100011mid {level6R}
yneuron neuron00100011 n00100011mid 0 level6Params 
R001000112 n00100011mid n00100011 {level6R}
R0010001101 n00100011 n001000110mid {level7R}
yneuron neuron001000110 n001000110mid 0 level7Params 
R0010001102 n001000110mid n001000110 {level7R}
R00100011001 n001000110 n0010001100mid {level8R}
yneuron neuron0010001100 n0010001100mid 0 level8Params 
R00100011002 n0010001100mid n0010001100 {level8R}
R001000110001 n0010001100 n00100011000mid {level9R}
yneuron neuron00100011000 n00100011000mid 0 level9Params 
R001000110002 n00100011000mid n00100011000 {level9R}
R001000110011 n0010001100 n00100011001mid {level9R}
yneuron neuron00100011001 n00100011001mid 0 level9Params 
R001000110012 n00100011001mid n00100011001 {level9R}
R00100011011 n001000110 n0010001101mid {level8R}
yneuron neuron0010001101 n0010001101mid 0 level8Params 
R00100011012 n0010001101mid n0010001101 {level8R}
R001000110101 n0010001101 n00100011010mid {level9R}
yneuron neuron00100011010 n00100011010mid 0 level9Params 
R001000110102 n00100011010mid n00100011010 {level9R}
R001000110111 n0010001101 n00100011011mid {level9R}
yneuron neuron00100011011 n00100011011mid 0 level9Params 
R001000110112 n00100011011mid n00100011011 {level9R}
R0010001111 n00100011 n001000111mid {level7R}
yneuron neuron001000111 n001000111mid 0 level7Params 
R0010001112 n001000111mid n001000111 {level7R}
R00100011101 n001000111 n0010001110mid {level8R}
yneuron neuron0010001110 n0010001110mid 0 level8Params 
R00100011102 n0010001110mid n0010001110 {level8R}
R001000111001 n0010001110 n00100011100mid {level9R}
yneuron neuron00100011100 n00100011100mid 0 level9Params 
R001000111002 n00100011100mid n00100011100 {level9R}
R001000111011 n0010001110 n00100011101mid {level9R}
yneuron neuron00100011101 n00100011101mid 0 level9Params 
R001000111012 n00100011101mid n00100011101 {level9R}
R00100011111 n001000111 n0010001111mid {level8R}
yneuron neuron0010001111 n0010001111mid 0 level8Params 
R00100011112 n0010001111mid n0010001111 {level8R}
R001000111101 n0010001111 n00100011110mid {level9R}
yneuron neuron00100011110 n00100011110mid 0 level9Params 
R001000111102 n00100011110mid n00100011110 {level9R}
R001000111111 n0010001111 n00100011111mid {level9R}
yneuron neuron00100011111 n00100011111mid 0 level9Params 
R001000111112 n00100011111mid n00100011111 {level9R}
R0010011 n00100 n001001mid {level4R}
yneuron neuron001001 n001001mid 0 level4Params 
R0010012 n001001mid n001001 {level4R}
R00100101 n001001 n0010010mid {level5R}
yneuron neuron0010010 n0010010mid 0 level5Params 
R00100102 n0010010mid n0010010 {level5R}
R001001001 n0010010 n00100100mid {level6R}
yneuron neuron00100100 n00100100mid 0 level6Params 
R001001002 n00100100mid n00100100 {level6R}
R0010010001 n00100100 n001001000mid {level7R}
yneuron neuron001001000 n001001000mid 0 level7Params 
R0010010002 n001001000mid n001001000 {level7R}
R00100100001 n001001000 n0010010000mid {level8R}
yneuron neuron0010010000 n0010010000mid 0 level8Params 
R00100100002 n0010010000mid n0010010000 {level8R}
R001001000001 n0010010000 n00100100000mid {level9R}
yneuron neuron00100100000 n00100100000mid 0 level9Params 
R001001000002 n00100100000mid n00100100000 {level9R}
R001001000011 n0010010000 n00100100001mid {level9R}
yneuron neuron00100100001 n00100100001mid 0 level9Params 
R001001000012 n00100100001mid n00100100001 {level9R}
R00100100011 n001001000 n0010010001mid {level8R}
yneuron neuron0010010001 n0010010001mid 0 level8Params 
R00100100012 n0010010001mid n0010010001 {level8R}
R001001000101 n0010010001 n00100100010mid {level9R}
yneuron neuron00100100010 n00100100010mid 0 level9Params 
R001001000102 n00100100010mid n00100100010 {level9R}
R001001000111 n0010010001 n00100100011mid {level9R}
yneuron neuron00100100011 n00100100011mid 0 level9Params 
R001001000112 n00100100011mid n00100100011 {level9R}
R0010010011 n00100100 n001001001mid {level7R}
yneuron neuron001001001 n001001001mid 0 level7Params 
R0010010012 n001001001mid n001001001 {level7R}
R00100100101 n001001001 n0010010010mid {level8R}
yneuron neuron0010010010 n0010010010mid 0 level8Params 
R00100100102 n0010010010mid n0010010010 {level8R}
R001001001001 n0010010010 n00100100100mid {level9R}
yneuron neuron00100100100 n00100100100mid 0 level9Params 
R001001001002 n00100100100mid n00100100100 {level9R}
R001001001011 n0010010010 n00100100101mid {level9R}
yneuron neuron00100100101 n00100100101mid 0 level9Params 
R001001001012 n00100100101mid n00100100101 {level9R}
R00100100111 n001001001 n0010010011mid {level8R}
yneuron neuron0010010011 n0010010011mid 0 level8Params 
R00100100112 n0010010011mid n0010010011 {level8R}
R001001001101 n0010010011 n00100100110mid {level9R}
yneuron neuron00100100110 n00100100110mid 0 level9Params 
R001001001102 n00100100110mid n00100100110 {level9R}
R001001001111 n0010010011 n00100100111mid {level9R}
yneuron neuron00100100111 n00100100111mid 0 level9Params 
R001001001112 n00100100111mid n00100100111 {level9R}
R001001011 n0010010 n00100101mid {level6R}
yneuron neuron00100101 n00100101mid 0 level6Params 
R001001012 n00100101mid n00100101 {level6R}
R0010010101 n00100101 n001001010mid {level7R}
yneuron neuron001001010 n001001010mid 0 level7Params 
R0010010102 n001001010mid n001001010 {level7R}
R00100101001 n001001010 n0010010100mid {level8R}
yneuron neuron0010010100 n0010010100mid 0 level8Params 
R00100101002 n0010010100mid n0010010100 {level8R}
R001001010001 n0010010100 n00100101000mid {level9R}
yneuron neuron00100101000 n00100101000mid 0 level9Params 
R001001010002 n00100101000mid n00100101000 {level9R}
R001001010011 n0010010100 n00100101001mid {level9R}
yneuron neuron00100101001 n00100101001mid 0 level9Params 
R001001010012 n00100101001mid n00100101001 {level9R}
R00100101011 n001001010 n0010010101mid {level8R}
yneuron neuron0010010101 n0010010101mid 0 level8Params 
R00100101012 n0010010101mid n0010010101 {level8R}
R001001010101 n0010010101 n00100101010mid {level9R}
yneuron neuron00100101010 n00100101010mid 0 level9Params 
R001001010102 n00100101010mid n00100101010 {level9R}
R001001010111 n0010010101 n00100101011mid {level9R}
yneuron neuron00100101011 n00100101011mid 0 level9Params 
R001001010112 n00100101011mid n00100101011 {level9R}
R0010010111 n00100101 n001001011mid {level7R}
yneuron neuron001001011 n001001011mid 0 level7Params 
R0010010112 n001001011mid n001001011 {level7R}
R00100101101 n001001011 n0010010110mid {level8R}
yneuron neuron0010010110 n0010010110mid 0 level8Params 
R00100101102 n0010010110mid n0010010110 {level8R}
R001001011001 n0010010110 n00100101100mid {level9R}
yneuron neuron00100101100 n00100101100mid 0 level9Params 
R001001011002 n00100101100mid n00100101100 {level9R}
R001001011011 n0010010110 n00100101101mid {level9R}
yneuron neuron00100101101 n00100101101mid 0 level9Params 
R001001011012 n00100101101mid n00100101101 {level9R}
R00100101111 n001001011 n0010010111mid {level8R}
yneuron neuron0010010111 n0010010111mid 0 level8Params 
R00100101112 n0010010111mid n0010010111 {level8R}
R001001011101 n0010010111 n00100101110mid {level9R}
yneuron neuron00100101110 n00100101110mid 0 level9Params 
R001001011102 n00100101110mid n00100101110 {level9R}
R001001011111 n0010010111 n00100101111mid {level9R}
yneuron neuron00100101111 n00100101111mid 0 level9Params 
R001001011112 n00100101111mid n00100101111 {level9R}
R00100111 n001001 n0010011mid {level5R}
yneuron neuron0010011 n0010011mid 0 level5Params 
R00100112 n0010011mid n0010011 {level5R}
R001001101 n0010011 n00100110mid {level6R}
yneuron neuron00100110 n00100110mid 0 level6Params 
R001001102 n00100110mid n00100110 {level6R}
R0010011001 n00100110 n001001100mid {level7R}
yneuron neuron001001100 n001001100mid 0 level7Params 
R0010011002 n001001100mid n001001100 {level7R}
R00100110001 n001001100 n0010011000mid {level8R}
yneuron neuron0010011000 n0010011000mid 0 level8Params 
R00100110002 n0010011000mid n0010011000 {level8R}
R001001100001 n0010011000 n00100110000mid {level9R}
yneuron neuron00100110000 n00100110000mid 0 level9Params 
R001001100002 n00100110000mid n00100110000 {level9R}
R001001100011 n0010011000 n00100110001mid {level9R}
yneuron neuron00100110001 n00100110001mid 0 level9Params 
R001001100012 n00100110001mid n00100110001 {level9R}
R00100110011 n001001100 n0010011001mid {level8R}
yneuron neuron0010011001 n0010011001mid 0 level8Params 
R00100110012 n0010011001mid n0010011001 {level8R}
R001001100101 n0010011001 n00100110010mid {level9R}
yneuron neuron00100110010 n00100110010mid 0 level9Params 
R001001100102 n00100110010mid n00100110010 {level9R}
R001001100111 n0010011001 n00100110011mid {level9R}
yneuron neuron00100110011 n00100110011mid 0 level9Params 
R001001100112 n00100110011mid n00100110011 {level9R}
R0010011011 n00100110 n001001101mid {level7R}
yneuron neuron001001101 n001001101mid 0 level7Params 
R0010011012 n001001101mid n001001101 {level7R}
R00100110101 n001001101 n0010011010mid {level8R}
yneuron neuron0010011010 n0010011010mid 0 level8Params 
R00100110102 n0010011010mid n0010011010 {level8R}
R001001101001 n0010011010 n00100110100mid {level9R}
yneuron neuron00100110100 n00100110100mid 0 level9Params 
R001001101002 n00100110100mid n00100110100 {level9R}
R001001101011 n0010011010 n00100110101mid {level9R}
yneuron neuron00100110101 n00100110101mid 0 level9Params 
R001001101012 n00100110101mid n00100110101 {level9R}
R00100110111 n001001101 n0010011011mid {level8R}
yneuron neuron0010011011 n0010011011mid 0 level8Params 
R00100110112 n0010011011mid n0010011011 {level8R}
R001001101101 n0010011011 n00100110110mid {level9R}
yneuron neuron00100110110 n00100110110mid 0 level9Params 
R001001101102 n00100110110mid n00100110110 {level9R}
R001001101111 n0010011011 n00100110111mid {level9R}
yneuron neuron00100110111 n00100110111mid 0 level9Params 
R001001101112 n00100110111mid n00100110111 {level9R}
R001001111 n0010011 n00100111mid {level6R}
yneuron neuron00100111 n00100111mid 0 level6Params 
R001001112 n00100111mid n00100111 {level6R}
R0010011101 n00100111 n001001110mid {level7R}
yneuron neuron001001110 n001001110mid 0 level7Params 
R0010011102 n001001110mid n001001110 {level7R}
R00100111001 n001001110 n0010011100mid {level8R}
yneuron neuron0010011100 n0010011100mid 0 level8Params 
R00100111002 n0010011100mid n0010011100 {level8R}
R001001110001 n0010011100 n00100111000mid {level9R}
yneuron neuron00100111000 n00100111000mid 0 level9Params 
R001001110002 n00100111000mid n00100111000 {level9R}
R001001110011 n0010011100 n00100111001mid {level9R}
yneuron neuron00100111001 n00100111001mid 0 level9Params 
R001001110012 n00100111001mid n00100111001 {level9R}
R00100111011 n001001110 n0010011101mid {level8R}
yneuron neuron0010011101 n0010011101mid 0 level8Params 
R00100111012 n0010011101mid n0010011101 {level8R}
R001001110101 n0010011101 n00100111010mid {level9R}
yneuron neuron00100111010 n00100111010mid 0 level9Params 
R001001110102 n00100111010mid n00100111010 {level9R}
R001001110111 n0010011101 n00100111011mid {level9R}
yneuron neuron00100111011 n00100111011mid 0 level9Params 
R001001110112 n00100111011mid n00100111011 {level9R}
R0010011111 n00100111 n001001111mid {level7R}
yneuron neuron001001111 n001001111mid 0 level7Params 
R0010011112 n001001111mid n001001111 {level7R}
R00100111101 n001001111 n0010011110mid {level8R}
yneuron neuron0010011110 n0010011110mid 0 level8Params 
R00100111102 n0010011110mid n0010011110 {level8R}
R001001111001 n0010011110 n00100111100mid {level9R}
yneuron neuron00100111100 n00100111100mid 0 level9Params 
R001001111002 n00100111100mid n00100111100 {level9R}
R001001111011 n0010011110 n00100111101mid {level9R}
yneuron neuron00100111101 n00100111101mid 0 level9Params 
R001001111012 n00100111101mid n00100111101 {level9R}
R00100111111 n001001111 n0010011111mid {level8R}
yneuron neuron0010011111 n0010011111mid 0 level8Params 
R00100111112 n0010011111mid n0010011111 {level8R}
R001001111101 n0010011111 n00100111110mid {level9R}
yneuron neuron00100111110 n00100111110mid 0 level9Params 
R001001111102 n00100111110mid n00100111110 {level9R}
R001001111111 n0010011111 n00100111111mid {level9R}
yneuron neuron00100111111 n00100111111mid 0 level9Params 
R001001111112 n00100111111mid n00100111111 {level9R}
R001011 n0010 n00101mid {level3R}
yneuron neuron00101 n00101mid 0 level3Params 
R001012 n00101mid n00101 {level3R}
R0010101 n00101 n001010mid {level4R}
yneuron neuron001010 n001010mid 0 level4Params 
R0010102 n001010mid n001010 {level4R}
R00101001 n001010 n0010100mid {level5R}
yneuron neuron0010100 n0010100mid 0 level5Params 
R00101002 n0010100mid n0010100 {level5R}
R001010001 n0010100 n00101000mid {level6R}
yneuron neuron00101000 n00101000mid 0 level6Params 
R001010002 n00101000mid n00101000 {level6R}
R0010100001 n00101000 n001010000mid {level7R}
yneuron neuron001010000 n001010000mid 0 level7Params 
R0010100002 n001010000mid n001010000 {level7R}
R00101000001 n001010000 n0010100000mid {level8R}
yneuron neuron0010100000 n0010100000mid 0 level8Params 
R00101000002 n0010100000mid n0010100000 {level8R}
R001010000001 n0010100000 n00101000000mid {level9R}
yneuron neuron00101000000 n00101000000mid 0 level9Params 
R001010000002 n00101000000mid n00101000000 {level9R}
R001010000011 n0010100000 n00101000001mid {level9R}
yneuron neuron00101000001 n00101000001mid 0 level9Params 
R001010000012 n00101000001mid n00101000001 {level9R}
R00101000011 n001010000 n0010100001mid {level8R}
yneuron neuron0010100001 n0010100001mid 0 level8Params 
R00101000012 n0010100001mid n0010100001 {level8R}
R001010000101 n0010100001 n00101000010mid {level9R}
yneuron neuron00101000010 n00101000010mid 0 level9Params 
R001010000102 n00101000010mid n00101000010 {level9R}
R001010000111 n0010100001 n00101000011mid {level9R}
yneuron neuron00101000011 n00101000011mid 0 level9Params 
R001010000112 n00101000011mid n00101000011 {level9R}
R0010100011 n00101000 n001010001mid {level7R}
yneuron neuron001010001 n001010001mid 0 level7Params 
R0010100012 n001010001mid n001010001 {level7R}
R00101000101 n001010001 n0010100010mid {level8R}
yneuron neuron0010100010 n0010100010mid 0 level8Params 
R00101000102 n0010100010mid n0010100010 {level8R}
R001010001001 n0010100010 n00101000100mid {level9R}
yneuron neuron00101000100 n00101000100mid 0 level9Params 
R001010001002 n00101000100mid n00101000100 {level9R}
R001010001011 n0010100010 n00101000101mid {level9R}
yneuron neuron00101000101 n00101000101mid 0 level9Params 
R001010001012 n00101000101mid n00101000101 {level9R}
R00101000111 n001010001 n0010100011mid {level8R}
yneuron neuron0010100011 n0010100011mid 0 level8Params 
R00101000112 n0010100011mid n0010100011 {level8R}
R001010001101 n0010100011 n00101000110mid {level9R}
yneuron neuron00101000110 n00101000110mid 0 level9Params 
R001010001102 n00101000110mid n00101000110 {level9R}
R001010001111 n0010100011 n00101000111mid {level9R}
yneuron neuron00101000111 n00101000111mid 0 level9Params 
R001010001112 n00101000111mid n00101000111 {level9R}
R001010011 n0010100 n00101001mid {level6R}
yneuron neuron00101001 n00101001mid 0 level6Params 
R001010012 n00101001mid n00101001 {level6R}
R0010100101 n00101001 n001010010mid {level7R}
yneuron neuron001010010 n001010010mid 0 level7Params 
R0010100102 n001010010mid n001010010 {level7R}
R00101001001 n001010010 n0010100100mid {level8R}
yneuron neuron0010100100 n0010100100mid 0 level8Params 
R00101001002 n0010100100mid n0010100100 {level8R}
R001010010001 n0010100100 n00101001000mid {level9R}
yneuron neuron00101001000 n00101001000mid 0 level9Params 
R001010010002 n00101001000mid n00101001000 {level9R}
R001010010011 n0010100100 n00101001001mid {level9R}
yneuron neuron00101001001 n00101001001mid 0 level9Params 
R001010010012 n00101001001mid n00101001001 {level9R}
R00101001011 n001010010 n0010100101mid {level8R}
yneuron neuron0010100101 n0010100101mid 0 level8Params 
R00101001012 n0010100101mid n0010100101 {level8R}
R001010010101 n0010100101 n00101001010mid {level9R}
yneuron neuron00101001010 n00101001010mid 0 level9Params 
R001010010102 n00101001010mid n00101001010 {level9R}
R001010010111 n0010100101 n00101001011mid {level9R}
yneuron neuron00101001011 n00101001011mid 0 level9Params 
R001010010112 n00101001011mid n00101001011 {level9R}
R0010100111 n00101001 n001010011mid {level7R}
yneuron neuron001010011 n001010011mid 0 level7Params 
R0010100112 n001010011mid n001010011 {level7R}
R00101001101 n001010011 n0010100110mid {level8R}
yneuron neuron0010100110 n0010100110mid 0 level8Params 
R00101001102 n0010100110mid n0010100110 {level8R}
R001010011001 n0010100110 n00101001100mid {level9R}
yneuron neuron00101001100 n00101001100mid 0 level9Params 
R001010011002 n00101001100mid n00101001100 {level9R}
R001010011011 n0010100110 n00101001101mid {level9R}
yneuron neuron00101001101 n00101001101mid 0 level9Params 
R001010011012 n00101001101mid n00101001101 {level9R}
R00101001111 n001010011 n0010100111mid {level8R}
yneuron neuron0010100111 n0010100111mid 0 level8Params 
R00101001112 n0010100111mid n0010100111 {level8R}
R001010011101 n0010100111 n00101001110mid {level9R}
yneuron neuron00101001110 n00101001110mid 0 level9Params 
R001010011102 n00101001110mid n00101001110 {level9R}
R001010011111 n0010100111 n00101001111mid {level9R}
yneuron neuron00101001111 n00101001111mid 0 level9Params 
R001010011112 n00101001111mid n00101001111 {level9R}
R00101011 n001010 n0010101mid {level5R}
yneuron neuron0010101 n0010101mid 0 level5Params 
R00101012 n0010101mid n0010101 {level5R}
R001010101 n0010101 n00101010mid {level6R}
yneuron neuron00101010 n00101010mid 0 level6Params 
R001010102 n00101010mid n00101010 {level6R}
R0010101001 n00101010 n001010100mid {level7R}
yneuron neuron001010100 n001010100mid 0 level7Params 
R0010101002 n001010100mid n001010100 {level7R}
R00101010001 n001010100 n0010101000mid {level8R}
yneuron neuron0010101000 n0010101000mid 0 level8Params 
R00101010002 n0010101000mid n0010101000 {level8R}
R001010100001 n0010101000 n00101010000mid {level9R}
yneuron neuron00101010000 n00101010000mid 0 level9Params 
R001010100002 n00101010000mid n00101010000 {level9R}
R001010100011 n0010101000 n00101010001mid {level9R}
yneuron neuron00101010001 n00101010001mid 0 level9Params 
R001010100012 n00101010001mid n00101010001 {level9R}
R00101010011 n001010100 n0010101001mid {level8R}
yneuron neuron0010101001 n0010101001mid 0 level8Params 
R00101010012 n0010101001mid n0010101001 {level8R}
R001010100101 n0010101001 n00101010010mid {level9R}
yneuron neuron00101010010 n00101010010mid 0 level9Params 
R001010100102 n00101010010mid n00101010010 {level9R}
R001010100111 n0010101001 n00101010011mid {level9R}
yneuron neuron00101010011 n00101010011mid 0 level9Params 
R001010100112 n00101010011mid n00101010011 {level9R}
R0010101011 n00101010 n001010101mid {level7R}
yneuron neuron001010101 n001010101mid 0 level7Params 
R0010101012 n001010101mid n001010101 {level7R}
R00101010101 n001010101 n0010101010mid {level8R}
yneuron neuron0010101010 n0010101010mid 0 level8Params 
R00101010102 n0010101010mid n0010101010 {level8R}
R001010101001 n0010101010 n00101010100mid {level9R}
yneuron neuron00101010100 n00101010100mid 0 level9Params 
R001010101002 n00101010100mid n00101010100 {level9R}
R001010101011 n0010101010 n00101010101mid {level9R}
yneuron neuron00101010101 n00101010101mid 0 level9Params 
R001010101012 n00101010101mid n00101010101 {level9R}
R00101010111 n001010101 n0010101011mid {level8R}
yneuron neuron0010101011 n0010101011mid 0 level8Params 
R00101010112 n0010101011mid n0010101011 {level8R}
R001010101101 n0010101011 n00101010110mid {level9R}
yneuron neuron00101010110 n00101010110mid 0 level9Params 
R001010101102 n00101010110mid n00101010110 {level9R}
R001010101111 n0010101011 n00101010111mid {level9R}
yneuron neuron00101010111 n00101010111mid 0 level9Params 
R001010101112 n00101010111mid n00101010111 {level9R}
R001010111 n0010101 n00101011mid {level6R}
yneuron neuron00101011 n00101011mid 0 level6Params 
R001010112 n00101011mid n00101011 {level6R}
R0010101101 n00101011 n001010110mid {level7R}
yneuron neuron001010110 n001010110mid 0 level7Params 
R0010101102 n001010110mid n001010110 {level7R}
R00101011001 n001010110 n0010101100mid {level8R}
yneuron neuron0010101100 n0010101100mid 0 level8Params 
R00101011002 n0010101100mid n0010101100 {level8R}
R001010110001 n0010101100 n00101011000mid {level9R}
yneuron neuron00101011000 n00101011000mid 0 level9Params 
R001010110002 n00101011000mid n00101011000 {level9R}
R001010110011 n0010101100 n00101011001mid {level9R}
yneuron neuron00101011001 n00101011001mid 0 level9Params 
R001010110012 n00101011001mid n00101011001 {level9R}
R00101011011 n001010110 n0010101101mid {level8R}
yneuron neuron0010101101 n0010101101mid 0 level8Params 
R00101011012 n0010101101mid n0010101101 {level8R}
R001010110101 n0010101101 n00101011010mid {level9R}
yneuron neuron00101011010 n00101011010mid 0 level9Params 
R001010110102 n00101011010mid n00101011010 {level9R}
R001010110111 n0010101101 n00101011011mid {level9R}
yneuron neuron00101011011 n00101011011mid 0 level9Params 
R001010110112 n00101011011mid n00101011011 {level9R}
R0010101111 n00101011 n001010111mid {level7R}
yneuron neuron001010111 n001010111mid 0 level7Params 
R0010101112 n001010111mid n001010111 {level7R}
R00101011101 n001010111 n0010101110mid {level8R}
yneuron neuron0010101110 n0010101110mid 0 level8Params 
R00101011102 n0010101110mid n0010101110 {level8R}
R001010111001 n0010101110 n00101011100mid {level9R}
yneuron neuron00101011100 n00101011100mid 0 level9Params 
R001010111002 n00101011100mid n00101011100 {level9R}
R001010111011 n0010101110 n00101011101mid {level9R}
yneuron neuron00101011101 n00101011101mid 0 level9Params 
R001010111012 n00101011101mid n00101011101 {level9R}
R00101011111 n001010111 n0010101111mid {level8R}
yneuron neuron0010101111 n0010101111mid 0 level8Params 
R00101011112 n0010101111mid n0010101111 {level8R}
R001010111101 n0010101111 n00101011110mid {level9R}
yneuron neuron00101011110 n00101011110mid 0 level9Params 
R001010111102 n00101011110mid n00101011110 {level9R}
R001010111111 n0010101111 n00101011111mid {level9R}
yneuron neuron00101011111 n00101011111mid 0 level9Params 
R001010111112 n00101011111mid n00101011111 {level9R}
R0010111 n00101 n001011mid {level4R}
yneuron neuron001011 n001011mid 0 level4Params 
R0010112 n001011mid n001011 {level4R}
R00101101 n001011 n0010110mid {level5R}
yneuron neuron0010110 n0010110mid 0 level5Params 
R00101102 n0010110mid n0010110 {level5R}
R001011001 n0010110 n00101100mid {level6R}
yneuron neuron00101100 n00101100mid 0 level6Params 
R001011002 n00101100mid n00101100 {level6R}
R0010110001 n00101100 n001011000mid {level7R}
yneuron neuron001011000 n001011000mid 0 level7Params 
R0010110002 n001011000mid n001011000 {level7R}
R00101100001 n001011000 n0010110000mid {level8R}
yneuron neuron0010110000 n0010110000mid 0 level8Params 
R00101100002 n0010110000mid n0010110000 {level8R}
R001011000001 n0010110000 n00101100000mid {level9R}
yneuron neuron00101100000 n00101100000mid 0 level9Params 
R001011000002 n00101100000mid n00101100000 {level9R}
R001011000011 n0010110000 n00101100001mid {level9R}
yneuron neuron00101100001 n00101100001mid 0 level9Params 
R001011000012 n00101100001mid n00101100001 {level9R}
R00101100011 n001011000 n0010110001mid {level8R}
yneuron neuron0010110001 n0010110001mid 0 level8Params 
R00101100012 n0010110001mid n0010110001 {level8R}
R001011000101 n0010110001 n00101100010mid {level9R}
yneuron neuron00101100010 n00101100010mid 0 level9Params 
R001011000102 n00101100010mid n00101100010 {level9R}
R001011000111 n0010110001 n00101100011mid {level9R}
yneuron neuron00101100011 n00101100011mid 0 level9Params 
R001011000112 n00101100011mid n00101100011 {level9R}
R0010110011 n00101100 n001011001mid {level7R}
yneuron neuron001011001 n001011001mid 0 level7Params 
R0010110012 n001011001mid n001011001 {level7R}
R00101100101 n001011001 n0010110010mid {level8R}
yneuron neuron0010110010 n0010110010mid 0 level8Params 
R00101100102 n0010110010mid n0010110010 {level8R}
R001011001001 n0010110010 n00101100100mid {level9R}
yneuron neuron00101100100 n00101100100mid 0 level9Params 
R001011001002 n00101100100mid n00101100100 {level9R}
R001011001011 n0010110010 n00101100101mid {level9R}
yneuron neuron00101100101 n00101100101mid 0 level9Params 
R001011001012 n00101100101mid n00101100101 {level9R}
R00101100111 n001011001 n0010110011mid {level8R}
yneuron neuron0010110011 n0010110011mid 0 level8Params 
R00101100112 n0010110011mid n0010110011 {level8R}
R001011001101 n0010110011 n00101100110mid {level9R}
yneuron neuron00101100110 n00101100110mid 0 level9Params 
R001011001102 n00101100110mid n00101100110 {level9R}
R001011001111 n0010110011 n00101100111mid {level9R}
yneuron neuron00101100111 n00101100111mid 0 level9Params 
R001011001112 n00101100111mid n00101100111 {level9R}
R001011011 n0010110 n00101101mid {level6R}
yneuron neuron00101101 n00101101mid 0 level6Params 
R001011012 n00101101mid n00101101 {level6R}
R0010110101 n00101101 n001011010mid {level7R}
yneuron neuron001011010 n001011010mid 0 level7Params 
R0010110102 n001011010mid n001011010 {level7R}
R00101101001 n001011010 n0010110100mid {level8R}
yneuron neuron0010110100 n0010110100mid 0 level8Params 
R00101101002 n0010110100mid n0010110100 {level8R}
R001011010001 n0010110100 n00101101000mid {level9R}
yneuron neuron00101101000 n00101101000mid 0 level9Params 
R001011010002 n00101101000mid n00101101000 {level9R}
R001011010011 n0010110100 n00101101001mid {level9R}
yneuron neuron00101101001 n00101101001mid 0 level9Params 
R001011010012 n00101101001mid n00101101001 {level9R}
R00101101011 n001011010 n0010110101mid {level8R}
yneuron neuron0010110101 n0010110101mid 0 level8Params 
R00101101012 n0010110101mid n0010110101 {level8R}
R001011010101 n0010110101 n00101101010mid {level9R}
yneuron neuron00101101010 n00101101010mid 0 level9Params 
R001011010102 n00101101010mid n00101101010 {level9R}
R001011010111 n0010110101 n00101101011mid {level9R}
yneuron neuron00101101011 n00101101011mid 0 level9Params 
R001011010112 n00101101011mid n00101101011 {level9R}
R0010110111 n00101101 n001011011mid {level7R}
yneuron neuron001011011 n001011011mid 0 level7Params 
R0010110112 n001011011mid n001011011 {level7R}
R00101101101 n001011011 n0010110110mid {level8R}
yneuron neuron0010110110 n0010110110mid 0 level8Params 
R00101101102 n0010110110mid n0010110110 {level8R}
R001011011001 n0010110110 n00101101100mid {level9R}
yneuron neuron00101101100 n00101101100mid 0 level9Params 
R001011011002 n00101101100mid n00101101100 {level9R}
R001011011011 n0010110110 n00101101101mid {level9R}
yneuron neuron00101101101 n00101101101mid 0 level9Params 
R001011011012 n00101101101mid n00101101101 {level9R}
R00101101111 n001011011 n0010110111mid {level8R}
yneuron neuron0010110111 n0010110111mid 0 level8Params 
R00101101112 n0010110111mid n0010110111 {level8R}
R001011011101 n0010110111 n00101101110mid {level9R}
yneuron neuron00101101110 n00101101110mid 0 level9Params 
R001011011102 n00101101110mid n00101101110 {level9R}
R001011011111 n0010110111 n00101101111mid {level9R}
yneuron neuron00101101111 n00101101111mid 0 level9Params 
R001011011112 n00101101111mid n00101101111 {level9R}
R00101111 n001011 n0010111mid {level5R}
yneuron neuron0010111 n0010111mid 0 level5Params 
R00101112 n0010111mid n0010111 {level5R}
R001011101 n0010111 n00101110mid {level6R}
yneuron neuron00101110 n00101110mid 0 level6Params 
R001011102 n00101110mid n00101110 {level6R}
R0010111001 n00101110 n001011100mid {level7R}
yneuron neuron001011100 n001011100mid 0 level7Params 
R0010111002 n001011100mid n001011100 {level7R}
R00101110001 n001011100 n0010111000mid {level8R}
yneuron neuron0010111000 n0010111000mid 0 level8Params 
R00101110002 n0010111000mid n0010111000 {level8R}
R001011100001 n0010111000 n00101110000mid {level9R}
yneuron neuron00101110000 n00101110000mid 0 level9Params 
R001011100002 n00101110000mid n00101110000 {level9R}
R001011100011 n0010111000 n00101110001mid {level9R}
yneuron neuron00101110001 n00101110001mid 0 level9Params 
R001011100012 n00101110001mid n00101110001 {level9R}
R00101110011 n001011100 n0010111001mid {level8R}
yneuron neuron0010111001 n0010111001mid 0 level8Params 
R00101110012 n0010111001mid n0010111001 {level8R}
R001011100101 n0010111001 n00101110010mid {level9R}
yneuron neuron00101110010 n00101110010mid 0 level9Params 
R001011100102 n00101110010mid n00101110010 {level9R}
R001011100111 n0010111001 n00101110011mid {level9R}
yneuron neuron00101110011 n00101110011mid 0 level9Params 
R001011100112 n00101110011mid n00101110011 {level9R}
R0010111011 n00101110 n001011101mid {level7R}
yneuron neuron001011101 n001011101mid 0 level7Params 
R0010111012 n001011101mid n001011101 {level7R}
R00101110101 n001011101 n0010111010mid {level8R}
yneuron neuron0010111010 n0010111010mid 0 level8Params 
R00101110102 n0010111010mid n0010111010 {level8R}
R001011101001 n0010111010 n00101110100mid {level9R}
yneuron neuron00101110100 n00101110100mid 0 level9Params 
R001011101002 n00101110100mid n00101110100 {level9R}
R001011101011 n0010111010 n00101110101mid {level9R}
yneuron neuron00101110101 n00101110101mid 0 level9Params 
R001011101012 n00101110101mid n00101110101 {level9R}
R00101110111 n001011101 n0010111011mid {level8R}
yneuron neuron0010111011 n0010111011mid 0 level8Params 
R00101110112 n0010111011mid n0010111011 {level8R}
R001011101101 n0010111011 n00101110110mid {level9R}
yneuron neuron00101110110 n00101110110mid 0 level9Params 
R001011101102 n00101110110mid n00101110110 {level9R}
R001011101111 n0010111011 n00101110111mid {level9R}
yneuron neuron00101110111 n00101110111mid 0 level9Params 
R001011101112 n00101110111mid n00101110111 {level9R}
R001011111 n0010111 n00101111mid {level6R}
yneuron neuron00101111 n00101111mid 0 level6Params 
R001011112 n00101111mid n00101111 {level6R}
R0010111101 n00101111 n001011110mid {level7R}
yneuron neuron001011110 n001011110mid 0 level7Params 
R0010111102 n001011110mid n001011110 {level7R}
R00101111001 n001011110 n0010111100mid {level8R}
yneuron neuron0010111100 n0010111100mid 0 level8Params 
R00101111002 n0010111100mid n0010111100 {level8R}
R001011110001 n0010111100 n00101111000mid {level9R}
yneuron neuron00101111000 n00101111000mid 0 level9Params 
R001011110002 n00101111000mid n00101111000 {level9R}
R001011110011 n0010111100 n00101111001mid {level9R}
yneuron neuron00101111001 n00101111001mid 0 level9Params 
R001011110012 n00101111001mid n00101111001 {level9R}
R00101111011 n001011110 n0010111101mid {level8R}
yneuron neuron0010111101 n0010111101mid 0 level8Params 
R00101111012 n0010111101mid n0010111101 {level8R}
R001011110101 n0010111101 n00101111010mid {level9R}
yneuron neuron00101111010 n00101111010mid 0 level9Params 
R001011110102 n00101111010mid n00101111010 {level9R}
R001011110111 n0010111101 n00101111011mid {level9R}
yneuron neuron00101111011 n00101111011mid 0 level9Params 
R001011110112 n00101111011mid n00101111011 {level9R}
R0010111111 n00101111 n001011111mid {level7R}
yneuron neuron001011111 n001011111mid 0 level7Params 
R0010111112 n001011111mid n001011111 {level7R}
R00101111101 n001011111 n0010111110mid {level8R}
yneuron neuron0010111110 n0010111110mid 0 level8Params 
R00101111102 n0010111110mid n0010111110 {level8R}
R001011111001 n0010111110 n00101111100mid {level9R}
yneuron neuron00101111100 n00101111100mid 0 level9Params 
R001011111002 n00101111100mid n00101111100 {level9R}
R001011111011 n0010111110 n00101111101mid {level9R}
yneuron neuron00101111101 n00101111101mid 0 level9Params 
R001011111012 n00101111101mid n00101111101 {level9R}
R00101111111 n001011111 n0010111111mid {level8R}
yneuron neuron0010111111 n0010111111mid 0 level8Params 
R00101111112 n0010111111mid n0010111111 {level8R}
R001011111101 n0010111111 n00101111110mid {level9R}
yneuron neuron00101111110 n00101111110mid 0 level9Params 
R001011111102 n00101111110mid n00101111110 {level9R}
R001011111111 n0010111111 n00101111111mid {level9R}
yneuron neuron00101111111 n00101111111mid 0 level9Params 
R001011111112 n00101111111mid n00101111111 {level9R}
R00111 n001 n0011mid {level2R}
yneuron neuron0011 n0011mid 0 level2Params 
R00112 n0011mid n0011 {level2R}
R001101 n0011 n00110mid {level3R}
yneuron neuron00110 n00110mid 0 level3Params 
R001102 n00110mid n00110 {level3R}
R0011001 n00110 n001100mid {level4R}
yneuron neuron001100 n001100mid 0 level4Params 
R0011002 n001100mid n001100 {level4R}
R00110001 n001100 n0011000mid {level5R}
yneuron neuron0011000 n0011000mid 0 level5Params 
R00110002 n0011000mid n0011000 {level5R}
R001100001 n0011000 n00110000mid {level6R}
yneuron neuron00110000 n00110000mid 0 level6Params 
R001100002 n00110000mid n00110000 {level6R}
R0011000001 n00110000 n001100000mid {level7R}
yneuron neuron001100000 n001100000mid 0 level7Params 
R0011000002 n001100000mid n001100000 {level7R}
R00110000001 n001100000 n0011000000mid {level8R}
yneuron neuron0011000000 n0011000000mid 0 level8Params 
R00110000002 n0011000000mid n0011000000 {level8R}
R001100000001 n0011000000 n00110000000mid {level9R}
yneuron neuron00110000000 n00110000000mid 0 level9Params 
R001100000002 n00110000000mid n00110000000 {level9R}
R001100000011 n0011000000 n00110000001mid {level9R}
yneuron neuron00110000001 n00110000001mid 0 level9Params 
R001100000012 n00110000001mid n00110000001 {level9R}
R00110000011 n001100000 n0011000001mid {level8R}
yneuron neuron0011000001 n0011000001mid 0 level8Params 
R00110000012 n0011000001mid n0011000001 {level8R}
R001100000101 n0011000001 n00110000010mid {level9R}
yneuron neuron00110000010 n00110000010mid 0 level9Params 
R001100000102 n00110000010mid n00110000010 {level9R}
R001100000111 n0011000001 n00110000011mid {level9R}
yneuron neuron00110000011 n00110000011mid 0 level9Params 
R001100000112 n00110000011mid n00110000011 {level9R}
R0011000011 n00110000 n001100001mid {level7R}
yneuron neuron001100001 n001100001mid 0 level7Params 
R0011000012 n001100001mid n001100001 {level7R}
R00110000101 n001100001 n0011000010mid {level8R}
yneuron neuron0011000010 n0011000010mid 0 level8Params 
R00110000102 n0011000010mid n0011000010 {level8R}
R001100001001 n0011000010 n00110000100mid {level9R}
yneuron neuron00110000100 n00110000100mid 0 level9Params 
R001100001002 n00110000100mid n00110000100 {level9R}
R001100001011 n0011000010 n00110000101mid {level9R}
yneuron neuron00110000101 n00110000101mid 0 level9Params 
R001100001012 n00110000101mid n00110000101 {level9R}
R00110000111 n001100001 n0011000011mid {level8R}
yneuron neuron0011000011 n0011000011mid 0 level8Params 
R00110000112 n0011000011mid n0011000011 {level8R}
R001100001101 n0011000011 n00110000110mid {level9R}
yneuron neuron00110000110 n00110000110mid 0 level9Params 
R001100001102 n00110000110mid n00110000110 {level9R}
R001100001111 n0011000011 n00110000111mid {level9R}
yneuron neuron00110000111 n00110000111mid 0 level9Params 
R001100001112 n00110000111mid n00110000111 {level9R}
R001100011 n0011000 n00110001mid {level6R}
yneuron neuron00110001 n00110001mid 0 level6Params 
R001100012 n00110001mid n00110001 {level6R}
R0011000101 n00110001 n001100010mid {level7R}
yneuron neuron001100010 n001100010mid 0 level7Params 
R0011000102 n001100010mid n001100010 {level7R}
R00110001001 n001100010 n0011000100mid {level8R}
yneuron neuron0011000100 n0011000100mid 0 level8Params 
R00110001002 n0011000100mid n0011000100 {level8R}
R001100010001 n0011000100 n00110001000mid {level9R}
yneuron neuron00110001000 n00110001000mid 0 level9Params 
R001100010002 n00110001000mid n00110001000 {level9R}
R001100010011 n0011000100 n00110001001mid {level9R}
yneuron neuron00110001001 n00110001001mid 0 level9Params 
R001100010012 n00110001001mid n00110001001 {level9R}
R00110001011 n001100010 n0011000101mid {level8R}
yneuron neuron0011000101 n0011000101mid 0 level8Params 
R00110001012 n0011000101mid n0011000101 {level8R}
R001100010101 n0011000101 n00110001010mid {level9R}
yneuron neuron00110001010 n00110001010mid 0 level9Params 
R001100010102 n00110001010mid n00110001010 {level9R}
R001100010111 n0011000101 n00110001011mid {level9R}
yneuron neuron00110001011 n00110001011mid 0 level9Params 
R001100010112 n00110001011mid n00110001011 {level9R}
R0011000111 n00110001 n001100011mid {level7R}
yneuron neuron001100011 n001100011mid 0 level7Params 
R0011000112 n001100011mid n001100011 {level7R}
R00110001101 n001100011 n0011000110mid {level8R}
yneuron neuron0011000110 n0011000110mid 0 level8Params 
R00110001102 n0011000110mid n0011000110 {level8R}
R001100011001 n0011000110 n00110001100mid {level9R}
yneuron neuron00110001100 n00110001100mid 0 level9Params 
R001100011002 n00110001100mid n00110001100 {level9R}
R001100011011 n0011000110 n00110001101mid {level9R}
yneuron neuron00110001101 n00110001101mid 0 level9Params 
R001100011012 n00110001101mid n00110001101 {level9R}
R00110001111 n001100011 n0011000111mid {level8R}
yneuron neuron0011000111 n0011000111mid 0 level8Params 
R00110001112 n0011000111mid n0011000111 {level8R}
R001100011101 n0011000111 n00110001110mid {level9R}
yneuron neuron00110001110 n00110001110mid 0 level9Params 
R001100011102 n00110001110mid n00110001110 {level9R}
R001100011111 n0011000111 n00110001111mid {level9R}
yneuron neuron00110001111 n00110001111mid 0 level9Params 
R001100011112 n00110001111mid n00110001111 {level9R}
R00110011 n001100 n0011001mid {level5R}
yneuron neuron0011001 n0011001mid 0 level5Params 
R00110012 n0011001mid n0011001 {level5R}
R001100101 n0011001 n00110010mid {level6R}
yneuron neuron00110010 n00110010mid 0 level6Params 
R001100102 n00110010mid n00110010 {level6R}
R0011001001 n00110010 n001100100mid {level7R}
yneuron neuron001100100 n001100100mid 0 level7Params 
R0011001002 n001100100mid n001100100 {level7R}
R00110010001 n001100100 n0011001000mid {level8R}
yneuron neuron0011001000 n0011001000mid 0 level8Params 
R00110010002 n0011001000mid n0011001000 {level8R}
R001100100001 n0011001000 n00110010000mid {level9R}
yneuron neuron00110010000 n00110010000mid 0 level9Params 
R001100100002 n00110010000mid n00110010000 {level9R}
R001100100011 n0011001000 n00110010001mid {level9R}
yneuron neuron00110010001 n00110010001mid 0 level9Params 
R001100100012 n00110010001mid n00110010001 {level9R}
R00110010011 n001100100 n0011001001mid {level8R}
yneuron neuron0011001001 n0011001001mid 0 level8Params 
R00110010012 n0011001001mid n0011001001 {level8R}
R001100100101 n0011001001 n00110010010mid {level9R}
yneuron neuron00110010010 n00110010010mid 0 level9Params 
R001100100102 n00110010010mid n00110010010 {level9R}
R001100100111 n0011001001 n00110010011mid {level9R}
yneuron neuron00110010011 n00110010011mid 0 level9Params 
R001100100112 n00110010011mid n00110010011 {level9R}
R0011001011 n00110010 n001100101mid {level7R}
yneuron neuron001100101 n001100101mid 0 level7Params 
R0011001012 n001100101mid n001100101 {level7R}
R00110010101 n001100101 n0011001010mid {level8R}
yneuron neuron0011001010 n0011001010mid 0 level8Params 
R00110010102 n0011001010mid n0011001010 {level8R}
R001100101001 n0011001010 n00110010100mid {level9R}
yneuron neuron00110010100 n00110010100mid 0 level9Params 
R001100101002 n00110010100mid n00110010100 {level9R}
R001100101011 n0011001010 n00110010101mid {level9R}
yneuron neuron00110010101 n00110010101mid 0 level9Params 
R001100101012 n00110010101mid n00110010101 {level9R}
R00110010111 n001100101 n0011001011mid {level8R}
yneuron neuron0011001011 n0011001011mid 0 level8Params 
R00110010112 n0011001011mid n0011001011 {level8R}
R001100101101 n0011001011 n00110010110mid {level9R}
yneuron neuron00110010110 n00110010110mid 0 level9Params 
R001100101102 n00110010110mid n00110010110 {level9R}
R001100101111 n0011001011 n00110010111mid {level9R}
yneuron neuron00110010111 n00110010111mid 0 level9Params 
R001100101112 n00110010111mid n00110010111 {level9R}
R001100111 n0011001 n00110011mid {level6R}
yneuron neuron00110011 n00110011mid 0 level6Params 
R001100112 n00110011mid n00110011 {level6R}
R0011001101 n00110011 n001100110mid {level7R}
yneuron neuron001100110 n001100110mid 0 level7Params 
R0011001102 n001100110mid n001100110 {level7R}
R00110011001 n001100110 n0011001100mid {level8R}
yneuron neuron0011001100 n0011001100mid 0 level8Params 
R00110011002 n0011001100mid n0011001100 {level8R}
R001100110001 n0011001100 n00110011000mid {level9R}
yneuron neuron00110011000 n00110011000mid 0 level9Params 
R001100110002 n00110011000mid n00110011000 {level9R}
R001100110011 n0011001100 n00110011001mid {level9R}
yneuron neuron00110011001 n00110011001mid 0 level9Params 
R001100110012 n00110011001mid n00110011001 {level9R}
R00110011011 n001100110 n0011001101mid {level8R}
yneuron neuron0011001101 n0011001101mid 0 level8Params 
R00110011012 n0011001101mid n0011001101 {level8R}
R001100110101 n0011001101 n00110011010mid {level9R}
yneuron neuron00110011010 n00110011010mid 0 level9Params 
R001100110102 n00110011010mid n00110011010 {level9R}
R001100110111 n0011001101 n00110011011mid {level9R}
yneuron neuron00110011011 n00110011011mid 0 level9Params 
R001100110112 n00110011011mid n00110011011 {level9R}
R0011001111 n00110011 n001100111mid {level7R}
yneuron neuron001100111 n001100111mid 0 level7Params 
R0011001112 n001100111mid n001100111 {level7R}
R00110011101 n001100111 n0011001110mid {level8R}
yneuron neuron0011001110 n0011001110mid 0 level8Params 
R00110011102 n0011001110mid n0011001110 {level8R}
R001100111001 n0011001110 n00110011100mid {level9R}
yneuron neuron00110011100 n00110011100mid 0 level9Params 
R001100111002 n00110011100mid n00110011100 {level9R}
R001100111011 n0011001110 n00110011101mid {level9R}
yneuron neuron00110011101 n00110011101mid 0 level9Params 
R001100111012 n00110011101mid n00110011101 {level9R}
R00110011111 n001100111 n0011001111mid {level8R}
yneuron neuron0011001111 n0011001111mid 0 level8Params 
R00110011112 n0011001111mid n0011001111 {level8R}
R001100111101 n0011001111 n00110011110mid {level9R}
yneuron neuron00110011110 n00110011110mid 0 level9Params 
R001100111102 n00110011110mid n00110011110 {level9R}
R001100111111 n0011001111 n00110011111mid {level9R}
yneuron neuron00110011111 n00110011111mid 0 level9Params 
R001100111112 n00110011111mid n00110011111 {level9R}
R0011011 n00110 n001101mid {level4R}
yneuron neuron001101 n001101mid 0 level4Params 
R0011012 n001101mid n001101 {level4R}
R00110101 n001101 n0011010mid {level5R}
yneuron neuron0011010 n0011010mid 0 level5Params 
R00110102 n0011010mid n0011010 {level5R}
R001101001 n0011010 n00110100mid {level6R}
yneuron neuron00110100 n00110100mid 0 level6Params 
R001101002 n00110100mid n00110100 {level6R}
R0011010001 n00110100 n001101000mid {level7R}
yneuron neuron001101000 n001101000mid 0 level7Params 
R0011010002 n001101000mid n001101000 {level7R}
R00110100001 n001101000 n0011010000mid {level8R}
yneuron neuron0011010000 n0011010000mid 0 level8Params 
R00110100002 n0011010000mid n0011010000 {level8R}
R001101000001 n0011010000 n00110100000mid {level9R}
yneuron neuron00110100000 n00110100000mid 0 level9Params 
R001101000002 n00110100000mid n00110100000 {level9R}
R001101000011 n0011010000 n00110100001mid {level9R}
yneuron neuron00110100001 n00110100001mid 0 level9Params 
R001101000012 n00110100001mid n00110100001 {level9R}
R00110100011 n001101000 n0011010001mid {level8R}
yneuron neuron0011010001 n0011010001mid 0 level8Params 
R00110100012 n0011010001mid n0011010001 {level8R}
R001101000101 n0011010001 n00110100010mid {level9R}
yneuron neuron00110100010 n00110100010mid 0 level9Params 
R001101000102 n00110100010mid n00110100010 {level9R}
R001101000111 n0011010001 n00110100011mid {level9R}
yneuron neuron00110100011 n00110100011mid 0 level9Params 
R001101000112 n00110100011mid n00110100011 {level9R}
R0011010011 n00110100 n001101001mid {level7R}
yneuron neuron001101001 n001101001mid 0 level7Params 
R0011010012 n001101001mid n001101001 {level7R}
R00110100101 n001101001 n0011010010mid {level8R}
yneuron neuron0011010010 n0011010010mid 0 level8Params 
R00110100102 n0011010010mid n0011010010 {level8R}
R001101001001 n0011010010 n00110100100mid {level9R}
yneuron neuron00110100100 n00110100100mid 0 level9Params 
R001101001002 n00110100100mid n00110100100 {level9R}
R001101001011 n0011010010 n00110100101mid {level9R}
yneuron neuron00110100101 n00110100101mid 0 level9Params 
R001101001012 n00110100101mid n00110100101 {level9R}
R00110100111 n001101001 n0011010011mid {level8R}
yneuron neuron0011010011 n0011010011mid 0 level8Params 
R00110100112 n0011010011mid n0011010011 {level8R}
R001101001101 n0011010011 n00110100110mid {level9R}
yneuron neuron00110100110 n00110100110mid 0 level9Params 
R001101001102 n00110100110mid n00110100110 {level9R}
R001101001111 n0011010011 n00110100111mid {level9R}
yneuron neuron00110100111 n00110100111mid 0 level9Params 
R001101001112 n00110100111mid n00110100111 {level9R}
R001101011 n0011010 n00110101mid {level6R}
yneuron neuron00110101 n00110101mid 0 level6Params 
R001101012 n00110101mid n00110101 {level6R}
R0011010101 n00110101 n001101010mid {level7R}
yneuron neuron001101010 n001101010mid 0 level7Params 
R0011010102 n001101010mid n001101010 {level7R}
R00110101001 n001101010 n0011010100mid {level8R}
yneuron neuron0011010100 n0011010100mid 0 level8Params 
R00110101002 n0011010100mid n0011010100 {level8R}
R001101010001 n0011010100 n00110101000mid {level9R}
yneuron neuron00110101000 n00110101000mid 0 level9Params 
R001101010002 n00110101000mid n00110101000 {level9R}
R001101010011 n0011010100 n00110101001mid {level9R}
yneuron neuron00110101001 n00110101001mid 0 level9Params 
R001101010012 n00110101001mid n00110101001 {level9R}
R00110101011 n001101010 n0011010101mid {level8R}
yneuron neuron0011010101 n0011010101mid 0 level8Params 
R00110101012 n0011010101mid n0011010101 {level8R}
R001101010101 n0011010101 n00110101010mid {level9R}
yneuron neuron00110101010 n00110101010mid 0 level9Params 
R001101010102 n00110101010mid n00110101010 {level9R}
R001101010111 n0011010101 n00110101011mid {level9R}
yneuron neuron00110101011 n00110101011mid 0 level9Params 
R001101010112 n00110101011mid n00110101011 {level9R}
R0011010111 n00110101 n001101011mid {level7R}
yneuron neuron001101011 n001101011mid 0 level7Params 
R0011010112 n001101011mid n001101011 {level7R}
R00110101101 n001101011 n0011010110mid {level8R}
yneuron neuron0011010110 n0011010110mid 0 level8Params 
R00110101102 n0011010110mid n0011010110 {level8R}
R001101011001 n0011010110 n00110101100mid {level9R}
yneuron neuron00110101100 n00110101100mid 0 level9Params 
R001101011002 n00110101100mid n00110101100 {level9R}
R001101011011 n0011010110 n00110101101mid {level9R}
yneuron neuron00110101101 n00110101101mid 0 level9Params 
R001101011012 n00110101101mid n00110101101 {level9R}
R00110101111 n001101011 n0011010111mid {level8R}
yneuron neuron0011010111 n0011010111mid 0 level8Params 
R00110101112 n0011010111mid n0011010111 {level8R}
R001101011101 n0011010111 n00110101110mid {level9R}
yneuron neuron00110101110 n00110101110mid 0 level9Params 
R001101011102 n00110101110mid n00110101110 {level9R}
R001101011111 n0011010111 n00110101111mid {level9R}
yneuron neuron00110101111 n00110101111mid 0 level9Params 
R001101011112 n00110101111mid n00110101111 {level9R}
R00110111 n001101 n0011011mid {level5R}
yneuron neuron0011011 n0011011mid 0 level5Params 
R00110112 n0011011mid n0011011 {level5R}
R001101101 n0011011 n00110110mid {level6R}
yneuron neuron00110110 n00110110mid 0 level6Params 
R001101102 n00110110mid n00110110 {level6R}
R0011011001 n00110110 n001101100mid {level7R}
yneuron neuron001101100 n001101100mid 0 level7Params 
R0011011002 n001101100mid n001101100 {level7R}
R00110110001 n001101100 n0011011000mid {level8R}
yneuron neuron0011011000 n0011011000mid 0 level8Params 
R00110110002 n0011011000mid n0011011000 {level8R}
R001101100001 n0011011000 n00110110000mid {level9R}
yneuron neuron00110110000 n00110110000mid 0 level9Params 
R001101100002 n00110110000mid n00110110000 {level9R}
R001101100011 n0011011000 n00110110001mid {level9R}
yneuron neuron00110110001 n00110110001mid 0 level9Params 
R001101100012 n00110110001mid n00110110001 {level9R}
R00110110011 n001101100 n0011011001mid {level8R}
yneuron neuron0011011001 n0011011001mid 0 level8Params 
R00110110012 n0011011001mid n0011011001 {level8R}
R001101100101 n0011011001 n00110110010mid {level9R}
yneuron neuron00110110010 n00110110010mid 0 level9Params 
R001101100102 n00110110010mid n00110110010 {level9R}
R001101100111 n0011011001 n00110110011mid {level9R}
yneuron neuron00110110011 n00110110011mid 0 level9Params 
R001101100112 n00110110011mid n00110110011 {level9R}
R0011011011 n00110110 n001101101mid {level7R}
yneuron neuron001101101 n001101101mid 0 level7Params 
R0011011012 n001101101mid n001101101 {level7R}
R00110110101 n001101101 n0011011010mid {level8R}
yneuron neuron0011011010 n0011011010mid 0 level8Params 
R00110110102 n0011011010mid n0011011010 {level8R}
R001101101001 n0011011010 n00110110100mid {level9R}
yneuron neuron00110110100 n00110110100mid 0 level9Params 
R001101101002 n00110110100mid n00110110100 {level9R}
R001101101011 n0011011010 n00110110101mid {level9R}
yneuron neuron00110110101 n00110110101mid 0 level9Params 
R001101101012 n00110110101mid n00110110101 {level9R}
R00110110111 n001101101 n0011011011mid {level8R}
yneuron neuron0011011011 n0011011011mid 0 level8Params 
R00110110112 n0011011011mid n0011011011 {level8R}
R001101101101 n0011011011 n00110110110mid {level9R}
yneuron neuron00110110110 n00110110110mid 0 level9Params 
R001101101102 n00110110110mid n00110110110 {level9R}
R001101101111 n0011011011 n00110110111mid {level9R}
yneuron neuron00110110111 n00110110111mid 0 level9Params 
R001101101112 n00110110111mid n00110110111 {level9R}
R001101111 n0011011 n00110111mid {level6R}
yneuron neuron00110111 n00110111mid 0 level6Params 
R001101112 n00110111mid n00110111 {level6R}
R0011011101 n00110111 n001101110mid {level7R}
yneuron neuron001101110 n001101110mid 0 level7Params 
R0011011102 n001101110mid n001101110 {level7R}
R00110111001 n001101110 n0011011100mid {level8R}
yneuron neuron0011011100 n0011011100mid 0 level8Params 
R00110111002 n0011011100mid n0011011100 {level8R}
R001101110001 n0011011100 n00110111000mid {level9R}
yneuron neuron00110111000 n00110111000mid 0 level9Params 
R001101110002 n00110111000mid n00110111000 {level9R}
R001101110011 n0011011100 n00110111001mid {level9R}
yneuron neuron00110111001 n00110111001mid 0 level9Params 
R001101110012 n00110111001mid n00110111001 {level9R}
R00110111011 n001101110 n0011011101mid {level8R}
yneuron neuron0011011101 n0011011101mid 0 level8Params 
R00110111012 n0011011101mid n0011011101 {level8R}
R001101110101 n0011011101 n00110111010mid {level9R}
yneuron neuron00110111010 n00110111010mid 0 level9Params 
R001101110102 n00110111010mid n00110111010 {level9R}
R001101110111 n0011011101 n00110111011mid {level9R}
yneuron neuron00110111011 n00110111011mid 0 level9Params 
R001101110112 n00110111011mid n00110111011 {level9R}
R0011011111 n00110111 n001101111mid {level7R}
yneuron neuron001101111 n001101111mid 0 level7Params 
R0011011112 n001101111mid n001101111 {level7R}
R00110111101 n001101111 n0011011110mid {level8R}
yneuron neuron0011011110 n0011011110mid 0 level8Params 
R00110111102 n0011011110mid n0011011110 {level8R}
R001101111001 n0011011110 n00110111100mid {level9R}
yneuron neuron00110111100 n00110111100mid 0 level9Params 
R001101111002 n00110111100mid n00110111100 {level9R}
R001101111011 n0011011110 n00110111101mid {level9R}
yneuron neuron00110111101 n00110111101mid 0 level9Params 
R001101111012 n00110111101mid n00110111101 {level9R}
R00110111111 n001101111 n0011011111mid {level8R}
yneuron neuron0011011111 n0011011111mid 0 level8Params 
R00110111112 n0011011111mid n0011011111 {level8R}
R001101111101 n0011011111 n00110111110mid {level9R}
yneuron neuron00110111110 n00110111110mid 0 level9Params 
R001101111102 n00110111110mid n00110111110 {level9R}
R001101111111 n0011011111 n00110111111mid {level9R}
yneuron neuron00110111111 n00110111111mid 0 level9Params 
R001101111112 n00110111111mid n00110111111 {level9R}
R001111 n0011 n00111mid {level3R}
yneuron neuron00111 n00111mid 0 level3Params 
R001112 n00111mid n00111 {level3R}
R0011101 n00111 n001110mid {level4R}
yneuron neuron001110 n001110mid 0 level4Params 
R0011102 n001110mid n001110 {level4R}
R00111001 n001110 n0011100mid {level5R}
yneuron neuron0011100 n0011100mid 0 level5Params 
R00111002 n0011100mid n0011100 {level5R}
R001110001 n0011100 n00111000mid {level6R}
yneuron neuron00111000 n00111000mid 0 level6Params 
R001110002 n00111000mid n00111000 {level6R}
R0011100001 n00111000 n001110000mid {level7R}
yneuron neuron001110000 n001110000mid 0 level7Params 
R0011100002 n001110000mid n001110000 {level7R}
R00111000001 n001110000 n0011100000mid {level8R}
yneuron neuron0011100000 n0011100000mid 0 level8Params 
R00111000002 n0011100000mid n0011100000 {level8R}
R001110000001 n0011100000 n00111000000mid {level9R}
yneuron neuron00111000000 n00111000000mid 0 level9Params 
R001110000002 n00111000000mid n00111000000 {level9R}
R001110000011 n0011100000 n00111000001mid {level9R}
yneuron neuron00111000001 n00111000001mid 0 level9Params 
R001110000012 n00111000001mid n00111000001 {level9R}
R00111000011 n001110000 n0011100001mid {level8R}
yneuron neuron0011100001 n0011100001mid 0 level8Params 
R00111000012 n0011100001mid n0011100001 {level8R}
R001110000101 n0011100001 n00111000010mid {level9R}
yneuron neuron00111000010 n00111000010mid 0 level9Params 
R001110000102 n00111000010mid n00111000010 {level9R}
R001110000111 n0011100001 n00111000011mid {level9R}
yneuron neuron00111000011 n00111000011mid 0 level9Params 
R001110000112 n00111000011mid n00111000011 {level9R}
R0011100011 n00111000 n001110001mid {level7R}
yneuron neuron001110001 n001110001mid 0 level7Params 
R0011100012 n001110001mid n001110001 {level7R}
R00111000101 n001110001 n0011100010mid {level8R}
yneuron neuron0011100010 n0011100010mid 0 level8Params 
R00111000102 n0011100010mid n0011100010 {level8R}
R001110001001 n0011100010 n00111000100mid {level9R}
yneuron neuron00111000100 n00111000100mid 0 level9Params 
R001110001002 n00111000100mid n00111000100 {level9R}
R001110001011 n0011100010 n00111000101mid {level9R}
yneuron neuron00111000101 n00111000101mid 0 level9Params 
R001110001012 n00111000101mid n00111000101 {level9R}
R00111000111 n001110001 n0011100011mid {level8R}
yneuron neuron0011100011 n0011100011mid 0 level8Params 
R00111000112 n0011100011mid n0011100011 {level8R}
R001110001101 n0011100011 n00111000110mid {level9R}
yneuron neuron00111000110 n00111000110mid 0 level9Params 
R001110001102 n00111000110mid n00111000110 {level9R}
R001110001111 n0011100011 n00111000111mid {level9R}
yneuron neuron00111000111 n00111000111mid 0 level9Params 
R001110001112 n00111000111mid n00111000111 {level9R}
R001110011 n0011100 n00111001mid {level6R}
yneuron neuron00111001 n00111001mid 0 level6Params 
R001110012 n00111001mid n00111001 {level6R}
R0011100101 n00111001 n001110010mid {level7R}
yneuron neuron001110010 n001110010mid 0 level7Params 
R0011100102 n001110010mid n001110010 {level7R}
R00111001001 n001110010 n0011100100mid {level8R}
yneuron neuron0011100100 n0011100100mid 0 level8Params 
R00111001002 n0011100100mid n0011100100 {level8R}
R001110010001 n0011100100 n00111001000mid {level9R}
yneuron neuron00111001000 n00111001000mid 0 level9Params 
R001110010002 n00111001000mid n00111001000 {level9R}
R001110010011 n0011100100 n00111001001mid {level9R}
yneuron neuron00111001001 n00111001001mid 0 level9Params 
R001110010012 n00111001001mid n00111001001 {level9R}
R00111001011 n001110010 n0011100101mid {level8R}
yneuron neuron0011100101 n0011100101mid 0 level8Params 
R00111001012 n0011100101mid n0011100101 {level8R}
R001110010101 n0011100101 n00111001010mid {level9R}
yneuron neuron00111001010 n00111001010mid 0 level9Params 
R001110010102 n00111001010mid n00111001010 {level9R}
R001110010111 n0011100101 n00111001011mid {level9R}
yneuron neuron00111001011 n00111001011mid 0 level9Params 
R001110010112 n00111001011mid n00111001011 {level9R}
R0011100111 n00111001 n001110011mid {level7R}
yneuron neuron001110011 n001110011mid 0 level7Params 
R0011100112 n001110011mid n001110011 {level7R}
R00111001101 n001110011 n0011100110mid {level8R}
yneuron neuron0011100110 n0011100110mid 0 level8Params 
R00111001102 n0011100110mid n0011100110 {level8R}
R001110011001 n0011100110 n00111001100mid {level9R}
yneuron neuron00111001100 n00111001100mid 0 level9Params 
R001110011002 n00111001100mid n00111001100 {level9R}
R001110011011 n0011100110 n00111001101mid {level9R}
yneuron neuron00111001101 n00111001101mid 0 level9Params 
R001110011012 n00111001101mid n00111001101 {level9R}
R00111001111 n001110011 n0011100111mid {level8R}
yneuron neuron0011100111 n0011100111mid 0 level8Params 
R00111001112 n0011100111mid n0011100111 {level8R}
R001110011101 n0011100111 n00111001110mid {level9R}
yneuron neuron00111001110 n00111001110mid 0 level9Params 
R001110011102 n00111001110mid n00111001110 {level9R}
R001110011111 n0011100111 n00111001111mid {level9R}
yneuron neuron00111001111 n00111001111mid 0 level9Params 
R001110011112 n00111001111mid n00111001111 {level9R}
R00111011 n001110 n0011101mid {level5R}
yneuron neuron0011101 n0011101mid 0 level5Params 
R00111012 n0011101mid n0011101 {level5R}
R001110101 n0011101 n00111010mid {level6R}
yneuron neuron00111010 n00111010mid 0 level6Params 
R001110102 n00111010mid n00111010 {level6R}
R0011101001 n00111010 n001110100mid {level7R}
yneuron neuron001110100 n001110100mid 0 level7Params 
R0011101002 n001110100mid n001110100 {level7R}
R00111010001 n001110100 n0011101000mid {level8R}
yneuron neuron0011101000 n0011101000mid 0 level8Params 
R00111010002 n0011101000mid n0011101000 {level8R}
R001110100001 n0011101000 n00111010000mid {level9R}
yneuron neuron00111010000 n00111010000mid 0 level9Params 
R001110100002 n00111010000mid n00111010000 {level9R}
R001110100011 n0011101000 n00111010001mid {level9R}
yneuron neuron00111010001 n00111010001mid 0 level9Params 
R001110100012 n00111010001mid n00111010001 {level9R}
R00111010011 n001110100 n0011101001mid {level8R}
yneuron neuron0011101001 n0011101001mid 0 level8Params 
R00111010012 n0011101001mid n0011101001 {level8R}
R001110100101 n0011101001 n00111010010mid {level9R}
yneuron neuron00111010010 n00111010010mid 0 level9Params 
R001110100102 n00111010010mid n00111010010 {level9R}
R001110100111 n0011101001 n00111010011mid {level9R}
yneuron neuron00111010011 n00111010011mid 0 level9Params 
R001110100112 n00111010011mid n00111010011 {level9R}
R0011101011 n00111010 n001110101mid {level7R}
yneuron neuron001110101 n001110101mid 0 level7Params 
R0011101012 n001110101mid n001110101 {level7R}
R00111010101 n001110101 n0011101010mid {level8R}
yneuron neuron0011101010 n0011101010mid 0 level8Params 
R00111010102 n0011101010mid n0011101010 {level8R}
R001110101001 n0011101010 n00111010100mid {level9R}
yneuron neuron00111010100 n00111010100mid 0 level9Params 
R001110101002 n00111010100mid n00111010100 {level9R}
R001110101011 n0011101010 n00111010101mid {level9R}
yneuron neuron00111010101 n00111010101mid 0 level9Params 
R001110101012 n00111010101mid n00111010101 {level9R}
R00111010111 n001110101 n0011101011mid {level8R}
yneuron neuron0011101011 n0011101011mid 0 level8Params 
R00111010112 n0011101011mid n0011101011 {level8R}
R001110101101 n0011101011 n00111010110mid {level9R}
yneuron neuron00111010110 n00111010110mid 0 level9Params 
R001110101102 n00111010110mid n00111010110 {level9R}
R001110101111 n0011101011 n00111010111mid {level9R}
yneuron neuron00111010111 n00111010111mid 0 level9Params 
R001110101112 n00111010111mid n00111010111 {level9R}
R001110111 n0011101 n00111011mid {level6R}
yneuron neuron00111011 n00111011mid 0 level6Params 
R001110112 n00111011mid n00111011 {level6R}
R0011101101 n00111011 n001110110mid {level7R}
yneuron neuron001110110 n001110110mid 0 level7Params 
R0011101102 n001110110mid n001110110 {level7R}
R00111011001 n001110110 n0011101100mid {level8R}
yneuron neuron0011101100 n0011101100mid 0 level8Params 
R00111011002 n0011101100mid n0011101100 {level8R}
R001110110001 n0011101100 n00111011000mid {level9R}
yneuron neuron00111011000 n00111011000mid 0 level9Params 
R001110110002 n00111011000mid n00111011000 {level9R}
R001110110011 n0011101100 n00111011001mid {level9R}
yneuron neuron00111011001 n00111011001mid 0 level9Params 
R001110110012 n00111011001mid n00111011001 {level9R}
R00111011011 n001110110 n0011101101mid {level8R}
yneuron neuron0011101101 n0011101101mid 0 level8Params 
R00111011012 n0011101101mid n0011101101 {level8R}
R001110110101 n0011101101 n00111011010mid {level9R}
yneuron neuron00111011010 n00111011010mid 0 level9Params 
R001110110102 n00111011010mid n00111011010 {level9R}
R001110110111 n0011101101 n00111011011mid {level9R}
yneuron neuron00111011011 n00111011011mid 0 level9Params 
R001110110112 n00111011011mid n00111011011 {level9R}
R0011101111 n00111011 n001110111mid {level7R}
yneuron neuron001110111 n001110111mid 0 level7Params 
R0011101112 n001110111mid n001110111 {level7R}
R00111011101 n001110111 n0011101110mid {level8R}
yneuron neuron0011101110 n0011101110mid 0 level8Params 
R00111011102 n0011101110mid n0011101110 {level8R}
R001110111001 n0011101110 n00111011100mid {level9R}
yneuron neuron00111011100 n00111011100mid 0 level9Params 
R001110111002 n00111011100mid n00111011100 {level9R}
R001110111011 n0011101110 n00111011101mid {level9R}
yneuron neuron00111011101 n00111011101mid 0 level9Params 
R001110111012 n00111011101mid n00111011101 {level9R}
R00111011111 n001110111 n0011101111mid {level8R}
yneuron neuron0011101111 n0011101111mid 0 level8Params 
R00111011112 n0011101111mid n0011101111 {level8R}
R001110111101 n0011101111 n00111011110mid {level9R}
yneuron neuron00111011110 n00111011110mid 0 level9Params 
R001110111102 n00111011110mid n00111011110 {level9R}
R001110111111 n0011101111 n00111011111mid {level9R}
yneuron neuron00111011111 n00111011111mid 0 level9Params 
R001110111112 n00111011111mid n00111011111 {level9R}
R0011111 n00111 n001111mid {level4R}
yneuron neuron001111 n001111mid 0 level4Params 
R0011112 n001111mid n001111 {level4R}
R00111101 n001111 n0011110mid {level5R}
yneuron neuron0011110 n0011110mid 0 level5Params 
R00111102 n0011110mid n0011110 {level5R}
R001111001 n0011110 n00111100mid {level6R}
yneuron neuron00111100 n00111100mid 0 level6Params 
R001111002 n00111100mid n00111100 {level6R}
R0011110001 n00111100 n001111000mid {level7R}
yneuron neuron001111000 n001111000mid 0 level7Params 
R0011110002 n001111000mid n001111000 {level7R}
R00111100001 n001111000 n0011110000mid {level8R}
yneuron neuron0011110000 n0011110000mid 0 level8Params 
R00111100002 n0011110000mid n0011110000 {level8R}
R001111000001 n0011110000 n00111100000mid {level9R}
yneuron neuron00111100000 n00111100000mid 0 level9Params 
R001111000002 n00111100000mid n00111100000 {level9R}
R001111000011 n0011110000 n00111100001mid {level9R}
yneuron neuron00111100001 n00111100001mid 0 level9Params 
R001111000012 n00111100001mid n00111100001 {level9R}
R00111100011 n001111000 n0011110001mid {level8R}
yneuron neuron0011110001 n0011110001mid 0 level8Params 
R00111100012 n0011110001mid n0011110001 {level8R}
R001111000101 n0011110001 n00111100010mid {level9R}
yneuron neuron00111100010 n00111100010mid 0 level9Params 
R001111000102 n00111100010mid n00111100010 {level9R}
R001111000111 n0011110001 n00111100011mid {level9R}
yneuron neuron00111100011 n00111100011mid 0 level9Params 
R001111000112 n00111100011mid n00111100011 {level9R}
R0011110011 n00111100 n001111001mid {level7R}
yneuron neuron001111001 n001111001mid 0 level7Params 
R0011110012 n001111001mid n001111001 {level7R}
R00111100101 n001111001 n0011110010mid {level8R}
yneuron neuron0011110010 n0011110010mid 0 level8Params 
R00111100102 n0011110010mid n0011110010 {level8R}
R001111001001 n0011110010 n00111100100mid {level9R}
yneuron neuron00111100100 n00111100100mid 0 level9Params 
R001111001002 n00111100100mid n00111100100 {level9R}
R001111001011 n0011110010 n00111100101mid {level9R}
yneuron neuron00111100101 n00111100101mid 0 level9Params 
R001111001012 n00111100101mid n00111100101 {level9R}
R00111100111 n001111001 n0011110011mid {level8R}
yneuron neuron0011110011 n0011110011mid 0 level8Params 
R00111100112 n0011110011mid n0011110011 {level8R}
R001111001101 n0011110011 n00111100110mid {level9R}
yneuron neuron00111100110 n00111100110mid 0 level9Params 
R001111001102 n00111100110mid n00111100110 {level9R}
R001111001111 n0011110011 n00111100111mid {level9R}
yneuron neuron00111100111 n00111100111mid 0 level9Params 
R001111001112 n00111100111mid n00111100111 {level9R}
R001111011 n0011110 n00111101mid {level6R}
yneuron neuron00111101 n00111101mid 0 level6Params 
R001111012 n00111101mid n00111101 {level6R}
R0011110101 n00111101 n001111010mid {level7R}
yneuron neuron001111010 n001111010mid 0 level7Params 
R0011110102 n001111010mid n001111010 {level7R}
R00111101001 n001111010 n0011110100mid {level8R}
yneuron neuron0011110100 n0011110100mid 0 level8Params 
R00111101002 n0011110100mid n0011110100 {level8R}
R001111010001 n0011110100 n00111101000mid {level9R}
yneuron neuron00111101000 n00111101000mid 0 level9Params 
R001111010002 n00111101000mid n00111101000 {level9R}
R001111010011 n0011110100 n00111101001mid {level9R}
yneuron neuron00111101001 n00111101001mid 0 level9Params 
R001111010012 n00111101001mid n00111101001 {level9R}
R00111101011 n001111010 n0011110101mid {level8R}
yneuron neuron0011110101 n0011110101mid 0 level8Params 
R00111101012 n0011110101mid n0011110101 {level8R}
R001111010101 n0011110101 n00111101010mid {level9R}
yneuron neuron00111101010 n00111101010mid 0 level9Params 
R001111010102 n00111101010mid n00111101010 {level9R}
R001111010111 n0011110101 n00111101011mid {level9R}
yneuron neuron00111101011 n00111101011mid 0 level9Params 
R001111010112 n00111101011mid n00111101011 {level9R}
R0011110111 n00111101 n001111011mid {level7R}
yneuron neuron001111011 n001111011mid 0 level7Params 
R0011110112 n001111011mid n001111011 {level7R}
R00111101101 n001111011 n0011110110mid {level8R}
yneuron neuron0011110110 n0011110110mid 0 level8Params 
R00111101102 n0011110110mid n0011110110 {level8R}
R001111011001 n0011110110 n00111101100mid {level9R}
yneuron neuron00111101100 n00111101100mid 0 level9Params 
R001111011002 n00111101100mid n00111101100 {level9R}
R001111011011 n0011110110 n00111101101mid {level9R}
yneuron neuron00111101101 n00111101101mid 0 level9Params 
R001111011012 n00111101101mid n00111101101 {level9R}
R00111101111 n001111011 n0011110111mid {level8R}
yneuron neuron0011110111 n0011110111mid 0 level8Params 
R00111101112 n0011110111mid n0011110111 {level8R}
R001111011101 n0011110111 n00111101110mid {level9R}
yneuron neuron00111101110 n00111101110mid 0 level9Params 
R001111011102 n00111101110mid n00111101110 {level9R}
R001111011111 n0011110111 n00111101111mid {level9R}
yneuron neuron00111101111 n00111101111mid 0 level9Params 
R001111011112 n00111101111mid n00111101111 {level9R}
R00111111 n001111 n0011111mid {level5R}
yneuron neuron0011111 n0011111mid 0 level5Params 
R00111112 n0011111mid n0011111 {level5R}
R001111101 n0011111 n00111110mid {level6R}
yneuron neuron00111110 n00111110mid 0 level6Params 
R001111102 n00111110mid n00111110 {level6R}
R0011111001 n00111110 n001111100mid {level7R}
yneuron neuron001111100 n001111100mid 0 level7Params 
R0011111002 n001111100mid n001111100 {level7R}
R00111110001 n001111100 n0011111000mid {level8R}
yneuron neuron0011111000 n0011111000mid 0 level8Params 
R00111110002 n0011111000mid n0011111000 {level8R}
R001111100001 n0011111000 n00111110000mid {level9R}
yneuron neuron00111110000 n00111110000mid 0 level9Params 
R001111100002 n00111110000mid n00111110000 {level9R}
R001111100011 n0011111000 n00111110001mid {level9R}
yneuron neuron00111110001 n00111110001mid 0 level9Params 
R001111100012 n00111110001mid n00111110001 {level9R}
R00111110011 n001111100 n0011111001mid {level8R}
yneuron neuron0011111001 n0011111001mid 0 level8Params 
R00111110012 n0011111001mid n0011111001 {level8R}
R001111100101 n0011111001 n00111110010mid {level9R}
yneuron neuron00111110010 n00111110010mid 0 level9Params 
R001111100102 n00111110010mid n00111110010 {level9R}
R001111100111 n0011111001 n00111110011mid {level9R}
yneuron neuron00111110011 n00111110011mid 0 level9Params 
R001111100112 n00111110011mid n00111110011 {level9R}
R0011111011 n00111110 n001111101mid {level7R}
yneuron neuron001111101 n001111101mid 0 level7Params 
R0011111012 n001111101mid n001111101 {level7R}
R00111110101 n001111101 n0011111010mid {level8R}
yneuron neuron0011111010 n0011111010mid 0 level8Params 
R00111110102 n0011111010mid n0011111010 {level8R}
R001111101001 n0011111010 n00111110100mid {level9R}
yneuron neuron00111110100 n00111110100mid 0 level9Params 
R001111101002 n00111110100mid n00111110100 {level9R}
R001111101011 n0011111010 n00111110101mid {level9R}
yneuron neuron00111110101 n00111110101mid 0 level9Params 
R001111101012 n00111110101mid n00111110101 {level9R}
R00111110111 n001111101 n0011111011mid {level8R}
yneuron neuron0011111011 n0011111011mid 0 level8Params 
R00111110112 n0011111011mid n0011111011 {level8R}
R001111101101 n0011111011 n00111110110mid {level9R}
yneuron neuron00111110110 n00111110110mid 0 level9Params 
R001111101102 n00111110110mid n00111110110 {level9R}
R001111101111 n0011111011 n00111110111mid {level9R}
yneuron neuron00111110111 n00111110111mid 0 level9Params 
R001111101112 n00111110111mid n00111110111 {level9R}
R001111111 n0011111 n00111111mid {level6R}
yneuron neuron00111111 n00111111mid 0 level6Params 
R001111112 n00111111mid n00111111 {level6R}
R0011111101 n00111111 n001111110mid {level7R}
yneuron neuron001111110 n001111110mid 0 level7Params 
R0011111102 n001111110mid n001111110 {level7R}
R00111111001 n001111110 n0011111100mid {level8R}
yneuron neuron0011111100 n0011111100mid 0 level8Params 
R00111111002 n0011111100mid n0011111100 {level8R}
R001111110001 n0011111100 n00111111000mid {level9R}
yneuron neuron00111111000 n00111111000mid 0 level9Params 
R001111110002 n00111111000mid n00111111000 {level9R}
R001111110011 n0011111100 n00111111001mid {level9R}
yneuron neuron00111111001 n00111111001mid 0 level9Params 
R001111110012 n00111111001mid n00111111001 {level9R}
R00111111011 n001111110 n0011111101mid {level8R}
yneuron neuron0011111101 n0011111101mid 0 level8Params 
R00111111012 n0011111101mid n0011111101 {level8R}
R001111110101 n0011111101 n00111111010mid {level9R}
yneuron neuron00111111010 n00111111010mid 0 level9Params 
R001111110102 n00111111010mid n00111111010 {level9R}
R001111110111 n0011111101 n00111111011mid {level9R}
yneuron neuron00111111011 n00111111011mid 0 level9Params 
R001111110112 n00111111011mid n00111111011 {level9R}
R0011111111 n00111111 n001111111mid {level7R}
yneuron neuron001111111 n001111111mid 0 level7Params 
R0011111112 n001111111mid n001111111 {level7R}
R00111111101 n001111111 n0011111110mid {level8R}
yneuron neuron0011111110 n0011111110mid 0 level8Params 
R00111111102 n0011111110mid n0011111110 {level8R}
R001111111001 n0011111110 n00111111100mid {level9R}
yneuron neuron00111111100 n00111111100mid 0 level9Params 
R001111111002 n00111111100mid n00111111100 {level9R}
R001111111011 n0011111110 n00111111101mid {level9R}
yneuron neuron00111111101 n00111111101mid 0 level9Params 
R001111111012 n00111111101mid n00111111101 {level9R}
R00111111111 n001111111 n0011111111mid {level8R}
yneuron neuron0011111111 n0011111111mid 0 level8Params 
R00111111112 n0011111111mid n0011111111 {level8R}
R001111111101 n0011111111 n00111111110mid {level9R}
yneuron neuron00111111110 n00111111110mid 0 level9Params 
R001111111102 n00111111110mid n00111111110 {level9R}
R001111111111 n0011111111 n00111111111mid {level9R}
yneuron neuron00111111111 n00111111111mid 0 level9Params 
R001111111112 n00111111111mid n00111111111 {level9R}

.print tran v(n0) 
*+ i(Iin) 
+ v(n00000000000) 

.end
