Baseline for subcircuit/expression tests
****************************************************************************
*
* Tests that expressions used in subcircuits work properly when using both
* local nodes and nodes from the .subckt line.
*
* This test simply puts the B source into a subcircuit, but with a chance that
* a subcircuit local node could be confused with the global node of the same
* name that is passed in to the subcircuit
*
****************************************************************************


V2 2 0 10V
R2 2 0 1
V3 3 0 100V
R3 3 0 1

XsubK1 1 2 3 4 SubK1

.subckt SubK1 S1 S2 S3 S4
B1 S4 0 V={V(S3)+V(S2)*V(3)}
R4 S4 0 1
V1 3 0 5V
R1 3 0 1
B2 S1 0 V={V(3)}
R2 S1 0 1
.ends

.print DC V(2) V(1) V(3) V(4)
.DC V2 0 10 1

.end