********************************************************
* Test that Xyce exits gracefully with a reasonable error
* message if the specified save file is in a subdirectory
* that does not exist.
*
* The contents of this netlist doesn't really matter.
* The .SAVE line is trying to write to a file in a 
* non-existent subdirectory.
*
*
*********************************************************
V1 1 0 SIN(0 1 1HZ)
R1 1 2 1
R2 2 0 2

.TRAN 0 1S
.PRINT TRAN V(2)

* attempting to write the Save file to a directory
.SAVE TYPE=IC FILE=bogo_dir/save.cir.ic

.END 
