Regression test to show proper transient RC circuit
********************************************************************************
* erkeite.  10/15/2007.
*
* This test is a simple test of .dcvolt.  It is nearly identical to the
* CAPACITOR/capacitor.cir test, except that it relies on .DCVOLT rather than
* IC= on the device instance line.  The result should be exactly the same.
* Similar to that test, this test compares directly to an analytic
* solution, rather than a numerically-generated gold standard.
*
* This version of the test uses the .DCVOLT form:  
*   .dcvolt v(node1)=val1  <v(node2)=val2> ...
*
*  Another, nearly identical test, IC_AND_NODESET/dcvolt_cap2.cir, is exactly
*  the same except that it uses the form:
*  .dcvolt node1 value1  <node2 value2>  <node3 value3> ...
*
********************************************************************************
.param V1=1.0
.dcvolt v(1)={V1}

c1 1 0 1uF 
R1 1 2 1K
v1 2 0 0V
.print tran v(1)
.tran 0 5ms
.options timeint reltol=1e-6 abstol=1e-6
.end

