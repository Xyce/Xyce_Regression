Multiple print HB lines --- baselne
* This test of a simple inverter circuit is use to produce the single
* print line baseline case for case 7 of the bug 538 SON test set.

.hb 1e5
.print hb_td file=foo1_bl {v(vout)+1.0} {v(in) +4.0}  {v(1) +4.0} ig(MP1) ig(MN1) is(MP1) id(MN1)  id(MP1)
.print hb_fd file=foo2_bl {v(vout)+1.0} {v(in) +4.0}  {v(1) +4.0} ig(MP1) ig(MN1) is(MP1) id(MN1)  id(MP1)

.options hbint numfreq=30 STARTUPPERIODS=2
.options linsol-hb type=aztecoo


VDDdev 	VDD	0	3V
RIN	IN	1	1K
*                   v1 v2   td  tr  tf   pw   per
*VIN1  1	0  5V PULSE (5V 0V 1.5us 5ns 5ns 1.5us 3us)
*VIN1  1	0  5V PULSE (5V 0V 1.5us 0.15us 0.15us 1.5us 3.3us)
VIN1 1 0 sin 0  3V 1e5 0 0

R1    VOUT  0  10K
C2    VOUT  0  0.1p
MN1   VOUT  IN 0 0 CD4012_NMOS L=5u W=175u
MP1   VOUT IN VDD VDD CD4012_PMOS L=5u W=270u
**************************************************************************
.MODEL cd4012_pmos PMOS (LEVEL=2)
**************************************************************************
.MODEL cd4012_nmos NMOS (
+ LEVEL = 2)
.END
