* Test various invalid .model statements
* See SRN Bug 2107 for more details.

.TRAN 0.5U 400ms
.PRINT TRAN v(3) v(2) 
VIN  1 0 PULSE(0 1 10U 1U 1U 100m)
R    2 1 1K
D1   3 2 D1N3940_short  
rload 3 0 1K

R2   4 1 1K
D2   4 5 D1N3940_UMP
rload2 5 0 1K

* .model statement must have at least three elements
.MODEL D1N3940_short

* .model statement lacks the closing parenthesis
.MODEL D1N3940_UMP D(
+ IS = 4E-10
+ RS = .105
+ N = 1.48
+ TT = 8E-7
+ CJO = 1.95E-11
+ VJ = .4
+ M = .38
+ EG = 1.36
+ XTI = -8
+ KF = 0
+ AF = 1
+ FC = .9
+ BV = 600
+ IBV = 1E-4

.END

