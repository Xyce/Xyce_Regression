irf130 test circuit
* This test tests the use of "options parser scale" 
*
* The point of this test is to make sure that if sampling 
* is applied to a scaled parameter, that it does the right 
* thing and applies the scaling every time it is updated.
*
* this version of the netlist is the reference version, so it does not use scale.
vd 3 1 0.5
vs 2 0 0
vg 4 0 10 pulse(0 10 300ns 50ns 50ns 400ns 1000ns)
vid 0 1 dc 0

m1 3 4 2 0 irf130 w=0.386e6u l='1.0e-6*agauss(2.5,0.25,1)'

.model irf130 nmos level=18
+ cv=1
+ cve=1
+ vto=3.5
+ rd= 0
+ rs= 0.005
+ lambda=0
+ m=3
+ sigma0=0
+ uo=230
+ vmax=4e4
+ delta=5
+ tox=50nm

.sampling useExpr=true

.options samples numsamples=10 seed=1923635719
+ outputs={i(vid)+0.5}
+ sample_type=lhs
+ stdoutput=false

.tran 0.5n 1u 0u 2n
.print tran precision=10 width=19 v(3) v(4) {i(vid)+0.5}

.options timeint reltol=1.0e-2 abstol=1.0e-7
.end

