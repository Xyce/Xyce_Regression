RAW File Output test for the Mutual Inductors.
************************************************************
* This test has two purposes:
*   1) Verify that the variable types (e.g., "current") and 
*      variable names are correct for the linear and
*      non-linear mutual inductors.  For the non-linear
*      mutual inductor, the m and r variables also appear and 
*      are listed as "voltage".
*
*   2) Verify that the data is actually correct for all of
*      the time-steps in the .RAW file output 
*
* The "gold" .RAW file output was generated by manually
* comparing that "gold" file with a .PRN file.  It was 
* generated for a limited set of fixed time-steps, so that
* a file comparison could be used to verify the test output's
* .RAW file against that "gold" .RAW file.
*
************************************************************  

*Linear mutual inductor
VS 1 0 SIN(0 169.7 60HZ)
R1 1 2 1K
R2 3 0 1K
L1 2 0 1mH
L2 3 0 1mH
K1 L1 L2 0.75

*Non-linear mutual inductor will be added later
Vprimary 0 node2 sin(0 115 60 0 0 0 )
xbr2 0 node2 node13 node14 bridge_rectifier2

.subckt bridge_rectifier2 pIn1 pIn2 sOut1 sOut2

Lprimary   pIn1 pIn2 495
Lsecondary node3 node4 34
Ktrans Lprimary Lsecondary 1.0 tMod
.model tMod CORE rvarscaling=1.0e6 factorms=1 MS=1.0e6 AREA=5.81

Rfeed node4 0 1000
Rtune node3 node5 0.1

dbridge1 sOut1  node5 dmod1
dbridge2 node5  sOut2 dmod1
dbridge3 sOut1  node4 dmod1
dbridge4 node4  sOut2 dmod1
.model dmod1 d CJ=1.0e-12 CJ0=1.0e-12

.ends

* simulation control
.OPTIONS OUTPUT INITIAL_INTERVAL=1ms
.TRAN 100US 25MS

* .PRINT statement is not actually used for .RAW output.
* It was included in the netslit so that the "gold" .RAW 
* file output could manually verified against a .PRN file
* during test development
.PRINT TRAN V(1) V(2) V(3) N(l1_branch) N(l2_branch) 
+ N(l:xbr2:primary_branch)  N(l:xbr2:secondary_branch)
+ V(node13) v(node14) v(2) I(vprimary) I(vs)
+ V(xbr2:node3) V(xbr2:node4) V(xbr2:node5)
+ N(xbr2:ymin!ktrans_m) N(xbr2:ymin!ktrans_r)
+ N(y:xbr2:min!ktrans_lprimary_branch) 
+ N(y:xbr2:min!ktrans_lsecondary_branch)
+ N(y:xbr2:min!ktrans_m) N(y:xbr2:min!ktrans_r)
+ N(ymil!k1_l1_branch) N(ymil!k1_l2_branch)


.END
