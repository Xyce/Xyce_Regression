Power test for S, SW and W devices (switches)
*
v1  1  0        PWL(0 0 1U 0 1.01U 5 2U 5 2.01U 0 3U 0 3.01U 5)
S1  2  1  3  0  VSW
W2  0  2  v3  ISW
v3  0  3        PWL (0 0 2U 0 2.01U 5)
r3  0  3        200
.MODEL VSW VSWITCH(RON=1 ROFF=1MEG VON=1 VOFF=0)
.MODEL ISW ISWITCH (ION=10mA IOFF=0mA RON=1 ROFF=1E6)

V4  4  0  PWL(0 0 1U 0 1.01U 5 2U 5 2.01U 0 3U 0 3.01U 5)
SW1 5  4  VSW ON CONTROL={V(3)}
SW2 0  5  ISW ON CONTROL={I(V3)} 

.options timeint method=trap
.options nonlin-tran rhstol=1.0e-7
.TRAN 0.02U 4U

* S1 and W2 should dissipate an equal amount of power.
* So, their individual power dissipation should also be "minus one-half" 
* of the power dissipation of V1.  Similar comments for SW1 and SW2 vs. V4.
.PRINT TRAN P(S1) W(S1) P(W2) W(W2) {V(2,1)*I(S1)} {V(0,2)*I(W2)} {-0.5*P(V1)} 
+ P(SW1) W(S1) P(SW2) W(SW2) {V(5,4)*I(SW1)} {V(0,5)*I(SW2)} {-0.5*P(V4)} 
+ V(1) V(2) I(S1) I(W2)
+ V(4) V(5) I(SW1) I(SW2)

.END
