Test "idvgh" from psp QA symmetric/nmos
*
* The PSP qa reference lists this test as:
*
*// Id-Vg @ Vs=0V, Vb=-1.0V, Vd=0.05 & 1.0V, SWIGATE=SWIMPACT=SWGIDL=1, SWJUNCAP=3
*test                        idvg0
*biases                      V(s)=0 V(b)=-1.0
*biasList                    V(d)=0.05,1.0
*biasSweep                   V(g)=-1.0,1.2,0.01
*outputs                     I(d) I(g) I(s) I(b)
*instanceParameters          W=10.0e-6 L=0.1e-6 AS=5e-12 AD=5e-12 PS=21e-6 PD=21e-6
*modelParameters             parameters/psp103_params
*modelParameters             SWIGATE=1 SWIMPACT=1 SWGIDL=1 SWJUNCAP=3
*
******
* PSP defines the drain, source, gate, and bulk currents as positive when they're into the 
* device, hence the goofy organization of these probe voltage sources.
*
*********

*idvg0 and idvgh share identical models and instances, only base bias is different.
.include "psp_nmos_idvg0.model"
M1 D G S B pspqan W=10.0e-6 L=0.1e-6 AS=5e-12 AD=5e-12 PS=21e-6 PD=21e-6

Vg G 0 DC 0v
Vd D 0 DC 0v
Vs S 0 DC 0v
Vb B 0 DC -1.0v

*Second transistor for finite differencing
Bdrain d2 0 V={V(d)}
Bgate g2 0  V={V(g)+((V(g)==0)?.00000001:(1e-8*abs(v(g))))}
Bsource s2 0 V={V(s)}
Bbulk b2 0 V={V(b)}

M2 D2 G2 S2 B2 pspqan W=10.0e-6 L=0.1e-6 AS=5e-12 AD=5e-12 PS=21e-6 PD=21e-6

.dc Vg -1 1.2 0.01  Vd LIST 0.05 1.0
.step TEMP LIST 27 -50 150
*COMP {N(M1:gm)-{((N(M2:ids)+N(M2:idedge)+N(M2:idb)-N(M2:igd))-(N(M1:ids)+N(M1:idedge)+N(M1:idb)-N(M1:igd)))/(V(g2)-V(g))}} abstol=1e-8
*COMP {((N(M2:ids)+N(M2:idedge)+N(M2:idb)-N(M2:igd))-(N(M1:ids)+N(M1:idedge)+N(M1:idb)-N(M1:igd)))/(V(g2)-V(g))} abstol=1e-8
* PSP "Ids" is only one term of the thing gm differentiates.
.print dc v(g) v(d) {N(M1:ids)+N(M1:idedge)+N(M1:idb)-N(M1:igd)}
+ {((N(M2:ids)+N(M2:idedge)+N(M2:idb)-N(M2:igd))-(N(M1:ids)+N(M1:idedge)+N(M1:idb)-N(M1:igd)))/(V(g2)-V(g))}
+ N(M1:gm)
+ {N(M1:gm)-{((N(M2:ids)+N(M2:idedge)+N(M2:idb)-N(M2:igd))-(N(M1:ids)+N(M1:idedge)+N(M1:idb)-N(M1:igd)))/(V(g2)-V(g))}}  N(M1:Vth) N(M1:Vds) N(M1:Vsb) N(M1:Vgs) N(M1:Vdss)
.end
