* Sensitivity of collector current to amplifier component
* This circuit was found  on page 298 of the book,
* "PSPICE and MATLAB for Electronics: An Integrated Approach" by John Okyere Attia.
*
* The relevant pages are excerpted in google books, and includes a printout of the
* PSPICE output.
*
.global_param VCCvalue=10V

VCC 4 0 DC {VCCvalue}
RB1 4 1 40k
RB2 1 0 10k
RE 2 0 1K
RC 5 3 6K
VM 4 5 DC 0; monitor collector current
Q1 3 1 2 Q2N2222 sw_et=0

.DC VCCvalue 1 10 0.4

.print dc v(4) I(VM)
.print sens v(4)


.SENS param=
+ Q2N2222:is,
+ Q2N2222:ibei,
+ Q2N2222:rci,
+ Q2N2222:mc,
+ Q2N2222:nf,
+ Q2N2222:tnom
+objfunc={I(VM)}

.options SENSITIVITY direct=1 adjoint=0  forcedevicefd=1  debuglevel=2

* VBIC model generated by sgp2vbic.pl from q2n2222 level 1 BJT model
.model q2n2222 npn
+ LEVEL=11  rcx=0.001 rci=0.0015 rbx=0.001 rbi=0 re=0.001 rb=0.001 rc=0.001
+ is=3.295e-14 nf=1 nr=1 fc=0.5 cje=0 pe=0.75 me=0.33 cjc=0 cjep=0 pc=0.75
+ mc=0.33 cjcp=0 ps=0.75 ms=0.001 ibei=3.295e-16 nei=1 iben=0 nen=1.5
+ ibci=3.295e-14 nci=1 ibcn=0 ncn=2 vef=134.605947186551 ver=6485118644.83438
+ ikf=0 ikr=0 tf=0 xtf=0 vtf=0 itf=0 tr=0 td=0 ea=1.11 eaie=1.11 eaic=1.11
+ eane=1.11 eanc=1.11 xis=3 xii=3 xin=3 kfn=0 afn=1 tnom=27
