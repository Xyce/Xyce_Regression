
* test for subcircuit instance parameters, when they refer to each other.
*
* this test also tests precedence rules for subcircuit parameters.   
* The resistor Rinside uses the parameter 'par3'.  It is defined in 3 places.  
* The one with highest priority is on the Xtest line.
*
.subckt simple in out PARAMS: par1=2.0 par2=2.0 par3='par1*par2*2.0'
.param par3=100.0
Rinside in out 'par3'
.ends

V1 1 0 1.0
R1 1 2 1.0
Xtest 2 0  simple par1=2.0 par2=3.0 par3='par1+par2'

.dc v1 1.0 1.0 1.0
.print dc v(1) {Xtest:Rinside:R}

