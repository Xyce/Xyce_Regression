Testing ill-formed .MEASURE lines
*********************************************************************
* Missing node specifier in I(), P() and W().    
* 
* See SON Bug 673
*
*
*
*
*
*********************************************************************
VS  1  0  SIN(0 1.0 1KHZ 0 0)
R1  1  0  100
.TRAN 0 1ms
.PRINT TRAN FORMAT=NOINDEX V(1) I(R1)

* bogo measure line that will cause a fatal error within
* the *makeOp() function in N_UTL_Op.C
.MEASURE TRAN MAX1 MAX I()
.MEASURE TRAN MAX1 MAX P()
.MEASURE TRAN MAX1 MAX W()

.END

