****************************************************
* Test Touchstone2 output using a 3-Port S-Parameter
* analysis.  This also tests:
* the cases where:
*
*   1) the ports have differing output impedances.
*
*   2) the .LIN line uses the default values, and hence
*      outputs Touchstone 2 format without generating
*      any warning messages.
*
* There is no .PRINT AC line.  So, there should
* not be any .AC output.
****************************************************

* RC ladder circuit
* Note that all ports (P devices) must use a common
* Reference Node, which is 0 here.
P1 1  0  port=1  z0=50
P2 12 0  port=2  z0=50
P3 5  0  port=3  Z0=100

C1 2 0 1e-2
Rgs 1 2 0.02

.subckt RCBlock IN OUT GND
R1 IN OUT 20
C1 IN OUT 1p
Cg1 OUT GND 1p
.ends

X1 2 3 0 RCBlock
X2 3 4 0 RCBlock
X3 4 5 0 RCBlock
X4 5 6 0 RCBlock
X5 6 7 0 RCBlock
X6 7 8 0 RCBlock
X7 8 9 0 RCBlock
X8 9 10 0 RCBlock
X9 10 11 0 RCBlock
X10 11 12 0 RCBlock

.AC DEC 10 10  1e5

* This .LIN line should use the defaults of FORMAT=TOUCHSTONE2
* and SPARCALC=1.  It explicitly sets LINTYPE=S.
.LIN LINTYPE=S

.END
