* Test syntax for function specified with .param keyword.
* Xyce functions were originally implemented with 
* the .func keyword, but some simulators specify 
* functions as a special type of .param.

* This test exercises multiple function params on the same line, 
* with a conventional parameter in the middle of the list, that has 
* a "naked" expression for its RHS.
*
* The old .func specification only allowed a single function per line.
*
* In this case the functions are NOT comma-separated, and the 
* functions have multiple arguments.  Also, in this case the parameter 
* "b" has parenthesis and commas as part of its specification of AGAUSS, 
* which is specified as a "naked" expression (ie, no single quotes or curly braces).
*
* This is a use case that potentially could confuse the parser, so it is a good test.
* Parens and commas can indicate (1) a separator between params 
* (but not in this case) and (2) function arguments (but not when 
* part of AGAUSS as in the case here).

.param a=1.0
.param ftest(x,y)={2*x+y}  b=agauss(12.0,1,1)  ftest2(x,y)={3*x+y}

v1 1 0 1.0
r1 1 2 {ftest(2.0,a)*b}
r2 2 0 {ftest2(2.0,a)*b}

.dc v1 1 1 1
.print dc v(1) v(2) {r1:r} {r2:r}

