module main;
initial $runXyceInSteps;
endmodule
