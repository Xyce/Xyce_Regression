*Test of parameter resolution
* This test used to pass Xyce 6.7 because of the early (and wrong)
* resolution that the pass 1 and pass MI used to make.  When bug 28
* was first fixed, the main netlist in this test case started to
* produce parameter resolution errors.  That's because it is a use
* case that had previously been untested in our test suite.

* That exposed limitations in the first approach to the bug 28 fix,
* requiring deeper modification.  This test case assures that we don't
* miss that sort of thing again.

* This netlist does not use the parameters at all, and serves as a baseline
* to which the main netlist in the test case can be compared, to make sure
* that it actually produces the CORRECT results when it resolves parameters.

.subckt transformer_v2 trans_start trans_end
.param pRHi = 0.34e-6
.param pL1 = 6.67e-6
.param pC1 = 2.4e-9
.param pCo = 28.9e-9
.param pL2 =4.65e-6
.param pC2 = 1.64e-15
.param pRLo = 0.233e-6
.param pRL1 = 47.6e-9
.param pRC1 = 0.26e-6
.param pRL2 = 0.2
.param pRC2 = 7.6

V_Meas_Trans_HV         TRANS_START     TRANS_HV        0
V_Meas_Trans_LV         TRANS_LV        TRANS_END       0

R_rhi        TRANS_HV    NODE1       pRHi
C1           NODE1       NODE3       pC1
RC1          NODE3       0           pRC1
L1           NODE1       NODE4       6.67e-6
RL1          NODE4       0           pRL1
Co           NODE1       NODE2       pCo
L2           NODE2       NODE5       4.65e-6
Ktrans       L1  L2  1.0
RL2          NODE5       0           pRL2
C2           NODE2       NODE6       pC2
RC2          NODE6       0           pRC2
RLo          NODE2       TRANS_LV    pRLo

.ends

xtest node1 node2 TRANSFORMER_V2 

r1 node1 0 100
r2 node2 0 100

vsrc node1 0 sin( 0 10.0 100k)

.tran 0 .1m
.print tran v(node1) v(node2)
.end

