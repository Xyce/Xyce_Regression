A test of the measure integral functionality
*******************************************************************************
*
* a few sources of different types
VS1  1  0  SIN(0 1.0 50HZ 0 0)
VP   2  0  PULSE( 0 100 0.2ms 0.2ms 0.2ms 1ms 2ms )
VS3  3  0  SIN(-0.5 1.0 250HZ 0 500)
VS4  4  0  SIN(0.5 -1.0 250HZ 0 500)

R1  1  0  100
R2  2  0  100
R3  3  0  100
R4  4  0  100

.TRAN 0  10ms
.PRINT TRAN FORMAT=NOINDEX V(1) V(2) V(3) V(4) V(1,0)

.measure tran intAll INTEGRAL v(1)
.measure tran int10All INTEGRAL v(1,0)
.measure tran intTop INTEG v(2)

* add TO-FROM modifiers
.measure tran sineHalfInterval Integ V(1) from=0 to=0.001

* mix in TDs before and after FROM value.
.measure tran sineTDbetween integ V(1) FROM=0 TO=0.005 TD=0.001
.measure tran sineTDbefore integ V(1) FROM=0.002 TO=0.005 TD=0.001

* these tests should return -1 and -100
.measure tran returnNegOne integ V(1) FROM=0.2e-3 TO=0.25e-3 TD=0.5e-3
.measure tran returnNeg100 integ V(1) FROM=0.2e-3 TO=0.25e-3 TD=0.5e-3 default_val=-100

* add tests for rise/fall/cross.  V3 and VS4 have a DC offset
* and are damped sinusoids
.measure tran intv3fall2 integ v(3) fall=2
.measure tran intv4rise1 integ v(4) rise=1
.measure tran intv3cross2 integ v(3) cross=2

* test LAST for rise/fall/cross
.measure tran int3falllast integ v(3) fall=last
.measure tran int4riselast integ v(4) rise=last
.measure tran int3crosslast integ v(3) cross=last

* test RFC_LEVEL keyword
.measure tran intv4Rise1RFClevel50 integral V(4) RFC_LEVEL=0.50 RISE=1
.measure tran intv4Fall1RFClevel50 integral V(4) RFC_LEVEL=0.50 FALL=1
.measure tran intv4Cross1RFClevel50 integral V(4) RFC_LEVEL=0.50 CROSS=1 

*test Failed measures for rise/fall/cross
.measure tran int3fallfail integ v(3) fall=25
.measure tran int4risefail integ v(4) rise=25
.measure tran intv3crossfail integ v(3) cross=25

.END

