Regression test to ensure that .STEP with .DATA can be applied to .param

.param testnorm={0.5K}
.param r1value={testnorm*2.0}

r2 1 0 7k
r1 1 2 {r1value}
v1 2 0 1000v

.dc v1 1000 1000 1
.print dc v(2) v(1)

.data eric
+ testnorm 
+ 0.5k 
+ 0.6k 
+ 0.7k
.enddata

.step data=eric

.end

