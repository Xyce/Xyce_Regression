Test for LIST capability in DC sweeps
*
* Eric Keiter, 9233.
* 8/29/04.
*
VT1 4 0 0V
R1  4 5 10
R2  5 0 5

.DC VT1 LIST  -17 12 188 5
.print DC V(4) V(5)

.END

