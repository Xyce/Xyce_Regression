************************************************
* T for warning for improperly formatted
* .ENDL line in a library file, that is still
* usable.
*
* See SON Bug 980 for more details.  Also this
* circuit is based on the example in the .LIB
* section of the Reference Guide.
************************************************

.LIB bogoLib2 high

V1 1 0 1
R1 1 2 {rval}

.DC V1 1 2 1
.PRINT DC V(1) V(2)

.END

