P-Channel Mosfet (Level 6) Circuit
************************************************************** 
VDD 2 0 DC 5V
R1 2 1 50K
R2 1 0 50K
RD 4 0 7.5K
VMON 3 4 0
M1 3 1 2 2 PFET L=10U W=160U
.MODEL PFET PMOS(LEVEL=6 KP=25U VTO=-0.8V)

.DC VDD 0 5 0.01
.PRINT DC V(2) I(VMON) V(2,3) V(2,1)
.END
