********************************************************
* Test FORMAT=GNUPLOT with .STEP.  This should 
* produce the same .prn file as FORMAT=STD, but with
* two blank lines before steps 1,2, ... N-1.  Note that
* first step is "step 0".  In this netlist, N is 4.
*******************************************************

V1 1 0 SIN(0 1 1)
R1 1 2 1
R2 2 0 1

* step over two variables
.STEP R1 1 2 1 
.STEP R2 3 4 1

.OPTIONS OUTPUT INITIAL_INTERVAL=0.01
.PRINT TRAN FORMAT=GNUPLOT R1:R R2:R V(1) V(2)
.TRAN 0 1

.END
