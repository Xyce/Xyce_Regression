branched cable simulation - rallpack 2 


.tran 0 0.25  
.options linsol type=klu
*.options timeint maxord=1
*.options output initial_interval=1.0e-3

* rallpack 2 calls for a steady current input.  But we need to use PULSE so
* that the current will be off during dcop calculation
Iin 0 n0 PULSE( 0 1.0e-10 1.0e-12 0.0 0.0 1.0e10 1.0e10)

* membrane properties (from rallpack2 README file)
* Ra = 1.0 ohms meter
* Rm = 4.0 ohms meter^2
* Cm = 0.01 F/m^2
* Em = -0.065 Volts
* confirmed that these are the same parameter values as for rallpack1

* axial resistance 1 ohms m
.param Ra = 1.0	; [ohm m]

* specific membrane capacitance 0.01 F/m^2 
.param memC = { 0.01 } ; [F/m^2]

* leak current has membrane resistivity of 4 ohms m^2, with reversal potential of -65mV
.param rm = { 4.0 }    ; [ohm m^2]
.param memG = { 1 / rm }                  ; [1/(ohm m^2)]
.param revE = -0.065                      ; [V]

* neuron model - this just specifies electrophysiological parameters; size parameters will vary
.model segParams neuron level=6 ionchannelmodel=passive cMem={memC}  gMem={memG} vRest={revE} R={Ra} N=1
 
  
yneuron neuron00 n0 n00 segParams L={3.20000e-05} A={8.00000e-06}
yneuron neuron000 n00 n000 segParams L={2.54000e-05} A={5.04000e-06}
yneuron neuron0000 n000 n0000 segParams L={2.01600e-05} A={3.17500e-06}
yneuron neuron00000 n0000 n00000 segParams L={1.60000e-05} A={2.00000e-06}
yneuron neuron000000 n00000 n000000 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0000000 n000000 n0000000 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00000000 n0000000 n00000000 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000000000 n00000000 n000000000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000000000 n000000000 n0000000000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000000000 n0000000000 n00000000000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000000001 n0000000000 n00000000001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000000001 n000000000 n0000000001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000000010 n0000000001 n00000000010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000000011 n0000000001 n00000000011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000000001 n00000000 n000000001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000000010 n000000001 n0000000010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000000100 n0000000010 n00000000100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000000101 n0000000010 n00000000101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000000011 n000000001 n0000000011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000000110 n0000000011 n00000000110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000000111 n0000000011 n00000000111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000001 n0000000 n00000001 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000000010 n00000001 n000000010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000000100 n000000010 n0000000100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000001000 n0000000100 n00000001000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000001001 n0000000100 n00000001001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000000101 n000000010 n0000000101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000001010 n0000000101 n00000001010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000001011 n0000000101 n00000001011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000000011 n00000001 n000000011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000000110 n000000011 n0000000110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000001100 n0000000110 n00000001100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000001101 n0000000110 n00000001101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000000111 n000000011 n0000000111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000001110 n0000000111 n00000001110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000001111 n0000000111 n00000001111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000001 n000000 n0000001 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00000010 n0000001 n00000010 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000000100 n00000010 n000000100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000001000 n000000100 n0000001000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000010000 n0000001000 n00000010000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000010001 n0000001000 n00000010001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000001001 n000000100 n0000001001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000010010 n0000001001 n00000010010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000010011 n0000001001 n00000010011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000000101 n00000010 n000000101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000001010 n000000101 n0000001010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000010100 n0000001010 n00000010100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000010101 n0000001010 n00000010101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000001011 n000000101 n0000001011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000010110 n0000001011 n00000010110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000010111 n0000001011 n00000010111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000011 n0000001 n00000011 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000000110 n00000011 n000000110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000001100 n000000110 n0000001100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000011000 n0000001100 n00000011000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000011001 n0000001100 n00000011001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000001101 n000000110 n0000001101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000011010 n0000001101 n00000011010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000011011 n0000001101 n00000011011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000000111 n00000011 n000000111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000001110 n000000111 n0000001110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000011100 n0000001110 n00000011100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000011101 n0000001110 n00000011101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000001111 n000000111 n0000001111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000011110 n0000001111 n00000011110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000011111 n0000001111 n00000011111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000001 n00000 n000001 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0000010 n000001 n0000010 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00000100 n0000010 n00000100 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000001000 n00000100 n000001000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000010000 n000001000 n0000010000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000100000 n0000010000 n00000100000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000100001 n0000010000 n00000100001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000010001 n000001000 n0000010001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000100010 n0000010001 n00000100010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000100011 n0000010001 n00000100011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000001001 n00000100 n000001001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000010010 n000001001 n0000010010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000100100 n0000010010 n00000100100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000100101 n0000010010 n00000100101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000010011 n000001001 n0000010011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000100110 n0000010011 n00000100110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000100111 n0000010011 n00000100111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000101 n0000010 n00000101 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000001010 n00000101 n000001010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000010100 n000001010 n0000010100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000101000 n0000010100 n00000101000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000101001 n0000010100 n00000101001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000010101 n000001010 n0000010101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000101010 n0000010101 n00000101010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000101011 n0000010101 n00000101011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000001011 n00000101 n000001011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000010110 n000001011 n0000010110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000101100 n0000010110 n00000101100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000101101 n0000010110 n00000101101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000010111 n000001011 n0000010111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000101110 n0000010111 n00000101110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000101111 n0000010111 n00000101111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000011 n000001 n0000011 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00000110 n0000011 n00000110 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000001100 n00000110 n000001100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000011000 n000001100 n0000011000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000110000 n0000011000 n00000110000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000110001 n0000011000 n00000110001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000011001 n000001100 n0000011001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000110010 n0000011001 n00000110010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000110011 n0000011001 n00000110011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000001101 n00000110 n000001101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000011010 n000001101 n0000011010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000110100 n0000011010 n00000110100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000110101 n0000011010 n00000110101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000011011 n000001101 n0000011011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000110110 n0000011011 n00000110110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000110111 n0000011011 n00000110111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000111 n0000011 n00000111 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000001110 n00000111 n000001110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000011100 n000001110 n0000011100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000111000 n0000011100 n00000111000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000111001 n0000011100 n00000111001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000011101 n000001110 n0000011101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000111010 n0000011101 n00000111010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000111011 n0000011101 n00000111011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000001111 n00000111 n000001111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000011110 n000001111 n0000011110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000111100 n0000011110 n00000111100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000111101 n0000011110 n00000111101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000011111 n000001111 n0000011111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00000111110 n0000011111 n00000111110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00000111111 n0000011111 n00000111111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001 n0000 n00001 segParams L={1.60000e-05} A={2.00000e-06}
yneuron neuron000010 n00001 n000010 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0000100 n000010 n0000100 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00001000 n0000100 n00001000 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000010000 n00001000 n000010000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000100000 n000010000 n0000100000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001000000 n0000100000 n00001000000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001000001 n0000100000 n00001000001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000100001 n000010000 n0000100001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001000010 n0000100001 n00001000010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001000011 n0000100001 n00001000011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000010001 n00001000 n000010001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000100010 n000010001 n0000100010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001000100 n0000100010 n00001000100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001000101 n0000100010 n00001000101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000100011 n000010001 n0000100011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001000110 n0000100011 n00001000110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001000111 n0000100011 n00001000111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001001 n0000100 n00001001 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000010010 n00001001 n000010010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000100100 n000010010 n0000100100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001001000 n0000100100 n00001001000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001001001 n0000100100 n00001001001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000100101 n000010010 n0000100101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001001010 n0000100101 n00001001010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001001011 n0000100101 n00001001011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000010011 n00001001 n000010011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000100110 n000010011 n0000100110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001001100 n0000100110 n00001001100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001001101 n0000100110 n00001001101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000100111 n000010011 n0000100111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001001110 n0000100111 n00001001110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001001111 n0000100111 n00001001111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000101 n000010 n0000101 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00001010 n0000101 n00001010 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000010100 n00001010 n000010100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000101000 n000010100 n0000101000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001010000 n0000101000 n00001010000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001010001 n0000101000 n00001010001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000101001 n000010100 n0000101001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001010010 n0000101001 n00001010010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001010011 n0000101001 n00001010011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000010101 n00001010 n000010101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000101010 n000010101 n0000101010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001010100 n0000101010 n00001010100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001010101 n0000101010 n00001010101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000101011 n000010101 n0000101011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001010110 n0000101011 n00001010110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001010111 n0000101011 n00001010111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001011 n0000101 n00001011 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000010110 n00001011 n000010110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000101100 n000010110 n0000101100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001011000 n0000101100 n00001011000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001011001 n0000101100 n00001011001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000101101 n000010110 n0000101101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001011010 n0000101101 n00001011010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001011011 n0000101101 n00001011011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000010111 n00001011 n000010111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000101110 n000010111 n0000101110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001011100 n0000101110 n00001011100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001011101 n0000101110 n00001011101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000101111 n000010111 n0000101111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001011110 n0000101111 n00001011110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001011111 n0000101111 n00001011111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000011 n00001 n000011 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0000110 n000011 n0000110 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00001100 n0000110 n00001100 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000011000 n00001100 n000011000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000110000 n000011000 n0000110000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001100000 n0000110000 n00001100000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001100001 n0000110000 n00001100001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000110001 n000011000 n0000110001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001100010 n0000110001 n00001100010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001100011 n0000110001 n00001100011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000011001 n00001100 n000011001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000110010 n000011001 n0000110010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001100100 n0000110010 n00001100100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001100101 n0000110010 n00001100101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000110011 n000011001 n0000110011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001100110 n0000110011 n00001100110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001100111 n0000110011 n00001100111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001101 n0000110 n00001101 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000011010 n00001101 n000011010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000110100 n000011010 n0000110100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001101000 n0000110100 n00001101000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001101001 n0000110100 n00001101001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000110101 n000011010 n0000110101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001101010 n0000110101 n00001101010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001101011 n0000110101 n00001101011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000011011 n00001101 n000011011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000110110 n000011011 n0000110110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001101100 n0000110110 n00001101100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001101101 n0000110110 n00001101101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000110111 n000011011 n0000110111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001101110 n0000110111 n00001101110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001101111 n0000110111 n00001101111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000111 n000011 n0000111 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00001110 n0000111 n00001110 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000011100 n00001110 n000011100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000111000 n000011100 n0000111000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001110000 n0000111000 n00001110000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001110001 n0000111000 n00001110001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000111001 n000011100 n0000111001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001110010 n0000111001 n00001110010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001110011 n0000111001 n00001110011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000011101 n00001110 n000011101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000111010 n000011101 n0000111010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001110100 n0000111010 n00001110100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001110101 n0000111010 n00001110101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000111011 n000011101 n0000111011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001110110 n0000111011 n00001110110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001110111 n0000111011 n00001110111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001111 n0000111 n00001111 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000011110 n00001111 n000011110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000111100 n000011110 n0000111100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001111000 n0000111100 n00001111000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001111001 n0000111100 n00001111001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000111101 n000011110 n0000111101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001111010 n0000111101 n00001111010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001111011 n0000111101 n00001111011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000011111 n00001111 n000011111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0000111110 n000011111 n0000111110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001111100 n0000111110 n00001111100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001111101 n0000111110 n00001111101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0000111111 n000011111 n0000111111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00001111110 n0000111111 n00001111110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00001111111 n0000111111 n00001111111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001 n000 n0001 segParams L={2.01600e-05} A={3.17500e-06}
yneuron neuron00010 n0001 n00010 segParams L={1.60000e-05} A={2.00000e-06}
yneuron neuron000100 n00010 n000100 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0001000 n000100 n0001000 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00010000 n0001000 n00010000 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000100000 n00010000 n000100000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001000000 n000100000 n0001000000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010000000 n0001000000 n00010000000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010000001 n0001000000 n00010000001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001000001 n000100000 n0001000001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010000010 n0001000001 n00010000010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010000011 n0001000001 n00010000011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000100001 n00010000 n000100001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001000010 n000100001 n0001000010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010000100 n0001000010 n00010000100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010000101 n0001000010 n00010000101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001000011 n000100001 n0001000011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010000110 n0001000011 n00010000110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010000111 n0001000011 n00010000111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010001 n0001000 n00010001 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000100010 n00010001 n000100010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001000100 n000100010 n0001000100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010001000 n0001000100 n00010001000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010001001 n0001000100 n00010001001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001000101 n000100010 n0001000101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010001010 n0001000101 n00010001010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010001011 n0001000101 n00010001011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000100011 n00010001 n000100011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001000110 n000100011 n0001000110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010001100 n0001000110 n00010001100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010001101 n0001000110 n00010001101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001000111 n000100011 n0001000111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010001110 n0001000111 n00010001110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010001111 n0001000111 n00010001111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001001 n000100 n0001001 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00010010 n0001001 n00010010 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000100100 n00010010 n000100100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001001000 n000100100 n0001001000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010010000 n0001001000 n00010010000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010010001 n0001001000 n00010010001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001001001 n000100100 n0001001001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010010010 n0001001001 n00010010010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010010011 n0001001001 n00010010011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000100101 n00010010 n000100101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001001010 n000100101 n0001001010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010010100 n0001001010 n00010010100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010010101 n0001001010 n00010010101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001001011 n000100101 n0001001011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010010110 n0001001011 n00010010110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010010111 n0001001011 n00010010111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010011 n0001001 n00010011 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000100110 n00010011 n000100110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001001100 n000100110 n0001001100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010011000 n0001001100 n00010011000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010011001 n0001001100 n00010011001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001001101 n000100110 n0001001101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010011010 n0001001101 n00010011010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010011011 n0001001101 n00010011011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000100111 n00010011 n000100111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001001110 n000100111 n0001001110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010011100 n0001001110 n00010011100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010011101 n0001001110 n00010011101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001001111 n000100111 n0001001111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010011110 n0001001111 n00010011110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010011111 n0001001111 n00010011111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000101 n00010 n000101 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0001010 n000101 n0001010 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00010100 n0001010 n00010100 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000101000 n00010100 n000101000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001010000 n000101000 n0001010000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010100000 n0001010000 n00010100000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010100001 n0001010000 n00010100001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001010001 n000101000 n0001010001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010100010 n0001010001 n00010100010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010100011 n0001010001 n00010100011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000101001 n00010100 n000101001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001010010 n000101001 n0001010010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010100100 n0001010010 n00010100100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010100101 n0001010010 n00010100101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001010011 n000101001 n0001010011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010100110 n0001010011 n00010100110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010100111 n0001010011 n00010100111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010101 n0001010 n00010101 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000101010 n00010101 n000101010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001010100 n000101010 n0001010100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010101000 n0001010100 n00010101000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010101001 n0001010100 n00010101001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001010101 n000101010 n0001010101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010101010 n0001010101 n00010101010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010101011 n0001010101 n00010101011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000101011 n00010101 n000101011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001010110 n000101011 n0001010110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010101100 n0001010110 n00010101100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010101101 n0001010110 n00010101101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001010111 n000101011 n0001010111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010101110 n0001010111 n00010101110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010101111 n0001010111 n00010101111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001011 n000101 n0001011 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00010110 n0001011 n00010110 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000101100 n00010110 n000101100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001011000 n000101100 n0001011000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010110000 n0001011000 n00010110000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010110001 n0001011000 n00010110001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001011001 n000101100 n0001011001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010110010 n0001011001 n00010110010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010110011 n0001011001 n00010110011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000101101 n00010110 n000101101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001011010 n000101101 n0001011010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010110100 n0001011010 n00010110100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010110101 n0001011010 n00010110101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001011011 n000101101 n0001011011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010110110 n0001011011 n00010110110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010110111 n0001011011 n00010110111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010111 n0001011 n00010111 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000101110 n00010111 n000101110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001011100 n000101110 n0001011100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010111000 n0001011100 n00010111000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010111001 n0001011100 n00010111001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001011101 n000101110 n0001011101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010111010 n0001011101 n00010111010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010111011 n0001011101 n00010111011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000101111 n00010111 n000101111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001011110 n000101111 n0001011110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010111100 n0001011110 n00010111100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010111101 n0001011110 n00010111101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001011111 n000101111 n0001011111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00010111110 n0001011111 n00010111110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00010111111 n0001011111 n00010111111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011 n0001 n00011 segParams L={1.60000e-05} A={2.00000e-06}
yneuron neuron000110 n00011 n000110 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0001100 n000110 n0001100 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00011000 n0001100 n00011000 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000110000 n00011000 n000110000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001100000 n000110000 n0001100000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011000000 n0001100000 n00011000000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011000001 n0001100000 n00011000001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001100001 n000110000 n0001100001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011000010 n0001100001 n00011000010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011000011 n0001100001 n00011000011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000110001 n00011000 n000110001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001100010 n000110001 n0001100010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011000100 n0001100010 n00011000100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011000101 n0001100010 n00011000101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001100011 n000110001 n0001100011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011000110 n0001100011 n00011000110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011000111 n0001100011 n00011000111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011001 n0001100 n00011001 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000110010 n00011001 n000110010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001100100 n000110010 n0001100100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011001000 n0001100100 n00011001000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011001001 n0001100100 n00011001001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001100101 n000110010 n0001100101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011001010 n0001100101 n00011001010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011001011 n0001100101 n00011001011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000110011 n00011001 n000110011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001100110 n000110011 n0001100110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011001100 n0001100110 n00011001100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011001101 n0001100110 n00011001101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001100111 n000110011 n0001100111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011001110 n0001100111 n00011001110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011001111 n0001100111 n00011001111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001101 n000110 n0001101 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00011010 n0001101 n00011010 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000110100 n00011010 n000110100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001101000 n000110100 n0001101000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011010000 n0001101000 n00011010000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011010001 n0001101000 n00011010001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001101001 n000110100 n0001101001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011010010 n0001101001 n00011010010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011010011 n0001101001 n00011010011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000110101 n00011010 n000110101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001101010 n000110101 n0001101010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011010100 n0001101010 n00011010100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011010101 n0001101010 n00011010101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001101011 n000110101 n0001101011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011010110 n0001101011 n00011010110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011010111 n0001101011 n00011010111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011011 n0001101 n00011011 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000110110 n00011011 n000110110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001101100 n000110110 n0001101100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011011000 n0001101100 n00011011000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011011001 n0001101100 n00011011001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001101101 n000110110 n0001101101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011011010 n0001101101 n00011011010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011011011 n0001101101 n00011011011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000110111 n00011011 n000110111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001101110 n000110111 n0001101110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011011100 n0001101110 n00011011100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011011101 n0001101110 n00011011101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001101111 n000110111 n0001101111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011011110 n0001101111 n00011011110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011011111 n0001101111 n00011011111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000111 n00011 n000111 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0001110 n000111 n0001110 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00011100 n0001110 n00011100 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000111000 n00011100 n000111000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001110000 n000111000 n0001110000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011100000 n0001110000 n00011100000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011100001 n0001110000 n00011100001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001110001 n000111000 n0001110001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011100010 n0001110001 n00011100010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011100011 n0001110001 n00011100011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000111001 n00011100 n000111001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001110010 n000111001 n0001110010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011100100 n0001110010 n00011100100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011100101 n0001110010 n00011100101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001110011 n000111001 n0001110011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011100110 n0001110011 n00011100110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011100111 n0001110011 n00011100111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011101 n0001110 n00011101 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000111010 n00011101 n000111010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001110100 n000111010 n0001110100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011101000 n0001110100 n00011101000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011101001 n0001110100 n00011101001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001110101 n000111010 n0001110101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011101010 n0001110101 n00011101010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011101011 n0001110101 n00011101011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000111011 n00011101 n000111011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001110110 n000111011 n0001110110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011101100 n0001110110 n00011101100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011101101 n0001110110 n00011101101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001110111 n000111011 n0001110111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011101110 n0001110111 n00011101110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011101111 n0001110111 n00011101111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001111 n000111 n0001111 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00011110 n0001111 n00011110 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000111100 n00011110 n000111100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001111000 n000111100 n0001111000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011110000 n0001111000 n00011110000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011110001 n0001111000 n00011110001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001111001 n000111100 n0001111001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011110010 n0001111001 n00011110010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011110011 n0001111001 n00011110011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000111101 n00011110 n000111101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001111010 n000111101 n0001111010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011110100 n0001111010 n00011110100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011110101 n0001111010 n00011110101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001111011 n000111101 n0001111011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011110110 n0001111011 n00011110110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011110111 n0001111011 n00011110111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011111 n0001111 n00011111 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron000111110 n00011111 n000111110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001111100 n000111110 n0001111100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011111000 n0001111100 n00011111000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011111001 n0001111100 n00011111001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001111101 n000111110 n0001111101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011111010 n0001111101 n00011111010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011111011 n0001111101 n00011111011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron000111111 n00011111 n000111111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0001111110 n000111111 n0001111110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011111100 n0001111110 n00011111100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011111101 n0001111110 n00011111101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0001111111 n000111111 n0001111111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00011111110 n0001111111 n00011111110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00011111111 n0001111111 n00011111111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001 n00 n001 segParams L={2.54000e-05} A={5.04000e-06}
yneuron neuron0010 n001 n0010 segParams L={2.01600e-05} A={3.17500e-06}
yneuron neuron00100 n0010 n00100 segParams L={1.60000e-05} A={2.00000e-06}
yneuron neuron001000 n00100 n001000 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0010000 n001000 n0010000 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00100000 n0010000 n00100000 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001000000 n00100000 n001000000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010000000 n001000000 n0010000000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100000000 n0010000000 n00100000000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100000001 n0010000000 n00100000001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010000001 n001000000 n0010000001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100000010 n0010000001 n00100000010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100000011 n0010000001 n00100000011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001000001 n00100000 n001000001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010000010 n001000001 n0010000010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100000100 n0010000010 n00100000100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100000101 n0010000010 n00100000101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010000011 n001000001 n0010000011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100000110 n0010000011 n00100000110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100000111 n0010000011 n00100000111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100001 n0010000 n00100001 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001000010 n00100001 n001000010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010000100 n001000010 n0010000100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100001000 n0010000100 n00100001000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100001001 n0010000100 n00100001001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010000101 n001000010 n0010000101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100001010 n0010000101 n00100001010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100001011 n0010000101 n00100001011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001000011 n00100001 n001000011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010000110 n001000011 n0010000110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100001100 n0010000110 n00100001100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100001101 n0010000110 n00100001101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010000111 n001000011 n0010000111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100001110 n0010000111 n00100001110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100001111 n0010000111 n00100001111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010001 n001000 n0010001 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00100010 n0010001 n00100010 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001000100 n00100010 n001000100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010001000 n001000100 n0010001000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100010000 n0010001000 n00100010000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100010001 n0010001000 n00100010001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010001001 n001000100 n0010001001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100010010 n0010001001 n00100010010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100010011 n0010001001 n00100010011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001000101 n00100010 n001000101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010001010 n001000101 n0010001010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100010100 n0010001010 n00100010100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100010101 n0010001010 n00100010101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010001011 n001000101 n0010001011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100010110 n0010001011 n00100010110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100010111 n0010001011 n00100010111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100011 n0010001 n00100011 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001000110 n00100011 n001000110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010001100 n001000110 n0010001100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100011000 n0010001100 n00100011000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100011001 n0010001100 n00100011001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010001101 n001000110 n0010001101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100011010 n0010001101 n00100011010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100011011 n0010001101 n00100011011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001000111 n00100011 n001000111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010001110 n001000111 n0010001110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100011100 n0010001110 n00100011100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100011101 n0010001110 n00100011101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010001111 n001000111 n0010001111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100011110 n0010001111 n00100011110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100011111 n0010001111 n00100011111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001001 n00100 n001001 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0010010 n001001 n0010010 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00100100 n0010010 n00100100 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001001000 n00100100 n001001000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010010000 n001001000 n0010010000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100100000 n0010010000 n00100100000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100100001 n0010010000 n00100100001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010010001 n001001000 n0010010001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100100010 n0010010001 n00100100010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100100011 n0010010001 n00100100011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001001001 n00100100 n001001001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010010010 n001001001 n0010010010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100100100 n0010010010 n00100100100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100100101 n0010010010 n00100100101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010010011 n001001001 n0010010011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100100110 n0010010011 n00100100110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100100111 n0010010011 n00100100111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100101 n0010010 n00100101 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001001010 n00100101 n001001010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010010100 n001001010 n0010010100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100101000 n0010010100 n00100101000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100101001 n0010010100 n00100101001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010010101 n001001010 n0010010101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100101010 n0010010101 n00100101010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100101011 n0010010101 n00100101011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001001011 n00100101 n001001011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010010110 n001001011 n0010010110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100101100 n0010010110 n00100101100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100101101 n0010010110 n00100101101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010010111 n001001011 n0010010111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100101110 n0010010111 n00100101110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100101111 n0010010111 n00100101111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010011 n001001 n0010011 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00100110 n0010011 n00100110 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001001100 n00100110 n001001100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010011000 n001001100 n0010011000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100110000 n0010011000 n00100110000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100110001 n0010011000 n00100110001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010011001 n001001100 n0010011001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100110010 n0010011001 n00100110010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100110011 n0010011001 n00100110011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001001101 n00100110 n001001101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010011010 n001001101 n0010011010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100110100 n0010011010 n00100110100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100110101 n0010011010 n00100110101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010011011 n001001101 n0010011011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100110110 n0010011011 n00100110110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100110111 n0010011011 n00100110111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100111 n0010011 n00100111 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001001110 n00100111 n001001110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010011100 n001001110 n0010011100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100111000 n0010011100 n00100111000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100111001 n0010011100 n00100111001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010011101 n001001110 n0010011101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100111010 n0010011101 n00100111010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100111011 n0010011101 n00100111011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001001111 n00100111 n001001111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010011110 n001001111 n0010011110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100111100 n0010011110 n00100111100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100111101 n0010011110 n00100111101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010011111 n001001111 n0010011111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00100111110 n0010011111 n00100111110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00100111111 n0010011111 n00100111111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101 n0010 n00101 segParams L={1.60000e-05} A={2.00000e-06}
yneuron neuron001010 n00101 n001010 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0010100 n001010 n0010100 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00101000 n0010100 n00101000 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001010000 n00101000 n001010000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010100000 n001010000 n0010100000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101000000 n0010100000 n00101000000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101000001 n0010100000 n00101000001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010100001 n001010000 n0010100001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101000010 n0010100001 n00101000010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101000011 n0010100001 n00101000011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001010001 n00101000 n001010001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010100010 n001010001 n0010100010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101000100 n0010100010 n00101000100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101000101 n0010100010 n00101000101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010100011 n001010001 n0010100011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101000110 n0010100011 n00101000110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101000111 n0010100011 n00101000111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101001 n0010100 n00101001 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001010010 n00101001 n001010010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010100100 n001010010 n0010100100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101001000 n0010100100 n00101001000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101001001 n0010100100 n00101001001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010100101 n001010010 n0010100101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101001010 n0010100101 n00101001010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101001011 n0010100101 n00101001011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001010011 n00101001 n001010011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010100110 n001010011 n0010100110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101001100 n0010100110 n00101001100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101001101 n0010100110 n00101001101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010100111 n001010011 n0010100111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101001110 n0010100111 n00101001110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101001111 n0010100111 n00101001111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010101 n001010 n0010101 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00101010 n0010101 n00101010 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001010100 n00101010 n001010100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010101000 n001010100 n0010101000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101010000 n0010101000 n00101010000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101010001 n0010101000 n00101010001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010101001 n001010100 n0010101001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101010010 n0010101001 n00101010010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101010011 n0010101001 n00101010011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001010101 n00101010 n001010101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010101010 n001010101 n0010101010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101010100 n0010101010 n00101010100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101010101 n0010101010 n00101010101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010101011 n001010101 n0010101011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101010110 n0010101011 n00101010110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101010111 n0010101011 n00101010111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101011 n0010101 n00101011 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001010110 n00101011 n001010110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010101100 n001010110 n0010101100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101011000 n0010101100 n00101011000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101011001 n0010101100 n00101011001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010101101 n001010110 n0010101101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101011010 n0010101101 n00101011010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101011011 n0010101101 n00101011011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001010111 n00101011 n001010111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010101110 n001010111 n0010101110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101011100 n0010101110 n00101011100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101011101 n0010101110 n00101011101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010101111 n001010111 n0010101111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101011110 n0010101111 n00101011110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101011111 n0010101111 n00101011111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001011 n00101 n001011 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0010110 n001011 n0010110 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00101100 n0010110 n00101100 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001011000 n00101100 n001011000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010110000 n001011000 n0010110000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101100000 n0010110000 n00101100000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101100001 n0010110000 n00101100001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010110001 n001011000 n0010110001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101100010 n0010110001 n00101100010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101100011 n0010110001 n00101100011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001011001 n00101100 n001011001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010110010 n001011001 n0010110010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101100100 n0010110010 n00101100100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101100101 n0010110010 n00101100101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010110011 n001011001 n0010110011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101100110 n0010110011 n00101100110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101100111 n0010110011 n00101100111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101101 n0010110 n00101101 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001011010 n00101101 n001011010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010110100 n001011010 n0010110100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101101000 n0010110100 n00101101000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101101001 n0010110100 n00101101001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010110101 n001011010 n0010110101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101101010 n0010110101 n00101101010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101101011 n0010110101 n00101101011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001011011 n00101101 n001011011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010110110 n001011011 n0010110110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101101100 n0010110110 n00101101100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101101101 n0010110110 n00101101101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010110111 n001011011 n0010110111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101101110 n0010110111 n00101101110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101101111 n0010110111 n00101101111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010111 n001011 n0010111 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00101110 n0010111 n00101110 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001011100 n00101110 n001011100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010111000 n001011100 n0010111000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101110000 n0010111000 n00101110000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101110001 n0010111000 n00101110001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010111001 n001011100 n0010111001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101110010 n0010111001 n00101110010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101110011 n0010111001 n00101110011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001011101 n00101110 n001011101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010111010 n001011101 n0010111010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101110100 n0010111010 n00101110100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101110101 n0010111010 n00101110101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010111011 n001011101 n0010111011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101110110 n0010111011 n00101110110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101110111 n0010111011 n00101110111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101111 n0010111 n00101111 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001011110 n00101111 n001011110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010111100 n001011110 n0010111100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101111000 n0010111100 n00101111000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101111001 n0010111100 n00101111001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010111101 n001011110 n0010111101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101111010 n0010111101 n00101111010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101111011 n0010111101 n00101111011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001011111 n00101111 n001011111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0010111110 n001011111 n0010111110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101111100 n0010111110 n00101111100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101111101 n0010111110 n00101111101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0010111111 n001011111 n0010111111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00101111110 n0010111111 n00101111110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00101111111 n0010111111 n00101111111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011 n001 n0011 segParams L={2.01600e-05} A={3.17500e-06}
yneuron neuron00110 n0011 n00110 segParams L={1.60000e-05} A={2.00000e-06}
yneuron neuron001100 n00110 n001100 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0011000 n001100 n0011000 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00110000 n0011000 n00110000 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001100000 n00110000 n001100000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011000000 n001100000 n0011000000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110000000 n0011000000 n00110000000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110000001 n0011000000 n00110000001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011000001 n001100000 n0011000001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110000010 n0011000001 n00110000010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110000011 n0011000001 n00110000011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001100001 n00110000 n001100001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011000010 n001100001 n0011000010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110000100 n0011000010 n00110000100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110000101 n0011000010 n00110000101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011000011 n001100001 n0011000011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110000110 n0011000011 n00110000110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110000111 n0011000011 n00110000111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110001 n0011000 n00110001 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001100010 n00110001 n001100010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011000100 n001100010 n0011000100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110001000 n0011000100 n00110001000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110001001 n0011000100 n00110001001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011000101 n001100010 n0011000101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110001010 n0011000101 n00110001010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110001011 n0011000101 n00110001011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001100011 n00110001 n001100011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011000110 n001100011 n0011000110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110001100 n0011000110 n00110001100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110001101 n0011000110 n00110001101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011000111 n001100011 n0011000111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110001110 n0011000111 n00110001110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110001111 n0011000111 n00110001111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011001 n001100 n0011001 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00110010 n0011001 n00110010 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001100100 n00110010 n001100100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011001000 n001100100 n0011001000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110010000 n0011001000 n00110010000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110010001 n0011001000 n00110010001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011001001 n001100100 n0011001001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110010010 n0011001001 n00110010010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110010011 n0011001001 n00110010011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001100101 n00110010 n001100101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011001010 n001100101 n0011001010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110010100 n0011001010 n00110010100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110010101 n0011001010 n00110010101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011001011 n001100101 n0011001011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110010110 n0011001011 n00110010110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110010111 n0011001011 n00110010111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110011 n0011001 n00110011 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001100110 n00110011 n001100110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011001100 n001100110 n0011001100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110011000 n0011001100 n00110011000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110011001 n0011001100 n00110011001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011001101 n001100110 n0011001101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110011010 n0011001101 n00110011010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110011011 n0011001101 n00110011011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001100111 n00110011 n001100111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011001110 n001100111 n0011001110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110011100 n0011001110 n00110011100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110011101 n0011001110 n00110011101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011001111 n001100111 n0011001111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110011110 n0011001111 n00110011110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110011111 n0011001111 n00110011111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001101 n00110 n001101 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0011010 n001101 n0011010 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00110100 n0011010 n00110100 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001101000 n00110100 n001101000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011010000 n001101000 n0011010000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110100000 n0011010000 n00110100000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110100001 n0011010000 n00110100001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011010001 n001101000 n0011010001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110100010 n0011010001 n00110100010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110100011 n0011010001 n00110100011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001101001 n00110100 n001101001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011010010 n001101001 n0011010010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110100100 n0011010010 n00110100100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110100101 n0011010010 n00110100101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011010011 n001101001 n0011010011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110100110 n0011010011 n00110100110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110100111 n0011010011 n00110100111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110101 n0011010 n00110101 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001101010 n00110101 n001101010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011010100 n001101010 n0011010100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110101000 n0011010100 n00110101000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110101001 n0011010100 n00110101001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011010101 n001101010 n0011010101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110101010 n0011010101 n00110101010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110101011 n0011010101 n00110101011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001101011 n00110101 n001101011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011010110 n001101011 n0011010110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110101100 n0011010110 n00110101100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110101101 n0011010110 n00110101101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011010111 n001101011 n0011010111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110101110 n0011010111 n00110101110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110101111 n0011010111 n00110101111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011011 n001101 n0011011 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00110110 n0011011 n00110110 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001101100 n00110110 n001101100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011011000 n001101100 n0011011000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110110000 n0011011000 n00110110000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110110001 n0011011000 n00110110001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011011001 n001101100 n0011011001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110110010 n0011011001 n00110110010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110110011 n0011011001 n00110110011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001101101 n00110110 n001101101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011011010 n001101101 n0011011010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110110100 n0011011010 n00110110100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110110101 n0011011010 n00110110101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011011011 n001101101 n0011011011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110110110 n0011011011 n00110110110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110110111 n0011011011 n00110110111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110111 n0011011 n00110111 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001101110 n00110111 n001101110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011011100 n001101110 n0011011100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110111000 n0011011100 n00110111000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110111001 n0011011100 n00110111001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011011101 n001101110 n0011011101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110111010 n0011011101 n00110111010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110111011 n0011011101 n00110111011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001101111 n00110111 n001101111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011011110 n001101111 n0011011110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110111100 n0011011110 n00110111100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110111101 n0011011110 n00110111101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011011111 n001101111 n0011011111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00110111110 n0011011111 n00110111110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00110111111 n0011011111 n00110111111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111 n0011 n00111 segParams L={1.60000e-05} A={2.00000e-06}
yneuron neuron001110 n00111 n001110 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0011100 n001110 n0011100 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00111000 n0011100 n00111000 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001110000 n00111000 n001110000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011100000 n001110000 n0011100000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111000000 n0011100000 n00111000000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111000001 n0011100000 n00111000001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011100001 n001110000 n0011100001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111000010 n0011100001 n00111000010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111000011 n0011100001 n00111000011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001110001 n00111000 n001110001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011100010 n001110001 n0011100010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111000100 n0011100010 n00111000100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111000101 n0011100010 n00111000101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011100011 n001110001 n0011100011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111000110 n0011100011 n00111000110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111000111 n0011100011 n00111000111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111001 n0011100 n00111001 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001110010 n00111001 n001110010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011100100 n001110010 n0011100100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111001000 n0011100100 n00111001000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111001001 n0011100100 n00111001001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011100101 n001110010 n0011100101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111001010 n0011100101 n00111001010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111001011 n0011100101 n00111001011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001110011 n00111001 n001110011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011100110 n001110011 n0011100110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111001100 n0011100110 n00111001100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111001101 n0011100110 n00111001101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011100111 n001110011 n0011100111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111001110 n0011100111 n00111001110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111001111 n0011100111 n00111001111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011101 n001110 n0011101 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00111010 n0011101 n00111010 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001110100 n00111010 n001110100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011101000 n001110100 n0011101000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111010000 n0011101000 n00111010000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111010001 n0011101000 n00111010001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011101001 n001110100 n0011101001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111010010 n0011101001 n00111010010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111010011 n0011101001 n00111010011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001110101 n00111010 n001110101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011101010 n001110101 n0011101010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111010100 n0011101010 n00111010100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111010101 n0011101010 n00111010101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011101011 n001110101 n0011101011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111010110 n0011101011 n00111010110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111010111 n0011101011 n00111010111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111011 n0011101 n00111011 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001110110 n00111011 n001110110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011101100 n001110110 n0011101100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111011000 n0011101100 n00111011000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111011001 n0011101100 n00111011001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011101101 n001110110 n0011101101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111011010 n0011101101 n00111011010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111011011 n0011101101 n00111011011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001110111 n00111011 n001110111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011101110 n001110111 n0011101110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111011100 n0011101110 n00111011100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111011101 n0011101110 n00111011101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011101111 n001110111 n0011101111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111011110 n0011101111 n00111011110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111011111 n0011101111 n00111011111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001111 n00111 n001111 segParams L={1.27000e-05} A={1.26000e-06}
yneuron neuron0011110 n001111 n0011110 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00111100 n0011110 n00111100 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001111000 n00111100 n001111000 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011110000 n001111000 n0011110000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111100000 n0011110000 n00111100000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111100001 n0011110000 n00111100001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011110001 n001111000 n0011110001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111100010 n0011110001 n00111100010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111100011 n0011110001 n00111100011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001111001 n00111100 n001111001 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011110010 n001111001 n0011110010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111100100 n0011110010 n00111100100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111100101 n0011110010 n00111100101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011110011 n001111001 n0011110011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111100110 n0011110011 n00111100110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111100111 n0011110011 n00111100111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111101 n0011110 n00111101 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001111010 n00111101 n001111010 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011110100 n001111010 n0011110100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111101000 n0011110100 n00111101000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111101001 n0011110100 n00111101001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011110101 n001111010 n0011110101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111101010 n0011110101 n00111101010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111101011 n0011110101 n00111101011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001111011 n00111101 n001111011 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011110110 n001111011 n0011110110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111101100 n0011110110 n00111101100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111101101 n0011110110 n00111101101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011110111 n001111011 n0011110111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111101110 n0011110111 n00111101110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111101111 n0011110111 n00111101111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011111 n001111 n0011111 segParams L={1.00800e-05} A={7.93500e-07}
yneuron neuron00111110 n0011111 n00111110 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001111100 n00111110 n001111100 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011111000 n001111100 n0011111000 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111110000 n0011111000 n00111110000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111110001 n0011111000 n00111110001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011111001 n001111100 n0011111001 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111110010 n0011111001 n00111110010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111110011 n0011111001 n00111110011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001111101 n00111110 n001111101 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011111010 n001111101 n0011111010 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111110100 n0011111010 n00111110100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111110101 n0011111010 n00111110101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011111011 n001111101 n0011111011 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111110110 n0011111011 n00111110110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111110111 n0011111011 n00111110111 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111111 n0011111 n00111111 segParams L={8.00000e-06} A={5.00000e-07}
yneuron neuron001111110 n00111111 n001111110 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011111100 n001111110 n0011111100 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111111000 n0011111100 n00111111000 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111111001 n0011111100 n00111111001 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011111101 n001111110 n0011111101 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111111010 n0011111101 n00111111010 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111111011 n0011111101 n00111111011 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron001111111 n00111111 n001111111 segParams L={6.35000e-06} A={3.15000e-07}
yneuron neuron0011111110 n001111111 n0011111110 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111111100 n0011111110 n00111111100 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111111101 n0011111110 n00111111101 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron0011111111 n001111111 n0011111111 segParams L={5.04000e-06} A={1.98500e-07}
yneuron neuron00111111110 n0011111111 n00111111110 segParams L={4.00000e-06} A={1.25000e-07}
yneuron neuron00111111111 n0011111111 n00111111111 segParams L={4.00000e-06} A={1.25000e-07}

.options output initial_interval=5.0e-5
.print tran  
+ v(n0) 
+ v(n00000000000) 

.end
