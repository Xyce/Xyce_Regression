Demonstration circuit for bug 889.
* This is a chain of 1 1-input CMOS inverters
* The NMOS and PMOS devices have their gates tied 
* together to form a CMOS inverter. VIN1, the input signal, is applied to a 1K
* resistor,RIN, which is connected to the gates of the inverter at node IN.

*
* erkeite:  12/10/2005
*
* This circuit is adapted from the lead_b3soi.cir test case.  
* However, as bug 889 is unrelated (somewhat) to lead currents, I've taken
* out all the lead current stuff.  Also, the original circuit had a bunch
* of resistors in the place of my vmon sources.  When I added these sources,
* (replacing the resistors), the circuit appeared to run all the way to the
* end, but in reality, the nonlinear solver very obviously failed on every
* solve, including the DCOP.
*
* In general, I can understand why the nonlinear solver would fail in 
* transient, but yet the time integrator would accept steps - there 
* are "soft failure" modes in place to handle that case in 
* transient.  For DCOP, however, this shouldn't happen.  
*

.tran 20ns 3us
.print tran v(in) v(vout)

.options timeint abstol=1.0e-5
.options nonlin maxstep=30

VDDdev 	VDD	0	4V
RIN	IN	1	1K
VIN1  1	0  0V PULSE (0V 4V 1.5us 5ns 5ns 1.5us 3.01us)
R1    VOUT  0  10K  
C2    VOUT  0  0.1p 
*IC=0V

* Note: the original version of this netlist included the above
* ic=0V statement.  However, the code has changed so that Xyce
* no longer ignores IC=0, as of Xyce 4.0.1.  In order to restore the 
* original behavior of the bug, this statement needed to be commented
* out.

vmon_nd   vout nd  0.0V
vmon_pd   vout pd  0.0V
vmon_ng   in   ng  0.0V
vmon_pg   in   pg  0.0V
vmon_ns   0    ns  0.0V
vmon_ps   vdd  ps  0.0V
vmon_ne   0    ne  0.0V
vmon_pe   0    pe  0.0V
vmon_nb   0    nb  0.0V
vmon_pb   0    pb  0.0V

MN1 nd ng ns ne nb  CMOSN L=0.258u W=19.585u
MP1 pd pg ps pe pb  CMOSP L=0.258u W=19.585u

.MODEL CMOSN NMOS (    LEVEL   = 10
+ soimod = 0
+ rgatemod = 1
+ mobmod = 2  capmod = 2
+ shmod = 1  igmod = 0  paramchk = 0 )
*
.MODEL CMOSP PMOS (   LEVEL   = 10
+ soimod = 0
+ rgatemod = 1
+ mobmod = 2  capmod = 2
+ shmod = 1  igmod = 0  paramchk = 0 )

.END
