Regression test for simple normal distribution sampling, .param version

.param testNorm={agauss(0.5K,0.05K,1)}
.param R1value={testNorm*2.0}

R2 1 0 7K
R1 1 2 {R1value}
v1 2 0 1000V

.dc v1 1000 1000 1

.sampling useExpr=true

.options samples numsamples=25000
+ outputs={R1:R},{V(1)}
+ sample_type=mc
+ stdoutput=true

.end

