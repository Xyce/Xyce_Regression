***************************************************************
* Calculate both the direct and adjoint sensitivities for
* the case of two objective functions and two parameters.
* This file has both a .PRINT AC and a .PRINT SENS line.
*
* The key points are:
*
*   1) the -o command line option should produce output from
* the .PRINT AC output.
*
*   2) there should be no output from the .PRINT SENS line.
*
*   3) the FILE= qualifier on the .PRINT AC line should have
*      no effect.
*
*   4) the other -o "features" for .PRINT AC are tested by ac.cir.
*
* See SON Bugs 911 and 1170 for more details.
***************************************************************

* Trivial high-pass filter

R2 c 0 1
R1 b c 1
C1 a b 1u
V1 a 0 DC 0V AC 1

.SENS OBJVARS=b,C PARAM=R1:R,c1:c
.options sensitivity direct=1 adjoint=1 stdoutput=1
.print AC file=acSensFoo vr(b) vi(b) vp(b) vm(b) R1:R C1:C
.PRINT SENS vr(b) vi(b) vp(b) vm(b) R1:R R2:R C1:C
.ac dec 5 100Hz 1e6

.end
