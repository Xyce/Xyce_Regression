*******************************************************
* Test of HB output with FILE= qualifiers.   
* See SON Bugs 652 and 701 for more details.
*
* Because we use VP and IP here, it is pretty essential that there be nontrivial
* power in frequencies other than the fundamental -- using a sinusoidal
* input source and only linear devices would have what is essentially
* roundoff error in all frequencies other than the fundamental.   This
* leads to platform-dependent failure when comparing the VP signal.
*
* Wwe're driving this circuit with a roughly square wave and making the 
* circuit slightly non-linear.  That produces nontrivial power in frequencies 
* other than the fundamental frequency.
* 

R1 1 0 1k
C1 1 0 1p
D1 2 1 D1N3940
.MODEL D1N3940 D (IS=4e-10 RS=.105 N=1.48 TT=8e-7 CJO=1.95E-11 VJ=.4 M=.38 EG=1.36 XTI=-8 KF=0 AF=1 FC=.9 BV=600 IBV=1e-4)
*            low high td tr  tf  pulsewidth    period
v1 2 0 pulse 1V 2V  0 1e-5 1e-5 {1/1e4/2-1e-5 } {1/1e4}

* Check the file names generated as "fallbacks" from 
* the .PRINT HB line.
.print HB FILE=hb_foo_csv FORMAT=CSV vr(1) vi(1)
.hb 1e4

.options hbint saveicdata=1 STARTUPPERIODS=2

.end

