* AC simulation for xyce
.options device temp=27
.subckt mysub c_x b_x e_x s_x
e_c c_v 0 c_x 0 1
v_c c_v c 0
f_c c_x 0 v_c   -0.01
e_b b_v 0 b_x 0 1
v_b b_v b 0
f_b b_x 0 v_b   -0.01
e_e e_v 0 e_x 0 1
v_e e_v e 0
f_e e_x 0 v_e   -0.01
e_s s_v 0 s_x 0 1
v_s s_v s 0
f_s s_x 0 v_s   -0.01
q1 c b e s mymodel
+ sw_et=0
+ m=100
.model mymodel npn level=12
+ IS=1e-16
+ IBEI=1e-18
+ IBEN=5e-15
+ IBCI=2e-17
+ IBCN=5e-15
+ ISP=1e-15
+ RCX=10
+ RCI=60
+ RBX=10
+ RBI=40
+ RE=2
+ RS=20
+ RBP=40
+ VEF=10
+ VER=4
+ IKF=2e-3
+ ITF=8e-2
+ XTF=20
+ IKR=2e-4
+ IKP=2e-4
+ CJE=1e-13
+ CJC=2e-14
+ CJEP=1e-13
+ CJCP=4e-13
+ VO=2
+ GAMM=2e-11
+ HRCF=2
+ QCO=1e-12
+ AVC1=2
+ AVC2=15
+ TF=10e-12
+ TR=100e-12
+ TD=2.0e-11
+ RTH=300
+ GMIN=0.0
.ends
v_c_b c_b 0 3
v_b_b b_b 0 0.7 ac 1
v_e_b e_b 0 0
v_s_b s_b 0 0
x_b c_b b_b e_b s_b mysub
.ac dec 10 1e6 1e10
.print ac
+ i(v_c_b)
+ i(v_b_b)
+ i(v_e_b)
+ i(v_s_b)
.end
