IRHC110 Test Circuit
*VD 1 0 DC 10
VD 1 0 DC 0
VS 4 0 0
VG 3 0 DC 0
VID 1 2 DC 0
M1 2 3 4 0 IRHC110 W=0.25 L=3u
.MODEL IRHC110 NMOS LEVEL=18
+ CV=1
+ CVE=1
+ VTO=4.0
+ RD= 0.12
+ RS= 0.055
+ LAMBDA=0.0
+ KAPPA=1e-3
+ NFS=3e11
+ M=3
+ SIGMA0=0
+ UO=700
+ TOX=100nm
+ NSUB=4.6e16
+ PHI=0.6
+ CBSO=2.65e-11
*
*.DC VG 0 8 0.5
.DC VD 0 10 1 VG 4 8 1
.PRINT DC V(1) V(3) V(2) I(VID)
.END

