module main;
initial $ADCStateTest;
endmodule
