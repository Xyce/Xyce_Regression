*********************************************************************
* This tests the error messages, from remeasure, that should occur
* if a TRAN or TRAN_CONT mode measure is included in a netlist that
* is doing a .DC analysis.
*
* See SON Bugs 889 and 1274 for more details.
*
*
*********************************************************************

vsrc1   1a 0 1
rload1a 1a 1b 0.1
rload1b 1b 0 1

.DC vsrc1 1 5 1
.print dc vsrc1:DCV0 v(1a) v(1b)

* Test what happens when a TRAN or TRAN_CONT measure is requested in a .DC netlist
* during remeasure
.MEASURE TRAN tranmax max v(1a)
.MEASURE TRAN_CONT tran_cont_when when v(1a)=2.5

.END


