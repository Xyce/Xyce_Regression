*Sample netlist for BSIM6
*Inverter Transient

.options timeint method=gear debuglevel=-100
.options device temp=25 debuglevel=-100

*.hdl "bsim6.va"
.include "modelcard_xyce.nmos"
.include "modelcard_xyce.pmos"

* --- Voltage Sources ---
vdd   supply  0 dc 1.0
VIN1 vi 0 PWL(0S 0V  7.0e-8 0V 0.1us 1.0V )

* --- Inverter Subcircuit ---
.subckt inverter vin vout vdd gnd
Mp1 vout vin vdd gnd pmos W=10u L=10u 
Mn1 vout vin gnd gnd nmos W=10u L=10u 
.ends

* --- Inverter ---
Xinv1  vi 1 supply 0 inverter
Xinv2  1 2 supply 0 inverter
Xinv3  2 3 supply 0 inverter
Xinv4  3 4 supply 0 inverter
Xinv5  4 vo supply 0 inverter

* --- Transient Analysis ---
.tran 2ns 1us

.print tran v(vi) v(1) v(2) v(3) v(4) v(vo) {ddt(v(vo))} 

.SENS objfunc={V(VO)}
+ param=
+ nmos:TOXE,
+ pmos:TOXE

.options SENSITIVITY adjoint=0 direct=1  forceDeviceFD=true

.print sens 

.end

