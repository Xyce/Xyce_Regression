Does .param work with functions?

.func foobar(x) {x*x}

.param foobie=3.1415926535
+ bletch={foobie*foobar(666)}

V1 1 0 1
R1 1 0 1
B1 2 0 V={foobie*foobar(V(1))}
R2 2 0 1
.DC V1 0 1 .1
.print DC V(1) V(2)
.end
