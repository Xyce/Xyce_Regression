* Xyce netlist for test of PSpice E-Source and 
* G-Source Table syntaxes

R2      2 0 1 
R3      3 0 1 
R4      4 0 1 
R5      5 0 1
R6      6 0 1
R7      7 0 1
R8      8 0 1
R9      9 0 1
R10    10 0 1 
R11    11 0 1
R12    12 0 1 
R13    13 0 1
R14    14 0 1 
R15    15 0 1
R16    16 0 1
R17    17 0 1
V1      1 0  SIN(0V 1V 1e6)

* All sources use the correct Xyce syntax
E2         2 0 TABLE {V(1, 0)} = (-2,-3) (2,3)
E3         3 0 TABLE {V(1, 0)} = (-2,-4) (2,4)
E4         4 0 TABLE {V(1, 0)} = (-2,-5) (2,5)
E5         5 0 TABLE {V(1, 0)} = (-2,-6) (2,6)
E6         6 0 TABLE {V(1, 0)} = (-2,-7) (2,7)
E7         7 0 TABLE {V(1, 0)} = (-2,-8) (2,8)
E8         8 0 TABLE {V(1, 0)} = (-2,-9) (2,9)
E9         9 0 TABLE {V(1, 0)} = (-2,-10) (2,10)

* repeat the subtests, but with G-sources
G10       10 0 TABLE {V(1, 0)} = (-2,-3) (2,3)
G11       11 0 TABLE {V(1, 0)} = (-2,-4) (2,4)
G12       12 0 TABLE {V(1, 0)} = (-2,-5) (2,5)
G13       13 0 TABLE {V(1, 0)} = (-2,-6) (2,6)
G14       14 0 TABLE {V(1, 0)} = (-2,-7) (2,7)
G15       15 0 TABLE {V(1, 0)} = (-2,-8) (2,8)
G16       16 0 TABLE {V(1, 0)} = (-2,-9) (2,9)
G17       17 0 TABLE {V(1, 0)} = (-2,-10) (2,10)

.TRAN 0 1U
.PRINT TRAN FORMAT=PROBE V(1) V(2) V(3) V(4) V(5)
+ V(6) V(7) V(8) V(9) V(10) V(11)
+ V(12) V(13) V(14) V(15) V(16) V(17)

.END
