*******************************************************************
* Xyce Gold Netlist
* Test voltage-controlled switch (S-device) and current-controlled
* switch (W-device).  Also test that XDM can handle cases where
* the device and model name are the same (e.g., VSW and VSW).
*
*******************************************************************

*Analysis directives
.TRAN 0.02U 4U
.PRINT TRAN FORMAT=PROBE W(V1) W(SVSW) W(WISW)

v1  1  0        PWL(0 0 1U 0 1.01U 5 2U 5 2.01U 0 3U 0 3.01U 5)
SVSW  2  1  3  0  VSW
R2  2  0 1
WISW  0  2  v3  ISW
v3  0  3        PWL (0 0 2U 0 2.01U 5)
r3  0  3        200
.MODEL VSW VSWITCH(RON=1 ROFF=1MEG VON=1 VOFF=0)
.MODEL ISW ISWITCH (ION=10mA IOFF=0mA RON=1 ROFF=1E6)

.TRAN 0.02U 4U

.END
