TEST OF A 1-BIT ADDER WITH SWITCHES
*
* Will add comments to this netlist at a later time. Regina Schells 6/1
*
.include bug_307_i.lib1
* MAIN CIRCUIT 
* 
X1 1 2 3 9 13 99 ONEBIT
RINA 1 0 1K
RINB 2 0 1K
RCIN 3 0 1K
RBIT0 9 0 1K
RCOUT 13 0 1K
VCC 99 0 5
VINA 1 0 PULSE(0 3 0 10N 10N 10N 50N)
VINB 2 0 PULSE(0 3 0 10N 10N 20N 100N)
VCIN 3 0 PULSE(0 3 100N 10N 10N 100N 200N)
.TRAN 0.5N 200N
.PRINT TRAN V(1) V(2) V(3) V(9) V(13)
.OPTIONS TIMEINT ABSTOL=1.0E-3 RELTOL=1.0E-3
.END   
