Capacitor Circuit Netlist - lower level.
********************************************************************************
c1 1 B 1uF IC=1
R1 A 1 1K

vconnect0000   A 0 1
vconnect0001   B 0 2

.options nonlin nox=1 
.options device debuglevel=-100
.options timeint reltol=1e-6 abstol=1e-6

.print tran v(1)
.tran 0 1ms

.END

