* Transient sensitivity example, pulse source, analytical version
**********************************************************************
.param cap=10u
.param res=1K

ipulse 0 1 pulse(1a 5a 1s 0.1s 0.4s 0.5s 2s)
r1 1 2 res
c1 2 0 cap
r2 2 3 res
c2 3 0 cap
r3 3 4 res
c3 4 0 cap
r4 4 0 res

.tran .1s 4s
.print tran v(1) v(2) v(3) v(4)

* Sensitivity commands
.print sens 
.SENS objfunc={V(4)} param=ipulse:v1,ipulse:v2,ipulse:td,ipulse:tr,ipulse:tf,ipulse:pw,ipulse:per
.options SENSITIVITY direct=1 adjoint=0  forceanalytic=true
.end
