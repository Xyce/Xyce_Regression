Test circuit for HB output through expressions

v1 a 0   sin  1  1 {SIG_FREQ} 
*v1 a 0 PULSE( 1V 5V 0  5n 5n {.5e-4-10n} 1e-4) AC 1
R1 a b 1k

d1 b 0 dmod

.model  dmod d

.options hbint numfreq=50   loadtimesources=0


.param SIG_PER=1e-5
.param SIG_FREQ={1/SIG_PER}

*v1 a 0 pulse(0 5 0 5n 5n {SIG_PER/2-10n} {SIG_PER})
*R1 a b 1
*R2 b 0 2
*C1 a b 1u

.hb 100kHz

.print hb V(B) {V(B)} VR(B) {VR(B)} VI(B) {VI(B)} VM(B) {VM(B)} VDB(B) {VDB(B)} VP(B) {VP(B)} 

.end
