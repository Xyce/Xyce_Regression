Basic diode circuit testing simple parameter use in model statement inside a
* subcircuit, with an expression on the call line

.param ISmant=100

XD1 1 0 DMODsub IS0={ISmant*1F} RS0=2K
V1 1 0 DC 5V

.subckt DMODsub 1 2 IS0=100mA RS0=2
D1 1 2 DMOD1
.model DMOD1 D (IS={IS0} RS={RS0})
.ends

.dc V1 0 5 1
.print DC v(1) I(v1)
.end
