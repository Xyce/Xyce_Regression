* curly braces for simple function calls
* Xyce netlist for corresponding HSPICE netlist.
* This tests XDM can correctly identify and put 
* curly braces around single functions in parameter 
* statements. This should also include removing 
* any delimiters embedded in the function call.
* See issue #154 in XDM gitlab.

.OPTIONS DEVICE TNOM=25

.PARAM 
+ P1=1.5 VAL3={sqrt(9)} VAL2={agauss(0,0,2*p1)} VAL1={max(1,3)}

Va 1 0 DC 0
R1 1 2 R=val1
R2 2 0 R=val2+val3
.DC LIN va 0 10 1


.PRINT DC FORMAT=PROBE v(1) v(2)
