Simple RC circuit
*
* Eric Keiter, SNL
*
* Tests simultaneous sweeps of frequency, magnitude and phase, using a
* data table to specify frequency, combined with expressions for magnitude 
* and phase.
*

.global_param mag={log10(freq)+1}
.global_param phase={0.1*mag}

Isrc 1 0 AC {mag} {phase} 
R1 1 0 1e3
C1 1 0 2e-6


.data table
+ freq
+  1.0e0
+  1.0e1
+  1.0e2
+  1.0e3
+  1.0e4
+  1.0e5
.enddata


.print ac 
+ {mag}
+ {phase}
+ {Isrc:acmag}
+ {Isrc:acphase}
+ v(1)

.AC data=table

.END
