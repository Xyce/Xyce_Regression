* Test N(), P(), W() with .FFT and .MEASURE FFT.
*
*************************************************

.TRAN 0 1
.OPTIONS FFT FFT_ACCURATE=1 FFTOUT=1

V1 1 0 1
R1 1 0 2

.FFT N(1) NP=8 WINDOW=HAMM FORMAT=UNORM
.FFT P(R1) NP=8 WINDOW=HANN FORMAT=UNORM
.FFT W(R1) NP=8 WINDOW=HANN FORMAT=UNORM

.MEASURE FFT ENOB ENOB N(1)
.MEASURE FFT THDPR1 THD P(R1)
.MEASURE FFT SFDRWR1 SFDR W(R1)

.PRINT TRAN N(1) P(R1) W(R1)

.END
