TEST A5_HS of subcircuit regression tests
* **********************************************************************
* A simple pair of MOSFET level 3 inverters
* The inverters are constructed from dissimilar mosfets, just for testing 
* purposes
*
* Test A5_HS uses a single inverter subcircuits with a model statement that 
* includes parameters from the subcircuit line. It also uses parameters for 
* the widths of the N and P mosfets.  By construction it should be identical
* to case A0
*
* This test case differs from test A4 only in the ordering of the subcircuit
* instances.  This case is meant to test whether the parser is appropriately
* resetting its context after handling the first instance with parameters.
*
*Note: ERK 10/22/09
* This test case differs from test A5 only in that the keyword PARAMS: has
* been removed, for Hspice compatibility, per bug 1733.
*
* Author:   $Author$
* Revision: $Revision$
* Date:     $Date$
*
* **********************************************************************

.subckt INV1 IN OUT VDD GND  WN=100u WP=200u VTON=1.679 VTOP=-1.6
MN1 OUT IN GND GND CD4012_NMOS L=5u W={WN}
MP1 OUT IN VDD VDD CD4012_PMOS L=5u W={WP}
***** original mosfets
.MODEL cd4012_nmos NMOS (
+ LEVEL = 3 UO = 190   VTO = {VTON}   TOX = 6E-08   NSUB = 8.601E+15
+ NSS = 0   RS = 13.21   RD = 11.59   RSH = 0   IS = 1E-14
+ VMAX = 4.206E+04 NFS=1E10  GAMMA=0.37 PHI=0.65 
+ XJ = 7.1E-06   LD = 8.6E-07   DELTA = 0   THETA = 0.0021   ETA = 0.057   KAPPA = 0.15
+ KP = 2.161E-05  L=5u W=175u
+ CBD=0.1P CBS=0.1P PB=0.81 CGSO=2P CGBO=4P CGDO=2P CJ=2E-4 MJ=0.5 CJSW=1E-9
+ MJSW=0.5 JS=1E-8 TPG=0 KF=1E-25 AF=1 FC=0.5 TNOM=27)
.MODEL cd4012_pmos PMOS (
+ LEVEL = 3  UO = 310  VTO = {VTOP}  TOX = 6E-08  NSUB = 5.701E+15
+ NSS = 0    VMAX = 5.374E+04   RS = 5.359   RD = 93.66   RSH = 0   IS = 1E-14
+ XJ = 7.9E-06   LD = 3E-08   DELTA = 0   THETA = 0.0278   ETA = 0.535   KAPPA = 0.643
+ KP = 1.711E-05 L=5u W=270u GAMMA=0.37 PHI=0.65 NFS=1E10
+ CBD=0.1P CBS=0.1P PB=0.81 CGSO=2P CGBO=4P CGDO=2P CJ=2E-4 MJ=0.5 CJSW=1E-9
+ MJSW=0.5 JS=1E-8 TPG=0 KF=1E-25 AF=1 FC=0.5 TNOM=27)
.ends


Xinv2 MID OUT VDD 0 INV1  WN=175u WP=270u VTON=1.0 VTOP=-1.0
Xinv1 IN MID VDD 0 INV1  WN=175u WP=270u 

VDDdev 	VDD	0	5V
RIN	IN	1	1K
VIN1  1	0  5V PULSE (5V 0V 1.5us 5ns 5ns 1.5us 3.01us)
R1    OUT  0  10K  
C2    OUT  0  0.1p

.tran 20ns 30us
.print tran PRECISION=10 WIDTH=19 v(out) v(in) v(1)


.end
