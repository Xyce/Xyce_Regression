Basic voltage divider circuit test of subcircuit usage
* Should produce results identical to Double_Resist_Control.
* Tests use of expressions involving function calls in params of subcircuit 
* *and* context issues 
* regarding those params.

.param R0=10k
.param R1=1k
.func R2(X)  {0.5*X}
XR1 1 2 Rsub PARAMS: R=R0
XR2 2 0 Rsub PARAMS: R={R2(R0)}
V1 1 0 DC 5V

.subckt Rsub 1 2 PARAMS: R=R1
R1 1 2 R
.ends

.dc V1 0 5 1
.print DC v(1) v(2) I(v1)
.end
