test of wodicka splines

b1 1 0 v={wodicka("sinewave.dat")}
r1 1 0 500
.tran 1us 10us

*COMP V(1) OFFSET=6
.print tran v(1)

.end
