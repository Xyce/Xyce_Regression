* Test of duplicate measure names in Xyce.  The first
* M1 and M2 definitions should be ignored and produce
* warning messages.  This test uses a mix of TRAN and
* TRAN_CONT measures, but it should not produce the
* <netlistName>.mt0 file since the TRAN mode M1
* definition is not used.  This also tests that
* PRINT=STDOUT works for a TRAN_CONT measure.
*
* See SON Bugs 1274 and 1300 for more details.
******************************************************
.TRAN 0 1
.PRINT TRAN V(1) V(2)

V1 1 0 PWL 0 0 0.5 1 1 0
R1 1 0 1

V2 2 0 PWL 0 1 0.5 0 1 1
R2 2 0 1

.MEASURE TRAN M1 MIN V(1)
.MEASURE TRAN_CONT M2 WHEN V(2)=0.2

.MEASURE TRAN_CONT M1 WHEN V(1)=0.3
.MEASURE TRAN_CONT M2 WHEN V(2)=0.4

* This should only send output to stdout
.MEASURE TRAN_CONT M3 WHEN V(1)=0.2 PRINT=STDOUT

.END
