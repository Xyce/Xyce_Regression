test multiplier

Vin 1 0 1.0
Rin 1 2 1.0

Xtest1 2 3 testA 
Xtest2 3 0 testA 

.subckt testA A B 
Xtest A B testB M=15
.ends

.subckt testB A B 
R1 A B 0.5 M=4
.ends

.DC Vin 1 1 1
.PRINT DC V(1) V(2) V(3) I(Vin)  { Xtest1:Xtest:R1:R } { Xtest2:Xtest:R1:R }

