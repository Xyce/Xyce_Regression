* This netlist is used to test the use of Xyce command line
* options, such as -o commandLine.prnOutput, in the
* Python initialize() method

V1 1 0 SIN(0 1 1)
R1 1 0 1

.TRAN 0 1
.PRINT TRAN V(1)

.MEASURE TRAN MAXV1 MAX V(1)

.END

