Test of synapse device

vin a1 0 1.0

.model synParams synapse alpha=1.1e6 beta=190 Tmax=1e-3 Vp=2e-3 Kp=5e-3 gmax=1e-10 Erev=0.0

ysynapse syn a1 a2  synParams

rload a2 0 100

.tran 0 1
.print tran v(a1) v(a2)
.end
