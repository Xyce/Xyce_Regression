Test error message capability when a mutual inductor references an undefined
*inductor

R1 1 2 1
L1 2 0 1
*L2 2 3 1
L3 2 0 1
V1 1 0 DC 1

K1 L1 L3 0.1
K2 L1 L3 0
K3 L1 L2 0

.DC V1 1 1 0.1
.end
