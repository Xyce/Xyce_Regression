* This netlist is used to test the getTimeStatePairsADC() 
* method for valid YADC names.  It also tests that the width 
* value on the instance line takes precedence over the width 
* value in the model card.

* Note: these WIDTH values will NOT be overwritten by the Python program.
* They will be used as set in device constructors.
YADC adc1 1 0 simpleADC R=1T WIDTH=2
YADC adc2 1 0 simpleADC R=1T
.model simpleADC ADC(settlingtime=50ns uppervoltagelimit=2 lowervoltagelimit=0 width=3)

v1 1 0 PWL 0 0 1e-4 2

* Limit the max. time step so that the simulation takes at
* least 1000 steps.  This is needed for the comparison of
* Python-generated timeArray and voltageArray in the .sh file.
.TRAN 0 1e-4 0 1e-7
.PRINT TRAN V(1) YADC!ADC1:WIDTH YADC!ADC2:WIDTH
.END

