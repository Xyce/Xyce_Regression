Regression test to show temperature-dependent capacitor behavior, using DTEMP

.param dtempParam=600

c1    1 0 CAP1 1uF IC=1 DTEMP={dtempParam}
r1    1 2 1K
v1 2 0 0V
.model CAP1 C ( TC1=1.77M TC2=-0.63U )

.options temp=27.0

.step dtempParam list 600 700 800

.print tran v(1)
.tran 0 5ms
.options timeint reltol=1e-6 abstol=1e-6
.END
