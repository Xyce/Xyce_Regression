A simple test case of a resistor with small resistance.  
* in this test node 'a' should be automatically removed and R1 removed.
* the result is a circuit with no devices.  check that.

* supernoding is off by default.  activate it
.options topology supernode=true
.options device zeroresistancetol=1e-10

* test case when resistance is lower than a given tolerance
R1 a 0 1e-12 

.TRAN 1us 5us
.print TRAN v(a)

.END
