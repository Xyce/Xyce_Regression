* Transient sensitivity example, PWL source, analytical version
.param cap=1u
.param res=1K

c1 1 0 cap
c2 2 0 cap
R1 1 3 res
R2 1 2 res

Vin 3 0 PWL(0 0 1ms 1 2ms -1 3ms -0.5 4ms 0.25 5ms 0.75 6ms 0.0  )

* Transient commands
.tran 0 10ms uic
.options timeint reltol=1e-6 abstol=1e-6


*comp V(2) offset=0.2
*comp V(2)_V0 offset=0.1
*comp V(2)_V1 offset=0.1
*comp V(2)_V2 offset=0.1
*comp V(2)_V3 offset=0.1
*comp V(2)_V4 offset=0.1
*comp V(2)_V5 offset=0.1
*comp V(2)_V6 offset=0.1

.print tran v(2)
+ V(2)_V0 
+ V(2)_V1 
+ V(2)_V2 
+ V(2)_V3 
+ V(2)_V4 
+ V(2)_V5 
+ V(2)_V6


.end

