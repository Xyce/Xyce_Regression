test of fast table, which has no breakpoints.

b1 1 0 v={fasttablefile("sinewave.dat")}
r1 1 0 500
.tran 1us 10us

*COMP V(1) OFFSET=6
.print tran v(1)

.end
