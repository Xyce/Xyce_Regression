* Operational Amplifier.  AC Analysis.
* BSIM3 testing, 3/16/96. 


.param m6w=2u
.param m6l=1u

*Operational Amplifier
M1 bias1 1 cm cm nmos w=10u l=1u
M2 bias2 in2 cm cm  nmos w=10u l=1u
M3 vdd bias1 bias1 vdd pmos w=2u l=1u
M4 bias2 bias1 vdd vdd pmos w=2u l=1u

m5 cm bias vss vss nmos w=2u l=1u
mbias bias bias vss vss nmos w=2u l=1u
rbias 0 bias 195k

* the "bogus" node is simply there to test out a bug.
*m6 8 bias vss vss  nmos w={m6w} l={m6l}
vbogus bogus vss 0.0
m6 8 bias vss bogus nmos w={m6w} l={m6l}
m7 8 bias2 vdd out nmos w=2u l=1u

Cfb bias2 8 2p

Vid 1 c 0 ac 0.1
eid in2 c 1 c -1
vic c 0 dc 0
vss1 vss 0 -5
Vdd1 vdd 0 5 

*AC analysis
.ac dec 10 1e2 100Meg 
.print ac v(8)

.sens objvars=8 param=m6:w,m6:l
.options sensitivity direct=0 adjoint=1  stdoutput=1  
*forcedevicefd=1
.print sens 
*+ format=tecplot

.model nmos nmos level=9 version=3.2.2
.model pmos pmos level=9 version=3.2.2

.end




