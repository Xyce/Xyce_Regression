Test of BSIM-CMG output variable feature
* This duplicates the gummel_n.cir test case, but adds gm computation
* and output of other output variables
*Sample netlist for BSIM-CMG
*Drain current symmetry for nmos

*.options nonlin abstol=1e-6 reltol=1e-6
.options device temp=25

.include "modelcard.nmos_xyce"

* --- Voltage Sources ---
vdrain drain 0 dc 0
esource source 0 drain 0 -1
vgate gate  0 dc 1.0
vbulk bulk 0 dc 0.0


* --- Transistor ---
M1 drain gate source bulk nmos1 TFIN=15n L=30n NFIN=10 NRS=1 NRD=1

* Second transistor for finite differencing
Bdrain drain2 0 V={V(drain)}
Bgate gate2 0  V={V(gate)+((V(gate)==0)?.00000001:(1e-8*abs(v(gate))))}
Bsource source2 0 V={V(source)}
Bbulk bulk2 0 V={V(bulk)}

M2 drain2 gate2 source2 bulk2 nmos1 TFIN=15n L=30n NFIN=10 NRS=1 NRD=1

* --- DC Analysis ---
.dc vdrain -0.1 0.1 0.001 vgate 0.0 1.0 0.2
*COMP {N(M1:gm)-{(N(M2:ids)-N(M1:ids))/(V(gate2)-V(gate))}} abstol=1e-9
*COMP {(N(M2:ids)-N(M1:ids))/(V(gate2)-V(gate))} abstol=1e-9
.print dc v(drain) v(gate) N(M1:ids) {(N(M2:ids)-N(M1:ids))/(V(gate2)-V(gate))} N(M1:gm) {N(M1:gm)-{(N(M2:ids)-N(M1:ids))/(V(gate2)-V(gate))}}  N(M1:Vth) N(M1:Vds) N(M1:Vbs) N(M1:Vgs) N(M1:Vdsat)

.end
