test multiplier

V1 1 0 PULSE (0v 5V 1us 10ns 10ns 1us 2us)
Xtest2 1 2 test  M=5
Rin 2 0 10k

.subckt test 1 2 
D1 1 2 DFOR 

.MODEL DFOR D
+ IS = 2.355E-14 N = 1.112 BV = 1000 IBV = 0.001
+ RS = 0.137 CJO = 2.993E-10 VJ = 0.5033 M = 0.3144
+ FC = 0.5 EG = 1.11 XTI = 3 TT = 1.7E-07
.ends

.tran 10ns 6us
.PRINT tran V(1) V(2) I(V1)  

