* Xyce netlist for testing SFFM V-Sources

ISFF1 15 0 DC 1A SFFM(0V 0.5A 20K 10 5K)
RSSF1 15 0 1
.TRAN 0 .5ms 0
.PRINT TRAN FORMAT=PROBE V(15)

.END
