********************************************************
* Test error messsage when .LIN analysis is requested
* but there are no port (P) devices in the netlist.
*
* See SON Bug 1202 for more details.
********************************************************

* Trivial high-pass filter
R1 b 0 2
C1 a b 1u
V1 a 0 DC 0V AC 1

.print AC vm(b)
.ac dec 5 100Hz 1e6

.LIN SPARCALC=1

.end

