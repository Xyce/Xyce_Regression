* Basic IV curves for EKV 2.6 NMOS

V1 g 0 1

v2 d1 0 1
vdmon d1 d 0

Mfoo d g 0 0 P L=.45u W=.8u AS=1e-12 AD=1e-12 PS=2e-6 PD=2e-6

* model card of absolutely no relation to a real device, just trying to
* use non-default parameters in reasonable ranges
.MODEL P PMOS (
+ LEVEL  = 260
+ TNOM = 27.00
+ COX = 4.379E-3
+ XJ = 22.53n
+ VTO =-570.6e-3
+ TCV =-1.194e-3
+ GAMMA = 670.7e-3
+ PHI = 450.0E-3
+ KP = 232.1e-6
+ BEX =-1.828
+ THETA=0
+ E0 = 42.216MEG
+ UCRIT = 3.146E6
+ UCEX=0.8
+ LAMBDA = 228.3e-3
+ DL =-60.86n
+ DW =-209.7n
+ WETA=2.001
+ LETA=264.6e-3
+ Q0 = 230e-6
+ LK=0.4e-6
+ IBA = 0.000
+ IBB = 300.0E6
+ IBBT = 800.0E-6
+ IBN = 1.000
+ RSH = 0.000
+ HDIF = 0.000
+ AVTO = 0.000
+ AKP = 1e-6
+)

.dc  v2 0 -3  -.01 v1 -3 -5 -.4
.print DC v(d1) v(g) ID(Mfoo)

