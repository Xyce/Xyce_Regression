* NMOS Id-Vd

.include modelcard.nmos

vg 1 0 1.2
vd 2 0 1.2
vb b 0 0.0

m1 2 1 0 b n1 W=10.0u L=0.09u NF=5

.dc vd 0.0 1.18 0.02 vg 0.2 1.2 0.2
.print dc v(2) v(1) i(vd)

.end

