Regression test for simple uniform distribution propagation via regression PCE
* The circuit is a simple voltage divider, so it has an analytic solution
* Also, the propagated mean, max and min can be computed analytically as well.
*
* Here is the results of that analytical analysis:
*
* analytical mean of R1 is 4.0e+3
* analytical max  of R1 is 2.0e+3
* analytical min  of R1 is 6.0e+3
*
* analytical mean of V1 is 600
*
* Analysis details:
*
* solution to voltage divider:  v(1) = V(2) * R2/(R1+R2)
*
* analytical mean of v(1) is: 1000 * 6/(4+6) = 1000 * 6/10 = 600
* analytical max  of v(1) is: 1000 * 6/(2+6) = 1000 * 6/8  = 750
* analytical min  of v(1) is: 1000 * 6/(6+6) = 1000 * 6/12 = 500
* analytical variance  of v(1) is: (max-min)^2/12.0 = (750-500)^2/12.0 = 5208.3333333333
* analytical stddev of v(1) is: sqrt(variance) = (750-500)/sqrt(12) = 72.1687836487
*
.global_param testNorm={aunif(2k,1k)}
.global_param R1value={testNorm*2.0}

R2 1 0 6K
R1 1 2 {R1value}
v1 2 0 1000V

.dc v1 1000 1000 1

.print dc format=tecplot v(1)

.result {v(1)}
*
.SAMPLING 
+ useExpr=true
*+ param=testNorm
*+ type=uniform
*+ lower_bounds=1k 
*+ upper_bounds=3k 

.options SAMPLES numsamples=10
+ regression_pce=true
+ order=5
+ outputs={v(1)}
+ sample_type=lhs
+ stdoutput=true
+ resample=true

.end

