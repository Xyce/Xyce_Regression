*Xyce netlist for testing G-sources syntaxes

.TRAN 0 1000ns
.PRINT TRAN FORMAT=PROBE V(N388954) V(N388906) V(N391734) V(N391678)
+ V(N392868) V(N392673) V(N393371) V(N393403)
+ V($G_CLK) V(2) V(3) V(4)

G_G1         N388906 0 N388954 N388948 2
R_R10        N388948 0 1
R_R11        N388906 0 1
V_V6         N388954 0  SIN(0V 1V 1e6 0 0 0)

* test the POLY form of the G-Source
R_R16        0 N391728 1
V_V9         N391734 0 SIN(0V 2V 1e6 0 0 0)
R_R17        0 N391678 1
G_G2         N391678 0 POLY(1) N391734 N391728 0.0 2

* test the VALUE form of the G-Source
G_G3         N392673 0 VALUE 2*V(N392868,0)
V_V10        N392475 0 1
R_R18        N392673 0 1 
V_V11        N392868 0 SIN(0V 1.5V 1e6 0 0 0)
R_R19        N392868 0 1

* test the TABLE form of the G-Source
R_R20         N393403 0  1 
G_G4          N393403 0 TABLE V(N393371,0) = (-1,-3) (1,3)
V_V12         N393371 0 SIN(0V 0.75V 1e6 0 0 0)

*Test of G-Source syntaxes with Global Node
RG1 $G_CLK 0 1
VG1 $G_CLK 0  SIN(0V 1V 1e6 0 0 0)

RG2  2 0 1
GG2  2 0 VALUE 2*V($G_CLK) 

RG3  3 0 1
GG3  3 0 VALUE 3*V($G_CLK) 

RG4  4 0 1
GG4  4 0 VALUE IF(((V($G_CLK) >= 0.8)&(V($G_CLK) >= 0.8)),3.5, 3.5)

.END