Test of netlist error.  
*
* The ojbfunc parameter is improperly formatted, so the code should emit an error message and gracefully exit.
*
* This is the same circuit as the one used in the twoObj.cir test.
*
.global_param VCCvalue=10V

VCC 4 0 DC {VCCvalue}
RB1 4 1 40k
RB2 1 0 10k
RE 2 0 1K
RC 5 3 6K
VM 4 5 DC 0; monitor collector current
Q1 3 1 2 Q2N2222
.model Q2N2222 NPN(BF=100 IS=3.295e-14 VA=200)

.options nonlin debuglevel=-100
.options device debuglevel=-100

.DC VCCvalue 1 10 0.2

* several of the sensitivities need offsets, as their computed values are
* near zero for the lower biases.
*comp  d_{v(3)*v(3)}/d_q2n2222:bf_adj offset=2.0e-6
*comp  d_{V(3)*V(3)}/d_Q2N2222:vaf_adj offset=1.0e-6
*comp  d_{v(3)*v(3)}/d_re:r_adj offset=-2.0e-9

.print dc v(4)
.print sens v(4)

.SENS param=
+ RB1:R,RB2:R,RE:R,RC:R,VM:DCV0,
+ Q2N2222:bf,
+ Q2N2222:is,
+ Q2N2222:nf,
+ Q2N2222:tnom,
+ Q2N2222:vaf
+objfunc={I(VM),V(3)*V(3)}

.op 

.options SENSITIVITY direct=0 adjoint=1  difference=forward  diagnosticfile=0 STDOUTPUT=1 debuglevel=-100 REUSEFACTORS=0

