
*Simulation of Checksum U74 OP AMP

.tran 1us 1ms 0 1ns

.print tran v(4)

*.options loca MAXNLITERS=200 MINSTEPSIZE=1e-12
.options nonlin searchmethod=1

*Voltage Source to OP Amplifier
V1 1 0 3.3

*OP Amplifier Passive Comp.
R1 3 3a 10k
R2 1 2 1.1M
R3 2 0 100
R4 3 4 1.1M
R5 4 5 10k
R6 5 0 1G
R7 3a 0 1k

C1 3 4 1n

D1 3a 0 1N4004
D2 0 3a 1N4004

*OP Amplifier
CB 1 0 0.1u
X1 2 3 1 0 4 LMV831

*CAP DUT
CDUT 3a 6 1.47u IC=0
RDUT 3a 6 7M
VCHR 0 6 50

* PINOUT ORDER +IN -IN +V -V OUT
* PINOUT ORDER 1 3 5 2 4
.SUBCKT LMV831 1 3 5 2 4
V120 28 58 362E-6
Q21 6 7 8 QLN
R633 9 10 2
R634 11 10 2
R635 7 12 1E3
R636 13 14 1E3
R637 15 5 5
R638 2 16 5
R640 17 18 400
R641 19 20 5
R642 8 21 5
D46 22 5 DD
D47 2 22 DD
D48 23 0 DIN
D49 24 0 DIN
I48 0 23 0.1E-3
I49 0 24 0.1E-3
E100 8 0 2 0 1
E101 20 0 5 0 1
D50 25 0 DVN
D51 26 0 DVN
I50 0 25 0.1E-3
I51 0 26 0.1E-3
E102 27 3 25 26 0.06
G37 28 3 23 24 2.4E-6
R643 2 5 1E6
E103 29 0 20 0 1
E104 30 0 8 0 1
E105 31 0 32 0 1
R644 29 33 1E5
R645 30 34 1E5
R646 31 35 1E5
R647 0 33 10
R648 0 34 10
R649 0 35 1E3
E106 36 1 35 0 -0.11
R650 37 38 1E3
R651 38 39 1E3
C106 29 33 0.2E-12
C107 30 34 1E-12
C108 31 35 7E-12
E107 40 36 34 0 -0.12
E108 41 40 33 0 0.28
E109 42 8 20 8 0.51
D52 17 20 DD
D53 8 17 DD
M56 43 44 16 16 NOUT L=3U W=1000U
M57 45 46 15 15 POUT L=3U W=1000U
M58 47 47 19 19 POUT L=3U W=1000U
M59 48 49 9 9 PIN L=3U W=460U
M60 50 51 11 11 PIN L=3U W=460U
M61 52 52 21 21 NOUT L=3U W=1000U
R652 53 46 100
R653 54 44 100
G38 17 42 55 42 0.2E-3
R654 42 17 1.8E8
C109 18 56 26E-12
R655 8 48 2E3
R656 8 50 2E3
C110 48 50 5E-12
C111 28 0 13E-12
C112 27 0 13E-12
C113 22 0 0.5E-12
D54 44 6 DD
D55 57 46 DD
Q22 57 14 20 QLP
M62 59 60 20 20 PIN L=6U W=500U
E110 39 0 28 0 1
E111 37 0 3 0 1
M63 60 60 20 20 PIN L=6U W=500U
V121 59 10 0.41
R657 22 45 15
R658 43 22 15
J5 61 28 61 JNC
J6 61 27 61 JNC
J7 27 62 27 JNC
J8 28 62 28 JNC
C114 28 63 0.1E-12
E112 64 42 50 48 1
R659 64 55 1E3
C115 55 42 11E-12
G39 65 42 17 42 -1E-3
G40 42 66 17 42 1E-3
G41 42 67 52 8 1E-3
G42 68 42 20 47 1E-3
D56 68 65 DD
D57 66 67 DD
R660 65 68 1E8
R661 67 66 1E8
R662 68 20 1E3
R663 8 67 1E3
E113 20 53 20 68 1
E114 54 8 67 8 1
R664 66 42 1E6
R665 67 42 1E6
R666 42 68 1E6
R667 42 65 1E6
G43 5 2 69 0 -2.5E-4
R668 40 41 1E9
R669 36 40 1E9
R670 1 36 1E9
R671 3 27 1E9
R672 42 55 1E9
R673 53 20 1E9
R674 8 54 1E9
R675 38 0 1E9
G44 60 8 70 0 140E-6
G45 47 52 70 0 5E-6
V125 70 0 1
I53 5 2 2.27E-4
L2 22 4 0.4E-9
R684 22 4 400
V127 20 61 0
V128 62 8 0.1
R685 47 20 1E8
R686 8 52 1E8
R687 16 44 1E8
R688 15 46 1E8
R689 0 69 1E9
R690 63 27 100
R691 51 27 1850
R692 49 58 1850
E121 20 13 5 15 2.2
E122 12 8 16 2 2.2
R715 60 20 1E12
E124 56 0 22 0 1
R717 17 56 3E8
C126 17 71 19E-12
R724 8 71 1E4
D58 72 73 DL
V144 73 0 3
R725 0 72 1E8
G53 27 0 72 0 15E-11
I66 27 0 0.2E-12
G54 28 0 72 0 15E-11
I67 28 0 0.2E-12
I68 0 74 1E-3
D59 74 0 DD
V146 74 69 0.6551
R726 0 69 1E6
E125 28 41 69 0 282E-6
R727 41 28 1E9
R729 0 70 1E12
E128 75 0 38 0 1
R730 75 32 1E5
R731 0 32 1E3
C127 75 32 7E-12
.MODEL DL D IS=0.95E-11 N=1.47 XTI=1.5
.MODEL DVN D KF=7E-13 IS=1E-16
.MODEL DD D
.MODEL DIN D
.MODEL QLN NPN
.MODEL QLP PNP
.MODEL JNC NJF
.MODEL POUT PMOS KP=200U VTO=-0.7
.MODEL NOUT NMOS KP=200U VTO=0.7
.MODEL PIN PMOS KP=200U VTO=-0.7
.ENDS
* END MODEL LMV831

.MODEL 1N4004 D (IS=5n RS=0 BV=200 IBV=5.00u CJO=4p M=0.333 N=2 EG=0.9)

.END
