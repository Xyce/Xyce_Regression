Test of different cap model types
VIN  1 0 PULSE(0 1 10U 1N 1N 30U)
R    1 2 1K
C1    3 0 CMODEL1 L=20U W=1U
C2    3 0 CMODEL2 L=20U W=1U
C3    3 0 {1*20U*1U*2}
VMON 2 3 0
.MODEL CMODEL1 C (CJ=1 C=2)
.MODEL CMODEL2 CAP (CJ=1 C=2)
.TRAN 1N 20U 
.PRINT TRAN  V(3) {I(VMON)*100.0+1.0} I(C1) I(C2) I(C3)
*.OPTIONS TIMEINT CONSTSTEP=1
.END
