Class AB Amplifier Circuit
********************************************************************************
* Tier No.: 3
* Directory/Circuit Name:SANDLER24/sandler24.cir
* Description:  The amplifer circuit netlist was developed by Steve Sandler to 
*       compare the validity of simulations using 3 different circuit simulation
*       tools.  The results were compared to measured data.
* Input: VIN=V(4)
* Output: V(4), V(6), V(11)
********************************************************************************
* NOTE: 7/30/02 Code enhancement to read E,F,G poly sources.
*       Updated netlist by replacing B sources with E,F,G sources from original
*       circuit. (RLS)
********************************************************************************
*
* MAIN CIRCUIT DEFINITION
*
VEE 1 0 -9
VCC 2 0 9
VIN 4 0 SIN 0 100M 1K
R1 4 5 1K
R2 5 11 22K
R_LOAD 11 0 50
R7 2 12 1K
R8 7 1 1K
R9 11 8 2.2
R10 9 11 2.2
Q5 2 12 9 QN2222A
Q7 1 7 8 QN2907A
D1 12 6 DN4148
D2 6 7 DN4148
X2 0 5 2 1 6 UA741T
*
* ANALYSIS AND OPTION STATEMENTS
*
.options timeint newdae=1
.options mpde IC=1 N2=11 oscsrc=VIN diff=1 wampde=1 oscout=4
.tran 1u 2m 
* These xyce_verify tolerances can be tighter, if the MPDE circuit
* is run with more fast time scale points. 
*COMP {v(11)+3.0} RELTOL=0.04
*COMP {v(6)+3.0} RELTOL=0.04
*COMP {v(4)+3.0} RELTOL=0.04
.print tran {v(4)+3.0}   {v(6)+3.0}  {v(11)+3.0}
*ALIAS  V(4)=IN  V(6)=PA_OUT V(11)=OUT
**********************************************************
* MODEL DEFINITIONS
.MODEL QN2222A NPN (IS=81.1F NF=1 BF=205 VAF=113 IKF=.5
+ ISE=10.6P NE=2 BR=4 NR=1 VAR=24 IKR=.225 RE=.343 RB=1.37
+ RC=.137 XTB=1.5 CJE=29.5P CJC=15.2P TF=397P TR=85N)
*   MOTOROLA 40 VOLT  .8 AMP  400 MHZ  SINPN  TRANSISTOR  04-11-1991
.MODEL QN2907A PNP (IS=381F NF=1 BF=154 VAF=139 IKF=.14
+ ISE=15.3P NE=2 BR=4 NR=1 VAR=20 IKR=.21 RE=.552 RB=2.21
+ RC=.221 XTB=1.5 CJE=15.6P CJC=20.8P TF=636P TR=63.7N)
*   60 VOLT  .6 AMP  250 MHZ  SIPNP  TRANSISTOR  04-11-1991
.MODEL DN4148 D(RS=.8 CJO=4PF IS=7E-09 N=2 VJ=.6V
+ TT=6E-09 M=.45 BV=100V)
***********************************************************
* SUBCIRCUIT DEFINITION
***********************************************************
.SUBCKT UA741T    1 2 3 4 5
*
C1   11 12 4.664E-12
C2    6  7 20.00E-12
DC    5 53 DX
DE   54  5 DX
DLP  90 91 DX
DLN  92 90 DX
DP    4  3 DX
*EGND 99 0 POLY(2) 3 0 4 0 0 0.5 0.5
*FB 7 99 POLY(5) VB VC VE VLP VLN 0 10.61E6 -10E6 10E6 10E6 -10E6
BGND 99 0 V={POLY(2) V(3) V(4) 0 0.5 0.5}
BB 7 99 I={POLY(5) I(VB) I(VC) I(VE) I(VLP) I(VLN) 0 10.61E6 -10E6 10E6 10E6 -10E6}
GA 6  0 11 12 137.7E-6
GCM 0  6 10 99 2.574E-9
IEE  10  4 DC 10.16E-6
*HLIM 90  0 VLIM 1K
BLIM 90 0 V={1E3 * I(VLIM)}
Q1   11  2 13 QX
Q2   12  1 14 QX
R2    6  9 100.0E3
RC1   3 11 7.957E3
RC2   3 12 7.957E3
RE1  13 10 2.740E3
RE2  14 10 2.740E3
REE  10 99 19.69E6
RO1   8  5 150
RO2   7 99 150
RP    3  4 18.11E3
VB    9  0 DC 0
VC 3 53 DC 2.600
VE   54  4 DC 2.600
VLIM  7  8 DC 0
VLP  91  0 DC 25
VLN   0 92 DC 25
.MODEL DX D(IS=800.0E-18)
.MODEL QX NPN(IS=800.0E-18 BF=62.50)
.ENDS
***********************************************************
.END

