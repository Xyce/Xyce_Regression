Test of BJT (Uniform Collector Doping) Photocurrent Model 
********************************************************************
* csradtckt1.cir
* Tier No.:  1
* Description:  
*
* Input:  Pulse representing radition dose level within the
*               model
* Output:       
* Circuit Elements: 
* Dose Rate:    
********************************************************************
* This netlist can be used to simulate at various rad levels by changing
* GRORDER (See note above).  The netlist include the basic MMBT2222 DC
* model parameters and the TF default and MMBT2222 model parameters
*------------------------------------------------------------------
*.options nonlin-tran reltol=1.0E-5 abstol=1.0E-6 deltaxtol=0.1 searchmethod=2
*+ maxsearchstep=10 maxstep=5000

Ib 3 0 DC -400E-6
VIB 3  8 0V
VC  4  0  2V
VIC 4  7  0V
VIE 9  0   0V
rxth dt 0 1e12
QNPN              7        8     9     dt   VND_0780

.MODEL VND_0780 
+ AFN=1.000
+ AJC=1.000m
+ AJE=1.000m
+ AJS=1.000m
+ ART=0.1
+ AVC1=Name
+ AVC2=Name
+ BFN=1.000
+ CBCO=0.000
+ CBEO=60.00f
+ CCSO=0
+ CJC=Name
+ CJCP=Name
+ CJE=Name
+ CJEP=0.000
+ CTH=0.000
+ DEAR=0
+ DTEMP=0
+ EA=1.529
+ EAIC=1.418
+ EAIE=1.533
+ EAIS=1.529
+ EANC=1.625
+ EANE=1.932
+ EANS=1.529
+ EAP=1.12
+ EBBE=0
+ FC=900.0m
+ GAMM=Name
+ HRCF=Name
+ IBBE=0.000001
+ IBCI=Name
+ IBCIP=0.000
+ IBCN=Name
+ IBCNP=0.000
+ IBEI=Name
+ IBEIP=0.000
+ IBEN=Name
+ IBENP=0.000
+ IKF=Name
+ IKP=Name
+ IKR=Name
+ IS=Name
+ ISP=Name
+ ISPMIN=0
+ ISRR=0.9247
+ ITF=0.000
+ KFN=0.000
+ MC=Name
+ ME=Name
+ MS=Name
+ NBBE=1
+ NCI=Name
+ NCIP=1.000
+ NCN=Name
+ NCNP=2.000
+ NEI=Name
+ NEN=Name
+ NF=Name
+ NFP=Name
+ NKF=0.5
+ NR=Name
+ PC=Name
+ PE=Name
+ PS=Name
+ QBM=0
+ QCO=Name
+ QTF=0.000
+ RBI=Name
+ RBP=1.000n
+ RBPMIN=0
+ RBX=Name
+ RCI=Name
+ RCX=Name
+ RE=Name
+ RS=Name
+ RTH=0.000
+ TAVC=0.000
+ TD=856.0f
+ TF=11.40p
+ TNBBE=0
+ TNF=-100.0u
+ TNOM=21.00
+ TR=11.40p
+ TVBBE1=0
+ TVBBE2=0
+ VBBE=7.7
+ VEF=0.000
+ VER=0.000
+ VO=Name
+ VRT=0
+ VTF=0.000
+ WBE=Name
+ WSP=1.000
+ XII=5.758
+ XIKF=0
+ XIN=1.903
+ XIS=3.834
+ XISR=0
+ XRB=0.000
+ XRBI=0
+ XRBP=0
+ XRBX=0
+ XRC=0.000
+ XRCI=0
+ XRCX=0
+ XRE=0.000
+ XRS=0.000
+ XTF=0.000
+ XVO=0.000

*.DC VB 0 1 1
*.DC Iecs 1e-4 1e-2 1e-4
.DC VC 0 10 0.25 Ib -5e-6 -100e-6 -10e-6
.PRINT DC   v(7) v(8) v(9) i(VIC) i(VIB) i(VIE)
*.TRAN 1.0E-5 .001 0.0 1.0E-5
*.PRINT TRAN FILE=csradtckt1b.prn v(1) v(3) v(4) v(5) v(6) v(10) i(VIC) i(VIB) i(VIE)
.END

