Test for DECADE capability in DC sweeps. Baseline
*
VT1 4 0 0V
R1  4 5 10
R2  5 0 5

.DC DEC VT1  0.1 100 4
.print DC V(4) V(5)

.END

