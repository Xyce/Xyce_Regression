Test of Function Handling in Expression Lib
********************************************************************************
* BUG 1085 was about the old expression library not being able to 
* handle .func names that started with "I" and had 2 characters.  It would
* confuse them with lead currents.
*
* This is the "reference" circuit, that does NOT include an I?-named .func
********************************************************************************
.func test(x,y) {y}
.func diff(x,y) {x-y}
.FUNC f(x,y,z) {diff(y,z)-4+test(z,x)**2}
VX  x  0  PWL(0 1v  1ms  2v  2ms  0v)
VY  y  0  PWL(0 2v  1ms  2v  2ms  0v)
VZ  z  0  PWL(0 3v  1ms  2v  2ms  1v)
BF  F  0  v = {f(v(x), v(y), v(z))}
RX  x  0  1M
RY  y  0  1M
RZ  z  0  1M
RF  f  0  1M
.TRAN 0.02MS 2MS
.PRINT TRAN v(x) v(y) v(z) v(f)
.END

