Simple RC circuit
**********************************************************************
*
* This circuit has the voltage source applied directly to the
* resistor, with the capacitor tied to ground.
*
**********************************************************************
Isrc 1 0 AC 1 0 sin(0 1 1e+5 0 0)
R1 1 0 {res}
C1 1 0 2e-6

.print ac v(1)  VR(1) VI(1) VM(1) VP(1) VDB(1)  {R1:R}

.global_param res=1e3

.data table
+ hertz  res
+ 1.00000000e+00	1.00000000e+00
+ 1.00000000e+01	1.00000000e+01
+ 1.00000000e+02	1.00000000e+02
+ 1.00000000e+03	1.00000000e+03
+ 1.00000000e+04	1.00000000e+04
+ 1.00000000e+05	1.00000000e+05
.enddata


*.AC DEC 10 1 1e5 
.AC data=table

.END
