* Test ERR, ERR1 and ERR2 measures.  This test is
* done via -remeasure because the measure values
* depend on the number of time-steps taken.
*
* See SON Bug 1278 for more details.
**************************************************

V3 3 0 2.5
R3 3 0 1

.TRAN 0 1
.PRINT TRAN V(1) V(2) V(3)

* Output the data at fixed time-steps, so that -remeasure
* gets a consistent answer on all platforms.
.OPTIONS OUTPUT INITIAL_INTERVAL=0.1

V1 1 0 PWL 0 0 1 5
R1 1 2 1
R2 2 0 3

.MEASURE TRAN ERR1MV1.5 ERR1 V(1) V(2) MINVAL=1.5
.MEASURE TRAN ERR1YMIN2.5 ERR1 V(1) V(3) YMIN=2.5
.MEASURE TRAN ERR1IGNOR2.5 ERR1 V(1) V(3) IGNOR=2.5
.MEASURE TRAN ERR1YMAX3.5 ERR1 V(1) V(3) YMAX=3.5
.MEASURE TRAN ERR1FT ERR1 {V(1)*V(1)} V(1) FROM=0.5 TO=0.8

.MEASURE TRAN ERR2MV1.5 ERR2 V(1) V(2) MINVAL=1.5
.MEASURE TRAN ERR2YMIN2.5 ERR2 V(1) V(3) YMIN=2.5
.MEASURE TRAN ERR2IGNOR2.5 ERR2 V(1) V(3) IGNOR=2.5
.MEASURE TRAN ERR2YMAX3.5 ERR2 V(1) V(3) YMAX=3.5
.MEASURE TRAN ERR2FT ERR2 {V(1)*V(1)} V(1) FROM=0.5 TO=0.8

.END
