* Xyce netlist for testing mixed current sources
.OPTIONS DEVICE TNOM=25

.TRAN  0 0.5ms 0
.PRINT TRAN FORMAT=PROBE V(1) V(2) I(R2)

IRAMP 1 0 EXP(0 0.2 2us 20us 40us 60us)
R1 1 2 100
R2 2 0 75

.END
