*Samle netlist for BSIM-MG
* Drain Noise Simulation 

**.option abstol=1e-6 reltol=1e-6 post ingold
*.options nonlin abstol=1e-6 reltol=1e-6
.options device temp=27

.include "modelcard.nmos_xyce_111"

* --- Voltage Sources ---
vds 1 0 dc 1v
vgs gate 0 dc 0.5v ac 1
vbs bulk 0 dc 0v

* --- Circuit ---
lbias 1 drain 1m
cload drain 2 1m
rload 2 0 1
M1 drain gate 0 bulk nmos1 TFIN=15n L=30n NFIN=10 NRS=1 NRD=1
M2 drain gate 0 bulk nmos1 TFIN=15n L=30n NFIN=10 NRS=1 NRD=1
M3 drain gate 0 bulk nmos1 TFIN=15n L=30n NFIN=10 NRS=1 NRD=1
M4 drain gate 0 bulk nmos1 TFIN=15n L=30n NFIN=10 NRS=1 NRD=1
M5 drain gate 0 bulk nmos1 TFIN=15n L=30n NFIN=10 NRS=1 NRD=1
M6 drain gate 0 bulk nmos1 TFIN=15n L=30n NFIN=10 NRS=1 NRD=1

* --- Analysis ---
.noise v(drain) vgs dec 11 1k 100g 1

.print noise inoise onoise

.end

