Power test for MOSFET Level 6
*
VDS 4 0  5V
VGS  1   0  pulse (0 1 1ns 1ns 1ns 1us 5us)
VMOND 4 3 0V
VMONS 0 2 0V
VMONG 1 1a 0
VMONB 0 6 0

M1 3 1a 2 6 CD4012_NMOS L=5u W=175u
.MODEL cd4012_nmos NMOS (
+ LEVEL = 6 UO = 190   VTO = 1.679  TOX = 6E-08   NSUB = 8.601E+15
+ NSS = 0     RS = 13.21   RD = 11.59   RSH = 0   IS = 1E-14
+ LD = 8.6E-07   L=5u W=175u lambda=0.02 GAMMA=0.37 PHI=0.65
+ CBD=0.1P CBS=0.1P PB=0.81 CGSO=2P CGBO=4P CGDO=2P CJ=2E-4 MJ=0.5 CJSW=1E-9
+ MJSW=0.5 JS=1E-8 TPG=0  FC=0.5 TNOM=27) 

.options timeint method=gear
.options nonlin-tran rhstol=1.0e-8
.tran 1ns 20us

* test that P(M1) and W(M1) are equal to the formula (Id*Vds + Ig*Vgs)
* and also equal to the combined power dissipation of the two
* source VDS and VGS.
.PRINT TRAN PRECISION=10 
+ P(M1) W(M1) {ID(M1)*V(4) + IG(M1)*V(1)} {-1*(P(VDS)+P(VGS))}
+ ID(M1) IG(M1) IS(M1) IB(M1) I(VDS) I(VGS) V(4) V(1) 

.END
