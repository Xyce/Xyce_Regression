***********************************************************
* AC test for .PRINT AC_IC without a .PRINT AC line.
* Netlist needs the .OP statement to get the AC_IC output.
* Also for "testing diversity", this netlist has the .OP
* statement before the .AC statement.
*
* Addresses SON Bug 942.
* *********************************************************

* Trivial high-pass filter
R1 b 0 2
C1 a b 1u
V1 a 0 DC 0V AC 1

.PRINT AC_IC R1:R vm(b)
.op
.ac dec 5 100Hz 1e6

.end
