Diode Circuit Netlist


VIN 1 0 PULSE ( 5 -1 0.05ms 100ns 100ns 0.1ms 0.2ms )
R1 1 2 2K
D1 3 0 DMOD
VMON 2 3 0

.global_param gpIS={100FA}
.param pIS={gpIS}

.step gpIS 100FA 150FA 10FA

.MODEL DMOD D (IS={pIS})
.TRAN 0 0.5ms
.options timeint reltol=1.0e-4
.PRINT TRAN I(VMON) V(3) {V(3)/I(VMON)}
*
.END
