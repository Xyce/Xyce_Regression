NPN Bipolar Circuit Netlist for MMBT2222LT, forward Gummels
************************************************************** 
VBB  6 0 0V
VMON1 6 1 0
VMON2 6 2 0
Q1 2 1 0 NBJT
.MODEL NBJT NPN (
+ IS=2.96E-14
+ BF=233.8
+ NF=1
+ ISE=2.30E-14
+ NE=1.780
+ VAF=2
+ IKF=0.340
*+ NK=0.5
+ NK=0.9

+ BR=1
+ NR=1
+ ISC=0
+ NC=2.0
+ VAR=100
+ IKR=1e99

* note that RB=RC for this problem (VBC=0)
+ RB=1.3
+ RC=1.3 
+ RE=0 )
.DC VBB 0.15 0.95 0.05
.PRINT DC V(6) I(VMON1) I(VMON2) 

.END
