
.tran 1ns 1ms
.print tran v(1)

r1   1   0   1
v3  $G_1  0  1

xg  $G_1 1  abc

.subckt abc $G_1 a
r2  $G_1 a 2
.ends

.end
