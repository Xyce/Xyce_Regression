* Test remeasure support for .DC analyses when the remeasured
* output file has a STEPNUM column.
*
**************************************************************

vsrc1   1a 0 1
rload1a 1a 1b 0.1
rload1b 1b 0 1

vsrc2   2a 0 1
rload2a 2a 1b 0.2

.DC vsrc1 1 16 2 vsrc2 2 5 3

.OPTIONS OUTPUT ADD_STEPNUM_COL=TRUE
.print dc vsrc1:DCV0 vsrc2:DCV0 v(1a) v(2a) v(1b)

* MAX measure
.measure dc maxv1b   max v(1b)

*MIN measure
.measure dc minv1b   min v(1b)

* PP measure
.measure dc ppv1b   pp v(1b)

.end
