** NMOSFET: Benchmarking Implementation of BSIM4.6.0 by Mohan V. Dunga 12/13/2006.

** Circuit Description **
m1 2 1 0 0 n1 L=0.09u W=10.0u rgeoMod=1
vgs 1 0 1.2 
vds 2 0 1.2

.dc vgs 0.0 1.18 0.02 vds 0.05 1.2 0.5 

.print dc v(1) v(2) i(vds)
*COMP i(vds) abstol=1e-5

.include modelcard.nmos
.end
