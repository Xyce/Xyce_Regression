* 51 stage Ring-Osc.

vin in out 2 pulse 2 0 0.1n 5n 1 1 1
vdd dd 0 1.0
*dc 0 pulse 0 2 0 1n 1 1 1
vss ss 0 dc 0
ve  sub  0 dc 0

xinv1 dd ss sub in out25 inv25 
xinv2 dd ss sub out25 out50 inv25
xinv5 dd ss sub out50 out inv1
xinv11 dd ss sub out buf inv1
cout  buf ss 1pF

xdum ss dum

*.option itl1=500 gmin=1e-15 itl4=10 
*.tran 0.2n 50n

.dc vdd 2 2 1

************************************
* **** Start Homotopy Setup ****
************************************
.options nonlin nlstrategy=0 searchmethod=0 
+ maxstep=50 maxsearchstep=20 continuation=1
 
.options loca stepper=1 stepcontrol=0
+ conparam=vdd
+ initialvalue=0.0 minvalue=-1.0 maxvalue=2.0
+ initialstepsize=0.02 minstepsize=0.02 maxstepsize=0.02 aggressiveness=1.0
+ maxsteps=5000 maxnliters=200
**********************************
* **** End Homotopy Setup ****
**********************************

.print dc v(in) v(out) 

.options device debuglevel=-5

*.include nmospd.mod
*.include pmospd.mod

.include nmos_3_2.mod
.include pmos_3_2.mod
.include lib.h
.end
