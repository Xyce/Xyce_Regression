Test IC formats (IC= vs. IC1= IC2= ) for U devices

*COMP v(sum1_out) reltol=0.02
*COMP v(carry1_out) reltol=0.02
*COMP v(sum2_out) reltol=0.02
*COMP v(carry2_out) reltol=0.02

* Analysis Commands
.options timeint reltol=1.0e-3
.tran 10ns 1us

* Analysis Commands
.options timeint reltol=1.0e-3
.tran 10ns 2us

* Sources
V1 in_1 0  PULSE ({V_HI} {V_LO} 100ns 20ns 20ns 80ns 200ns)
V2 in_2 0  PULSE ({V_HI} {V_LO} 100ns 20ns 20ns 180ns 400ns)
V3 carry_in 0  PULSE ({V_HI} {V_LO} 100ns 20ns 20ns 380ns 800ns)

* Output
.print tran PRECISION=10 WIDTH=19 v(in_1) v(in_2) v(carry_in) v(sum1_out)
+ v(carry1_out) v(sum2_out) v(carry2_out)

* Digital power and reference node
V4 dig_pn 0 3 

* Set digital default parameters:
.param R1HI=5 R1LO=200 R0HI=200 R0LO=5 RIN=1000 R1=100
.param SW=5.e-9  CAPOUT=1.e-12  CAPIN=1.e-12
.param V_LO=0 V_REF=0 V_HI=3

UADD1 ADD dig_pn 0 in_1 in_2 carry_in sum1_out carry1_out DMOD IC=FALSE,FALSE
UADD2 ADD dig_pn 0 in_1 in_2 carry_in sum2_out carry2_out DMOD IC1=FALSE IC2=FALSE

R1 sum1_out 0 100K
R2 carry1_out 0 100K
R3 sum2_out 0 100K
R4 carry2_out 0 100K

.model DMOD DIG ( CLO=CAPOUT  CHI=CAPOUT
+ S0RLO=R0LO  S0RHI=R0HI  S0TSW=SW
+ S0VLO=-1  S0VHI=1.8
+ S1RLO=R1LO  S1RHI=R1HI  S1TSW=SW
+ S1VLO=1  S1VHI=3
+ RLOAD=RIN   CLOAD=CAPIN
+ DELAY=20ns )

.end
