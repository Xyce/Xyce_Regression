level=1 diode circuit
*
R 1 2 0.0001
V2 2 0 0.21
V1 3 0 0.0
D2 1 3 DA

.MODEL DA D (RS=6.5e-05 IS=1.0e-09 N=1.037)

.print DC width=22 v(2) I(V1)  
.print SENS width=22 v(2) I(V1)  
.SENS objfunc={I(V1)} param=DA:RS,DA:IS
.options SENSITIVITY DAKOTAFILE=0  adjoint=1 direct=0  STDOUTPUT=0

.DC V2 0.005 2.0 0.005

.END

