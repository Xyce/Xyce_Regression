Test of global params in VSRC combined with no source stepping

.global_param dvdd = '1.8'

V1 1 0 'dvdd'
R1 1 2 1.0
R2 2 0 2.0

.DC R1 1.0 1.0 1.0
.PRINT dc V(2)
.end