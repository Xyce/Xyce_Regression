ram2k.sp SPICE FILE
.model nenh nmos
+ level = 2
+   vto = 0.761   kp = 3.843e-05   gamma = 0.639243
+   phi = 0.31
+
+   cgso = 3.54e-10   cgdo = 3.54e-10
+   rsh = 66   cj = 0.000343
+   mj = 1.067   cjsw = 1.83e-10   mjsw = 0.195
+   tox = 2.41e-08   nsub = 1.066e+16
+   nss = 3e+10   nfs = 4.55168e+12   tpg = 1
+   xj = 9e-07   ld = -1.68e-07   uo = 790
+   ucrit = 174667   uexp = 0.0461235
+   vmax = 177269   neff = 4.6883
+
+   delta = 0
.model penh pmos
+ level = 2
+   vto = -0.79   kp = 1.601e-05   gamma = 0.618101
+   phi = 0.541111
+
+   cgso = 4.01e-10   cgdo = 4.01e-10
+   rsh = 165   cj = 0.000499
+   mj = 0.341   cjsw = 2.34e-10   mjsw = 0.307
+   tox = 2.41e-08   nsub = 6.57544e+16
+   nss = 3e+10   nfs = 1.66844e+11   tpg = -1
+   xj = 1.12799e-07   ld = -1.38e-07   uo = 235
+   ucrit = 637449   uexp = 0.0888696
+   vmax = 63253.3   neff = 0.64354
+
+   delta = 0
m0 3 5 4 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m1 3 6 4 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m2 3 7 4 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m3 3 8 4 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m4 9 5 10 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=4.54e-12 ps=1.54e-05 pd=9.35e-06 
+ nrs=1.78 nrd=1.03 
m5 9 6 10 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=4.54e-12 ps=1.54e-05 pd=9.35e-06 
+ nrs=1.78 nrd=1.03 
m6 9 7 10 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=4.54e-12 ps=1.54e-05 pd=9.35e-06 
+ nrs=1.78 nrd=1.03 
m7 9 8 10 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=4.54e-12 ps=1.54e-05 pd=9.35e-06 
+ nrs=1.78 nrd=1.03 
m8 11 5 12 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=5.23e-12 ps=1.355e-05 pd=1.027e-05 
+ nrs=1.52 nrd=1.19 
m9 11 6 12 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=5.23e-12 ps=1.355e-05 pd=1.027e-05 
+ nrs=1.52 nrd=1.19 
m10 11 7 12 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=5.23e-12 ps=1.355e-05 pd=1.027e-05 
+ nrs=1.52 nrd=1.19 
m11 11 8 12 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=5.23e-12 ps=1.355e-05 pd=1.027e-05 
+ nrs=1.52 nrd=1.19 
m12 13 5 14 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.68e-12 ad=4.54e-12 ps=1.493e-05 pd=9.35e-06 
+ nrs=1.74 nrd=1.03 
m13 13 6 14 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.68e-12 ad=4.54e-12 ps=1.493e-05 pd=9.35e-06 
+ nrs=1.74 nrd=1.03 
m14 13 7 14 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.68e-12 ad=4.54e-12 ps=1.493e-05 pd=9.35e-06 
+ nrs=1.74 nrd=1.03 
m15 13 8 14 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.68e-12 ad=4.54e-12 ps=1.493e-05 pd=9.35e-06 
+ nrs=1.74 nrd=1.03 
m16 15 6 16 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m17 15 5 16 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m18 15 7 16 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m19 15 17 16 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m20 18 5 19 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m21 18 6 19 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m22 18 7 19 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m23 18 17 19 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m24 20 5 21 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.15e-12 ad=5.23e-12 ps=1.145e-05 pd=1.027e-05 
+ nrs=1.39 nrd=1.19 
m25 20 6 21 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.15e-12 ad=5.23e-12 ps=1.145e-05 pd=1.027e-05 
+ nrs=1.39 nrd=1.19 
m26 20 7 21 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.15e-12 ad=5.23e-12 ps=1.145e-05 pd=1.027e-05 
+ nrs=1.39 nrd=1.19 
m27 20 17 21 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.15e-12 ad=5.23e-12 ps=1.145e-05 pd=1.027e-05 
+ nrs=1.39 nrd=1.19 
m28 22 5 23 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m29 22 6 23 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m30 22 7 23 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m31 22 17 23 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m32 24 5 25 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m33 24 6 25 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m34 24 8 25 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m35 24 26 25 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m36 27 5 28 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m37 27 6 28 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m38 27 8 28 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m39 27 26 28 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m40 29 5 30 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m41 29 6 30 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m42 29 8 30 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m43 29 26 30 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m44 31 5 32 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.68e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m45 31 6 32 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.68e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m46 31 8 32 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.68e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m47 31 26 32 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.68e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m48 33 5 34 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m49 33 6 34 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m50 33 26 34 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m51 33 17 34 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m52 35 5 36 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m53 35 6 36 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m54 35 26 36 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m55 35 17 36 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m56 37 5 38 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m57 37 6 38 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m58 37 26 38 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m59 37 17 38 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m60 39 5 40 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m61 39 6 40 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m62 39 26 40 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m63 39 17 40 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m64 41 5 42 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.21e-12 ad=6.21e-12 ps=1.031e-05 pd=1.213e-05 
+ nrs=1.18 nrd=1.41 
m65 41 7 42 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.21e-12 ad=6.21e-12 ps=1.031e-05 pd=1.213e-05 
+ nrs=1.18 nrd=1.41 
m66 41 43 42 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.21e-12 ad=6.21e-12 ps=1.031e-05 pd=1.213e-05 
+ nrs=1.18 nrd=1.41 
m67 41 8 42 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.21e-12 ad=6.21e-12 ps=1.031e-05 pd=1.213e-05 
+ nrs=1.18 nrd=1.41 
m68 44 5 45 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m69 44 7 45 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m70 44 43 45 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m71 44 8 45 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m72 46 5 47 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m73 46 7 47 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m74 46 43 47 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m75 46 8 47 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m76 48 5 49 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=3.88e-12 ps=1.167e-05 pd=8.5e-06 
+ nrs=1.37 nrd=0.88 
m77 48 7 49 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=3.88e-12 ps=1.167e-05 pd=8.5e-06 
+ nrs=1.37 nrd=0.88 
m78 48 43 49 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=3.88e-12 ps=1.167e-05 pd=8.5e-06 
+ nrs=1.37 nrd=0.88 
m79 48 8 49 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=3.88e-12 ps=1.167e-05 pd=8.5e-06 
+ nrs=1.37 nrd=0.88 
m80 50 5 51 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m81 50 7 51 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m82 50 43 51 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m83 50 17 51 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m84 52 5 53 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m85 52 7 53 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m86 52 43 53 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m87 52 17 53 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m88 54 5 55 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m89 54 7 55 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m90 54 43 55 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m91 54 17 55 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m92 56 5 57 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m93 56 7 57 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m94 56 43 57 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m95 56 17 57 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m96 58 5 59 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=2.94e-12 ps=1.088e-05 pd=6.18e-06 
+ nrs=1.21 nrd=0.67 
m97 58 43 59 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=2.94e-12 ps=1.088e-05 pd=6.18e-06 
+ nrs=1.21 nrd=0.67 
m98 58 8 59 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=2.94e-12 ps=1.088e-05 pd=6.18e-06 
+ nrs=1.21 nrd=0.67 
m99 58 26 59 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=2.94e-12 ps=1.088e-05 pd=6.18e-06 
+ nrs=1.21 nrd=0.67 
m100 60 5 61 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m101 60 43 61 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m102 60 8 61 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m103 60 26 61 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m104 62 5 63 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m105 62 43 63 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m106 62 8 63 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m107 62 26 63 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m108 64 5 65 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m109 64 43 65 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m110 64 8 65 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m111 64 26 65 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m112 66 5 67 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m113 66 43 67 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m114 66 26 67 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m115 66 17 67 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m116 68 5 69 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=4.28e-12 ps=1.213e-05 pd=9.16e-06 
+ nrs=1.41 nrd=0.97 
m117 68 43 69 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=4.28e-12 ps=1.213e-05 pd=9.16e-06 
+ nrs=1.41 nrd=0.97 
m118 68 26 69 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=4.28e-12 ps=1.213e-05 pd=9.16e-06 
+ nrs=1.41 nrd=0.97 
m119 68 17 69 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=4.28e-12 ps=1.213e-05 pd=9.16e-06 
+ nrs=1.41 nrd=0.97 
m120 70 5 71 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m121 70 43 71 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m122 70 26 71 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m123 70 17 71 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m124 72 5 73 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m125 72 43 73 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m126 72 26 73 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m127 72 17 73 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m128 74 6 75 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m129 74 76 75 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m130 74 7 75 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m131 74 8 75 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m132 77 6 78 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m133 77 76 78 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m134 77 7 78 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m135 77 8 78 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m136 79 6 80 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=8.98e-06 
+ nrs=1.03 nrd=1.19 
m137 79 76 80 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=8.98e-06 
+ nrs=1.03 nrd=1.19 
m138 79 7 80 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=8.98e-06 
+ nrs=1.03 nrd=1.19 
m139 79 8 80 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=8.98e-06 
+ nrs=1.03 nrd=1.19 
m140 81 6 82 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m141 81 76 82 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m142 81 7 82 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m143 81 8 82 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m144 83 6 84 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m145 83 76 84 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m146 83 7 84 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m147 83 17 84 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m148 85 6 86 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m149 85 76 86 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m150 85 7 86 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m151 85 17 86 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m152 87 6 88 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m153 87 76 88 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m154 87 7 88 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m155 87 17 88 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m156 89 6 90 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.72e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.3 nrd=1.03 
m157 89 76 90 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.72e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.3 nrd=1.03 
m158 89 7 90 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.72e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.3 nrd=1.03 
m159 89 17 90 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.72e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.3 nrd=1.03 
m160 91 6 92 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m161 91 76 92 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m162 91 8 92 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m163 91 26 92 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m164 93 6 94 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m165 93 76 94 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m166 93 8 94 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m167 93 26 94 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m168 95 6 96 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m169 95 76 96 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m170 95 8 96 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m171 95 26 96 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m172 97 6 98 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m173 97 76 98 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m174 97 8 98 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m175 97 26 98 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m176 99 6 100 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m177 99 76 100 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m178 99 26 100 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m179 99 17 100 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m180 101 6 102 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m181 101 76 102 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m182 101 26 102 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m183 101 17 102 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m184 103 6 104 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m185 103 76 104 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m186 103 26 104 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m187 103 17 104 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m188 105 6 106 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m189 105 76 106 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m190 105 26 106 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m191 105 17 106 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m192 107 76 108 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m193 107 7 108 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m194 107 43 108 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m195 107 8 108 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m196 109 76 110 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.155e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m197 109 7 110 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.155e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m198 109 43 110 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.155e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m199 109 8 110 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.155e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m200 111 76 112 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m201 111 7 112 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m202 111 43 112 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m203 111 8 112 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m204 113 76 114 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m205 113 7 114 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m206 113 43 114 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m207 113 8 114 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m208 115 76 116 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m209 115 7 116 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m210 115 43 116 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m211 115 17 116 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m212 117 76 118 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m213 117 7 118 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m214 117 43 118 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m215 117 17 118 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m216 119 76 120 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.81e-12 ad=6.21e-12 ps=8.5e-06 pd=1.213e-05 
+ nrs=1.09 nrd=1.41 
m217 119 7 120 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.81e-12 ad=6.21e-12 ps=8.5e-06 pd=1.213e-05 
+ nrs=1.09 nrd=1.41 
m218 119 43 120 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.81e-12 ad=6.21e-12 ps=8.5e-06 pd=1.213e-05 
+ nrs=1.09 nrd=1.41 
m219 119 17 120 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.81e-12 ad=6.21e-12 ps=8.5e-06 pd=1.213e-05 
+ nrs=1.09 nrd=1.41 
m220 121 76 122 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m221 121 7 122 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m222 121 43 122 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m223 121 17 122 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m224 123 76 124 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m225 123 43 124 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m226 123 8 124 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m227 123 26 124 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m228 125 76 126 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=2.67e-12 ps=1.213e-05 pd=5.92e-06 
+ nrs=1.41 nrd=0.61 
m229 125 43 126 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=2.67e-12 ps=1.213e-05 pd=5.92e-06 
+ nrs=1.41 nrd=0.61 
m230 125 8 126 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=2.67e-12 ps=1.213e-05 pd=5.92e-06 
+ nrs=1.41 nrd=0.61 
m231 125 26 126 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=2.67e-12 ps=1.213e-05 pd=5.92e-06 
+ nrs=1.41 nrd=0.61 
m232 127 76 128 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m233 127 43 128 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m234 127 8 128 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m235 127 26 128 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m236 129 76 130 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m237 129 43 130 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m238 129 8 130 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m239 129 26 130 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m240 131 76 132 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m241 131 43 132 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m242 131 26 132 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m243 131 17 132 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m244 133 76 134 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m245 133 43 134 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m246 133 26 134 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m247 133 17 134 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m248 135 76 136 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m249 135 43 136 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m250 135 26 136 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m251 135 17 136 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m252 137 76 138 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m253 137 43 138 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m254 137 26 138 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m255 137 17 138 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m256 1 140 139 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m257 141 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m258 1 140 142 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m259 143 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m260 1 140 144 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m261 145 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m262 1 140 146 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=9.8e-12 ps=1.734e-05 pd=1.68e-05 
+ nrs=0.95 nrd=0.56 
m263 147 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=9.8e-12 ad=1.678e-11 ps=1.68e-05 pd=1.734e-05 
+ nrs=0.56 nrd=0.95 
m264 1 5 76 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m265 1 6 43 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m266 1 7 26 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m267 1 8 17 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m268 1 149 148 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m269 1 151 150 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m270 152 153 139 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.277e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=1.05 
m271 154 153 141 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m272 155 156 142 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m273 157 156 143 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m274 158 159 144 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m275 160 159 145 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m276 161 162 146 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m277 163 162 147 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.089e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.99 
m278 0 164 152 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m279 0 165 154 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m280 0 164 155 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m281 0 165 157 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m282 0 164 158 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m283 0 165 160 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m284 0 164 161 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m285 0 165 163 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m286 0 5 76 0 nenh l=1.1e-06 w=9.1e-06 
+ as=2.709e-11 ad=1.078e-11 ps=2.848e-05 pd=2.38e-05 
+ nrs=0.33 nrd=0.13 
m287 0 6 43 0 nenh l=1.1e-06 w=9.1e-06 
+ as=2.709e-11 ad=1.078e-11 ps=2.848e-05 pd=2.38e-05 
+ nrs=0.33 nrd=0.13 
m288 0 7 26 0 nenh l=1.1e-06 w=9.1e-06 
+ as=2.709e-11 ad=1.078e-11 ps=2.848e-05 pd=2.38e-05 
+ nrs=0.33 nrd=0.13 
m289 0 8 17 0 nenh l=1.1e-06 w=1.05e-05 
+ as=3.125e-11 ad=1.47e-11 ps=3.287e-05 pd=2.66e-05 
+ nrs=0.28 nrd=0.13 
m290 0 149 148 0 nenh l=1.1e-06 w=1.05e-05 
+ as=3.125e-11 ad=1.47e-11 ps=3.287e-05 pd=2.66e-05 
+ nrs=0.28 nrd=0.13 
m291 0 151 150 0 nenh l=1.1e-06 w=1.05e-05 
+ as=3.125e-11 ad=1.47e-11 ps=3.287e-05 pd=2.66e-05 
+ nrs=0.28 nrd=0.13 
m292 166 167 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m293 166 167 0 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=2.917e-11 ps=2.1e-05 pd=3.068e-05 
+ nrs=0.07 nrd=0.3 
m294 168 169 0 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=2.917e-11 ps=2.1e-05 pd=3.068e-05 
+ nrs=0.07 nrd=0.3 
m295 170 169 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=1.19e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m296 162 171 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m297 162 171 0 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=2.917e-11 ps=2.1e-05 pd=3.068e-05 
+ nrs=0.07 nrd=0.3 
m298 0 172 168 0 nenh l=1.1e-06 w=9.8e-06 
+ as=2.917e-11 ad=6.86e-12 ps=3.068e-05 pd=2.1e-05 
+ nrs=0.3 nrd=0.07 
m299 168 172 170 1 penh l=1.1e-06 w=1.05e-05 
+ as=8.33e-12 ad=7.35e-12 ps=2.52e-05 pd=1.19e-05 
+ nrs=0.08 nrd=0.07 
m300 1 167 173 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m301 174 167 173 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=6.86e-12 ps=1.12e-05 pd=2.1e-05 
+ nrs=0.07 nrd=0.07 
m302 175 1 174 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=6.86e-12 ps=1.12e-05 pd=1.12e-05 
+ nrs=0.07 nrd=0.07 
m303 1 167 171 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m304 176 167 171 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=6.86e-12 ps=1.12e-05 pd=2.1e-05 
+ nrs=0.07 nrd=0.07 
m305 0 165 164 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m306 0 177 165 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m307 178 165 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=4.2e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m308 177 140 178 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=4.2e-06 
+ nrs=0.25 nrd=0.25 
m309 179 172 177 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m310 0 180 179 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m311 181 179 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=7e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m312 0 182 181 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m313 180 183 181 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m314 184 185 180 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m315 156 173 0 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=2.917e-11 ps=2.1e-05 pd=3.068e-05 
+ nrs=0.07 nrd=0.3 
m316 156 173 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m317 173 1 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m318 0 168 175 0 nenh l=1.1e-06 w=9.8e-06 
+ as=2.917e-11 ad=6.86e-12 ps=3.068e-05 pd=1.12e-05 
+ nrs=0.3 nrd=0.07 
m319 186 187 176 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=6.86e-12 ps=1.12e-05 pd=1.12e-05 
+ nrs=0.07 nrd=0.07 
m320 171 187 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m321 0 168 186 0 nenh l=1.1e-06 w=9.8e-06 
+ as=2.917e-11 ad=6.86e-12 ps=3.068e-05 pd=1.12e-05 
+ nrs=0.3 nrd=0.07 
m322 1 168 173 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m323 1 165 164 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m324 1 177 165 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m325 188 165 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=2.94e-12 ad=1.678e-11 ps=5.6e-06 pd=1.734e-05 
+ nrs=0.17 nrd=0.95 
m326 177 172 188 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=2.94e-12 ps=1.4e-05 pd=5.6e-06 
+ nrs=0.28 nrd=0.17 
m327 179 140 177 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m328 1 180 179 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.4e-05 
+ nrs=0.95 nrd=0.28 
m329 189 179 1 1 penh l=1.1e-06 w=8.4e-06 
+ as=5.88e-12 ad=3.355e-11 ps=9.8e-06 pd=3.468e-05 
+ nrs=0.08 nrd=0.48 
m330 181 182 189 1 penh l=1.1e-06 w=8.4e-06 
+ as=9.8e-12 ad=5.88e-12 ps=2.613e-05 pd=9.8e-06 
+ nrs=0.14 nrd=0.08 
m331 1 168 171 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m332 180 185 181 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.307e-05 
+ nrs=0.28 nrd=0.28 
m333 184 183 180 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.54e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m334 190 168 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m335 191 168 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m336 0 190 153 0 nenh l=1.1e-06 w=9.8e-06 
+ as=2.917e-11 ad=6.86e-12 ps=3.068e-05 pd=2.1e-05 
+ nrs=0.3 nrd=0.07 
m337 1 190 153 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m338 1 1 190 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m339 192 168 0 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=2.917e-11 ps=1.12e-05 pd=3.068e-05 
+ nrs=0.07 nrd=0.3 
m340 193 168 0 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=2.917e-11 ps=1.12e-05 pd=3.068e-05 
+ nrs=0.07 nrd=0.3 
m341 1 187 191 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m342 194 1 192 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=6.86e-12 ps=1.12e-05 pd=1.12e-05 
+ nrs=0.07 nrd=0.07 
m343 190 166 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m344 190 166 194 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=6.86e-12 ps=2.1e-05 pd=1.12e-05 
+ nrs=0.07 nrd=0.07 
m345 195 187 193 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=6.86e-12 ps=1.12e-05 pd=1.12e-05 
+ nrs=0.07 nrd=0.07 
m346 191 166 195 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=6.86e-12 ps=2.1e-05 pd=1.12e-05 
+ nrs=0.07 nrd=0.07 
m347 191 166 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m348 1 191 159 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m349 0 191 159 0 nenh l=1.1e-06 w=9.8e-06 
+ as=2.917e-11 ad=6.86e-12 ps=3.068e-05 pd=2.1e-05 
+ nrs=0.3 nrd=0.07 
m350 0 187 1 0 nenh l=1.1e-06 w=9.8e-06 
+ as=2.917e-11 ad=6.86e-12 ps=3.068e-05 pd=2.1e-05 
+ nrs=0.3 nrd=0.07 
m351 1 187 1 1 penh l=1.1e-06 w=1.54e-05 
+ as=6.151e-11 ad=6.151e-11 ps=6.359e-05 pd=6.359e-05 
+ nrs=0.26 nrd=0.26 
m352 1 140 196 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m353 197 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m354 1 140 198 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m355 199 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m356 1 140 200 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m357 201 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m358 1 140 202 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=9.8e-12 ps=1.734e-05 pd=1.68e-05 
+ nrs=0.95 nrd=0.56 
m359 203 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=9.8e-12 ad=1.678e-11 ps=1.68e-05 pd=1.734e-05 
+ nrs=0.56 nrd=0.95 
m360 204 153 196 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.277e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=1.05 
m361 205 153 197 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m362 206 156 198 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m363 207 156 199 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m364 208 159 200 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m365 209 159 201 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m366 210 162 202 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m367 211 162 203 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.089e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.99 
m368 0 212 204 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m369 0 213 205 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m370 0 212 206 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m371 0 213 207 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m372 0 212 208 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m373 0 213 209 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m374 0 212 210 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m375 0 213 211 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m376 0 213 212 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m377 0 214 213 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m378 215 213 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=4.2e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m379 214 140 215 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=4.2e-06 
+ nrs=0.25 nrd=0.25 
m380 216 172 214 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m381 0 217 216 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m382 218 216 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=7e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m383 0 182 218 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m384 217 183 218 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m385 219 185 217 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m386 1 213 212 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m387 1 214 213 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m388 220 213 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=2.94e-12 ad=1.678e-11 ps=5.6e-06 pd=1.734e-05 
+ nrs=0.17 nrd=0.95 
m389 214 172 220 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=2.94e-12 ps=1.4e-05 pd=5.6e-06 
+ nrs=0.28 nrd=0.17 
m390 216 140 214 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m391 1 217 216 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.4e-05 
+ nrs=0.95 nrd=0.28 
m392 221 216 1 1 penh l=1.1e-06 w=8.4e-06 
+ as=5.88e-12 ad=3.355e-11 ps=9.8e-06 pd=3.468e-05 
+ nrs=0.08 nrd=0.48 
m393 218 182 221 1 penh l=1.1e-06 w=8.4e-06 
+ as=9.8e-12 ad=5.88e-12 ps=2.613e-05 pd=9.8e-06 
+ nrs=0.14 nrd=0.08 
m394 217 185 218 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.307e-05 
+ nrs=0.28 nrd=0.28 
m395 219 183 217 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.54e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m396 1 140 222 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m397 223 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m398 1 140 224 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m399 225 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m400 1 140 226 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m401 227 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m402 1 140 228 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=9.8e-12 ps=1.734e-05 pd=1.68e-05 
+ nrs=0.95 nrd=0.56 
m403 229 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=9.8e-12 ad=1.678e-11 ps=1.68e-05 pd=1.734e-05 
+ nrs=0.56 nrd=0.95 
m404 230 153 222 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.277e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=1.05 
m405 231 153 223 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m406 232 156 224 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m407 233 156 225 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m408 234 159 226 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m409 235 159 227 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m410 236 162 228 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m411 237 162 229 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.089e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.99 
m412 0 238 230 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m413 0 239 231 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m414 0 238 232 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m415 0 239 233 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m416 0 238 234 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m417 0 239 235 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m418 0 238 236 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m419 0 239 237 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m420 0 239 238 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m421 0 240 239 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m422 241 239 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=4.2e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m423 240 140 241 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=4.2e-06 
+ nrs=0.25 nrd=0.25 
m424 242 172 240 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m425 0 243 242 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m426 244 242 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=7e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m427 0 182 244 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m428 243 183 244 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m429 245 185 243 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m430 1 239 238 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m431 1 240 239 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m432 246 239 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=2.94e-12 ad=1.678e-11 ps=5.6e-06 pd=1.734e-05 
+ nrs=0.17 nrd=0.95 
m433 240 172 246 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=2.94e-12 ps=1.4e-05 pd=5.6e-06 
+ nrs=0.28 nrd=0.17 
m434 242 140 240 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m435 1 243 242 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.4e-05 
+ nrs=0.95 nrd=0.28 
m436 247 242 1 1 penh l=1.1e-06 w=8.4e-06 
+ as=5.88e-12 ad=3.355e-11 ps=9.8e-06 pd=3.468e-05 
+ nrs=0.08 nrd=0.48 
m437 244 182 247 1 penh l=1.1e-06 w=8.4e-06 
+ as=9.8e-12 ad=5.88e-12 ps=2.613e-05 pd=9.8e-06 
+ nrs=0.14 nrd=0.08 
m438 243 185 244 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.307e-05 
+ nrs=0.28 nrd=0.28 
m439 245 183 243 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.54e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m440 1 140 248 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m441 249 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m442 1 140 250 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m443 251 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m444 1 140 252 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m445 253 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m446 1 140 254 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=9.8e-12 ps=1.734e-05 pd=1.68e-05 
+ nrs=0.95 nrd=0.56 
m447 255 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=9.8e-12 ad=1.678e-11 ps=1.68e-05 pd=1.734e-05 
+ nrs=0.56 nrd=0.95 
m448 256 153 248 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.277e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=1.05 
m449 257 153 249 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m450 258 156 250 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m451 259 156 251 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m452 260 159 252 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m453 261 159 253 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m454 262 162 254 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m455 263 162 255 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.089e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.99 
m456 0 264 256 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m457 0 265 257 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m458 0 264 258 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m459 0 265 259 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m460 0 264 260 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m461 0 265 261 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m462 0 264 262 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m463 0 265 263 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m464 0 265 264 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m465 0 266 265 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m466 267 265 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=4.2e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m467 266 140 267 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=4.2e-06 
+ nrs=0.25 nrd=0.25 
m468 268 172 266 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m469 0 269 268 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m470 270 268 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=7e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m471 0 182 270 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m472 269 183 270 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m473 271 185 269 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m474 1 265 264 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m475 1 266 265 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m476 272 265 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=2.94e-12 ad=1.678e-11 ps=5.6e-06 pd=1.734e-05 
+ nrs=0.17 nrd=0.95 
m477 266 172 272 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=2.94e-12 ps=1.4e-05 pd=5.6e-06 
+ nrs=0.28 nrd=0.17 
m478 268 140 266 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m479 1 269 268 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.4e-05 
+ nrs=0.95 nrd=0.28 
m480 273 268 1 1 penh l=1.1e-06 w=8.4e-06 
+ as=5.88e-12 ad=3.355e-11 ps=9.8e-06 pd=3.468e-05 
+ nrs=0.08 nrd=0.48 
m481 270 182 273 1 penh l=1.1e-06 w=8.4e-06 
+ as=9.8e-12 ad=5.88e-12 ps=2.613e-05 pd=9.8e-06 
+ nrs=0.14 nrd=0.08 
m482 269 185 270 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.307e-05 
+ nrs=0.28 nrd=0.28 
m483 271 183 269 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.54e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m484 1 140 274 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m485 275 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m486 1 140 276 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m487 277 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m488 1 140 278 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m489 279 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m490 1 140 280 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=9.8e-12 ps=1.734e-05 pd=1.68e-05 
+ nrs=0.95 nrd=0.56 
m491 281 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=9.8e-12 ad=1.678e-11 ps=1.68e-05 pd=1.734e-05 
+ nrs=0.56 nrd=0.95 
m492 282 153 274 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.277e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=1.05 
m493 283 153 275 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m494 284 156 276 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m495 285 156 277 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m496 286 159 278 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m497 287 159 279 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m498 288 162 280 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m499 289 162 281 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.089e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.99 
m500 0 290 282 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m501 0 291 283 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m502 0 290 284 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m503 0 291 285 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m504 0 290 286 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m505 0 291 287 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m506 0 290 288 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m507 0 291 289 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m508 0 291 290 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m509 0 292 291 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m510 293 291 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=4.2e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m511 292 140 293 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=4.2e-06 
+ nrs=0.25 nrd=0.25 
m512 294 172 292 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m513 0 295 294 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m514 296 294 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=7e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m515 0 182 296 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m516 295 183 296 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m517 297 185 295 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m518 1 291 290 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m519 1 292 291 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m520 298 291 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=2.94e-12 ad=1.678e-11 ps=5.6e-06 pd=1.734e-05 
+ nrs=0.17 nrd=0.95 
m521 292 172 298 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=2.94e-12 ps=1.4e-05 pd=5.6e-06 
+ nrs=0.28 nrd=0.17 
m522 294 140 292 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m523 1 295 294 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.4e-05 
+ nrs=0.95 nrd=0.28 
m524 299 294 1 1 penh l=1.1e-06 w=8.4e-06 
+ as=5.88e-12 ad=3.355e-11 ps=9.8e-06 pd=3.468e-05 
+ nrs=0.08 nrd=0.48 
m525 296 182 299 1 penh l=1.1e-06 w=8.4e-06 
+ as=9.8e-12 ad=5.88e-12 ps=2.613e-05 pd=9.8e-06 
+ nrs=0.14 nrd=0.08 
m526 295 185 296 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.307e-05 
+ nrs=0.28 nrd=0.28 
m527 297 183 295 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.54e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m528 1 140 300 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m529 301 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m530 1 140 302 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m531 303 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m532 1 140 304 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m533 305 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m534 1 140 306 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=9.8e-12 ps=1.734e-05 pd=1.68e-05 
+ nrs=0.95 nrd=0.56 
m535 307 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=9.8e-12 ad=1.678e-11 ps=1.68e-05 pd=1.734e-05 
+ nrs=0.56 nrd=0.95 
m536 308 153 300 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.277e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=1.05 
m537 309 153 301 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m538 310 156 302 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m539 311 156 303 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m540 312 159 304 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m541 313 159 305 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m542 314 162 306 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m543 315 162 307 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.089e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.99 
m544 0 316 308 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m545 0 317 309 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m546 0 316 310 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m547 0 317 311 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m548 0 316 312 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m549 0 317 313 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m550 0 316 314 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m551 0 317 315 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m552 0 317 316 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m553 0 318 317 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m554 319 317 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=4.2e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m555 318 140 319 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=4.2e-06 
+ nrs=0.25 nrd=0.25 
m556 320 172 318 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m557 0 321 320 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m558 322 320 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=7e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m559 0 182 322 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m560 321 183 322 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m561 323 185 321 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m562 1 317 316 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m563 1 318 317 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m564 324 317 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=2.94e-12 ad=1.678e-11 ps=5.6e-06 pd=1.734e-05 
+ nrs=0.17 nrd=0.95 
m565 318 172 324 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=2.94e-12 ps=1.4e-05 pd=5.6e-06 
+ nrs=0.28 nrd=0.17 
m566 320 140 318 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m567 1 321 320 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.4e-05 
+ nrs=0.95 nrd=0.28 
m568 325 320 1 1 penh l=1.1e-06 w=8.4e-06 
+ as=5.88e-12 ad=3.355e-11 ps=9.8e-06 pd=3.468e-05 
+ nrs=0.08 nrd=0.48 
m569 322 182 325 1 penh l=1.1e-06 w=8.4e-06 
+ as=9.8e-12 ad=5.88e-12 ps=2.613e-05 pd=9.8e-06 
+ nrs=0.14 nrd=0.08 
m570 321 185 322 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.307e-05 
+ nrs=0.28 nrd=0.28 
m571 323 183 321 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.54e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m572 1 140 326 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m573 327 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m574 1 140 328 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m575 329 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m576 1 140 330 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m577 331 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m578 1 140 332 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=9.8e-12 ps=1.734e-05 pd=1.68e-05 
+ nrs=0.95 nrd=0.56 
m579 333 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=9.8e-12 ad=1.678e-11 ps=1.68e-05 pd=1.734e-05 
+ nrs=0.56 nrd=0.95 
m580 334 153 326 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.277e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=1.05 
m581 335 153 327 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m582 336 156 328 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m583 337 156 329 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m584 338 159 330 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m585 339 159 331 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m586 340 162 332 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m587 341 162 333 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.089e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.99 
m588 0 342 334 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m589 0 343 335 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m590 0 342 336 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m591 0 343 337 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m592 0 342 338 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m593 0 343 339 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m594 0 342 340 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m595 0 343 341 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m596 0 343 342 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m597 0 344 343 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m598 345 343 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=4.2e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m599 344 140 345 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=4.2e-06 
+ nrs=0.25 nrd=0.25 
m600 346 172 344 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m601 0 347 346 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m602 348 346 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=7e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m603 0 182 348 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m604 347 183 348 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m605 349 185 347 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m606 1 343 342 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m607 1 344 343 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m608 350 343 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=2.94e-12 ad=1.678e-11 ps=5.6e-06 pd=1.734e-05 
+ nrs=0.17 nrd=0.95 
m609 344 172 350 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=2.94e-12 ps=1.4e-05 pd=5.6e-06 
+ nrs=0.28 nrd=0.17 
m610 346 140 344 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m611 1 347 346 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.4e-05 
+ nrs=0.95 nrd=0.28 
m612 351 346 1 1 penh l=1.1e-06 w=8.4e-06 
+ as=5.88e-12 ad=3.355e-11 ps=9.8e-06 pd=3.468e-05 
+ nrs=0.08 nrd=0.48 
m613 348 182 351 1 penh l=1.1e-06 w=8.4e-06 
+ as=9.8e-12 ad=5.88e-12 ps=2.613e-05 pd=9.8e-06 
+ nrs=0.14 nrd=0.08 
m614 347 185 348 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.307e-05 
+ nrs=0.28 nrd=0.28 
m615 349 183 347 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.54e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m616 1 140 352 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m617 353 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m618 1 140 354 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m619 355 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m620 1 140 356 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=1.274e-11 ps=1.734e-05 pd=1.82e-05 
+ nrs=0.95 nrd=0.72 
m621 357 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.274e-11 ad=1.678e-11 ps=1.82e-05 pd=1.734e-05 
+ nrs=0.72 nrd=0.95 
m622 1 140 358 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=9.8e-12 ps=1.734e-05 pd=1.68e-05 
+ nrs=0.95 nrd=0.56 
m623 359 140 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=9.8e-12 ad=1.678e-11 ps=1.68e-05 pd=1.734e-05 
+ nrs=0.56 nrd=0.95 
m624 360 153 352 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.277e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=1.05 
m625 361 153 353 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m626 362 156 354 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m627 363 156 355 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m628 364 159 356 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.901e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.93 
m629 365 159 357 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m630 366 162 358 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.524e-11 ps=7e-06 pd=3.814e-05 
+ nrs=0.12 nrd=0.81 
m631 367 162 359 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=3.089e-11 ps=7e-06 pd=3.993e-05 
+ nrs=0.12 nrd=0.99 
m632 0 368 360 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m633 0 369 361 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m634 0 368 362 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m635 0 369 363 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m636 0 368 364 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m637 0 369 365 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m638 0 368 366 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m639 0 369 367 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=7e-06 
+ nrs=0.53 nrd=0.12 
m640 0 369 368 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m641 0 370 369 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m642 371 369 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=4.2e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m643 370 140 371 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=4.2e-06 
+ nrs=0.25 nrd=0.25 
m644 372 172 370 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m645 0 373 372 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m646 374 372 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=8.33e-12 ps=7e-06 pd=8.76e-06 
+ nrs=0.25 nrd=1.06 
m647 0 182 374 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=1.96e-12 ps=8.76e-06 pd=7e-06 
+ nrs=1.06 nrd=0.25 
m648 373 183 374 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m649 375 185 373 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=1.96e-12 ps=7e-06 pd=7e-06 
+ nrs=0.25 nrd=0.25 
m650 1 369 368 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m651 1 370 369 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.54e-05 
+ nrs=0.95 nrd=0.28 
m652 376 369 1 1 penh l=1.1e-06 w=4.2e-06 
+ as=2.94e-12 ad=1.678e-11 ps=5.6e-06 pd=1.734e-05 
+ nrs=0.17 nrd=0.95 
m653 370 172 376 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=2.94e-12 ps=1.4e-05 pd=5.6e-06 
+ nrs=0.28 nrd=0.17 
m654 372 140 370 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m655 1 373 372 1 penh l=1.1e-06 w=4.2e-06 
+ as=1.678e-11 ad=4.9e-12 ps=1.734e-05 pd=1.4e-05 
+ nrs=0.95 nrd=0.28 
m656 377 372 1 1 penh l=1.1e-06 w=8.4e-06 
+ as=5.88e-12 ad=3.355e-11 ps=9.8e-06 pd=3.468e-05 
+ nrs=0.08 nrd=0.48 
m657 374 182 377 1 penh l=1.1e-06 w=8.4e-06 
+ as=9.8e-12 ad=5.88e-12 ps=2.613e-05 pd=9.8e-06 
+ nrs=0.14 nrd=0.08 
m658 373 185 374 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.4e-05 pd=1.307e-05 
+ nrs=0.28 nrd=0.28 
m659 375 183 373 1 penh l=1.1e-06 w=4.2e-06 
+ as=4.9e-12 ad=4.9e-12 ps=1.54e-05 pd=1.4e-05 
+ nrs=0.28 nrd=0.28 
m660 378 132 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m661 379 185 378 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m662 1 140 132 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m663 380 379 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m664 380 379 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m665 131 149 132 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m666 131 151 132 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m667 131 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.13e-12 ad=8.33e-12 ps=1.451e-05 pd=8.76e-06 
+ nrs=0.91 nrd=1.06 
m668 381 380 379 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m669 0 140 381 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m670 1 140 379 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m671 382 383 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m672 384 140 382 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m673 1 384 383 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m674 0 384 383 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m675 384 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m676 133 149 134 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m677 385 133 384 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m678 0 140 134 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=7.13e-12 ps=8.76e-06 pd=1.451e-05 
+ nrs=1.06 nrd=0.91 
m679 0 185 385 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m680 133 150 134 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m681 1 140 133 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m682 136 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m683 386 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m684 387 136 386 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m685 388 387 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m686 388 387 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m687 135 151 136 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m688 135 148 136 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m689 135 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.13e-12 ad=8.33e-12 ps=1.451e-05 pd=8.76e-06 
+ nrs=0.91 nrd=1.06 
m690 389 388 387 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m691 1 140 387 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m692 0 140 389 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m693 390 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m694 391 392 390 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m695 391 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m696 1 391 392 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m697 0 391 392 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m698 0 140 138 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=7.13e-12 ps=8.76e-06 pd=1.451e-05 
+ nrs=1.06 nrd=0.91 
m699 393 137 391 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m700 137 148 138 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m701 137 150 138 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m702 0 185 393 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m703 1 140 137 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m704 394 124 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m705 395 185 394 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m706 1 140 124 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m707 396 395 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m708 396 395 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m709 123 149 124 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m710 123 151 124 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m711 123 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.13e-12 ad=8.33e-12 ps=1.451e-05 pd=8.76e-06 
+ nrs=0.91 nrd=1.06 
m712 397 396 395 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m713 0 140 397 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m714 1 140 395 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m715 398 399 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m716 400 140 398 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m717 1 400 399 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m718 0 400 399 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m719 400 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m720 125 149 126 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=2.67e-12 ps=1.213e-05 pd=5.92e-06 
+ nrs=1.41 nrd=0.61 
m721 401 125 400 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m722 0 140 126 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=3.56e-12 ps=8.76e-06 pd=7.89e-06 
+ nrs=1.06 nrd=0.45 
m723 0 185 401 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m724 125 150 126 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=2.67e-12 ps=1.213e-05 pd=5.92e-06 
+ nrs=1.41 nrd=0.61 
m725 1 140 125 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m726 128 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m727 402 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m728 403 128 402 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m729 404 403 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m730 404 403 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m731 127 151 128 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m732 127 148 128 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m733 127 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.13e-12 ad=8.33e-12 ps=1.451e-05 pd=8.76e-06 
+ nrs=0.91 nrd=1.06 
m734 405 404 403 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m735 1 140 403 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m736 0 140 405 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m737 406 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m738 407 408 406 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m739 407 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m740 1 407 408 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m741 0 407 408 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m742 0 140 130 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=7.13e-12 ps=8.76e-06 pd=1.451e-05 
+ nrs=1.06 nrd=0.91 
m743 409 129 407 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m744 129 148 130 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m745 129 150 130 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m746 0 185 409 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m747 1 140 129 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m748 410 116 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m749 411 185 410 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m750 1 140 116 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m751 412 411 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m752 412 411 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m753 115 149 116 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m754 115 151 116 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m755 115 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.13e-12 ad=8.33e-12 ps=1.451e-05 pd=8.76e-06 
+ nrs=0.91 nrd=1.06 
m756 413 412 411 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m757 0 140 413 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m758 1 140 411 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m759 414 415 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m760 416 140 414 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m761 1 416 415 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m762 0 416 415 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m763 416 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m764 117 149 118 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m765 417 117 416 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m766 0 140 118 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=7.13e-12 ps=8.76e-06 pd=1.451e-05 
+ nrs=1.06 nrd=0.91 
m767 0 185 417 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m768 117 150 118 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m769 1 140 117 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m770 120 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m771 418 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m772 419 120 418 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m773 420 419 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m774 420 419 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m775 119 151 120 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.81e-12 ad=6.21e-12 ps=8.5e-06 pd=1.213e-05 
+ nrs=1.09 nrd=1.41 
m776 119 148 120 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.81e-12 ad=6.21e-12 ps=8.5e-06 pd=1.213e-05 
+ nrs=1.09 nrd=1.41 
m777 119 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.41e-12 ad=8.33e-12 ps=1.133e-05 pd=8.76e-06 
+ nrs=0.82 nrd=1.06 
m778 421 420 419 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m779 1 140 419 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m780 0 140 421 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m781 422 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m782 423 424 422 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m783 423 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m784 1 423 424 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m785 0 423 424 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m786 0 140 122 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=7.13e-12 ps=8.76e-06 pd=1.451e-05 
+ nrs=1.06 nrd=0.91 
m787 425 121 423 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m788 121 148 122 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m789 121 150 122 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m790 0 185 425 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m791 1 140 121 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m792 426 108 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m793 427 185 426 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m794 1 140 108 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m795 428 427 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m796 428 427 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m797 107 149 108 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m798 107 151 108 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m799 107 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.13e-12 ad=8.33e-12 ps=1.451e-05 pd=8.76e-06 
+ nrs=0.91 nrd=1.06 
m800 429 428 427 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m801 0 140 429 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m802 1 140 427 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m803 430 431 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m804 432 140 430 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m805 1 432 431 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m806 0 432 431 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m807 432 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m808 109 149 110 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.155e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m809 433 109 432 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m810 0 140 110 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=7.13e-12 ps=8.76e-06 pd=1.451e-05 
+ nrs=1.06 nrd=0.91 
m811 0 185 433 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m812 109 150 110 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.155e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m813 1 140 109 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m814 112 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m815 434 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m816 435 112 434 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m817 436 435 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m818 436 435 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m819 111 151 112 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m820 111 148 112 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m821 111 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.13e-12 ad=8.33e-12 ps=1.451e-05 pd=8.76e-06 
+ nrs=0.91 nrd=1.06 
m822 437 436 435 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m823 1 140 435 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m824 0 140 437 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m825 438 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m826 439 440 438 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m827 439 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m828 1 439 440 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m829 0 439 440 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m830 0 140 114 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=7.13e-12 ps=8.76e-06 pd=1.451e-05 
+ nrs=1.06 nrd=0.91 
m831 441 113 439 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m832 113 148 114 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m833 113 150 114 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m834 0 185 441 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m835 1 140 113 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m836 442 100 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m837 443 185 442 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m838 1 140 100 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m839 444 443 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m840 444 443 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m841 99 149 100 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m842 99 151 100 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m843 99 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.91e-12 ad=8.33e-12 ps=1.807e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m844 445 444 443 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m845 0 140 445 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m846 1 140 443 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m847 446 447 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m848 448 140 446 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m849 1 448 447 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m850 0 448 447 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m851 448 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m852 101 149 102 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m853 449 101 448 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m854 0 140 102 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.91e-12 ps=8.76e-06 pd=1.807e-05 
+ nrs=1.06 nrd=1.14 
m855 0 185 449 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m856 101 150 102 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m857 1 140 101 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m858 104 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m859 450 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m860 451 104 450 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m861 452 451 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m862 452 451 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m863 103 151 104 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m864 103 148 104 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m865 103 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.06e-12 ad=8.33e-12 ps=1.247e-05 pd=8.76e-06 
+ nrs=0.77 nrd=1.06 
m866 453 452 451 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m867 1 140 451 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m868 0 140 453 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m869 454 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m870 455 456 454 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m871 455 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m872 1 455 456 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m873 0 455 456 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m874 0 140 106 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=6.06e-12 ps=8.76e-06 pd=1.247e-05 
+ nrs=1.06 nrd=0.77 
m875 457 105 455 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m876 105 148 106 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m877 105 150 106 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m878 0 185 457 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m879 1 140 105 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m880 458 92 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m881 459 185 458 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m882 1 140 92 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m883 460 459 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m884 460 459 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m885 91 149 92 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m886 91 151 92 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m887 91 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.91e-12 ad=8.33e-12 ps=1.807e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m888 461 460 459 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m889 0 140 461 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m890 1 140 459 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m891 462 463 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m892 464 140 462 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m893 1 464 463 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m894 0 464 463 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m895 464 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m896 93 149 94 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m897 465 93 464 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m898 0 140 94 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=6.06e-12 ps=8.76e-06 pd=1.247e-05 
+ nrs=1.06 nrd=0.77 
m899 0 185 465 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m900 93 150 94 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m901 1 140 93 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m902 96 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m903 466 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m904 467 96 466 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m905 468 467 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m906 468 467 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m907 95 151 96 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m908 95 148 96 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m909 95 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.06e-12 ad=8.33e-12 ps=1.247e-05 pd=8.76e-06 
+ nrs=0.77 nrd=1.06 
m910 469 468 467 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m911 1 140 467 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m912 0 140 469 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m913 470 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m914 471 472 470 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m915 471 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m916 1 471 472 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m917 0 471 472 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m918 0 140 98 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=6.06e-12 ps=8.76e-06 pd=1.247e-05 
+ nrs=1.06 nrd=0.77 
m919 473 97 471 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m920 97 148 98 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m921 97 150 98 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m922 0 185 473 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m923 1 140 97 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m924 474 84 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m925 475 185 474 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m926 1 140 84 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m927 476 475 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m928 476 475 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m929 83 149 84 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m930 83 151 84 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m931 83 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.06e-12 ad=8.33e-12 ps=1.247e-05 pd=8.76e-06 
+ nrs=0.77 nrd=1.06 
m932 477 476 475 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m933 0 140 477 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m934 1 140 475 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m935 478 479 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m936 480 140 478 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m937 1 480 479 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m938 0 480 479 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m939 480 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m940 85 149 86 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m941 481 85 480 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m942 0 140 86 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=6.06e-12 ps=8.76e-06 pd=1.247e-05 
+ nrs=1.06 nrd=0.77 
m943 0 185 481 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m944 85 150 86 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m945 1 140 85 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m946 88 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m947 482 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m948 483 88 482 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m949 484 483 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m950 484 483 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m951 87 151 88 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m952 87 148 88 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m953 87 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.06e-12 ad=8.33e-12 ps=1.247e-05 pd=8.76e-06 
+ nrs=0.77 nrd=1.06 
m954 485 484 483 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m955 1 140 483 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m956 0 140 485 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m957 486 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m958 487 488 486 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m959 487 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m960 1 487 488 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m961 0 487 488 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m962 0 140 90 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=6.06e-12 ps=8.76e-06 pd=1.247e-05 
+ nrs=1.06 nrd=0.77 
m963 489 89 487 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m964 89 148 90 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.72e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.3 nrd=1.03 
m965 89 150 90 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.72e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.3 nrd=1.03 
m966 0 185 489 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m967 1 140 89 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m968 490 75 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m969 491 185 490 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m970 1 140 75 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=1.078e-11 ps=3.179e-05 pd=3.36e-05 
+ nrs=0.52 nrd=0.18 
m971 492 491 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m972 492 491 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m973 74 149 75 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m974 74 151 75 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m975 74 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.91e-12 ad=8.33e-12 ps=1.807e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m976 493 492 491 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m977 0 140 493 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m978 1 140 491 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m979 494 495 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m980 496 140 494 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m981 1 496 495 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m982 0 496 495 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m983 496 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m984 77 149 78 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m985 497 77 496 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m986 0 140 78 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=6.06e-12 ps=8.76e-06 pd=1.247e-05 
+ nrs=1.06 nrd=0.77 
m987 0 185 497 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m988 77 150 78 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m989 1 140 77 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m990 80 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m991 498 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m992 499 80 498 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m993 500 499 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m994 500 499 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m995 79 151 80 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=8.98e-06 
+ nrs=1.03 nrd=1.19 
m996 79 148 80 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=8.98e-06 
+ nrs=1.03 nrd=1.19 
m997 79 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.06e-12 ad=8.33e-12 ps=1.247e-05 pd=8.76e-06 
+ nrs=0.77 nrd=1.06 
m998 501 500 499 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m999 1 140 499 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1000 0 140 501 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1001 502 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1002 503 504 502 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1003 503 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m1004 1 503 504 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1005 0 503 504 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1006 0 140 82 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=6.06e-12 ps=8.76e-06 pd=1.247e-05 
+ nrs=1.06 nrd=0.77 
m1007 505 81 503 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1008 81 148 82 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m1009 81 150 82 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m1010 0 185 505 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1011 1 140 81 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m1012 506 67 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1013 507 185 506 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1014 1 140 67 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m1015 508 507 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1016 508 507 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1017 66 149 67 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m1018 66 151 67 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m1019 66 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.13e-12 ad=8.33e-12 ps=1.451e-05 pd=8.76e-06 
+ nrs=0.91 nrd=1.06 
m1020 509 508 507 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1021 0 140 509 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1022 1 140 507 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1023 510 511 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1024 512 140 510 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1025 1 512 511 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1026 0 512 511 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1027 512 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m1028 68 149 69 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=4.28e-12 ps=1.213e-05 pd=9.16e-06 
+ nrs=1.41 nrd=0.97 
m1029 513 68 512 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1030 0 140 69 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=5.7e-12 ps=8.76e-06 pd=1.222e-05 
+ nrs=1.06 nrd=0.73 
m1031 0 185 513 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1032 68 150 69 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=4.28e-12 ps=1.213e-05 pd=9.16e-06 
+ nrs=1.41 nrd=0.97 
m1033 1 140 68 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m1034 71 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m1035 514 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1036 515 71 514 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1037 516 515 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1038 516 515 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1039 70 151 71 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m1040 70 148 71 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m1041 70 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.13e-12 ad=8.33e-12 ps=1.451e-05 pd=8.76e-06 
+ nrs=0.91 nrd=1.06 
m1042 517 516 515 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1043 1 140 515 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1044 0 140 517 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1045 518 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1046 519 520 518 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1047 519 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m1048 1 519 520 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1049 0 519 520 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1050 0 140 73 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=7.13e-12 ps=8.76e-06 pd=1.451e-05 
+ nrs=1.06 nrd=0.91 
m1051 521 72 519 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1052 72 148 73 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m1053 72 150 73 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m1054 0 185 521 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1055 1 140 72 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m1056 522 59 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1057 523 185 522 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1058 1 140 59 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m1059 524 523 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1060 524 523 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1061 58 149 59 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=2.94e-12 ps=1.088e-05 pd=6.18e-06 
+ nrs=1.21 nrd=0.67 
m1062 58 151 59 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=2.94e-12 ps=1.088e-05 pd=6.18e-06 
+ nrs=1.21 nrd=0.67 
m1063 58 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.13e-12 ad=8.33e-12 ps=1.451e-05 pd=8.76e-06 
+ nrs=0.91 nrd=1.06 
m1064 525 524 523 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1065 0 140 525 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1066 1 140 523 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1067 526 527 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1068 528 140 526 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1069 1 528 527 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1070 0 528 527 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1071 528 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m1072 60 149 61 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m1073 529 60 528 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1074 0 140 61 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=7.13e-12 ps=8.76e-06 pd=1.451e-05 
+ nrs=1.06 nrd=0.91 
m1075 0 185 529 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1076 60 150 61 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m1077 1 140 60 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m1078 63 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m1079 530 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1080 531 63 530 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1081 532 531 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1082 532 531 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1083 62 151 63 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m1084 62 148 63 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m1085 62 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.13e-12 ad=8.33e-12 ps=1.451e-05 pd=8.76e-06 
+ nrs=0.91 nrd=1.06 
m1086 533 532 531 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1087 1 140 531 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1088 0 140 533 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1089 534 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1090 535 536 534 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1091 535 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m1092 1 535 536 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1093 0 535 536 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1094 0 140 65 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=7.13e-12 ps=8.76e-06 pd=1.451e-05 
+ nrs=1.06 nrd=0.91 
m1095 537 64 535 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1096 64 148 65 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m1097 64 150 65 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m1098 0 185 537 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1099 1 140 64 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m1100 538 51 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1101 539 185 538 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1102 1 140 51 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m1103 540 539 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1104 540 539 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1105 50 149 51 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m1106 50 151 51 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m1107 50 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.13e-12 ad=8.33e-12 ps=1.451e-05 pd=8.76e-06 
+ nrs=0.91 nrd=1.06 
m1108 541 540 539 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1109 0 140 541 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1110 1 140 539 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1111 542 543 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1112 544 140 542 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1113 1 544 543 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1114 0 544 543 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1115 544 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m1116 52 149 53 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m1117 545 52 544 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1118 0 140 53 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=7.13e-12 ps=8.76e-06 pd=1.451e-05 
+ nrs=1.06 nrd=0.91 
m1119 0 185 545 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1120 52 150 53 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m1121 1 140 52 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m1122 55 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m1123 546 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1124 547 55 546 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1125 548 547 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1126 548 547 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1127 54 151 55 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m1128 54 148 55 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m1129 54 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.13e-12 ad=8.33e-12 ps=1.451e-05 pd=8.76e-06 
+ nrs=0.91 nrd=1.06 
m1130 549 548 547 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1131 1 140 547 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1132 0 140 549 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1133 550 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1134 551 552 550 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1135 551 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m1136 1 551 552 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1137 0 551 552 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1138 0 140 57 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=7.13e-12 ps=8.76e-06 pd=1.451e-05 
+ nrs=1.06 nrd=0.91 
m1139 553 56 551 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1140 56 148 57 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m1141 56 150 57 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=5.35e-12 ps=1.167e-05 pd=1.088e-05 
+ nrs=1.37 nrd=1.21 
m1142 0 185 553 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1143 1 140 56 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m1144 554 42 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1145 555 185 554 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1146 1 140 42 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m1147 556 555 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1148 556 555 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1149 41 149 42 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.21e-12 ad=6.21e-12 ps=1.031e-05 pd=1.213e-05 
+ nrs=1.18 nrd=1.41 
m1150 41 151 42 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.21e-12 ad=6.21e-12 ps=1.031e-05 pd=1.213e-05 
+ nrs=1.18 nrd=1.41 
m1151 41 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.95e-12 ad=8.33e-12 ps=1.375e-05 pd=8.76e-06 
+ nrs=0.89 nrd=1.06 
m1152 557 556 555 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1153 0 140 557 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1154 1 140 555 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1155 558 559 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1156 560 140 558 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1157 1 560 559 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1158 0 560 559 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1159 560 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m1160 44 149 45 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m1161 561 44 560 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1162 0 140 45 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=7.13e-12 ps=8.76e-06 pd=1.451e-05 
+ nrs=1.06 nrd=0.91 
m1163 0 185 561 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1164 44 150 45 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.21e-12 ad=5.35e-12 ps=1.213e-05 pd=1.088e-05 
+ nrs=1.41 nrd=1.21 
m1165 1 140 44 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m1166 47 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m1167 562 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1168 563 47 562 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1169 564 563 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1170 564 563 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1171 46 151 47 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m1172 46 148 47 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.35e-12 ad=6.21e-12 ps=1.088e-05 pd=1.213e-05 
+ nrs=1.21 nrd=1.41 
m1173 46 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=7.13e-12 ad=8.33e-12 ps=1.451e-05 pd=8.76e-06 
+ nrs=0.91 nrd=1.06 
m1174 565 564 563 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1175 1 140 563 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1176 0 140 565 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1177 566 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1178 567 568 566 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1179 567 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m1180 1 567 568 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1181 0 567 568 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1182 0 140 49 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=5.17e-12 ps=8.76e-06 pd=1.133e-05 
+ nrs=1.06 nrd=0.66 
m1183 569 48 567 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1184 48 148 49 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=3.88e-12 ps=1.167e-05 pd=8.5e-06 
+ nrs=1.37 nrd=0.88 
m1185 48 150 49 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.04e-12 ad=3.88e-12 ps=1.167e-05 pd=8.5e-06 
+ nrs=1.37 nrd=0.88 
m1186 0 185 569 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1187 1 140 48 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m1188 570 34 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1189 571 185 570 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1190 1 140 34 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m1191 572 571 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1192 572 571 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1193 33 149 34 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m1194 33 151 34 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m1195 33 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.91e-12 ad=8.33e-12 ps=1.807e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1196 573 572 571 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1197 0 140 573 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1198 1 140 571 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1199 574 575 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1200 576 140 574 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1201 1 576 575 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1202 0 576 575 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1203 576 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m1204 35 149 36 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m1205 577 35 576 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1206 0 140 36 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.91e-12 ps=8.76e-06 pd=1.807e-05 
+ nrs=1.06 nrd=1.14 
m1207 0 185 577 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1208 35 150 36 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m1209 1 140 35 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m1210 38 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m1211 578 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1212 579 38 578 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1213 580 579 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1214 580 579 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1215 37 151 38 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m1216 37 148 38 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m1217 37 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.06e-12 ad=8.33e-12 ps=1.247e-05 pd=8.76e-06 
+ nrs=0.77 nrd=1.06 
m1218 581 580 579 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1219 1 140 579 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1220 0 140 581 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1221 582 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1222 583 584 582 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1223 583 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m1224 1 583 584 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1225 0 583 584 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1226 0 140 40 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=6.06e-12 ps=8.76e-06 pd=1.247e-05 
+ nrs=1.06 nrd=0.77 
m1227 585 39 583 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1228 39 148 40 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m1229 39 150 40 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m1230 0 185 585 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1231 1 140 39 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m1232 586 25 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1233 587 185 586 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1234 1 140 25 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m1235 588 587 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1236 588 587 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1237 24 149 25 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m1238 24 151 25 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m1239 24 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.91e-12 ad=8.33e-12 ps=1.807e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1240 589 588 587 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1241 0 140 589 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1242 1 140 587 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1243 590 591 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1244 592 140 590 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1245 1 592 591 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1246 0 592 591 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1247 592 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m1248 27 149 28 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m1249 593 27 592 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1250 0 140 28 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.91e-12 ps=8.76e-06 pd=1.807e-05 
+ nrs=1.06 nrd=1.14 
m1251 0 185 593 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1252 27 150 28 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=6.68e-12 ps=1.54e-05 pd=1.355e-05 
+ nrs=1.78 nrd=1.52 
m1253 1 140 27 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m1254 30 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m1255 594 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1256 595 30 594 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1257 596 595 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1258 596 595 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1259 29 151 30 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m1260 29 148 30 0 nenh l=1.1e-06 w=2.1e-06 
+ as=4.54e-12 ad=5.23e-12 ps=9.35e-06 pd=1.027e-05 
+ nrs=1.03 nrd=1.19 
m1261 29 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=6.06e-12 ad=8.33e-12 ps=1.247e-05 pd=8.76e-06 
+ nrs=0.77 nrd=1.06 
m1262 597 596 595 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1263 1 140 595 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1264 0 140 597 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1265 598 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1266 599 600 598 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1267 599 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m1268 1 599 600 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1269 0 599 600 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1270 0 140 32 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=6.06e-12 ps=8.76e-06 pd=1.247e-05 
+ nrs=1.06 nrd=0.77 
m1271 601 31 599 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1272 31 148 32 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.68e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m1273 31 150 32 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.68e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m1274 0 185 601 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1275 1 140 31 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m1276 602 16 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1277 603 185 602 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1278 1 140 16 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=1.078e-11 ps=3.179e-05 pd=3.36e-05 
+ nrs=0.52 nrd=0.18 
m1279 604 603 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1280 604 603 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1281 15 149 16 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m1282 15 151 16 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m1283 15 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.91e-12 ad=8.33e-12 ps=1.807e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1284 605 604 603 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1285 0 140 605 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1286 1 140 603 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1287 606 607 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1288 608 140 606 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1289 1 608 607 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1290 0 608 607 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1291 608 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=6.86e-12 ad=2.796e-11 ps=2.1e-05 pd=2.89e-05 
+ nrs=0.14 nrd=0.57 
m1292 18 149 19 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m1293 609 18 608 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1294 0 140 19 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=6.06e-12 ps=8.76e-06 pd=1.247e-05 
+ nrs=1.06 nrd=0.77 
m1295 0 185 609 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1296 18 150 19 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.23e-12 ad=4.54e-12 ps=1.027e-05 pd=9.35e-06 
+ nrs=1.19 nrd=1.03 
m1297 1 140 18 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=7.35e-12 ps=3.179e-05 pd=2.24e-05 
+ nrs=0.52 nrd=0.12 
m1298 21 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m1299 610 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1300 611 21 610 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1301 612 611 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1302 612 611 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1303 20 151 21 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.15e-12 ad=5.23e-12 ps=1.145e-05 pd=1.027e-05 
+ nrs=1.39 nrd=1.19 
m1304 20 148 21 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.15e-12 ad=5.23e-12 ps=1.145e-05 pd=1.027e-05 
+ nrs=1.39 nrd=1.19 
m1305 20 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.2e-12 ad=8.33e-12 ps=1.527e-05 pd=8.76e-06 
+ nrs=1.05 nrd=1.06 
m1306 613 612 611 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1307 1 140 611 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1308 0 140 613 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1309 614 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1310 615 616 614 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1311 615 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m1312 1 615 616 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1313 0 615 616 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1314 0 140 23 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=6.06e-12 ps=8.76e-06 pd=1.247e-05 
+ nrs=1.06 nrd=0.77 
m1315 617 22 615 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1316 22 148 23 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m1317 22 150 23 0 nenh l=1.1e-06 w=2.1e-06 
+ as=5.06e-12 ad=4.54e-12 ps=9.8e-06 pd=9.35e-06 
+ nrs=1.15 nrd=1.03 
m1318 0 185 617 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1319 1 140 22 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=5.39e-12 ps=3.179e-05 pd=1.68e-05 
+ nrs=0.52 nrd=0.09 
m1320 618 4 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1321 1 140 4 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=1.078e-11 ps=3.179e-05 pd=3.36e-05 
+ nrs=0.52 nrd=0.18 
m1322 619 185 618 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1323 620 619 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1324 620 619 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1325 3 149 4 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m1326 3 151 4 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=7.84e-12 ps=1.355e-05 pd=1.54e-05 
+ nrs=1.52 nrd=1.78 
m1327 621 620 619 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1328 3 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.91e-12 ad=8.33e-12 ps=1.807e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1329 1 140 619 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1330 0 140 621 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1331 622 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1332 623 624 622 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1333 1 623 624 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1334 0 623 624 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1335 623 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m1336 9 149 10 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=4.54e-12 ps=1.54e-05 pd=9.35e-06 
+ nrs=1.78 nrd=1.03 
m1337 625 9 623 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1338 0 140 10 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=6.06e-12 ps=8.76e-06 pd=1.247e-05 
+ nrs=1.06 nrd=0.77 
m1339 0 185 625 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1340 9 150 10 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.84e-12 ad=4.54e-12 ps=1.54e-05 pd=9.35e-06 
+ nrs=1.78 nrd=1.03 
m1341 1 140 9 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=1.078e-11 ps=3.179e-05 pd=3.36e-05 
+ nrs=0.52 nrd=0.18 
m1342 12 140 1 1 penh l=1.1e-06 w=7.7e-06 
+ as=7.35e-12 ad=3.076e-11 ps=2.24e-05 pd=3.179e-05 
+ nrs=0.12 nrd=0.52 
m1343 626 185 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1344 627 12 626 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1345 628 627 1 1 penh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=2.237e-11 ps=1.26e-05 pd=2.312e-05 
+ nrs=0.12 nrd=0.71 
m1346 628 627 0 0 nenh l=1.1e-06 w=5.6e-06 
+ as=3.92e-12 ad=1.667e-11 ps=1.26e-05 pd=1.753e-05 
+ nrs=0.12 nrd=0.53 
m1347 11 151 12 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=5.23e-12 ps=1.355e-05 pd=1.027e-05 
+ nrs=1.52 nrd=1.19 
m1348 11 148 12 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.68e-12 ad=5.23e-12 ps=1.355e-05 pd=1.027e-05 
+ nrs=1.52 nrd=1.19 
m1349 1 140 627 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=4.9e-12 ps=2.89e-05 pd=1.54e-05 
+ nrs=0.57 nrd=0.1 
m1350 11 140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.91e-12 ad=8.33e-12 ps=1.807e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1351 629 628 627 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1352 0 140 629 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1353 630 140 0 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=6.25e-12 ps=3.5e-06 pd=6.57e-06 
+ nrs=0.33 nrd=1.42 
m1354 631 632 630 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=5.6e-06 pd=3.5e-06 
+ nrs=0.33 nrd=0.33 
m1355 1 631 632 1 penh l=1.1e-06 w=5.6e-06 
+ as=2.237e-11 ad=3.92e-12 ps=2.312e-05 pd=1.26e-05 
+ nrs=0.71 nrd=0.12 
m1356 0 631 632 0 nenh l=1.1e-06 w=5.6e-06 
+ as=1.667e-11 ad=3.92e-12 ps=1.753e-05 pd=1.26e-05 
+ nrs=0.53 nrd=0.12 
m1357 631 140 1 1 penh l=1.1e-06 w=7e-06 
+ as=4.9e-12 ad=2.796e-11 ps=1.54e-05 pd=2.89e-05 
+ nrs=0.1 nrd=0.57 
m1358 0 140 14 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=6.06e-12 ps=8.76e-06 pd=1.247e-05 
+ nrs=1.06 nrd=0.77 
m1359 13 148 14 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.68e-12 ad=4.54e-12 ps=1.493e-05 pd=9.35e-06 
+ nrs=1.74 nrd=1.03 
m1360 633 13 631 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.47e-12 ad=1.47e-12 ps=3.5e-06 pd=5.6e-06 
+ nrs=0.33 nrd=0.33 
m1361 13 150 14 0 nenh l=1.1e-06 w=2.1e-06 
+ as=7.68e-12 ad=4.54e-12 ps=1.493e-05 pd=9.35e-06 
+ nrs=1.74 nrd=1.03 
m1362 0 185 633 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.25e-12 ad=1.47e-12 ps=6.57e-06 pd=3.5e-06 
+ nrs=1.42 nrd=0.33 
m1363 1 140 13 1 penh l=1.1e-06 w=7.7e-06 
+ as=3.076e-11 ad=1.078e-11 ps=3.179e-05 pd=3.36e-05 
+ nrs=0.52 nrd=0.18 
m1364 1 635 634 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1365 635 634 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m1366 1 637 636 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1367 637 636 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1368 1 639 638 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1369 639 638 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1370 1 641 640 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m1371 641 640 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1372 0 635 634 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1373 635 634 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1374 0 637 636 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1375 637 636 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1376 0 639 638 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1377 639 638 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1378 0 641 640 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1379 641 640 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1380 196 380 634 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m1381 197 380 635 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1382 198 380 636 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1383 199 380 637 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1384 200 380 638 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1385 201 380 639 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1386 202 380 640 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1387 203 380 641 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m1388 642 383 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m1389 643 383 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1390 644 383 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1391 645 383 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1392 646 383 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1393 647 383 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1394 648 383 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1395 649 383 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m1396 0 643 642 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1397 643 642 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1398 0 645 644 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1399 645 644 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1400 0 647 646 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1401 647 646 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1402 0 649 648 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1403 649 648 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1404 1 643 642 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1405 643 642 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1406 1 645 644 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1407 645 644 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1408 1 651 650 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1409 651 650 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m1410 1 653 652 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1411 653 652 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1412 1 647 646 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1413 647 646 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1414 1 649 648 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1415 649 648 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1416 1 655 654 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1417 655 654 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1418 1 657 656 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m1419 657 656 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1420 0 651 650 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1421 651 650 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1422 0 653 652 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1423 653 652 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1424 0 655 654 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1425 655 654 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1426 0 657 656 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1427 657 656 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1428 196 388 650 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m1429 197 388 651 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1430 198 388 652 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1431 199 388 653 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1432 200 388 654 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1433 201 388 655 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1434 202 388 656 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1435 203 388 657 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m1436 658 392 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m1437 659 392 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1438 660 392 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1439 661 392 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1440 662 392 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1441 663 392 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1442 664 392 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1443 665 392 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m1444 0 659 658 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1445 659 658 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1446 0 661 660 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1447 661 660 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1448 0 663 662 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1449 663 662 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1450 0 665 664 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1451 665 664 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1452 1 659 658 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1453 659 658 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1454 1 661 660 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1455 661 660 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1456 1 663 662 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1457 663 662 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1458 1 665 664 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1459 665 664 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1460 1 667 666 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1461 667 666 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m1462 1 669 668 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1463 669 668 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1464 1 671 670 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1465 671 670 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1466 1 673 672 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m1467 673 672 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1468 0 667 666 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1469 667 666 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1470 0 669 668 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1471 669 668 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1472 0 671 670 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1473 671 670 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1474 0 673 672 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1475 673 672 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1476 196 396 666 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m1477 197 396 667 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1478 198 396 668 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1479 199 396 669 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1480 200 396 670 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1481 201 396 671 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1482 202 396 672 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1483 203 396 673 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m1484 674 399 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m1485 675 399 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1486 676 399 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1487 677 399 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1488 678 399 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1489 679 399 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1490 680 399 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1491 681 399 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m1492 0 675 674 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1493 675 674 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1494 0 677 676 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1495 677 676 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1496 0 679 678 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1497 679 678 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1498 0 681 680 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1499 681 680 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1500 1 675 674 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1501 675 674 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1502 1 677 676 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1503 677 676 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1504 1 683 682 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1505 683 682 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m1506 1 685 684 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1507 685 684 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1508 1 679 678 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1509 679 678 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1510 1 681 680 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1511 681 680 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1512 1 687 686 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1513 687 686 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1514 1 689 688 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m1515 689 688 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1516 0 683 682 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1517 683 682 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1518 0 685 684 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1519 685 684 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1520 0 687 686 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1521 687 686 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1522 0 689 688 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1523 689 688 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1524 196 404 682 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m1525 197 404 683 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1526 198 404 684 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1527 199 404 685 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1528 200 404 686 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1529 201 404 687 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1530 202 404 688 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1531 203 404 689 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m1532 690 408 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m1533 691 408 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1534 692 408 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1535 693 408 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1536 694 408 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1537 695 408 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1538 696 408 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1539 697 408 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m1540 0 691 690 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1541 691 690 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1542 0 693 692 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1543 693 692 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1544 0 695 694 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1545 695 694 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1546 0 697 696 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1547 697 696 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1548 1 691 690 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1549 691 690 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1550 1 693 692 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1551 693 692 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1552 1 695 694 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1553 695 694 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1554 1 697 696 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1555 697 696 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1556 1 699 698 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1557 699 698 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m1558 1 701 700 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1559 701 700 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1560 1 703 702 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1561 703 702 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1562 1 705 704 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m1563 705 704 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1564 0 699 698 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1565 699 698 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1566 0 701 700 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1567 701 700 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1568 0 703 702 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1569 703 702 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1570 0 705 704 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1571 705 704 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1572 196 412 698 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m1573 197 412 699 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1574 198 412 700 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1575 199 412 701 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1576 200 412 702 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1577 201 412 703 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1578 202 412 704 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1579 203 412 705 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m1580 706 415 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m1581 707 415 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1582 708 415 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1583 709 415 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1584 710 415 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1585 711 415 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1586 712 415 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1587 713 415 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m1588 0 707 706 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1589 707 706 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1590 0 709 708 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1591 709 708 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1592 0 711 710 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1593 711 710 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1594 0 713 712 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1595 713 712 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1596 1 707 706 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1597 707 706 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1598 1 709 708 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1599 709 708 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1600 1 715 714 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1601 715 714 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m1602 1 717 716 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1603 717 716 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1604 1 711 710 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1605 711 710 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1606 1 713 712 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1607 713 712 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1608 1 719 718 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1609 719 718 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1610 1 721 720 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m1611 721 720 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1612 0 715 714 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1613 715 714 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1614 0 717 716 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1615 717 716 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1616 0 719 718 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1617 719 718 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1618 0 721 720 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1619 721 720 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1620 196 420 714 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m1621 197 420 715 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1622 198 420 716 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1623 199 420 717 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1624 200 420 718 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1625 201 420 719 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1626 202 420 720 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1627 203 420 721 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m1628 722 424 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m1629 723 424 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1630 724 424 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1631 725 424 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1632 726 424 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1633 727 424 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1634 728 424 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1635 729 424 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m1636 0 723 722 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1637 723 722 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1638 0 725 724 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1639 725 724 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1640 0 727 726 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1641 727 726 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1642 0 729 728 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1643 729 728 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1644 1 723 722 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1645 723 722 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1646 1 725 724 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1647 725 724 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1648 1 727 726 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1649 727 726 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1650 1 729 728 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1651 729 728 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1652 1 731 730 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1653 731 730 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m1654 1 733 732 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1655 733 732 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1656 1 735 734 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1657 735 734 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1658 1 737 736 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m1659 737 736 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1660 0 731 730 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1661 731 730 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1662 0 733 732 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1663 733 732 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1664 0 735 734 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1665 735 734 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1666 0 737 736 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1667 737 736 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1668 196 428 730 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m1669 197 428 731 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1670 198 428 732 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1671 199 428 733 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1672 200 428 734 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1673 201 428 735 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1674 202 428 736 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1675 203 428 737 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m1676 738 431 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m1677 739 431 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1678 740 431 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1679 741 431 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1680 742 431 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1681 743 431 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1682 744 431 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1683 745 431 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m1684 0 739 738 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1685 739 738 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1686 0 741 740 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1687 741 740 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1688 0 743 742 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1689 743 742 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1690 0 745 744 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1691 745 744 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1692 1 739 738 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1693 739 738 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1694 1 741 740 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1695 741 740 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1696 1 747 746 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1697 747 746 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m1698 1 749 748 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1699 749 748 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1700 1 743 742 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1701 743 742 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1702 1 745 744 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1703 745 744 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1704 1 751 750 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1705 751 750 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1706 1 753 752 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m1707 753 752 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1708 0 747 746 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1709 747 746 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1710 0 749 748 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1711 749 748 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1712 0 751 750 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1713 751 750 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1714 0 753 752 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1715 753 752 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1716 196 436 746 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m1717 197 436 747 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1718 198 436 748 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1719 199 436 749 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1720 200 436 750 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1721 201 436 751 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1722 202 436 752 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1723 203 436 753 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m1724 754 440 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m1725 755 440 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1726 756 440 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1727 757 440 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1728 758 440 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1729 759 440 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1730 760 440 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1731 761 440 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m1732 0 755 754 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1733 755 754 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1734 0 757 756 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1735 757 756 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1736 0 759 758 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1737 759 758 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1738 0 761 760 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1739 761 760 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1740 1 755 754 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1741 755 754 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1742 1 757 756 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1743 757 756 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1744 1 759 758 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1745 759 758 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1746 1 761 760 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1747 761 760 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1748 1 763 762 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1749 763 762 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m1750 1 765 764 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1751 765 764 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1752 1 767 766 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1753 767 766 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1754 1 769 768 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m1755 769 768 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1756 0 763 762 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1757 763 762 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1758 0 765 764 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1759 765 764 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1760 0 767 766 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1761 767 766 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1762 0 769 768 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1763 769 768 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1764 196 444 762 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m1765 197 444 763 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1766 198 444 764 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1767 199 444 765 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1768 200 444 766 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1769 201 444 767 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1770 202 444 768 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1771 203 444 769 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m1772 770 447 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m1773 771 447 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1774 772 447 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1775 773 447 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1776 774 447 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1777 775 447 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1778 776 447 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1779 777 447 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m1780 0 771 770 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1781 771 770 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1782 0 773 772 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1783 773 772 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1784 0 775 774 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1785 775 774 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1786 0 777 776 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1787 777 776 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1788 1 771 770 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1789 771 770 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1790 1 773 772 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1791 773 772 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1792 1 779 778 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1793 779 778 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m1794 1 781 780 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1795 781 780 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1796 1 775 774 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1797 775 774 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1798 1 777 776 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1799 777 776 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1800 1 783 782 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1801 783 782 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1802 1 785 784 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m1803 785 784 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1804 0 779 778 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1805 779 778 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1806 0 781 780 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1807 781 780 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1808 0 783 782 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1809 783 782 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1810 0 785 784 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1811 785 784 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1812 196 452 778 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m1813 197 452 779 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1814 198 452 780 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1815 199 452 781 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1816 200 452 782 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1817 201 452 783 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1818 202 452 784 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1819 203 452 785 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m1820 786 456 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m1821 787 456 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1822 788 456 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1823 789 456 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1824 790 456 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1825 791 456 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1826 792 456 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1827 793 456 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m1828 0 787 786 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1829 787 786 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1830 0 789 788 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1831 789 788 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1832 0 791 790 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1833 791 790 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1834 0 793 792 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1835 793 792 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1836 1 787 786 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1837 787 786 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1838 1 789 788 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1839 789 788 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1840 1 791 790 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1841 791 790 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1842 1 793 792 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1843 793 792 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1844 1 795 794 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1845 795 794 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m1846 1 797 796 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1847 797 796 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1848 1 799 798 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1849 799 798 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1850 1 801 800 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m1851 801 800 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1852 0 795 794 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1853 795 794 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1854 0 797 796 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1855 797 796 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1856 0 799 798 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1857 799 798 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1858 0 801 800 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1859 801 800 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1860 196 460 794 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m1861 197 460 795 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1862 198 460 796 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1863 199 460 797 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1864 200 460 798 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1865 201 460 799 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1866 202 460 800 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1867 203 460 801 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m1868 802 463 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m1869 803 463 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1870 804 463 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1871 805 463 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1872 806 463 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1873 807 463 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1874 808 463 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1875 809 463 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m1876 0 803 802 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1877 803 802 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1878 0 805 804 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1879 805 804 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1880 0 807 806 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1881 807 806 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1882 0 809 808 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1883 809 808 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1884 1 803 802 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1885 803 802 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1886 1 805 804 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1887 805 804 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1888 1 811 810 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1889 811 810 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m1890 1 813 812 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1891 813 812 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1892 1 807 806 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1893 807 806 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1894 1 809 808 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1895 809 808 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1896 1 815 814 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1897 815 814 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1898 1 817 816 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m1899 817 816 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1900 0 811 810 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1901 811 810 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1902 0 813 812 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1903 813 812 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1904 0 815 814 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1905 815 814 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1906 0 817 816 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1907 817 816 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1908 196 468 810 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m1909 197 468 811 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1910 198 468 812 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1911 199 468 813 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1912 200 468 814 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1913 201 468 815 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1914 202 468 816 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1915 203 468 817 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m1916 818 472 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m1917 819 472 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1918 820 472 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1919 821 472 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1920 822 472 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1921 823 472 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1922 824 472 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1923 825 472 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m1924 0 819 818 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1925 819 818 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1926 0 821 820 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1927 821 820 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1928 0 823 822 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1929 823 822 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1930 0 825 824 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1931 825 824 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1932 1 819 818 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1933 819 818 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1934 1 821 820 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1935 821 820 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1936 1 823 822 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1937 823 822 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1938 1 825 824 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1939 825 824 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1940 1 827 826 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1941 827 826 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m1942 1 829 828 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1943 829 828 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1944 1 831 830 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1945 831 830 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1946 1 833 832 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m1947 833 832 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1948 0 827 826 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1949 827 826 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1950 0 829 828 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1951 829 828 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1952 0 831 830 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1953 831 830 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1954 0 833 832 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1955 833 832 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1956 196 476 826 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m1957 197 476 827 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1958 198 476 828 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1959 199 476 829 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1960 200 476 830 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m1961 201 476 831 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m1962 202 476 832 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m1963 203 476 833 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m1964 834 479 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m1965 835 479 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1966 836 479 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1967 837 479 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1968 838 479 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m1969 839 479 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m1970 840 479 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m1971 841 479 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m1972 0 835 834 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1973 835 834 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1974 0 837 836 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1975 837 836 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1976 0 839 838 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1977 839 838 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1978 0 841 840 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m1979 841 840 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m1980 1 835 834 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1981 835 834 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1982 1 837 836 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1983 837 836 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1984 1 843 842 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1985 843 842 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m1986 1 845 844 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1987 845 844 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1988 1 839 838 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1989 839 838 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1990 1 841 840 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1991 841 840 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1992 1 847 846 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m1993 847 846 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1994 1 849 848 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m1995 849 848 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m1996 0 843 842 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1997 843 842 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m1998 0 845 844 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m1999 845 844 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2000 0 847 846 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2001 847 846 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2002 0 849 848 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2003 849 848 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2004 196 484 842 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2005 197 484 843 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2006 198 484 844 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2007 199 484 845 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2008 200 484 846 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2009 201 484 847 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2010 202 484 848 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2011 203 484 849 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2012 850 488 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2013 851 488 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2014 852 488 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2015 853 488 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2016 854 488 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2017 855 488 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2018 856 488 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2019 857 488 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2020 0 851 850 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2021 851 850 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2022 0 853 852 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2023 853 852 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2024 0 855 854 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2025 855 854 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2026 0 857 856 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2027 857 856 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2028 1 851 850 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2029 851 850 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2030 1 853 852 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2031 853 852 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2032 1 855 854 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2033 855 854 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2034 1 857 856 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2035 857 856 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2036 1 859 858 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2037 859 858 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2038 1 861 860 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2039 861 860 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2040 1 863 862 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2041 863 862 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2042 1 865 864 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2043 865 864 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2044 0 859 858 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2045 859 858 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2046 0 861 860 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2047 861 860 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2048 0 863 862 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2049 863 862 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2050 0 865 864 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2051 865 864 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2052 196 492 858 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2053 197 492 859 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2054 198 492 860 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2055 199 492 861 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2056 200 492 862 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2057 201 492 863 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2058 202 492 864 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2059 203 492 865 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2060 866 495 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2061 867 495 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2062 868 495 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2063 869 495 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2064 870 495 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2065 871 495 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2066 872 495 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2067 873 495 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2068 0 867 866 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2069 867 866 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2070 0 869 868 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2071 869 868 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2072 0 871 870 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2073 871 870 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2074 0 873 872 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2075 873 872 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2076 1 867 866 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2077 867 866 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2078 1 869 868 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2079 869 868 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2080 1 875 874 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2081 875 874 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2082 1 877 876 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2083 877 876 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2084 1 871 870 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2085 871 870 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2086 1 873 872 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2087 873 872 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2088 1 879 878 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2089 879 878 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2090 1 881 880 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2091 881 880 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2092 0 875 874 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2093 875 874 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2094 0 877 876 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2095 877 876 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2096 0 879 878 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2097 879 878 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2098 0 881 880 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2099 881 880 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2100 196 500 874 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2101 197 500 875 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2102 198 500 876 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2103 199 500 877 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2104 200 500 878 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2105 201 500 879 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2106 202 500 880 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2107 203 500 881 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2108 882 504 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2109 883 504 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2110 884 504 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2111 885 504 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2112 886 504 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2113 887 504 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2114 888 504 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2115 889 504 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2116 0 883 882 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2117 883 882 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2118 0 885 884 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2119 885 884 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2120 0 887 886 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2121 887 886 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2122 0 889 888 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2123 889 888 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2124 1 883 882 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2125 883 882 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2126 1 885 884 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2127 885 884 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2128 1 887 886 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2129 887 886 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2130 1 889 888 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2131 889 888 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2132 1 891 890 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2133 891 890 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2134 1 893 892 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2135 893 892 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2136 1 895 894 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2137 895 894 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2138 1 897 896 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2139 897 896 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2140 0 891 890 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2141 891 890 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2142 0 893 892 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2143 893 892 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2144 0 895 894 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2145 895 894 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2146 0 897 896 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2147 897 896 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2148 196 508 890 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2149 197 508 891 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2150 198 508 892 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2151 199 508 893 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2152 200 508 894 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2153 201 508 895 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2154 202 508 896 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2155 203 508 897 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2156 898 511 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2157 899 511 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2158 900 511 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2159 901 511 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2160 902 511 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2161 903 511 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2162 904 511 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2163 905 511 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2164 0 899 898 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2165 899 898 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2166 0 901 900 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2167 901 900 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2168 0 903 902 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2169 903 902 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2170 0 905 904 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2171 905 904 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2172 1 899 898 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2173 899 898 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2174 1 901 900 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2175 901 900 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2176 1 907 906 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2177 907 906 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2178 1 909 908 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2179 909 908 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2180 1 903 902 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2181 903 902 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2182 1 905 904 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2183 905 904 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2184 1 911 910 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2185 911 910 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2186 1 913 912 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2187 913 912 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2188 0 907 906 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2189 907 906 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2190 0 909 908 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2191 909 908 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2192 0 911 910 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2193 911 910 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2194 0 913 912 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2195 913 912 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2196 196 516 906 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2197 197 516 907 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2198 198 516 908 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2199 199 516 909 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2200 200 516 910 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2201 201 516 911 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2202 202 516 912 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2203 203 516 913 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2204 914 520 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2205 915 520 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2206 916 520 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2207 917 520 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2208 918 520 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2209 919 520 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2210 920 520 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2211 921 520 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2212 0 915 914 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2213 915 914 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2214 0 917 916 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2215 917 916 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2216 0 919 918 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2217 919 918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2218 0 921 920 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2219 921 920 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2220 1 915 914 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2221 915 914 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2222 1 917 916 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2223 917 916 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2224 1 919 918 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2225 919 918 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2226 1 921 920 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2227 921 920 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2228 1 923 922 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2229 923 922 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2230 1 925 924 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2231 925 924 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2232 1 927 926 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2233 927 926 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2234 1 929 928 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2235 929 928 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2236 0 923 922 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2237 923 922 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2238 0 925 924 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2239 925 924 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2240 0 927 926 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2241 927 926 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2242 0 929 928 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2243 929 928 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2244 196 524 922 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2245 197 524 923 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2246 198 524 924 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2247 199 524 925 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2248 200 524 926 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2249 201 524 927 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2250 202 524 928 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2251 203 524 929 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2252 930 527 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2253 931 527 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2254 932 527 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2255 933 527 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2256 934 527 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2257 935 527 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2258 936 527 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2259 937 527 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2260 0 931 930 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2261 931 930 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2262 0 933 932 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2263 933 932 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2264 0 935 934 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2265 935 934 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2266 0 937 936 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2267 937 936 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2268 1 931 930 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2269 931 930 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2270 1 933 932 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2271 933 932 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2272 1 939 938 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2273 939 938 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2274 1 941 940 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2275 941 940 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2276 1 935 934 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2277 935 934 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2278 1 937 936 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2279 937 936 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2280 1 943 942 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2281 943 942 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2282 1 945 944 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2283 945 944 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2284 0 939 938 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2285 939 938 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2286 0 941 940 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2287 941 940 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2288 0 943 942 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2289 943 942 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2290 0 945 944 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2291 945 944 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2292 196 532 938 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2293 197 532 939 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2294 198 532 940 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2295 199 532 941 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2296 200 532 942 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2297 201 532 943 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2298 202 532 944 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2299 203 532 945 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2300 946 536 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2301 947 536 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2302 948 536 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2303 949 536 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2304 950 536 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2305 951 536 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2306 952 536 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2307 953 536 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2308 0 947 946 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2309 947 946 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2310 0 949 948 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2311 949 948 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2312 0 951 950 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2313 951 950 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2314 0 953 952 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2315 953 952 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2316 1 947 946 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2317 947 946 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2318 1 949 948 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2319 949 948 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2320 1 951 950 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2321 951 950 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2322 1 953 952 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2323 953 952 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2324 1 955 954 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2325 955 954 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2326 1 957 956 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2327 957 956 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2328 1 959 958 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2329 959 958 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2330 1 961 960 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2331 961 960 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2332 0 955 954 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2333 955 954 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2334 0 957 956 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2335 957 956 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2336 0 959 958 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2337 959 958 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2338 0 961 960 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2339 961 960 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2340 196 540 954 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2341 197 540 955 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2342 198 540 956 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2343 199 540 957 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2344 200 540 958 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2345 201 540 959 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2346 202 540 960 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2347 203 540 961 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2348 962 543 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2349 963 543 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2350 964 543 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2351 965 543 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2352 966 543 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2353 967 543 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2354 968 543 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2355 969 543 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2356 0 963 962 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2357 963 962 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2358 0 965 964 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2359 965 964 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2360 0 967 966 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2361 967 966 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2362 0 969 968 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2363 969 968 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2364 1 963 962 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2365 963 962 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2366 1 965 964 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2367 965 964 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2368 1 971 970 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2369 971 970 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2370 1 973 972 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2371 973 972 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2372 1 967 966 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2373 967 966 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2374 1 969 968 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2375 969 968 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2376 1 975 974 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2377 975 974 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2378 1 977 976 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2379 977 976 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2380 0 971 970 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2381 971 970 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2382 0 973 972 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2383 973 972 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2384 0 975 974 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2385 975 974 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2386 0 977 976 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2387 977 976 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2388 196 548 970 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2389 197 548 971 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2390 198 548 972 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2391 199 548 973 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2392 200 548 974 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2393 201 548 975 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2394 202 548 976 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2395 203 548 977 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2396 978 552 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2397 979 552 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2398 980 552 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2399 981 552 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2400 982 552 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2401 983 552 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2402 984 552 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2403 985 552 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2404 0 979 978 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2405 979 978 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2406 0 981 980 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2407 981 980 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2408 0 983 982 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2409 983 982 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2410 0 985 984 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2411 985 984 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2412 1 979 978 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2413 979 978 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2414 1 981 980 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2415 981 980 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2416 1 983 982 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2417 983 982 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2418 1 985 984 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2419 985 984 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2420 1 987 986 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2421 987 986 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2422 1 989 988 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2423 989 988 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2424 1 991 990 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2425 991 990 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2426 1 993 992 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2427 993 992 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2428 0 987 986 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2429 987 986 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2430 0 989 988 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2431 989 988 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2432 0 991 990 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2433 991 990 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2434 0 993 992 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2435 993 992 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2436 196 556 986 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2437 197 556 987 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2438 198 556 988 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2439 199 556 989 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2440 200 556 990 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2441 201 556 991 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2442 202 556 992 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2443 203 556 993 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2444 994 559 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2445 995 559 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2446 996 559 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2447 997 559 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2448 998 559 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2449 999 559 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2450 1000 559 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2451 1001 559 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2452 0 995 994 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2453 995 994 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2454 0 997 996 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2455 997 996 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2456 0 999 998 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2457 999 998 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2458 0 1001 1000 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2459 1001 1000 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2460 1 995 994 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2461 995 994 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2462 1 997 996 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2463 997 996 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2464 1 1003 1002 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2465 1003 1002 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2466 1 1005 1004 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2467 1005 1004 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2468 1 999 998 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2469 999 998 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2470 1 1001 1000 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2471 1001 1000 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2472 1 1007 1006 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2473 1007 1006 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2474 1 1009 1008 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2475 1009 1008 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2476 0 1003 1002 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2477 1003 1002 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2478 0 1005 1004 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2479 1005 1004 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2480 0 1007 1006 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2481 1007 1006 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2482 0 1009 1008 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2483 1009 1008 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2484 196 564 1002 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2485 197 564 1003 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2486 198 564 1004 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2487 199 564 1005 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2488 200 564 1006 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2489 201 564 1007 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2490 202 564 1008 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2491 203 564 1009 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2492 1010 568 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2493 1011 568 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2494 1012 568 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2495 1013 568 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2496 1014 568 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2497 1015 568 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2498 1016 568 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2499 1017 568 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2500 0 1011 1010 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2501 1011 1010 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2502 0 1013 1012 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2503 1013 1012 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2504 0 1015 1014 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2505 1015 1014 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2506 0 1017 1016 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2507 1017 1016 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2508 1 1011 1010 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2509 1011 1010 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2510 1 1013 1012 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2511 1013 1012 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2512 1 1015 1014 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2513 1015 1014 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2514 1 1017 1016 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2515 1017 1016 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2516 1 1019 1018 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2517 1019 1018 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2518 1 1021 1020 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2519 1021 1020 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2520 1 1023 1022 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2521 1023 1022 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2522 1 1025 1024 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2523 1025 1024 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2524 0 1019 1018 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2525 1019 1018 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2526 0 1021 1020 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2527 1021 1020 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2528 0 1023 1022 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2529 1023 1022 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2530 0 1025 1024 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2531 1025 1024 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2532 196 572 1018 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2533 197 572 1019 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2534 198 572 1020 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2535 199 572 1021 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2536 200 572 1022 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2537 201 572 1023 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2538 202 572 1024 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2539 203 572 1025 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2540 1026 575 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2541 1027 575 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2542 1028 575 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2543 1029 575 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2544 1030 575 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2545 1031 575 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2546 1032 575 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2547 1033 575 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2548 0 1027 1026 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2549 1027 1026 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2550 0 1029 1028 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2551 1029 1028 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2552 0 1031 1030 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2553 1031 1030 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2554 0 1033 1032 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2555 1033 1032 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2556 1 1027 1026 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2557 1027 1026 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2558 1 1029 1028 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2559 1029 1028 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2560 1 1035 1034 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2561 1035 1034 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2562 1 1037 1036 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2563 1037 1036 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2564 1 1031 1030 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2565 1031 1030 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2566 1 1033 1032 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2567 1033 1032 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2568 1 1039 1038 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2569 1039 1038 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2570 1 1041 1040 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2571 1041 1040 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2572 0 1035 1034 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2573 1035 1034 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2574 0 1037 1036 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2575 1037 1036 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2576 0 1039 1038 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2577 1039 1038 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2578 0 1041 1040 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2579 1041 1040 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2580 196 580 1034 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2581 197 580 1035 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2582 198 580 1036 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2583 199 580 1037 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2584 200 580 1038 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2585 201 580 1039 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2586 202 580 1040 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2587 203 580 1041 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2588 1042 584 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2589 1043 584 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2590 1044 584 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2591 1045 584 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2592 1046 584 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2593 1047 584 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2594 1048 584 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2595 1049 584 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2596 0 1043 1042 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2597 1043 1042 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2598 0 1045 1044 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2599 1045 1044 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2600 0 1047 1046 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2601 1047 1046 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2602 0 1049 1048 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2603 1049 1048 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2604 1 1043 1042 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2605 1043 1042 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2606 1 1045 1044 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2607 1045 1044 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2608 1 1047 1046 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2609 1047 1046 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2610 1 1049 1048 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2611 1049 1048 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2612 1 1051 1050 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2613 1051 1050 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2614 1 1053 1052 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2615 1053 1052 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2616 1 1055 1054 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2617 1055 1054 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2618 1 1057 1056 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2619 1057 1056 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2620 0 1051 1050 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2621 1051 1050 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2622 0 1053 1052 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2623 1053 1052 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2624 0 1055 1054 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2625 1055 1054 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2626 0 1057 1056 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2627 1057 1056 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2628 196 588 1050 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2629 197 588 1051 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2630 198 588 1052 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2631 199 588 1053 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2632 200 588 1054 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2633 201 588 1055 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2634 202 588 1056 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2635 203 588 1057 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2636 1058 591 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2637 1059 591 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2638 1060 591 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2639 1061 591 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2640 1062 591 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2641 1063 591 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2642 1064 591 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2643 1065 591 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2644 0 1059 1058 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2645 1059 1058 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2646 0 1061 1060 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2647 1061 1060 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2648 0 1063 1062 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2649 1063 1062 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2650 0 1065 1064 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2651 1065 1064 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2652 1 1059 1058 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2653 1059 1058 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2654 1 1061 1060 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2655 1061 1060 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2656 1 1067 1066 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2657 1067 1066 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2658 1 1069 1068 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2659 1069 1068 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2660 1 1063 1062 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2661 1063 1062 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2662 1 1065 1064 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2663 1065 1064 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2664 1 1071 1070 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2665 1071 1070 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2666 1 1073 1072 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2667 1073 1072 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2668 0 1067 1066 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2669 1067 1066 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2670 0 1069 1068 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2671 1069 1068 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2672 0 1071 1070 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2673 1071 1070 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2674 0 1073 1072 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2675 1073 1072 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2676 196 596 1066 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2677 197 596 1067 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2678 198 596 1068 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2679 199 596 1069 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2680 200 596 1070 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2681 201 596 1071 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2682 202 596 1072 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2683 203 596 1073 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2684 1074 600 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2685 1075 600 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2686 1076 600 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2687 1077 600 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2688 1078 600 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2689 1079 600 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2690 1080 600 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2691 1081 600 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2692 0 1075 1074 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2693 1075 1074 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2694 0 1077 1076 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2695 1077 1076 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2696 0 1079 1078 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2697 1079 1078 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2698 0 1081 1080 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2699 1081 1080 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2700 1 1075 1074 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2701 1075 1074 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2702 1 1077 1076 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2703 1077 1076 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2704 1 1079 1078 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2705 1079 1078 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2706 1 1081 1080 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2707 1081 1080 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2708 1 1083 1082 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2709 1083 1082 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2710 1 1085 1084 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2711 1085 1084 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2712 1 1087 1086 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2713 1087 1086 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2714 1 1089 1088 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2715 1089 1088 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2716 0 1083 1082 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2717 1083 1082 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2718 0 1085 1084 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2719 1085 1084 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2720 0 1087 1086 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2721 1087 1086 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2722 0 1089 1088 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2723 1089 1088 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2724 196 604 1082 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2725 197 604 1083 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2726 198 604 1084 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2727 199 604 1085 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2728 200 604 1086 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2729 201 604 1087 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2730 202 604 1088 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2731 203 604 1089 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2732 1090 607 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2733 1091 607 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2734 1092 607 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2735 1093 607 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2736 1094 607 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2737 1095 607 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2738 1096 607 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2739 1097 607 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2740 0 1091 1090 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2741 1091 1090 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2742 0 1093 1092 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2743 1093 1092 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2744 0 1095 1094 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2745 1095 1094 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2746 0 1097 1096 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2747 1097 1096 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2748 1 1091 1090 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2749 1091 1090 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2750 1 1093 1092 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2751 1093 1092 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2752 1 1099 1098 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2753 1099 1098 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2754 1 1101 1100 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2755 1101 1100 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2756 1 1095 1094 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2757 1095 1094 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2758 1 1097 1096 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2759 1097 1096 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2760 1 1103 1102 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2761 1103 1102 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2762 1 1105 1104 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2763 1105 1104 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2764 0 1099 1098 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2765 1099 1098 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2766 0 1101 1100 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2767 1101 1100 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2768 0 1103 1102 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2769 1103 1102 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2770 0 1105 1104 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2771 1105 1104 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2772 196 612 1098 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2773 197 612 1099 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2774 198 612 1100 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2775 199 612 1101 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2776 200 612 1102 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2777 201 612 1103 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2778 202 612 1104 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2779 203 612 1105 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2780 1106 616 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2781 1107 616 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2782 1108 616 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2783 1109 616 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2784 1110 616 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2785 1111 616 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2786 1112 616 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2787 1113 616 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2788 0 1107 1106 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2789 1107 1106 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2790 0 1109 1108 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2791 1109 1108 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2792 0 1111 1110 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2793 1111 1110 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2794 0 1113 1112 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2795 1113 1112 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2796 1 1107 1106 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2797 1107 1106 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2798 1 1109 1108 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2799 1109 1108 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2800 1 1111 1110 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2801 1111 1110 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2802 1 1113 1112 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2803 1113 1112 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2804 1 1115 1114 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2805 1115 1114 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2806 1 1117 1116 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2807 1117 1116 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2808 1 1119 1118 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2809 1119 1118 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2810 1 1121 1120 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2811 1121 1120 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2812 0 1115 1114 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2813 1115 1114 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2814 0 1117 1116 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2815 1117 1116 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2816 0 1119 1118 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2817 1119 1118 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2818 0 1121 1120 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2819 1121 1120 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2820 196 620 1114 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2821 197 620 1115 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2822 198 620 1116 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2823 199 620 1117 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2824 200 620 1118 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2825 201 620 1119 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2826 202 620 1120 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2827 203 620 1121 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2828 1122 624 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2829 1123 624 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2830 1124 624 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2831 1125 624 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2832 1126 624 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2833 1127 624 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2834 1128 624 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2835 1129 624 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2836 0 1123 1122 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2837 1123 1122 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2838 0 1125 1124 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2839 1125 1124 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2840 0 1127 1126 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2841 1127 1126 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2842 0 1129 1128 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2843 1129 1128 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2844 1 1123 1122 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2845 1123 1122 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2846 1 1125 1124 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2847 1125 1124 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2848 1 1131 1130 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2849 1131 1130 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2850 1 1133 1132 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2851 1133 1132 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2852 1 1127 1126 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2853 1127 1126 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2854 1 1129 1128 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2855 1129 1128 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2856 1 1135 1134 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2857 1135 1134 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2858 1 1137 1136 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2859 1137 1136 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2860 0 1131 1130 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2861 1131 1130 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2862 0 1133 1132 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2863 1133 1132 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2864 0 1135 1134 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2865 1135 1134 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2866 0 1137 1136 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2867 1137 1136 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2868 196 628 1130 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2869 197 628 1131 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2870 198 628 1132 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2871 199 628 1133 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2872 200 628 1134 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2873 201 628 1135 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2874 202 628 1136 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2875 203 628 1137 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2876 1138 632 196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2877 1139 632 197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2878 1140 632 198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2879 1141 632 199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2880 1142 632 200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2881 1143 632 201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2882 1144 632 202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2883 1145 632 203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2884 0 1139 1138 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2885 1139 1138 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2886 0 1141 1140 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2887 1141 1140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2888 0 1143 1142 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2889 1143 1142 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2890 0 1145 1144 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2891 1145 1144 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2892 1 1139 1138 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2893 1139 1138 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2894 1 1141 1140 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2895 1141 1140 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2896 1 1143 1142 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2897 1143 1142 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2898 1 1145 1144 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2899 1145 1144 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2900 1 1147 1146 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2901 1147 1146 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2902 1 1149 1148 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2903 1149 1148 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2904 1 1151 1150 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2905 1151 1150 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2906 1 1153 1152 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2907 1153 1152 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2908 0 1147 1146 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2909 1147 1146 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2910 0 1149 1148 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2911 1149 1148 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2912 0 1151 1150 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2913 1151 1150 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2914 0 1153 1152 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2915 1153 1152 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2916 222 380 1146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2917 223 380 1147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2918 224 380 1148 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2919 225 380 1149 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2920 226 380 1150 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2921 227 380 1151 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2922 228 380 1152 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2923 229 380 1153 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2924 1154 383 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2925 1155 383 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2926 1156 383 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2927 1157 383 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2928 1158 383 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2929 1159 383 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2930 1160 383 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2931 1161 383 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2932 0 1155 1154 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2933 1155 1154 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2934 0 1157 1156 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2935 1157 1156 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2936 0 1159 1158 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2937 1159 1158 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2938 0 1161 1160 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2939 1161 1160 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2940 1 1155 1154 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2941 1155 1154 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2942 1 1157 1156 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2943 1157 1156 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2944 1 1163 1162 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2945 1163 1162 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2946 1 1165 1164 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2947 1165 1164 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2948 1 1159 1158 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2949 1159 1158 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2950 1 1161 1160 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2951 1161 1160 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2952 1 1167 1166 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2953 1167 1166 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2954 1 1169 1168 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m2955 1169 1168 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2956 0 1163 1162 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2957 1163 1162 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2958 0 1165 1164 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2959 1165 1164 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2960 0 1167 1166 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2961 1167 1166 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2962 0 1169 1168 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2963 1169 1168 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2964 222 388 1162 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m2965 223 388 1163 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2966 224 388 1164 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2967 225 388 1165 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2968 226 388 1166 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m2969 227 388 1167 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m2970 228 388 1168 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m2971 229 388 1169 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m2972 1170 392 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m2973 1171 392 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2974 1172 392 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2975 1173 392 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2976 1174 392 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m2977 1175 392 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m2978 1176 392 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m2979 1177 392 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m2980 0 1171 1170 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2981 1171 1170 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2982 0 1173 1172 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m2983 1173 1172 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m2984 0 1175 1174 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2985 1175 1174 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2986 0 1177 1176 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m2987 1177 1176 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m2988 1 1171 1170 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2989 1171 1170 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2990 1 1173 1172 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2991 1173 1172 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2992 1 1175 1174 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2993 1175 1174 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2994 1 1177 1176 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2995 1177 1176 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m2996 1 1179 1178 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2997 1179 1178 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m2998 1 1181 1180 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m2999 1181 1180 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3000 1 1183 1182 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3001 1183 1182 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3002 1 1185 1184 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3003 1185 1184 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3004 0 1179 1178 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3005 1179 1178 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3006 0 1181 1180 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3007 1181 1180 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3008 0 1183 1182 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3009 1183 1182 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3010 0 1185 1184 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3011 1185 1184 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3012 222 396 1178 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3013 223 396 1179 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3014 224 396 1180 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3015 225 396 1181 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3016 226 396 1182 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3017 227 396 1183 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3018 228 396 1184 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3019 229 396 1185 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3020 1186 399 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3021 1187 399 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3022 1188 399 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3023 1189 399 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3024 1190 399 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3025 1191 399 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3026 1192 399 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3027 1193 399 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3028 0 1187 1186 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3029 1187 1186 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3030 0 1189 1188 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3031 1189 1188 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3032 0 1191 1190 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3033 1191 1190 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3034 0 1193 1192 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3035 1193 1192 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3036 1 1187 1186 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3037 1187 1186 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3038 1 1189 1188 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3039 1189 1188 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3040 1 1195 1194 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3041 1195 1194 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3042 1 1197 1196 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3043 1197 1196 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3044 1 1191 1190 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3045 1191 1190 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3046 1 1193 1192 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3047 1193 1192 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3048 1 1199 1198 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3049 1199 1198 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3050 1 1201 1200 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3051 1201 1200 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3052 0 1195 1194 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3053 1195 1194 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3054 0 1197 1196 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3055 1197 1196 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3056 0 1199 1198 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3057 1199 1198 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3058 0 1201 1200 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3059 1201 1200 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3060 222 404 1194 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3061 223 404 1195 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3062 224 404 1196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3063 225 404 1197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3064 226 404 1198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3065 227 404 1199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3066 228 404 1200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3067 229 404 1201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3068 1202 408 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3069 1203 408 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3070 1204 408 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3071 1205 408 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3072 1206 408 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3073 1207 408 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3074 1208 408 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3075 1209 408 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3076 0 1203 1202 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3077 1203 1202 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3078 0 1205 1204 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3079 1205 1204 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3080 0 1207 1206 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3081 1207 1206 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3082 0 1209 1208 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3083 1209 1208 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3084 1 1203 1202 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3085 1203 1202 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3086 1 1205 1204 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3087 1205 1204 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3088 1 1207 1206 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3089 1207 1206 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3090 1 1209 1208 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3091 1209 1208 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3092 1 1211 1210 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3093 1211 1210 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3094 1 1213 1212 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3095 1213 1212 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3096 1 1215 1214 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3097 1215 1214 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3098 1 1217 1216 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3099 1217 1216 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3100 0 1211 1210 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3101 1211 1210 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3102 0 1213 1212 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3103 1213 1212 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3104 0 1215 1214 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3105 1215 1214 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3106 0 1217 1216 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3107 1217 1216 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3108 222 412 1210 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3109 223 412 1211 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3110 224 412 1212 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3111 225 412 1213 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3112 226 412 1214 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3113 227 412 1215 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3114 228 412 1216 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3115 229 412 1217 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3116 1218 415 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3117 1219 415 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3118 1220 415 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3119 1221 415 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3120 1222 415 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3121 1223 415 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3122 1224 415 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3123 1225 415 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3124 0 1219 1218 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3125 1219 1218 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3126 0 1221 1220 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3127 1221 1220 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3128 0 1223 1222 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3129 1223 1222 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3130 0 1225 1224 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3131 1225 1224 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3132 1 1219 1218 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3133 1219 1218 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3134 1 1221 1220 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3135 1221 1220 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3136 1 1227 1226 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3137 1227 1226 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3138 1 1229 1228 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3139 1229 1228 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3140 1 1223 1222 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3141 1223 1222 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3142 1 1225 1224 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3143 1225 1224 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3144 1 1231 1230 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3145 1231 1230 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3146 1 1233 1232 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3147 1233 1232 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3148 0 1227 1226 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3149 1227 1226 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3150 0 1229 1228 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3151 1229 1228 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3152 0 1231 1230 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3153 1231 1230 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3154 0 1233 1232 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3155 1233 1232 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3156 222 420 1226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3157 223 420 1227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3158 224 420 1228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3159 225 420 1229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3160 226 420 1230 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3161 227 420 1231 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3162 228 420 1232 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3163 229 420 1233 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3164 1234 424 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3165 1235 424 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3166 1236 424 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3167 1237 424 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3168 1238 424 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3169 1239 424 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3170 1240 424 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3171 1241 424 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3172 0 1235 1234 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3173 1235 1234 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3174 0 1237 1236 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3175 1237 1236 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3176 0 1239 1238 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3177 1239 1238 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3178 0 1241 1240 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3179 1241 1240 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3180 1 1235 1234 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3181 1235 1234 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3182 1 1237 1236 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3183 1237 1236 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3184 1 1239 1238 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3185 1239 1238 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3186 1 1241 1240 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3187 1241 1240 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3188 1 1243 1242 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3189 1243 1242 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3190 1 1245 1244 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3191 1245 1244 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3192 1 1247 1246 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3193 1247 1246 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3194 1 1249 1248 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3195 1249 1248 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3196 0 1243 1242 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3197 1243 1242 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3198 0 1245 1244 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3199 1245 1244 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3200 0 1247 1246 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3201 1247 1246 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3202 0 1249 1248 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3203 1249 1248 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3204 222 428 1242 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3205 223 428 1243 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3206 224 428 1244 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3207 225 428 1245 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3208 226 428 1246 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3209 227 428 1247 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3210 228 428 1248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3211 229 428 1249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3212 1250 431 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3213 1251 431 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3214 1252 431 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3215 1253 431 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3216 1254 431 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3217 1255 431 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3218 1256 431 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3219 1257 431 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3220 0 1251 1250 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3221 1251 1250 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3222 0 1253 1252 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3223 1253 1252 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3224 0 1255 1254 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3225 1255 1254 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3226 0 1257 1256 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3227 1257 1256 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3228 1 1251 1250 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3229 1251 1250 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3230 1 1253 1252 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3231 1253 1252 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3232 1 1259 1258 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3233 1259 1258 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3234 1 1261 1260 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3235 1261 1260 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3236 1 1255 1254 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3237 1255 1254 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3238 1 1257 1256 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3239 1257 1256 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3240 1 1263 1262 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3241 1263 1262 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3242 1 1265 1264 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3243 1265 1264 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3244 0 1259 1258 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3245 1259 1258 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3246 0 1261 1260 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3247 1261 1260 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3248 0 1263 1262 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3249 1263 1262 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3250 0 1265 1264 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3251 1265 1264 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3252 222 436 1258 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3253 223 436 1259 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3254 224 436 1260 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3255 225 436 1261 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3256 226 436 1262 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3257 227 436 1263 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3258 228 436 1264 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3259 229 436 1265 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3260 1266 440 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3261 1267 440 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3262 1268 440 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3263 1269 440 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3264 1270 440 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3265 1271 440 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3266 1272 440 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3267 1273 440 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3268 0 1267 1266 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3269 1267 1266 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3270 0 1269 1268 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3271 1269 1268 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3272 0 1271 1270 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3273 1271 1270 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3274 0 1273 1272 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3275 1273 1272 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3276 1 1267 1266 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3277 1267 1266 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3278 1 1269 1268 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3279 1269 1268 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3280 1 1271 1270 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3281 1271 1270 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3282 1 1273 1272 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3283 1273 1272 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3284 1 1275 1274 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3285 1275 1274 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3286 1 1277 1276 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3287 1277 1276 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3288 1 1279 1278 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3289 1279 1278 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3290 1 1281 1280 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3291 1281 1280 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3292 0 1275 1274 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3293 1275 1274 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3294 0 1277 1276 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3295 1277 1276 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3296 0 1279 1278 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3297 1279 1278 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3298 0 1281 1280 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3299 1281 1280 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3300 222 444 1274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3301 223 444 1275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3302 224 444 1276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3303 225 444 1277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3304 226 444 1278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3305 227 444 1279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3306 228 444 1280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3307 229 444 1281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3308 1282 447 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3309 1283 447 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3310 1284 447 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3311 1285 447 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3312 1286 447 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3313 1287 447 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3314 1288 447 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3315 1289 447 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3316 0 1283 1282 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3317 1283 1282 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3318 0 1285 1284 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3319 1285 1284 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3320 0 1287 1286 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3321 1287 1286 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3322 0 1289 1288 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3323 1289 1288 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3324 1 1283 1282 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3325 1283 1282 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3326 1 1285 1284 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3327 1285 1284 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3328 1 1291 1290 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3329 1291 1290 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3330 1 1293 1292 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3331 1293 1292 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3332 1 1287 1286 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3333 1287 1286 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3334 1 1289 1288 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3335 1289 1288 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3336 1 1295 1294 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3337 1295 1294 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3338 1 1297 1296 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3339 1297 1296 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3340 0 1291 1290 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3341 1291 1290 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3342 0 1293 1292 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3343 1293 1292 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3344 0 1295 1294 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3345 1295 1294 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3346 0 1297 1296 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3347 1297 1296 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3348 222 452 1290 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3349 223 452 1291 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3350 224 452 1292 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3351 225 452 1293 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3352 226 452 1294 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3353 227 452 1295 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3354 228 452 1296 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3355 229 452 1297 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3356 1298 456 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3357 1299 456 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3358 1300 456 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3359 1301 456 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3360 1302 456 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3361 1303 456 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3362 1304 456 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3363 1305 456 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3364 0 1299 1298 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3365 1299 1298 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3366 0 1301 1300 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3367 1301 1300 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3368 0 1303 1302 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3369 1303 1302 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3370 0 1305 1304 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3371 1305 1304 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3372 1 1299 1298 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3373 1299 1298 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3374 1 1301 1300 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3375 1301 1300 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3376 1 1303 1302 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3377 1303 1302 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3378 1 1305 1304 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3379 1305 1304 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3380 1 1307 1306 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3381 1307 1306 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3382 1 1309 1308 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3383 1309 1308 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3384 1 1311 1310 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3385 1311 1310 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3386 1 1313 1312 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3387 1313 1312 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3388 0 1307 1306 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3389 1307 1306 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3390 0 1309 1308 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3391 1309 1308 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3392 0 1311 1310 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3393 1311 1310 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3394 0 1313 1312 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3395 1313 1312 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3396 222 460 1306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3397 223 460 1307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3398 224 460 1308 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3399 225 460 1309 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3400 226 460 1310 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3401 227 460 1311 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3402 228 460 1312 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3403 229 460 1313 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3404 1314 463 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3405 1315 463 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3406 1316 463 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3407 1317 463 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3408 1318 463 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3409 1319 463 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3410 1320 463 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3411 1321 463 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3412 0 1315 1314 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3413 1315 1314 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3414 0 1317 1316 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3415 1317 1316 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3416 0 1319 1318 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3417 1319 1318 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3418 0 1321 1320 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3419 1321 1320 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3420 1 1315 1314 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3421 1315 1314 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3422 1 1317 1316 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3423 1317 1316 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3424 1 1323 1322 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3425 1323 1322 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3426 1 1325 1324 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3427 1325 1324 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3428 1 1319 1318 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3429 1319 1318 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3430 1 1321 1320 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3431 1321 1320 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3432 1 1327 1326 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3433 1327 1326 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3434 1 1329 1328 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3435 1329 1328 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3436 0 1323 1322 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3437 1323 1322 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3438 0 1325 1324 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3439 1325 1324 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3440 0 1327 1326 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3441 1327 1326 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3442 0 1329 1328 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3443 1329 1328 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3444 222 468 1322 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3445 223 468 1323 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3446 224 468 1324 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3447 225 468 1325 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3448 226 468 1326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3449 227 468 1327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3450 228 468 1328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3451 229 468 1329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3452 1330 472 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3453 1331 472 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3454 1332 472 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3455 1333 472 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3456 1334 472 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3457 1335 472 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3458 1336 472 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3459 1337 472 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3460 0 1331 1330 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3461 1331 1330 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3462 0 1333 1332 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3463 1333 1332 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3464 0 1335 1334 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3465 1335 1334 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3466 0 1337 1336 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3467 1337 1336 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3468 1 1331 1330 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3469 1331 1330 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3470 1 1333 1332 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3471 1333 1332 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3472 1 1335 1334 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3473 1335 1334 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3474 1 1337 1336 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3475 1337 1336 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3476 1 1339 1338 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3477 1339 1338 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3478 1 1341 1340 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3479 1341 1340 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3480 1 1343 1342 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3481 1343 1342 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3482 1 1345 1344 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3483 1345 1344 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3484 0 1339 1338 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3485 1339 1338 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3486 0 1341 1340 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3487 1341 1340 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3488 0 1343 1342 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3489 1343 1342 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3490 0 1345 1344 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3491 1345 1344 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3492 222 476 1338 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3493 223 476 1339 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3494 224 476 1340 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3495 225 476 1341 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3496 226 476 1342 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3497 227 476 1343 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3498 228 476 1344 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3499 229 476 1345 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3500 1346 479 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3501 1347 479 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3502 1348 479 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3503 1349 479 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3504 1350 479 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3505 1351 479 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3506 1352 479 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3507 1353 479 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3508 0 1347 1346 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3509 1347 1346 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3510 0 1349 1348 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3511 1349 1348 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3512 0 1351 1350 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3513 1351 1350 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3514 0 1353 1352 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3515 1353 1352 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3516 1 1347 1346 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3517 1347 1346 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3518 1 1349 1348 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3519 1349 1348 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3520 1 1355 1354 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3521 1355 1354 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3522 1 1357 1356 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3523 1357 1356 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3524 1 1351 1350 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3525 1351 1350 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3526 1 1353 1352 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3527 1353 1352 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3528 1 1359 1358 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3529 1359 1358 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3530 1 1361 1360 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3531 1361 1360 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3532 0 1355 1354 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3533 1355 1354 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3534 0 1357 1356 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3535 1357 1356 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3536 0 1359 1358 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3537 1359 1358 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3538 0 1361 1360 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3539 1361 1360 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3540 222 484 1354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3541 223 484 1355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3542 224 484 1356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3543 225 484 1357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3544 226 484 1358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3545 227 484 1359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3546 228 484 1360 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3547 229 484 1361 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3548 1362 488 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3549 1363 488 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3550 1364 488 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3551 1365 488 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3552 1366 488 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3553 1367 488 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3554 1368 488 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3555 1369 488 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3556 0 1363 1362 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3557 1363 1362 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3558 0 1365 1364 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3559 1365 1364 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3560 0 1367 1366 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3561 1367 1366 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3562 0 1369 1368 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3563 1369 1368 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3564 1 1363 1362 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3565 1363 1362 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3566 1 1365 1364 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3567 1365 1364 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3568 1 1367 1366 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3569 1367 1366 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3570 1 1369 1368 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3571 1369 1368 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3572 1 1371 1370 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3573 1371 1370 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3574 1 1373 1372 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3575 1373 1372 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3576 1 1375 1374 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3577 1375 1374 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3578 1 1377 1376 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3579 1377 1376 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3580 0 1371 1370 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3581 1371 1370 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3582 0 1373 1372 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3583 1373 1372 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3584 0 1375 1374 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3585 1375 1374 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3586 0 1377 1376 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3587 1377 1376 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3588 222 492 1370 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3589 223 492 1371 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3590 224 492 1372 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3591 225 492 1373 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3592 226 492 1374 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3593 227 492 1375 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3594 228 492 1376 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3595 229 492 1377 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3596 1378 495 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3597 1379 495 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3598 1380 495 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3599 1381 495 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3600 1382 495 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3601 1383 495 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3602 1384 495 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3603 1385 495 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3604 0 1379 1378 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3605 1379 1378 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3606 0 1381 1380 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3607 1381 1380 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3608 0 1383 1382 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3609 1383 1382 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3610 0 1385 1384 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3611 1385 1384 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3612 1 1379 1378 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3613 1379 1378 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3614 1 1381 1380 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3615 1381 1380 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3616 1 1387 1386 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3617 1387 1386 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3618 1 1389 1388 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3619 1389 1388 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3620 1 1383 1382 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3621 1383 1382 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3622 1 1385 1384 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3623 1385 1384 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3624 1 1391 1390 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3625 1391 1390 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3626 1 1393 1392 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3627 1393 1392 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3628 0 1387 1386 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3629 1387 1386 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3630 0 1389 1388 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3631 1389 1388 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3632 0 1391 1390 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3633 1391 1390 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3634 0 1393 1392 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3635 1393 1392 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3636 222 500 1386 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3637 223 500 1387 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3638 224 500 1388 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3639 225 500 1389 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3640 226 500 1390 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3641 227 500 1391 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3642 228 500 1392 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3643 229 500 1393 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3644 1394 504 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3645 1395 504 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3646 1396 504 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3647 1397 504 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3648 1398 504 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3649 1399 504 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3650 1400 504 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3651 1401 504 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3652 0 1395 1394 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3653 1395 1394 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3654 0 1397 1396 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3655 1397 1396 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3656 0 1399 1398 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3657 1399 1398 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3658 0 1401 1400 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3659 1401 1400 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3660 1 1395 1394 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3661 1395 1394 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3662 1 1397 1396 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3663 1397 1396 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3664 1 1399 1398 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3665 1399 1398 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3666 1 1401 1400 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3667 1401 1400 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3668 1 1403 1402 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3669 1403 1402 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3670 1 1405 1404 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3671 1405 1404 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3672 1 1407 1406 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3673 1407 1406 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3674 1 1409 1408 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3675 1409 1408 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3676 0 1403 1402 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3677 1403 1402 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3678 0 1405 1404 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3679 1405 1404 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3680 0 1407 1406 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3681 1407 1406 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3682 0 1409 1408 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3683 1409 1408 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3684 222 508 1402 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3685 223 508 1403 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3686 224 508 1404 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3687 225 508 1405 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3688 226 508 1406 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3689 227 508 1407 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3690 228 508 1408 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3691 229 508 1409 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3692 1410 511 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3693 1411 511 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3694 1412 511 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3695 1413 511 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3696 1414 511 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3697 1415 511 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3698 1416 511 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3699 1417 511 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3700 0 1411 1410 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3701 1411 1410 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3702 0 1413 1412 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3703 1413 1412 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3704 0 1415 1414 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3705 1415 1414 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3706 0 1417 1416 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3707 1417 1416 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3708 1 1411 1410 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3709 1411 1410 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3710 1 1413 1412 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3711 1413 1412 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3712 1 1419 1418 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3713 1419 1418 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3714 1 1421 1420 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3715 1421 1420 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3716 1 1415 1414 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3717 1415 1414 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3718 1 1417 1416 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3719 1417 1416 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3720 1 1423 1422 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3721 1423 1422 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3722 1 1425 1424 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3723 1425 1424 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3724 0 1419 1418 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3725 1419 1418 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3726 0 1421 1420 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3727 1421 1420 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3728 0 1423 1422 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3729 1423 1422 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3730 0 1425 1424 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3731 1425 1424 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3732 222 516 1418 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3733 223 516 1419 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3734 224 516 1420 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3735 225 516 1421 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3736 226 516 1422 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3737 227 516 1423 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3738 228 516 1424 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3739 229 516 1425 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3740 1426 520 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3741 1427 520 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3742 1428 520 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3743 1429 520 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3744 1430 520 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3745 1431 520 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3746 1432 520 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3747 1433 520 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3748 0 1427 1426 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3749 1427 1426 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3750 0 1429 1428 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3751 1429 1428 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3752 0 1431 1430 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3753 1431 1430 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3754 0 1433 1432 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3755 1433 1432 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3756 1 1427 1426 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3757 1427 1426 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3758 1 1429 1428 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3759 1429 1428 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3760 1 1431 1430 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3761 1431 1430 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3762 1 1433 1432 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3763 1433 1432 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3764 1 1435 1434 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3765 1435 1434 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3766 1 1437 1436 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3767 1437 1436 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3768 1 1439 1438 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3769 1439 1438 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3770 1 1441 1440 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3771 1441 1440 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3772 0 1435 1434 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3773 1435 1434 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3774 0 1437 1436 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3775 1437 1436 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3776 0 1439 1438 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3777 1439 1438 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3778 0 1441 1440 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3779 1441 1440 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3780 222 524 1434 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3781 223 524 1435 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3782 224 524 1436 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3783 225 524 1437 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3784 226 524 1438 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3785 227 524 1439 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3786 228 524 1440 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3787 229 524 1441 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3788 1442 527 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3789 1443 527 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3790 1444 527 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3791 1445 527 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3792 1446 527 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3793 1447 527 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3794 1448 527 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3795 1449 527 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3796 0 1443 1442 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3797 1443 1442 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3798 0 1445 1444 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3799 1445 1444 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3800 0 1447 1446 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3801 1447 1446 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3802 0 1449 1448 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3803 1449 1448 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3804 1 1443 1442 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3805 1443 1442 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3806 1 1445 1444 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3807 1445 1444 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3808 1 1451 1450 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3809 1451 1450 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3810 1 1453 1452 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3811 1453 1452 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3812 1 1447 1446 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3813 1447 1446 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3814 1 1449 1448 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3815 1449 1448 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3816 1 1455 1454 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3817 1455 1454 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3818 1 1457 1456 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3819 1457 1456 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3820 0 1451 1450 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3821 1451 1450 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3822 0 1453 1452 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3823 1453 1452 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3824 0 1455 1454 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3825 1455 1454 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3826 0 1457 1456 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3827 1457 1456 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3828 222 532 1450 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3829 223 532 1451 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3830 224 532 1452 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3831 225 532 1453 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3832 226 532 1454 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3833 227 532 1455 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3834 228 532 1456 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3835 229 532 1457 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3836 1458 536 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3837 1459 536 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3838 1460 536 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3839 1461 536 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3840 1462 536 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3841 1463 536 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3842 1464 536 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3843 1465 536 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3844 0 1459 1458 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3845 1459 1458 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3846 0 1461 1460 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3847 1461 1460 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3848 0 1463 1462 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3849 1463 1462 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3850 0 1465 1464 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3851 1465 1464 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3852 1 1459 1458 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3853 1459 1458 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3854 1 1461 1460 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3855 1461 1460 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3856 1 1463 1462 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3857 1463 1462 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3858 1 1465 1464 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3859 1465 1464 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3860 1 1467 1466 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3861 1467 1466 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3862 1 1469 1468 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3863 1469 1468 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3864 1 1471 1470 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3865 1471 1470 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3866 1 1473 1472 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3867 1473 1472 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3868 0 1467 1466 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3869 1467 1466 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3870 0 1469 1468 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3871 1469 1468 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3872 0 1471 1470 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3873 1471 1470 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3874 0 1473 1472 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3875 1473 1472 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3876 222 540 1466 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3877 223 540 1467 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3878 224 540 1468 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3879 225 540 1469 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3880 226 540 1470 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3881 227 540 1471 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3882 228 540 1472 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3883 229 540 1473 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3884 1474 543 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3885 1475 543 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3886 1476 543 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3887 1477 543 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3888 1478 543 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3889 1479 543 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3890 1480 543 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3891 1481 543 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3892 0 1475 1474 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3893 1475 1474 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3894 0 1477 1476 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3895 1477 1476 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3896 0 1479 1478 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3897 1479 1478 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3898 0 1481 1480 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3899 1481 1480 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3900 1 1475 1474 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3901 1475 1474 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3902 1 1477 1476 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3903 1477 1476 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3904 1 1483 1482 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3905 1483 1482 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3906 1 1485 1484 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3907 1485 1484 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3908 1 1479 1478 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3909 1479 1478 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3910 1 1481 1480 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3911 1481 1480 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3912 1 1487 1486 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3913 1487 1486 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3914 1 1489 1488 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3915 1489 1488 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3916 0 1483 1482 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3917 1483 1482 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3918 0 1485 1484 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3919 1485 1484 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3920 0 1487 1486 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3921 1487 1486 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3922 0 1489 1488 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3923 1489 1488 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3924 222 548 1482 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3925 223 548 1483 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3926 224 548 1484 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3927 225 548 1485 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3928 226 548 1486 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3929 227 548 1487 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3930 228 548 1488 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3931 229 548 1489 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3932 1490 552 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3933 1491 552 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3934 1492 552 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3935 1493 552 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3936 1494 552 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3937 1495 552 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3938 1496 552 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3939 1497 552 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3940 0 1491 1490 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3941 1491 1490 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3942 0 1493 1492 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3943 1493 1492 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3944 0 1495 1494 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3945 1495 1494 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3946 0 1497 1496 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3947 1497 1496 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3948 1 1491 1490 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3949 1491 1490 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3950 1 1493 1492 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3951 1493 1492 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3952 1 1495 1494 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3953 1495 1494 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3954 1 1497 1496 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3955 1497 1496 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3956 1 1499 1498 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3957 1499 1498 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m3958 1 1501 1500 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3959 1501 1500 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3960 1 1503 1502 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3961 1503 1502 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3962 1 1505 1504 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m3963 1505 1504 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3964 0 1499 1498 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3965 1499 1498 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3966 0 1501 1500 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3967 1501 1500 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3968 0 1503 1502 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3969 1503 1502 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3970 0 1505 1504 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3971 1505 1504 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3972 222 556 1498 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m3973 223 556 1499 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3974 224 556 1500 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3975 225 556 1501 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3976 226 556 1502 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m3977 227 556 1503 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m3978 228 556 1504 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m3979 229 556 1505 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m3980 1506 559 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m3981 1507 559 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3982 1508 559 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3983 1509 559 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3984 1510 559 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m3985 1511 559 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m3986 1512 559 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m3987 1513 559 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m3988 0 1507 1506 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3989 1507 1506 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3990 0 1509 1508 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m3991 1509 1508 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m3992 0 1511 1510 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3993 1511 1510 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3994 0 1513 1512 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m3995 1513 1512 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m3996 1 1507 1506 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3997 1507 1506 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m3998 1 1509 1508 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m3999 1509 1508 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4000 1 1515 1514 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4001 1515 1514 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4002 1 1517 1516 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4003 1517 1516 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4004 1 1511 1510 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4005 1511 1510 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4006 1 1513 1512 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4007 1513 1512 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4008 1 1519 1518 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4009 1519 1518 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4010 1 1521 1520 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4011 1521 1520 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4012 0 1515 1514 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4013 1515 1514 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4014 0 1517 1516 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4015 1517 1516 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4016 0 1519 1518 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4017 1519 1518 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4018 0 1521 1520 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4019 1521 1520 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4020 222 564 1514 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4021 223 564 1515 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4022 224 564 1516 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4023 225 564 1517 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4024 226 564 1518 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4025 227 564 1519 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4026 228 564 1520 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4027 229 564 1521 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4028 1522 568 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4029 1523 568 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4030 1524 568 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4031 1525 568 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4032 1526 568 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4033 1527 568 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4034 1528 568 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4035 1529 568 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4036 0 1523 1522 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4037 1523 1522 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4038 0 1525 1524 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4039 1525 1524 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4040 0 1527 1526 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4041 1527 1526 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4042 0 1529 1528 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4043 1529 1528 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4044 1 1523 1522 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4045 1523 1522 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4046 1 1525 1524 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4047 1525 1524 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4048 1 1527 1526 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4049 1527 1526 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4050 1 1529 1528 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4051 1529 1528 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4052 1 1531 1530 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4053 1531 1530 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4054 1 1533 1532 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4055 1533 1532 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4056 1 1535 1534 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4057 1535 1534 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4058 1 1537 1536 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4059 1537 1536 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4060 0 1531 1530 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4061 1531 1530 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4062 0 1533 1532 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4063 1533 1532 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4064 0 1535 1534 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4065 1535 1534 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4066 0 1537 1536 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4067 1537 1536 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4068 222 572 1530 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4069 223 572 1531 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4070 224 572 1532 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4071 225 572 1533 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4072 226 572 1534 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4073 227 572 1535 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4074 228 572 1536 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4075 229 572 1537 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4076 1538 575 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4077 1539 575 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4078 1540 575 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4079 1541 575 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4080 1542 575 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4081 1543 575 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4082 1544 575 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4083 1545 575 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4084 0 1539 1538 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4085 1539 1538 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4086 0 1541 1540 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4087 1541 1540 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4088 0 1543 1542 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4089 1543 1542 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4090 0 1545 1544 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4091 1545 1544 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4092 1 1539 1538 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4093 1539 1538 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4094 1 1541 1540 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4095 1541 1540 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4096 1 1547 1546 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4097 1547 1546 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4098 1 1549 1548 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4099 1549 1548 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4100 1 1543 1542 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4101 1543 1542 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4102 1 1545 1544 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4103 1545 1544 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4104 1 1551 1550 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4105 1551 1550 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4106 1 1553 1552 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4107 1553 1552 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4108 0 1547 1546 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4109 1547 1546 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4110 0 1549 1548 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4111 1549 1548 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4112 0 1551 1550 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4113 1551 1550 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4114 0 1553 1552 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4115 1553 1552 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4116 222 580 1546 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4117 223 580 1547 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4118 224 580 1548 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4119 225 580 1549 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4120 226 580 1550 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4121 227 580 1551 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4122 228 580 1552 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4123 229 580 1553 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4124 1554 584 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4125 1555 584 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4126 1556 584 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4127 1557 584 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4128 1558 584 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4129 1559 584 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4130 1560 584 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4131 1561 584 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4132 0 1555 1554 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4133 1555 1554 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4134 0 1557 1556 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4135 1557 1556 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4136 0 1559 1558 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4137 1559 1558 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4138 0 1561 1560 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4139 1561 1560 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4140 1 1555 1554 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4141 1555 1554 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4142 1 1557 1556 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4143 1557 1556 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4144 1 1559 1558 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4145 1559 1558 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4146 1 1561 1560 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4147 1561 1560 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4148 1 1563 1562 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4149 1563 1562 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4150 1 1565 1564 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4151 1565 1564 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4152 1 1567 1566 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4153 1567 1566 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4154 1 1569 1568 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4155 1569 1568 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4156 0 1563 1562 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4157 1563 1562 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4158 0 1565 1564 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4159 1565 1564 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4160 0 1567 1566 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4161 1567 1566 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4162 0 1569 1568 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4163 1569 1568 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4164 222 588 1562 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4165 223 588 1563 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4166 224 588 1564 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4167 225 588 1565 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4168 226 588 1566 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4169 227 588 1567 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4170 228 588 1568 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4171 229 588 1569 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4172 1570 591 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4173 1571 591 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4174 1572 591 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4175 1573 591 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4176 1574 591 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4177 1575 591 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4178 1576 591 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4179 1577 591 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4180 0 1571 1570 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4181 1571 1570 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4182 0 1573 1572 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4183 1573 1572 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4184 0 1575 1574 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4185 1575 1574 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4186 0 1577 1576 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4187 1577 1576 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4188 1 1571 1570 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4189 1571 1570 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4190 1 1573 1572 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4191 1573 1572 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4192 1 1579 1578 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4193 1579 1578 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4194 1 1581 1580 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4195 1581 1580 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4196 1 1575 1574 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4197 1575 1574 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4198 1 1577 1576 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4199 1577 1576 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4200 1 1583 1582 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4201 1583 1582 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4202 1 1585 1584 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4203 1585 1584 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4204 0 1579 1578 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4205 1579 1578 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4206 0 1581 1580 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4207 1581 1580 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4208 0 1583 1582 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4209 1583 1582 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4210 0 1585 1584 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4211 1585 1584 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4212 222 596 1578 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4213 223 596 1579 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4214 224 596 1580 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4215 225 596 1581 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4216 226 596 1582 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4217 227 596 1583 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4218 228 596 1584 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4219 229 596 1585 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4220 1586 600 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4221 1587 600 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4222 1588 600 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4223 1589 600 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4224 1590 600 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4225 1591 600 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4226 1592 600 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4227 1593 600 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4228 0 1587 1586 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4229 1587 1586 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4230 0 1589 1588 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4231 1589 1588 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4232 0 1591 1590 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4233 1591 1590 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4234 0 1593 1592 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4235 1593 1592 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4236 1 1587 1586 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4237 1587 1586 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4238 1 1589 1588 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4239 1589 1588 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4240 1 1591 1590 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4241 1591 1590 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4242 1 1593 1592 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4243 1593 1592 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4244 1 1595 1594 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4245 1595 1594 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4246 1 1597 1596 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4247 1597 1596 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4248 1 1599 1598 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4249 1599 1598 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4250 1 1601 1600 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4251 1601 1600 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4252 0 1595 1594 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4253 1595 1594 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4254 0 1597 1596 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4255 1597 1596 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4256 0 1599 1598 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4257 1599 1598 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4258 0 1601 1600 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4259 1601 1600 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4260 222 604 1594 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4261 223 604 1595 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4262 224 604 1596 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4263 225 604 1597 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4264 226 604 1598 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4265 227 604 1599 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4266 228 604 1600 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4267 229 604 1601 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4268 1602 607 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4269 1603 607 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4270 1604 607 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4271 1605 607 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4272 1606 607 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4273 1607 607 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4274 1608 607 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4275 1609 607 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4276 0 1603 1602 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4277 1603 1602 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4278 0 1605 1604 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4279 1605 1604 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4280 0 1607 1606 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4281 1607 1606 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4282 0 1609 1608 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4283 1609 1608 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4284 1 1603 1602 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4285 1603 1602 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4286 1 1605 1604 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4287 1605 1604 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4288 1 1611 1610 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4289 1611 1610 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4290 1 1613 1612 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4291 1613 1612 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4292 1 1607 1606 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4293 1607 1606 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4294 1 1609 1608 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4295 1609 1608 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4296 1 1615 1614 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4297 1615 1614 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4298 1 1617 1616 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4299 1617 1616 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4300 0 1611 1610 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4301 1611 1610 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4302 0 1613 1612 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4303 1613 1612 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4304 0 1615 1614 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4305 1615 1614 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4306 0 1617 1616 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4307 1617 1616 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4308 222 612 1610 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4309 223 612 1611 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4310 224 612 1612 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4311 225 612 1613 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4312 226 612 1614 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4313 227 612 1615 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4314 228 612 1616 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4315 229 612 1617 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4316 1618 616 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4317 1619 616 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4318 1620 616 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4319 1621 616 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4320 1622 616 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4321 1623 616 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4322 1624 616 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4323 1625 616 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4324 0 1619 1618 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4325 1619 1618 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4326 0 1621 1620 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4327 1621 1620 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4328 0 1623 1622 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4329 1623 1622 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4330 0 1625 1624 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4331 1625 1624 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4332 1 1619 1618 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4333 1619 1618 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4334 1 1621 1620 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4335 1621 1620 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4336 1 1623 1622 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4337 1623 1622 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4338 1 1625 1624 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4339 1625 1624 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4340 1 1627 1626 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4341 1627 1626 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4342 1 1629 1628 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4343 1629 1628 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4344 1 1631 1630 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4345 1631 1630 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4346 1 1633 1632 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4347 1633 1632 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4348 0 1627 1626 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4349 1627 1626 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4350 0 1629 1628 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4351 1629 1628 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4352 0 1631 1630 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4353 1631 1630 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4354 0 1633 1632 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4355 1633 1632 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4356 222 620 1626 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4357 223 620 1627 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4358 224 620 1628 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4359 225 620 1629 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4360 226 620 1630 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4361 227 620 1631 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4362 228 620 1632 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4363 229 620 1633 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4364 1634 624 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4365 1635 624 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4366 1636 624 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4367 1637 624 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4368 1638 624 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4369 1639 624 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4370 1640 624 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4371 1641 624 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4372 0 1635 1634 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4373 1635 1634 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4374 0 1637 1636 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4375 1637 1636 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4376 0 1639 1638 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4377 1639 1638 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4378 0 1641 1640 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4379 1641 1640 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4380 1 1635 1634 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4381 1635 1634 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4382 1 1637 1636 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4383 1637 1636 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4384 1 1643 1642 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4385 1643 1642 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4386 1 1645 1644 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4387 1645 1644 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4388 1 1639 1638 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4389 1639 1638 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4390 1 1641 1640 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4391 1641 1640 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4392 1 1647 1646 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4393 1647 1646 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4394 1 1649 1648 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4395 1649 1648 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4396 0 1643 1642 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4397 1643 1642 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4398 0 1645 1644 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4399 1645 1644 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4400 0 1647 1646 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4401 1647 1646 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4402 0 1649 1648 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4403 1649 1648 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4404 222 628 1642 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4405 223 628 1643 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4406 224 628 1644 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4407 225 628 1645 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4408 226 628 1646 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4409 227 628 1647 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4410 228 628 1648 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4411 229 628 1649 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4412 1650 632 222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4413 1651 632 223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4414 1652 632 224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4415 1653 632 225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4416 1654 632 226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4417 1655 632 227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4418 1656 632 228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4419 1657 632 229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4420 0 1651 1650 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4421 1651 1650 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4422 0 1653 1652 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4423 1653 1652 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4424 0 1655 1654 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4425 1655 1654 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4426 0 1657 1656 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4427 1657 1656 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4428 1 1651 1650 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4429 1651 1650 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4430 1 1653 1652 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4431 1653 1652 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4432 1 1655 1654 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4433 1655 1654 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4434 1 1657 1656 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4435 1657 1656 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4436 1 1659 1658 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4437 1659 1658 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4438 1 1661 1660 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4439 1661 1660 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4440 1 1663 1662 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4441 1663 1662 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4442 1 1665 1664 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4443 1665 1664 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4444 0 1659 1658 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4445 1659 1658 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4446 0 1661 1660 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4447 1661 1660 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4448 0 1663 1662 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4449 1663 1662 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4450 0 1665 1664 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4451 1665 1664 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4452 248 380 1658 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4453 249 380 1659 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4454 250 380 1660 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4455 251 380 1661 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4456 252 380 1662 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4457 253 380 1663 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4458 254 380 1664 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4459 255 380 1665 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4460 1666 383 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4461 1667 383 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4462 1668 383 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4463 1669 383 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4464 1670 383 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4465 1671 383 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4466 1672 383 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4467 1673 383 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4468 0 1667 1666 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4469 1667 1666 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4470 0 1669 1668 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4471 1669 1668 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4472 0 1671 1670 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4473 1671 1670 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4474 0 1673 1672 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4475 1673 1672 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4476 1 1667 1666 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4477 1667 1666 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4478 1 1669 1668 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4479 1669 1668 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4480 1 1675 1674 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4481 1675 1674 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4482 1 1677 1676 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4483 1677 1676 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4484 1 1671 1670 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4485 1671 1670 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4486 1 1673 1672 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4487 1673 1672 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4488 1 1679 1678 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4489 1679 1678 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4490 1 1681 1680 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4491 1681 1680 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4492 0 1675 1674 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4493 1675 1674 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4494 0 1677 1676 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4495 1677 1676 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4496 0 1679 1678 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4497 1679 1678 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4498 0 1681 1680 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4499 1681 1680 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4500 248 388 1674 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4501 249 388 1675 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4502 250 388 1676 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4503 251 388 1677 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4504 252 388 1678 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4505 253 388 1679 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4506 254 388 1680 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4507 255 388 1681 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4508 1682 392 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4509 1683 392 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4510 1684 392 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4511 1685 392 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4512 1686 392 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4513 1687 392 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4514 1688 392 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4515 1689 392 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4516 0 1683 1682 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4517 1683 1682 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4518 0 1685 1684 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4519 1685 1684 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4520 0 1687 1686 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4521 1687 1686 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4522 0 1689 1688 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4523 1689 1688 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4524 1 1683 1682 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4525 1683 1682 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4526 1 1685 1684 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4527 1685 1684 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4528 1 1687 1686 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4529 1687 1686 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4530 1 1689 1688 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4531 1689 1688 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4532 1 1691 1690 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4533 1691 1690 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4534 1 1693 1692 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4535 1693 1692 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4536 1 1695 1694 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4537 1695 1694 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4538 1 1697 1696 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4539 1697 1696 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4540 0 1691 1690 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4541 1691 1690 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4542 0 1693 1692 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4543 1693 1692 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4544 0 1695 1694 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4545 1695 1694 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4546 0 1697 1696 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4547 1697 1696 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4548 248 396 1690 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4549 249 396 1691 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4550 250 396 1692 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4551 251 396 1693 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4552 252 396 1694 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4553 253 396 1695 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4554 254 396 1696 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4555 255 396 1697 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4556 1698 399 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4557 1699 399 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4558 1700 399 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4559 1701 399 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4560 1702 399 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4561 1703 399 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4562 1704 399 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4563 1705 399 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4564 0 1699 1698 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4565 1699 1698 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4566 0 1701 1700 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4567 1701 1700 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4568 0 1703 1702 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4569 1703 1702 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4570 0 1705 1704 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4571 1705 1704 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4572 1 1699 1698 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4573 1699 1698 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4574 1 1701 1700 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4575 1701 1700 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4576 1 1707 1706 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4577 1707 1706 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4578 1 1709 1708 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4579 1709 1708 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4580 1 1703 1702 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4581 1703 1702 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4582 1 1705 1704 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4583 1705 1704 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4584 1 1711 1710 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4585 1711 1710 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4586 1 1713 1712 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4587 1713 1712 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4588 0 1707 1706 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4589 1707 1706 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4590 0 1709 1708 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4591 1709 1708 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4592 0 1711 1710 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4593 1711 1710 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4594 0 1713 1712 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4595 1713 1712 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4596 248 404 1706 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4597 249 404 1707 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4598 250 404 1708 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4599 251 404 1709 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4600 252 404 1710 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4601 253 404 1711 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4602 254 404 1712 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4603 255 404 1713 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4604 1714 408 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4605 1715 408 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4606 1716 408 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4607 1717 408 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4608 1718 408 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4609 1719 408 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4610 1720 408 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4611 1721 408 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4612 0 1715 1714 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4613 1715 1714 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4614 0 1717 1716 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4615 1717 1716 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4616 0 1719 1718 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4617 1719 1718 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4618 0 1721 1720 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4619 1721 1720 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4620 1 1715 1714 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4621 1715 1714 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4622 1 1717 1716 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4623 1717 1716 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4624 1 1719 1718 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4625 1719 1718 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4626 1 1721 1720 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4627 1721 1720 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4628 1 1723 1722 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4629 1723 1722 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4630 1 1725 1724 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4631 1725 1724 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4632 1 1727 1726 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4633 1727 1726 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4634 1 1729 1728 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4635 1729 1728 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4636 0 1723 1722 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4637 1723 1722 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4638 0 1725 1724 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4639 1725 1724 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4640 0 1727 1726 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4641 1727 1726 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4642 0 1729 1728 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4643 1729 1728 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4644 248 412 1722 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4645 249 412 1723 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4646 250 412 1724 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4647 251 412 1725 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4648 252 412 1726 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4649 253 412 1727 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4650 254 412 1728 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4651 255 412 1729 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4652 1730 415 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4653 1731 415 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4654 1732 415 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4655 1733 415 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4656 1734 415 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4657 1735 415 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4658 1736 415 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4659 1737 415 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4660 0 1731 1730 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4661 1731 1730 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4662 0 1733 1732 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4663 1733 1732 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4664 0 1735 1734 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4665 1735 1734 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4666 0 1737 1736 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4667 1737 1736 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4668 1 1731 1730 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4669 1731 1730 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4670 1 1733 1732 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4671 1733 1732 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4672 1 1739 1738 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4673 1739 1738 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4674 1 1741 1740 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4675 1741 1740 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4676 1 1735 1734 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4677 1735 1734 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4678 1 1737 1736 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4679 1737 1736 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4680 1 1743 1742 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4681 1743 1742 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4682 1 1745 1744 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4683 1745 1744 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4684 0 1739 1738 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4685 1739 1738 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4686 0 1741 1740 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4687 1741 1740 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4688 0 1743 1742 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4689 1743 1742 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4690 0 1745 1744 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4691 1745 1744 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4692 248 420 1738 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4693 249 420 1739 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4694 250 420 1740 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4695 251 420 1741 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4696 252 420 1742 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4697 253 420 1743 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4698 254 420 1744 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4699 255 420 1745 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4700 1746 424 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4701 1747 424 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4702 1748 424 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4703 1749 424 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4704 1750 424 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4705 1751 424 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4706 1752 424 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4707 1753 424 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4708 0 1747 1746 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4709 1747 1746 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4710 0 1749 1748 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4711 1749 1748 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4712 0 1751 1750 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4713 1751 1750 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4714 0 1753 1752 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4715 1753 1752 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4716 1 1747 1746 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4717 1747 1746 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4718 1 1749 1748 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4719 1749 1748 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4720 1 1751 1750 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4721 1751 1750 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4722 1 1753 1752 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4723 1753 1752 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4724 1 1755 1754 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4725 1755 1754 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4726 1 1757 1756 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4727 1757 1756 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4728 1 1759 1758 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4729 1759 1758 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4730 1 1761 1760 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4731 1761 1760 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4732 0 1755 1754 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4733 1755 1754 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4734 0 1757 1756 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4735 1757 1756 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4736 0 1759 1758 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4737 1759 1758 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4738 0 1761 1760 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4739 1761 1760 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4740 248 428 1754 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4741 249 428 1755 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4742 250 428 1756 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4743 251 428 1757 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4744 252 428 1758 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4745 253 428 1759 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4746 254 428 1760 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4747 255 428 1761 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4748 1762 431 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4749 1763 431 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4750 1764 431 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4751 1765 431 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4752 1766 431 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4753 1767 431 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4754 1768 431 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4755 1769 431 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4756 0 1763 1762 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4757 1763 1762 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4758 0 1765 1764 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4759 1765 1764 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4760 0 1767 1766 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4761 1767 1766 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4762 0 1769 1768 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4763 1769 1768 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4764 1 1763 1762 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4765 1763 1762 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4766 1 1765 1764 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4767 1765 1764 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4768 1 1771 1770 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4769 1771 1770 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4770 1 1773 1772 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4771 1773 1772 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4772 1 1767 1766 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4773 1767 1766 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4774 1 1769 1768 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4775 1769 1768 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4776 1 1775 1774 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4777 1775 1774 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4778 1 1777 1776 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4779 1777 1776 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4780 0 1771 1770 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4781 1771 1770 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4782 0 1773 1772 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4783 1773 1772 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4784 0 1775 1774 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4785 1775 1774 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4786 0 1777 1776 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4787 1777 1776 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4788 248 436 1770 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4789 249 436 1771 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4790 250 436 1772 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4791 251 436 1773 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4792 252 436 1774 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4793 253 436 1775 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4794 254 436 1776 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4795 255 436 1777 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4796 1778 440 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4797 1779 440 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4798 1780 440 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4799 1781 440 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4800 1782 440 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4801 1783 440 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4802 1784 440 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4803 1785 440 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4804 0 1779 1778 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4805 1779 1778 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4806 0 1781 1780 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4807 1781 1780 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4808 0 1783 1782 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4809 1783 1782 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4810 0 1785 1784 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4811 1785 1784 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4812 1 1779 1778 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4813 1779 1778 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4814 1 1781 1780 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4815 1781 1780 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4816 1 1783 1782 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4817 1783 1782 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4818 1 1785 1784 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4819 1785 1784 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4820 1 1787 1786 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4821 1787 1786 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4822 1 1789 1788 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4823 1789 1788 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4824 1 1791 1790 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4825 1791 1790 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4826 1 1793 1792 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4827 1793 1792 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4828 0 1787 1786 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4829 1787 1786 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4830 0 1789 1788 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4831 1789 1788 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4832 0 1791 1790 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4833 1791 1790 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4834 0 1793 1792 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4835 1793 1792 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4836 248 444 1786 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4837 249 444 1787 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4838 250 444 1788 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4839 251 444 1789 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4840 252 444 1790 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4841 253 444 1791 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4842 254 444 1792 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4843 255 444 1793 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4844 1794 447 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4845 1795 447 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4846 1796 447 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4847 1797 447 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4848 1798 447 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4849 1799 447 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4850 1800 447 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4851 1801 447 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4852 0 1795 1794 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4853 1795 1794 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4854 0 1797 1796 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4855 1797 1796 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4856 0 1799 1798 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4857 1799 1798 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4858 0 1801 1800 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4859 1801 1800 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4860 1 1795 1794 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4861 1795 1794 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4862 1 1797 1796 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4863 1797 1796 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4864 1 1803 1802 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4865 1803 1802 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4866 1 1805 1804 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4867 1805 1804 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4868 1 1799 1798 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4869 1799 1798 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4870 1 1801 1800 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4871 1801 1800 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4872 1 1807 1806 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4873 1807 1806 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4874 1 1809 1808 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4875 1809 1808 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4876 0 1803 1802 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4877 1803 1802 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4878 0 1805 1804 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4879 1805 1804 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4880 0 1807 1806 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4881 1807 1806 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4882 0 1809 1808 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4883 1809 1808 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4884 248 452 1802 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4885 249 452 1803 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4886 250 452 1804 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4887 251 452 1805 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4888 252 452 1806 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4889 253 452 1807 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4890 254 452 1808 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4891 255 452 1809 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4892 1810 456 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4893 1811 456 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4894 1812 456 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4895 1813 456 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4896 1814 456 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4897 1815 456 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4898 1816 456 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4899 1817 456 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4900 0 1811 1810 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4901 1811 1810 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4902 0 1813 1812 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4903 1813 1812 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4904 0 1815 1814 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4905 1815 1814 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4906 0 1817 1816 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4907 1817 1816 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4908 1 1811 1810 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4909 1811 1810 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4910 1 1813 1812 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4911 1813 1812 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4912 1 1815 1814 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4913 1815 1814 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4914 1 1817 1816 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4915 1817 1816 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4916 1 1819 1818 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4917 1819 1818 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4918 1 1821 1820 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4919 1821 1820 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4920 1 1823 1822 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4921 1823 1822 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4922 1 1825 1824 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4923 1825 1824 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4924 0 1819 1818 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4925 1819 1818 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4926 0 1821 1820 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4927 1821 1820 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4928 0 1823 1822 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4929 1823 1822 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4930 0 1825 1824 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4931 1825 1824 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4932 248 460 1818 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4933 249 460 1819 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4934 250 460 1820 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4935 251 460 1821 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4936 252 460 1822 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4937 253 460 1823 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4938 254 460 1824 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4939 255 460 1825 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4940 1826 463 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4941 1827 463 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4942 1828 463 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4943 1829 463 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4944 1830 463 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4945 1831 463 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4946 1832 463 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4947 1833 463 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4948 0 1827 1826 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4949 1827 1826 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4950 0 1829 1828 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4951 1829 1828 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4952 0 1831 1830 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4953 1831 1830 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4954 0 1833 1832 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4955 1833 1832 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4956 1 1827 1826 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4957 1827 1826 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4958 1 1829 1828 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4959 1829 1828 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4960 1 1835 1834 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4961 1835 1834 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m4962 1 1837 1836 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4963 1837 1836 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4964 1 1831 1830 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4965 1831 1830 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4966 1 1833 1832 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4967 1833 1832 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4968 1 1839 1838 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m4969 1839 1838 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4970 1 1841 1840 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m4971 1841 1840 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m4972 0 1835 1834 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4973 1835 1834 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4974 0 1837 1836 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4975 1837 1836 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4976 0 1839 1838 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4977 1839 1838 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4978 0 1841 1840 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m4979 1841 1840 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m4980 248 468 1834 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m4981 249 468 1835 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4982 250 468 1836 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4983 251 468 1837 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4984 252 468 1838 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m4985 253 468 1839 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m4986 254 468 1840 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m4987 255 468 1841 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m4988 1842 472 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m4989 1843 472 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4990 1844 472 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4991 1845 472 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4992 1846 472 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m4993 1847 472 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m4994 1848 472 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m4995 1849 472 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m4996 0 1843 1842 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4997 1843 1842 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m4998 0 1845 1844 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m4999 1845 1844 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5000 0 1847 1846 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5001 1847 1846 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5002 0 1849 1848 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5003 1849 1848 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5004 1 1843 1842 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5005 1843 1842 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5006 1 1845 1844 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5007 1845 1844 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5008 1 1847 1846 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5009 1847 1846 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5010 1 1849 1848 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5011 1849 1848 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5012 1 1851 1850 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5013 1851 1850 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5014 1 1853 1852 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5015 1853 1852 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5016 1 1855 1854 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5017 1855 1854 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5018 1 1857 1856 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5019 1857 1856 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5020 0 1851 1850 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5021 1851 1850 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5022 0 1853 1852 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5023 1853 1852 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5024 0 1855 1854 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5025 1855 1854 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5026 0 1857 1856 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5027 1857 1856 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5028 248 476 1850 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5029 249 476 1851 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5030 250 476 1852 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5031 251 476 1853 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5032 252 476 1854 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5033 253 476 1855 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5034 254 476 1856 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5035 255 476 1857 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5036 1858 479 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5037 1859 479 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5038 1860 479 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5039 1861 479 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5040 1862 479 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5041 1863 479 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5042 1864 479 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5043 1865 479 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5044 0 1859 1858 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5045 1859 1858 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5046 0 1861 1860 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5047 1861 1860 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5048 0 1863 1862 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5049 1863 1862 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5050 0 1865 1864 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5051 1865 1864 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5052 1 1859 1858 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5053 1859 1858 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5054 1 1861 1860 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5055 1861 1860 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5056 1 1867 1866 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5057 1867 1866 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5058 1 1869 1868 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5059 1869 1868 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5060 1 1863 1862 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5061 1863 1862 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5062 1 1865 1864 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5063 1865 1864 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5064 1 1871 1870 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5065 1871 1870 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5066 1 1873 1872 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5067 1873 1872 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5068 0 1867 1866 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5069 1867 1866 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5070 0 1869 1868 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5071 1869 1868 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5072 0 1871 1870 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5073 1871 1870 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5074 0 1873 1872 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5075 1873 1872 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5076 248 484 1866 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5077 249 484 1867 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5078 250 484 1868 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5079 251 484 1869 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5080 252 484 1870 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5081 253 484 1871 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5082 254 484 1872 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5083 255 484 1873 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5084 1874 488 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5085 1875 488 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5086 1876 488 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5087 1877 488 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5088 1878 488 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5089 1879 488 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5090 1880 488 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5091 1881 488 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5092 0 1875 1874 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5093 1875 1874 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5094 0 1877 1876 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5095 1877 1876 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5096 0 1879 1878 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5097 1879 1878 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5098 0 1881 1880 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5099 1881 1880 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5100 1 1875 1874 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5101 1875 1874 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5102 1 1877 1876 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5103 1877 1876 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5104 1 1879 1878 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5105 1879 1878 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5106 1 1881 1880 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5107 1881 1880 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5108 1 1883 1882 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5109 1883 1882 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5110 1 1885 1884 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5111 1885 1884 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5112 1 1887 1886 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5113 1887 1886 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5114 1 1889 1888 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5115 1889 1888 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5116 0 1883 1882 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5117 1883 1882 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5118 0 1885 1884 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5119 1885 1884 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5120 0 1887 1886 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5121 1887 1886 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5122 0 1889 1888 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5123 1889 1888 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5124 248 492 1882 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5125 249 492 1883 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5126 250 492 1884 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5127 251 492 1885 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5128 252 492 1886 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5129 253 492 1887 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5130 254 492 1888 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5131 255 492 1889 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5132 1890 495 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5133 1891 495 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5134 1892 495 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5135 1893 495 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5136 1894 495 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5137 1895 495 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5138 1896 495 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5139 1897 495 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5140 0 1891 1890 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5141 1891 1890 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5142 0 1893 1892 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5143 1893 1892 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5144 0 1895 1894 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5145 1895 1894 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5146 0 1897 1896 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5147 1897 1896 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5148 1 1891 1890 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5149 1891 1890 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5150 1 1893 1892 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5151 1893 1892 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5152 1 1899 1898 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5153 1899 1898 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5154 1 1901 1900 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5155 1901 1900 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5156 1 1895 1894 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5157 1895 1894 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5158 1 1897 1896 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5159 1897 1896 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5160 1 1903 1902 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5161 1903 1902 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5162 1 1905 1904 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5163 1905 1904 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5164 0 1899 1898 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5165 1899 1898 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5166 0 1901 1900 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5167 1901 1900 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5168 0 1903 1902 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5169 1903 1902 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5170 0 1905 1904 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5171 1905 1904 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5172 248 500 1898 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5173 249 500 1899 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5174 250 500 1900 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5175 251 500 1901 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5176 252 500 1902 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5177 253 500 1903 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5178 254 500 1904 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5179 255 500 1905 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5180 1906 504 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5181 1907 504 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5182 1908 504 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5183 1909 504 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5184 1910 504 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5185 1911 504 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5186 1912 504 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5187 1913 504 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5188 0 1907 1906 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5189 1907 1906 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5190 0 1909 1908 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5191 1909 1908 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5192 0 1911 1910 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5193 1911 1910 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5194 0 1913 1912 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5195 1913 1912 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5196 1 1907 1906 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5197 1907 1906 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5198 1 1909 1908 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5199 1909 1908 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5200 1 1911 1910 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5201 1911 1910 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5202 1 1913 1912 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5203 1913 1912 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5204 1 1915 1914 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5205 1915 1914 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5206 1 1917 1916 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5207 1917 1916 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5208 1 1919 1918 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5209 1919 1918 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5210 1 1921 1920 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5211 1921 1920 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5212 0 1915 1914 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5213 1915 1914 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5214 0 1917 1916 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5215 1917 1916 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5216 0 1919 1918 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5217 1919 1918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5218 0 1921 1920 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5219 1921 1920 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5220 248 508 1914 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5221 249 508 1915 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5222 250 508 1916 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5223 251 508 1917 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5224 252 508 1918 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5225 253 508 1919 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5226 254 508 1920 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5227 255 508 1921 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5228 1922 511 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5229 1923 511 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5230 1924 511 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5231 1925 511 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5232 1926 511 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5233 1927 511 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5234 1928 511 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5235 1929 511 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5236 0 1923 1922 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5237 1923 1922 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5238 0 1925 1924 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5239 1925 1924 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5240 0 1927 1926 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5241 1927 1926 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5242 0 1929 1928 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5243 1929 1928 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5244 1 1923 1922 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5245 1923 1922 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5246 1 1925 1924 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5247 1925 1924 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5248 1 1931 1930 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5249 1931 1930 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5250 1 1933 1932 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5251 1933 1932 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5252 1 1927 1926 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5253 1927 1926 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5254 1 1929 1928 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5255 1929 1928 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5256 1 1935 1934 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5257 1935 1934 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5258 1 1937 1936 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5259 1937 1936 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5260 0 1931 1930 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5261 1931 1930 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5262 0 1933 1932 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5263 1933 1932 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5264 0 1935 1934 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5265 1935 1934 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5266 0 1937 1936 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5267 1937 1936 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5268 248 516 1930 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5269 249 516 1931 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5270 250 516 1932 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5271 251 516 1933 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5272 252 516 1934 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5273 253 516 1935 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5274 254 516 1936 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5275 255 516 1937 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5276 1938 520 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5277 1939 520 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5278 1940 520 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5279 1941 520 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5280 1942 520 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5281 1943 520 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5282 1944 520 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5283 1945 520 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5284 0 1939 1938 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5285 1939 1938 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5286 0 1941 1940 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5287 1941 1940 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5288 0 1943 1942 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5289 1943 1942 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5290 0 1945 1944 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5291 1945 1944 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5292 1 1939 1938 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5293 1939 1938 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5294 1 1941 1940 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5295 1941 1940 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5296 1 1943 1942 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5297 1943 1942 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5298 1 1945 1944 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5299 1945 1944 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5300 1 1947 1946 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5301 1947 1946 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5302 1 1949 1948 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5303 1949 1948 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5304 1 1951 1950 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5305 1951 1950 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5306 1 1953 1952 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5307 1953 1952 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5308 0 1947 1946 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5309 1947 1946 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5310 0 1949 1948 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5311 1949 1948 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5312 0 1951 1950 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5313 1951 1950 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5314 0 1953 1952 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5315 1953 1952 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5316 248 524 1946 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5317 249 524 1947 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5318 250 524 1948 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5319 251 524 1949 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5320 252 524 1950 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5321 253 524 1951 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5322 254 524 1952 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5323 255 524 1953 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5324 1954 527 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5325 1955 527 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5326 1956 527 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5327 1957 527 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5328 1958 527 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5329 1959 527 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5330 1960 527 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5331 1961 527 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5332 0 1955 1954 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5333 1955 1954 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5334 0 1957 1956 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5335 1957 1956 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5336 0 1959 1958 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5337 1959 1958 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5338 0 1961 1960 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5339 1961 1960 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5340 1 1955 1954 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5341 1955 1954 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5342 1 1957 1956 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5343 1957 1956 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5344 1 1963 1962 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5345 1963 1962 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5346 1 1965 1964 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5347 1965 1964 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5348 1 1959 1958 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5349 1959 1958 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5350 1 1961 1960 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5351 1961 1960 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5352 1 1967 1966 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5353 1967 1966 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5354 1 1969 1968 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5355 1969 1968 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5356 0 1963 1962 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5357 1963 1962 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5358 0 1965 1964 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5359 1965 1964 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5360 0 1967 1966 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5361 1967 1966 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5362 0 1969 1968 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5363 1969 1968 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5364 248 532 1962 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5365 249 532 1963 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5366 250 532 1964 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5367 251 532 1965 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5368 252 532 1966 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5369 253 532 1967 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5370 254 532 1968 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5371 255 532 1969 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5372 1970 536 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5373 1971 536 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5374 1972 536 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5375 1973 536 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5376 1974 536 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5377 1975 536 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5378 1976 536 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5379 1977 536 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5380 0 1971 1970 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5381 1971 1970 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5382 0 1973 1972 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5383 1973 1972 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5384 0 1975 1974 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5385 1975 1974 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5386 0 1977 1976 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5387 1977 1976 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5388 1 1971 1970 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5389 1971 1970 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5390 1 1973 1972 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5391 1973 1972 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5392 1 1975 1974 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5393 1975 1974 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5394 1 1977 1976 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5395 1977 1976 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5396 1 1979 1978 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5397 1979 1978 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5398 1 1981 1980 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5399 1981 1980 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5400 1 1983 1982 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5401 1983 1982 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5402 1 1985 1984 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5403 1985 1984 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5404 0 1979 1978 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5405 1979 1978 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5406 0 1981 1980 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5407 1981 1980 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5408 0 1983 1982 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5409 1983 1982 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5410 0 1985 1984 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5411 1985 1984 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5412 248 540 1978 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5413 249 540 1979 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5414 250 540 1980 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5415 251 540 1981 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5416 252 540 1982 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5417 253 540 1983 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5418 254 540 1984 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5419 255 540 1985 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5420 1986 543 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5421 1987 543 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5422 1988 543 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5423 1989 543 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5424 1990 543 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5425 1991 543 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5426 1992 543 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5427 1993 543 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5428 0 1987 1986 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5429 1987 1986 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5430 0 1989 1988 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5431 1989 1988 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5432 0 1991 1990 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5433 1991 1990 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5434 0 1993 1992 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5435 1993 1992 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5436 1 1987 1986 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5437 1987 1986 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5438 1 1989 1988 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5439 1989 1988 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5440 1 1995 1994 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5441 1995 1994 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5442 1 1997 1996 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5443 1997 1996 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5444 1 1991 1990 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5445 1991 1990 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5446 1 1993 1992 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5447 1993 1992 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5448 1 1999 1998 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5449 1999 1998 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5450 1 2001 2000 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5451 2001 2000 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5452 0 1995 1994 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5453 1995 1994 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5454 0 1997 1996 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5455 1997 1996 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5456 0 1999 1998 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5457 1999 1998 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5458 0 2001 2000 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5459 2001 2000 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5460 248 548 1994 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5461 249 548 1995 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5462 250 548 1996 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5463 251 548 1997 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5464 252 548 1998 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5465 253 548 1999 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5466 254 548 2000 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5467 255 548 2001 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5468 2002 552 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5469 2003 552 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5470 2004 552 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5471 2005 552 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5472 2006 552 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5473 2007 552 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5474 2008 552 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5475 2009 552 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5476 0 2003 2002 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5477 2003 2002 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5478 0 2005 2004 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5479 2005 2004 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5480 0 2007 2006 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5481 2007 2006 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5482 0 2009 2008 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5483 2009 2008 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5484 1 2003 2002 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5485 2003 2002 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5486 1 2005 2004 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5487 2005 2004 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5488 1 2007 2006 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5489 2007 2006 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5490 1 2009 2008 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5491 2009 2008 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5492 1 2011 2010 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5493 2011 2010 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5494 1 2013 2012 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5495 2013 2012 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5496 1 2015 2014 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5497 2015 2014 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5498 1 2017 2016 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5499 2017 2016 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5500 0 2011 2010 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5501 2011 2010 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5502 0 2013 2012 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5503 2013 2012 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5504 0 2015 2014 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5505 2015 2014 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5506 0 2017 2016 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5507 2017 2016 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5508 248 556 2010 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5509 249 556 2011 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5510 250 556 2012 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5511 251 556 2013 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5512 252 556 2014 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5513 253 556 2015 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5514 254 556 2016 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5515 255 556 2017 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5516 2018 559 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5517 2019 559 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5518 2020 559 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5519 2021 559 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5520 2022 559 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5521 2023 559 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5522 2024 559 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5523 2025 559 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5524 0 2019 2018 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5525 2019 2018 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5526 0 2021 2020 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5527 2021 2020 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5528 0 2023 2022 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5529 2023 2022 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5530 0 2025 2024 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5531 2025 2024 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5532 1 2019 2018 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5533 2019 2018 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5534 1 2021 2020 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5535 2021 2020 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5536 1 2027 2026 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5537 2027 2026 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5538 1 2029 2028 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5539 2029 2028 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5540 1 2023 2022 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5541 2023 2022 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5542 1 2025 2024 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5543 2025 2024 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5544 1 2031 2030 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5545 2031 2030 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5546 1 2033 2032 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5547 2033 2032 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5548 0 2027 2026 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5549 2027 2026 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5550 0 2029 2028 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5551 2029 2028 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5552 0 2031 2030 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5553 2031 2030 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5554 0 2033 2032 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5555 2033 2032 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5556 248 564 2026 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5557 249 564 2027 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5558 250 564 2028 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5559 251 564 2029 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5560 252 564 2030 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5561 253 564 2031 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5562 254 564 2032 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5563 255 564 2033 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5564 2034 568 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5565 2035 568 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5566 2036 568 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5567 2037 568 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5568 2038 568 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5569 2039 568 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5570 2040 568 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5571 2041 568 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5572 0 2035 2034 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5573 2035 2034 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5574 0 2037 2036 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5575 2037 2036 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5576 0 2039 2038 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5577 2039 2038 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5578 0 2041 2040 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5579 2041 2040 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5580 1 2035 2034 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5581 2035 2034 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5582 1 2037 2036 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5583 2037 2036 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5584 1 2039 2038 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5585 2039 2038 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5586 1 2041 2040 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5587 2041 2040 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5588 1 2043 2042 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5589 2043 2042 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5590 1 2045 2044 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5591 2045 2044 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5592 1 2047 2046 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5593 2047 2046 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5594 1 2049 2048 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5595 2049 2048 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5596 0 2043 2042 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5597 2043 2042 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5598 0 2045 2044 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5599 2045 2044 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5600 0 2047 2046 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5601 2047 2046 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5602 0 2049 2048 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5603 2049 2048 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5604 248 572 2042 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5605 249 572 2043 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5606 250 572 2044 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5607 251 572 2045 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5608 252 572 2046 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5609 253 572 2047 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5610 254 572 2048 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5611 255 572 2049 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5612 2050 575 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5613 2051 575 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5614 2052 575 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5615 2053 575 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5616 2054 575 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5617 2055 575 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5618 2056 575 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5619 2057 575 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5620 0 2051 2050 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5621 2051 2050 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5622 0 2053 2052 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5623 2053 2052 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5624 0 2055 2054 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5625 2055 2054 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5626 0 2057 2056 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5627 2057 2056 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5628 1 2051 2050 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5629 2051 2050 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5630 1 2053 2052 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5631 2053 2052 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5632 1 2059 2058 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5633 2059 2058 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5634 1 2061 2060 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5635 2061 2060 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5636 1 2055 2054 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5637 2055 2054 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5638 1 2057 2056 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5639 2057 2056 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5640 1 2063 2062 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5641 2063 2062 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5642 1 2065 2064 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5643 2065 2064 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5644 0 2059 2058 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5645 2059 2058 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5646 0 2061 2060 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5647 2061 2060 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5648 0 2063 2062 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5649 2063 2062 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5650 0 2065 2064 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5651 2065 2064 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5652 248 580 2058 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5653 249 580 2059 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5654 250 580 2060 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5655 251 580 2061 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5656 252 580 2062 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5657 253 580 2063 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5658 254 580 2064 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5659 255 580 2065 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5660 2066 584 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5661 2067 584 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5662 2068 584 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5663 2069 584 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5664 2070 584 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5665 2071 584 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5666 2072 584 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5667 2073 584 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5668 0 2067 2066 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5669 2067 2066 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5670 0 2069 2068 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5671 2069 2068 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5672 0 2071 2070 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5673 2071 2070 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5674 0 2073 2072 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5675 2073 2072 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5676 1 2067 2066 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5677 2067 2066 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5678 1 2069 2068 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5679 2069 2068 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5680 1 2071 2070 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5681 2071 2070 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5682 1 2073 2072 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5683 2073 2072 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5684 1 2075 2074 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5685 2075 2074 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5686 1 2077 2076 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5687 2077 2076 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5688 1 2079 2078 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5689 2079 2078 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5690 1 2081 2080 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5691 2081 2080 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5692 0 2075 2074 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5693 2075 2074 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5694 0 2077 2076 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5695 2077 2076 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5696 0 2079 2078 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5697 2079 2078 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5698 0 2081 2080 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5699 2081 2080 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5700 248 588 2074 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5701 249 588 2075 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5702 250 588 2076 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5703 251 588 2077 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5704 252 588 2078 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5705 253 588 2079 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5706 254 588 2080 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5707 255 588 2081 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5708 2082 591 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5709 2083 591 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5710 2084 591 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5711 2085 591 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5712 2086 591 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5713 2087 591 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5714 2088 591 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5715 2089 591 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5716 0 2083 2082 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5717 2083 2082 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5718 0 2085 2084 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5719 2085 2084 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5720 0 2087 2086 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5721 2087 2086 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5722 0 2089 2088 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5723 2089 2088 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5724 1 2083 2082 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5725 2083 2082 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5726 1 2085 2084 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5727 2085 2084 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5728 1 2091 2090 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5729 2091 2090 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5730 1 2093 2092 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5731 2093 2092 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5732 1 2087 2086 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5733 2087 2086 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5734 1 2089 2088 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5735 2089 2088 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5736 1 2095 2094 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5737 2095 2094 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5738 1 2097 2096 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5739 2097 2096 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5740 0 2091 2090 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5741 2091 2090 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5742 0 2093 2092 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5743 2093 2092 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5744 0 2095 2094 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5745 2095 2094 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5746 0 2097 2096 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5747 2097 2096 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5748 248 596 2090 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5749 249 596 2091 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5750 250 596 2092 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5751 251 596 2093 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5752 252 596 2094 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5753 253 596 2095 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5754 254 596 2096 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5755 255 596 2097 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5756 2098 600 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5757 2099 600 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5758 2100 600 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5759 2101 600 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5760 2102 600 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5761 2103 600 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5762 2104 600 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5763 2105 600 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5764 0 2099 2098 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5765 2099 2098 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5766 0 2101 2100 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5767 2101 2100 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5768 0 2103 2102 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5769 2103 2102 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5770 0 2105 2104 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5771 2105 2104 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5772 1 2099 2098 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5773 2099 2098 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5774 1 2101 2100 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5775 2101 2100 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5776 1 2103 2102 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5777 2103 2102 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5778 1 2105 2104 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5779 2105 2104 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5780 1 2107 2106 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5781 2107 2106 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5782 1 2109 2108 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5783 2109 2108 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5784 1 2111 2110 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5785 2111 2110 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5786 1 2113 2112 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5787 2113 2112 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5788 0 2107 2106 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5789 2107 2106 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5790 0 2109 2108 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5791 2109 2108 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5792 0 2111 2110 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5793 2111 2110 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5794 0 2113 2112 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5795 2113 2112 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5796 248 604 2106 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5797 249 604 2107 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5798 250 604 2108 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5799 251 604 2109 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5800 252 604 2110 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5801 253 604 2111 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5802 254 604 2112 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5803 255 604 2113 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5804 2114 607 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5805 2115 607 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5806 2116 607 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5807 2117 607 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5808 2118 607 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5809 2119 607 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5810 2120 607 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5811 2121 607 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5812 0 2115 2114 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5813 2115 2114 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5814 0 2117 2116 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5815 2117 2116 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5816 0 2119 2118 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5817 2119 2118 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5818 0 2121 2120 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5819 2121 2120 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5820 1 2115 2114 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5821 2115 2114 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5822 1 2117 2116 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5823 2117 2116 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5824 1 2123 2122 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5825 2123 2122 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5826 1 2125 2124 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5827 2125 2124 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5828 1 2119 2118 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5829 2119 2118 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5830 1 2121 2120 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5831 2121 2120 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5832 1 2127 2126 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5833 2127 2126 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5834 1 2129 2128 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5835 2129 2128 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5836 0 2123 2122 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5837 2123 2122 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5838 0 2125 2124 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5839 2125 2124 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5840 0 2127 2126 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5841 2127 2126 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5842 0 2129 2128 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5843 2129 2128 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5844 248 612 2122 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5845 249 612 2123 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5846 250 612 2124 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5847 251 612 2125 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5848 252 612 2126 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5849 253 612 2127 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5850 254 612 2128 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5851 255 612 2129 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5852 2130 616 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5853 2131 616 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5854 2132 616 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5855 2133 616 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5856 2134 616 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5857 2135 616 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5858 2136 616 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5859 2137 616 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5860 0 2131 2130 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5861 2131 2130 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5862 0 2133 2132 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5863 2133 2132 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5864 0 2135 2134 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5865 2135 2134 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5866 0 2137 2136 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5867 2137 2136 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5868 1 2131 2130 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5869 2131 2130 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5870 1 2133 2132 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5871 2133 2132 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5872 1 2135 2134 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5873 2135 2134 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5874 1 2137 2136 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5875 2137 2136 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5876 1 2139 2138 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5877 2139 2138 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5878 1 2141 2140 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5879 2141 2140 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5880 1 2143 2142 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5881 2143 2142 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5882 1 2145 2144 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5883 2145 2144 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5884 0 2139 2138 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5885 2139 2138 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5886 0 2141 2140 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5887 2141 2140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5888 0 2143 2142 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5889 2143 2142 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5890 0 2145 2144 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5891 2145 2144 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5892 248 620 2138 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5893 249 620 2139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5894 250 620 2140 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5895 251 620 2141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5896 252 620 2142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5897 253 620 2143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5898 254 620 2144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5899 255 620 2145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5900 2146 624 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5901 2147 624 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5902 2148 624 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5903 2149 624 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5904 2150 624 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5905 2151 624 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5906 2152 624 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5907 2153 624 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5908 0 2147 2146 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5909 2147 2146 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5910 0 2149 2148 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5911 2149 2148 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5912 0 2151 2150 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5913 2151 2150 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5914 0 2153 2152 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5915 2153 2152 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5916 1 2147 2146 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5917 2147 2146 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5918 1 2149 2148 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5919 2149 2148 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5920 1 2155 2154 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5921 2155 2154 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5922 1 2157 2156 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5923 2157 2156 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5924 1 2151 2150 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5925 2151 2150 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5926 1 2153 2152 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5927 2153 2152 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5928 1 2159 2158 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5929 2159 2158 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5930 1 2161 2160 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5931 2161 2160 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5932 0 2155 2154 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5933 2155 2154 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5934 0 2157 2156 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5935 2157 2156 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5936 0 2159 2158 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5937 2159 2158 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5938 0 2161 2160 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5939 2161 2160 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5940 248 628 2154 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5941 249 628 2155 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5942 250 628 2156 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5943 251 628 2157 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5944 252 628 2158 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5945 253 628 2159 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5946 254 628 2160 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5947 255 628 2161 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5948 2162 632 248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5949 2163 632 249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5950 2164 632 250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5951 2165 632 251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5952 2166 632 252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m5953 2167 632 253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5954 2168 632 254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5955 2169 632 255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m5956 0 2163 2162 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5957 2163 2162 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5958 0 2165 2164 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5959 2165 2164 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5960 0 2167 2166 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5961 2167 2166 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5962 0 2169 2168 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5963 2169 2168 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5964 1 2163 2162 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5965 2163 2162 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5966 1 2165 2164 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5967 2165 2164 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5968 1 2167 2166 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5969 2167 2166 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5970 1 2169 2168 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5971 2169 2168 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5972 1 2171 2170 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5973 2171 2170 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m5974 1 2173 2172 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5975 2173 2172 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5976 1 2175 2174 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m5977 2175 2174 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5978 1 2177 2176 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m5979 2177 2176 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m5980 0 2171 2170 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5981 2171 2170 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5982 0 2173 2172 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m5983 2173 2172 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m5984 0 2175 2174 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5985 2175 2174 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5986 0 2177 2176 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m5987 2177 2176 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m5988 274 380 2170 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m5989 275 380 2171 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5990 276 380 2172 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5991 277 380 2173 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5992 278 380 2174 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m5993 279 380 2175 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m5994 280 380 2176 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m5995 281 380 2177 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m5996 2178 383 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m5997 2179 383 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m5998 2180 383 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m5999 2181 383 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6000 2182 383 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6001 2183 383 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6002 2184 383 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6003 2185 383 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6004 0 2179 2178 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6005 2179 2178 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6006 0 2181 2180 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6007 2181 2180 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6008 0 2183 2182 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6009 2183 2182 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6010 0 2185 2184 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6011 2185 2184 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6012 1 2179 2178 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6013 2179 2178 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6014 1 2181 2180 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6015 2181 2180 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6016 1 2187 2186 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6017 2187 2186 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6018 1 2189 2188 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6019 2189 2188 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6020 1 2183 2182 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6021 2183 2182 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6022 1 2185 2184 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6023 2185 2184 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6024 1 2191 2190 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6025 2191 2190 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6026 1 2193 2192 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6027 2193 2192 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6028 0 2187 2186 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6029 2187 2186 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6030 0 2189 2188 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6031 2189 2188 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6032 0 2191 2190 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6033 2191 2190 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6034 0 2193 2192 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6035 2193 2192 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6036 274 388 2186 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6037 275 388 2187 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6038 276 388 2188 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6039 277 388 2189 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6040 278 388 2190 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6041 279 388 2191 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6042 280 388 2192 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6043 281 388 2193 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6044 2194 392 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6045 2195 392 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6046 2196 392 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6047 2197 392 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6048 2198 392 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6049 2199 392 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6050 2200 392 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6051 2201 392 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6052 0 2195 2194 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6053 2195 2194 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6054 0 2197 2196 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6055 2197 2196 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6056 0 2199 2198 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6057 2199 2198 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6058 0 2201 2200 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6059 2201 2200 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6060 1 2195 2194 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6061 2195 2194 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6062 1 2197 2196 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6063 2197 2196 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6064 1 2199 2198 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6065 2199 2198 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6066 1 2201 2200 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6067 2201 2200 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6068 1 2203 2202 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6069 2203 2202 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6070 1 2205 2204 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6071 2205 2204 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6072 1 2207 2206 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6073 2207 2206 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6074 1 2209 2208 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6075 2209 2208 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6076 0 2203 2202 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6077 2203 2202 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6078 0 2205 2204 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6079 2205 2204 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6080 0 2207 2206 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6081 2207 2206 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6082 0 2209 2208 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6083 2209 2208 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6084 274 396 2202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6085 275 396 2203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6086 276 396 2204 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6087 277 396 2205 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6088 278 396 2206 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6089 279 396 2207 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6090 280 396 2208 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6091 281 396 2209 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6092 2210 399 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6093 2211 399 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6094 2212 399 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6095 2213 399 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6096 2214 399 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6097 2215 399 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6098 2216 399 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6099 2217 399 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6100 0 2211 2210 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6101 2211 2210 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6102 0 2213 2212 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6103 2213 2212 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6104 0 2215 2214 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6105 2215 2214 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6106 0 2217 2216 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6107 2217 2216 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6108 1 2211 2210 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6109 2211 2210 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6110 1 2213 2212 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6111 2213 2212 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6112 1 2219 2218 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6113 2219 2218 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6114 1 2221 2220 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6115 2221 2220 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6116 1 2215 2214 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6117 2215 2214 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6118 1 2217 2216 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6119 2217 2216 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6120 1 2223 2222 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6121 2223 2222 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6122 1 2225 2224 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6123 2225 2224 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6124 0 2219 2218 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6125 2219 2218 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6126 0 2221 2220 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6127 2221 2220 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6128 0 2223 2222 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6129 2223 2222 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6130 0 2225 2224 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6131 2225 2224 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6132 274 404 2218 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6133 275 404 2219 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6134 276 404 2220 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6135 277 404 2221 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6136 278 404 2222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6137 279 404 2223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6138 280 404 2224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6139 281 404 2225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6140 2226 408 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6141 2227 408 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6142 2228 408 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6143 2229 408 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6144 2230 408 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6145 2231 408 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6146 2232 408 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6147 2233 408 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6148 0 2227 2226 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6149 2227 2226 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6150 0 2229 2228 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6151 2229 2228 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6152 0 2231 2230 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6153 2231 2230 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6154 0 2233 2232 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6155 2233 2232 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6156 1 2227 2226 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6157 2227 2226 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6158 1 2229 2228 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6159 2229 2228 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6160 1 2231 2230 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6161 2231 2230 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6162 1 2233 2232 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6163 2233 2232 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6164 1 2235 2234 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6165 2235 2234 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6166 1 2237 2236 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6167 2237 2236 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6168 1 2239 2238 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6169 2239 2238 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6170 1 2241 2240 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6171 2241 2240 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6172 0 2235 2234 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6173 2235 2234 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6174 0 2237 2236 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6175 2237 2236 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6176 0 2239 2238 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6177 2239 2238 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6178 0 2241 2240 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6179 2241 2240 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6180 274 412 2234 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6181 275 412 2235 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6182 276 412 2236 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6183 277 412 2237 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6184 278 412 2238 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6185 279 412 2239 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6186 280 412 2240 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6187 281 412 2241 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6188 2242 415 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6189 2243 415 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6190 2244 415 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6191 2245 415 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6192 2246 415 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6193 2247 415 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6194 2248 415 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6195 2249 415 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6196 0 2243 2242 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6197 2243 2242 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6198 0 2245 2244 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6199 2245 2244 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6200 0 2247 2246 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6201 2247 2246 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6202 0 2249 2248 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6203 2249 2248 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6204 1 2243 2242 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6205 2243 2242 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6206 1 2245 2244 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6207 2245 2244 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6208 1 2251 2250 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6209 2251 2250 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6210 1 2253 2252 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6211 2253 2252 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6212 1 2247 2246 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6213 2247 2246 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6214 1 2249 2248 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6215 2249 2248 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6216 1 2255 2254 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6217 2255 2254 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6218 1 2257 2256 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6219 2257 2256 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6220 0 2251 2250 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6221 2251 2250 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6222 0 2253 2252 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6223 2253 2252 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6224 0 2255 2254 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6225 2255 2254 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6226 0 2257 2256 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6227 2257 2256 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6228 274 420 2250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6229 275 420 2251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6230 276 420 2252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6231 277 420 2253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6232 278 420 2254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6233 279 420 2255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6234 280 420 2256 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6235 281 420 2257 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6236 2258 424 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6237 2259 424 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6238 2260 424 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6239 2261 424 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6240 2262 424 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6241 2263 424 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6242 2264 424 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6243 2265 424 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6244 0 2259 2258 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6245 2259 2258 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6246 0 2261 2260 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6247 2261 2260 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6248 0 2263 2262 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6249 2263 2262 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6250 0 2265 2264 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6251 2265 2264 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6252 1 2259 2258 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6253 2259 2258 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6254 1 2261 2260 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6255 2261 2260 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6256 1 2263 2262 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6257 2263 2262 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6258 1 2265 2264 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6259 2265 2264 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6260 1 2267 2266 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6261 2267 2266 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6262 1 2269 2268 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6263 2269 2268 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6264 1 2271 2270 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6265 2271 2270 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6266 1 2273 2272 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6267 2273 2272 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6268 0 2267 2266 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6269 2267 2266 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6270 0 2269 2268 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6271 2269 2268 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6272 0 2271 2270 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6273 2271 2270 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6274 0 2273 2272 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6275 2273 2272 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6276 274 428 2266 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6277 275 428 2267 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6278 276 428 2268 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6279 277 428 2269 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6280 278 428 2270 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6281 279 428 2271 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6282 280 428 2272 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6283 281 428 2273 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6284 2274 431 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6285 2275 431 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6286 2276 431 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6287 2277 431 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6288 2278 431 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6289 2279 431 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6290 2280 431 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6291 2281 431 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6292 0 2275 2274 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6293 2275 2274 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6294 0 2277 2276 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6295 2277 2276 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6296 0 2279 2278 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6297 2279 2278 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6298 0 2281 2280 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6299 2281 2280 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6300 1 2275 2274 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6301 2275 2274 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6302 1 2277 2276 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6303 2277 2276 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6304 1 2283 2282 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6305 2283 2282 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6306 1 2285 2284 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6307 2285 2284 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6308 1 2279 2278 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6309 2279 2278 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6310 1 2281 2280 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6311 2281 2280 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6312 1 2287 2286 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6313 2287 2286 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6314 1 2289 2288 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6315 2289 2288 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6316 0 2283 2282 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6317 2283 2282 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6318 0 2285 2284 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6319 2285 2284 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6320 0 2287 2286 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6321 2287 2286 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6322 0 2289 2288 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6323 2289 2288 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6324 274 436 2282 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6325 275 436 2283 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6326 276 436 2284 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6327 277 436 2285 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6328 278 436 2286 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6329 279 436 2287 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6330 280 436 2288 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6331 281 436 2289 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6332 2290 440 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6333 2291 440 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6334 2292 440 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6335 2293 440 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6336 2294 440 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6337 2295 440 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6338 2296 440 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6339 2297 440 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6340 0 2291 2290 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6341 2291 2290 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6342 0 2293 2292 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6343 2293 2292 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6344 0 2295 2294 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6345 2295 2294 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6346 0 2297 2296 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6347 2297 2296 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6348 1 2291 2290 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6349 2291 2290 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6350 1 2293 2292 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6351 2293 2292 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6352 1 2295 2294 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6353 2295 2294 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6354 1 2297 2296 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6355 2297 2296 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6356 1 2299 2298 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6357 2299 2298 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6358 1 2301 2300 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6359 2301 2300 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6360 1 2303 2302 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6361 2303 2302 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6362 1 2305 2304 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6363 2305 2304 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6364 0 2299 2298 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6365 2299 2298 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6366 0 2301 2300 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6367 2301 2300 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6368 0 2303 2302 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6369 2303 2302 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6370 0 2305 2304 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6371 2305 2304 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6372 274 444 2298 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6373 275 444 2299 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6374 276 444 2300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6375 277 444 2301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6376 278 444 2302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6377 279 444 2303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6378 280 444 2304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6379 281 444 2305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6380 2306 447 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6381 2307 447 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6382 2308 447 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6383 2309 447 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6384 2310 447 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6385 2311 447 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6386 2312 447 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6387 2313 447 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6388 0 2307 2306 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6389 2307 2306 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6390 0 2309 2308 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6391 2309 2308 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6392 0 2311 2310 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6393 2311 2310 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6394 0 2313 2312 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6395 2313 2312 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6396 1 2307 2306 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6397 2307 2306 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6398 1 2309 2308 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6399 2309 2308 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6400 1 2315 2314 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6401 2315 2314 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6402 1 2317 2316 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6403 2317 2316 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6404 1 2311 2310 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6405 2311 2310 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6406 1 2313 2312 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6407 2313 2312 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6408 1 2319 2318 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6409 2319 2318 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6410 1 2321 2320 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6411 2321 2320 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6412 0 2315 2314 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6413 2315 2314 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6414 0 2317 2316 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6415 2317 2316 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6416 0 2319 2318 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6417 2319 2318 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6418 0 2321 2320 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6419 2321 2320 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6420 274 452 2314 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6421 275 452 2315 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6422 276 452 2316 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6423 277 452 2317 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6424 278 452 2318 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6425 279 452 2319 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6426 280 452 2320 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6427 281 452 2321 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6428 2322 456 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6429 2323 456 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6430 2324 456 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6431 2325 456 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6432 2326 456 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6433 2327 456 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6434 2328 456 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6435 2329 456 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6436 0 2323 2322 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6437 2323 2322 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6438 0 2325 2324 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6439 2325 2324 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6440 0 2327 2326 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6441 2327 2326 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6442 0 2329 2328 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6443 2329 2328 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6444 1 2323 2322 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6445 2323 2322 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6446 1 2325 2324 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6447 2325 2324 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6448 1 2327 2326 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6449 2327 2326 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6450 1 2329 2328 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6451 2329 2328 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6452 1 2331 2330 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6453 2331 2330 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6454 1 2333 2332 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6455 2333 2332 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6456 1 2335 2334 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6457 2335 2334 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6458 1 2337 2336 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6459 2337 2336 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6460 0 2331 2330 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6461 2331 2330 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6462 0 2333 2332 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6463 2333 2332 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6464 0 2335 2334 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6465 2335 2334 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6466 0 2337 2336 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6467 2337 2336 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6468 274 460 2330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6469 275 460 2331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6470 276 460 2332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6471 277 460 2333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6472 278 460 2334 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6473 279 460 2335 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6474 280 460 2336 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6475 281 460 2337 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6476 2338 463 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6477 2339 463 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6478 2340 463 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6479 2341 463 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6480 2342 463 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6481 2343 463 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6482 2344 463 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6483 2345 463 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6484 0 2339 2338 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6485 2339 2338 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6486 0 2341 2340 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6487 2341 2340 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6488 0 2343 2342 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6489 2343 2342 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6490 0 2345 2344 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6491 2345 2344 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6492 1 2339 2338 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6493 2339 2338 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6494 1 2341 2340 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6495 2341 2340 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6496 1 2347 2346 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6497 2347 2346 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6498 1 2349 2348 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6499 2349 2348 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6500 1 2343 2342 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6501 2343 2342 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6502 1 2345 2344 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6503 2345 2344 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6504 1 2351 2350 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6505 2351 2350 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6506 1 2353 2352 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6507 2353 2352 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6508 0 2347 2346 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6509 2347 2346 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6510 0 2349 2348 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6511 2349 2348 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6512 0 2351 2350 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6513 2351 2350 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6514 0 2353 2352 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6515 2353 2352 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6516 274 468 2346 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6517 275 468 2347 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6518 276 468 2348 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6519 277 468 2349 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6520 278 468 2350 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6521 279 468 2351 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6522 280 468 2352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6523 281 468 2353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6524 2354 472 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6525 2355 472 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6526 2356 472 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6527 2357 472 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6528 2358 472 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6529 2359 472 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6530 2360 472 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6531 2361 472 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6532 0 2355 2354 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6533 2355 2354 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6534 0 2357 2356 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6535 2357 2356 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6536 0 2359 2358 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6537 2359 2358 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6538 0 2361 2360 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6539 2361 2360 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6540 1 2355 2354 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6541 2355 2354 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6542 1 2357 2356 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6543 2357 2356 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6544 1 2359 2358 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6545 2359 2358 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6546 1 2361 2360 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6547 2361 2360 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6548 1 2363 2362 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6549 2363 2362 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6550 1 2365 2364 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6551 2365 2364 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6552 1 2367 2366 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6553 2367 2366 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6554 1 2369 2368 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6555 2369 2368 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6556 0 2363 2362 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6557 2363 2362 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6558 0 2365 2364 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6559 2365 2364 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6560 0 2367 2366 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6561 2367 2366 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6562 0 2369 2368 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6563 2369 2368 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6564 274 476 2362 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6565 275 476 2363 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6566 276 476 2364 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6567 277 476 2365 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6568 278 476 2366 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6569 279 476 2367 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6570 280 476 2368 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6571 281 476 2369 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6572 2370 479 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6573 2371 479 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6574 2372 479 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6575 2373 479 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6576 2374 479 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6577 2375 479 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6578 2376 479 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6579 2377 479 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6580 0 2371 2370 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6581 2371 2370 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6582 0 2373 2372 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6583 2373 2372 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6584 0 2375 2374 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6585 2375 2374 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6586 0 2377 2376 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6587 2377 2376 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6588 1 2371 2370 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6589 2371 2370 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6590 1 2373 2372 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6591 2373 2372 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6592 1 2379 2378 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6593 2379 2378 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6594 1 2381 2380 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6595 2381 2380 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6596 1 2375 2374 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6597 2375 2374 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6598 1 2377 2376 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6599 2377 2376 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6600 1 2383 2382 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6601 2383 2382 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6602 1 2385 2384 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6603 2385 2384 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6604 0 2379 2378 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6605 2379 2378 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6606 0 2381 2380 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6607 2381 2380 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6608 0 2383 2382 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6609 2383 2382 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6610 0 2385 2384 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6611 2385 2384 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6612 274 484 2378 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6613 275 484 2379 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6614 276 484 2380 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6615 277 484 2381 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6616 278 484 2382 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6617 279 484 2383 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6618 280 484 2384 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6619 281 484 2385 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6620 2386 488 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6621 2387 488 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6622 2388 488 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6623 2389 488 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6624 2390 488 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6625 2391 488 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6626 2392 488 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6627 2393 488 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6628 0 2387 2386 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6629 2387 2386 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6630 0 2389 2388 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6631 2389 2388 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6632 0 2391 2390 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6633 2391 2390 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6634 0 2393 2392 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6635 2393 2392 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6636 1 2387 2386 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6637 2387 2386 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6638 1 2389 2388 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6639 2389 2388 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6640 1 2391 2390 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6641 2391 2390 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6642 1 2393 2392 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6643 2393 2392 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6644 1 2395 2394 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6645 2395 2394 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6646 1 2397 2396 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6647 2397 2396 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6648 1 2399 2398 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6649 2399 2398 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6650 1 2401 2400 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6651 2401 2400 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6652 0 2395 2394 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6653 2395 2394 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6654 0 2397 2396 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6655 2397 2396 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6656 0 2399 2398 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6657 2399 2398 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6658 0 2401 2400 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6659 2401 2400 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6660 274 492 2394 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6661 275 492 2395 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6662 276 492 2396 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6663 277 492 2397 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6664 278 492 2398 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6665 279 492 2399 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6666 280 492 2400 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6667 281 492 2401 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6668 2402 495 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6669 2403 495 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6670 2404 495 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6671 2405 495 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6672 2406 495 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6673 2407 495 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6674 2408 495 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6675 2409 495 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6676 0 2403 2402 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6677 2403 2402 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6678 0 2405 2404 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6679 2405 2404 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6680 0 2407 2406 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6681 2407 2406 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6682 0 2409 2408 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6683 2409 2408 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6684 1 2403 2402 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6685 2403 2402 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6686 1 2405 2404 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6687 2405 2404 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6688 1 2411 2410 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6689 2411 2410 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6690 1 2413 2412 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6691 2413 2412 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6692 1 2407 2406 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6693 2407 2406 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6694 1 2409 2408 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6695 2409 2408 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6696 1 2415 2414 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6697 2415 2414 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6698 1 2417 2416 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6699 2417 2416 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6700 0 2411 2410 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6701 2411 2410 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6702 0 2413 2412 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6703 2413 2412 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6704 0 2415 2414 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6705 2415 2414 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6706 0 2417 2416 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6707 2417 2416 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6708 274 500 2410 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6709 275 500 2411 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6710 276 500 2412 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6711 277 500 2413 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6712 278 500 2414 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6713 279 500 2415 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6714 280 500 2416 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6715 281 500 2417 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6716 2418 504 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6717 2419 504 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6718 2420 504 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6719 2421 504 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6720 2422 504 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6721 2423 504 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6722 2424 504 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6723 2425 504 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6724 0 2419 2418 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6725 2419 2418 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6726 0 2421 2420 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6727 2421 2420 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6728 0 2423 2422 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6729 2423 2422 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6730 0 2425 2424 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6731 2425 2424 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6732 1 2419 2418 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6733 2419 2418 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6734 1 2421 2420 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6735 2421 2420 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6736 1 2423 2422 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6737 2423 2422 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6738 1 2425 2424 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6739 2425 2424 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6740 1 2427 2426 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6741 2427 2426 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6742 1 2429 2428 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6743 2429 2428 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6744 1 2431 2430 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6745 2431 2430 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6746 1 2433 2432 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6747 2433 2432 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6748 0 2427 2426 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6749 2427 2426 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6750 0 2429 2428 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6751 2429 2428 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6752 0 2431 2430 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6753 2431 2430 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6754 0 2433 2432 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6755 2433 2432 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6756 274 508 2426 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6757 275 508 2427 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6758 276 508 2428 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6759 277 508 2429 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6760 278 508 2430 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6761 279 508 2431 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6762 280 508 2432 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6763 281 508 2433 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6764 2434 511 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6765 2435 511 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6766 2436 511 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6767 2437 511 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6768 2438 511 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6769 2439 511 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6770 2440 511 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6771 2441 511 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6772 0 2435 2434 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6773 2435 2434 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6774 0 2437 2436 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6775 2437 2436 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6776 0 2439 2438 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6777 2439 2438 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6778 0 2441 2440 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6779 2441 2440 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6780 1 2435 2434 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6781 2435 2434 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6782 1 2437 2436 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6783 2437 2436 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6784 1 2443 2442 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6785 2443 2442 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6786 1 2445 2444 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6787 2445 2444 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6788 1 2439 2438 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6789 2439 2438 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6790 1 2441 2440 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6791 2441 2440 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6792 1 2447 2446 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6793 2447 2446 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6794 1 2449 2448 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6795 2449 2448 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6796 0 2443 2442 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6797 2443 2442 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6798 0 2445 2444 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6799 2445 2444 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6800 0 2447 2446 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6801 2447 2446 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6802 0 2449 2448 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6803 2449 2448 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6804 274 516 2442 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6805 275 516 2443 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6806 276 516 2444 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6807 277 516 2445 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6808 278 516 2446 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6809 279 516 2447 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6810 280 516 2448 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6811 281 516 2449 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6812 2450 520 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6813 2451 520 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6814 2452 520 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6815 2453 520 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6816 2454 520 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6817 2455 520 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6818 2456 520 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6819 2457 520 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6820 0 2451 2450 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6821 2451 2450 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6822 0 2453 2452 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6823 2453 2452 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6824 0 2455 2454 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6825 2455 2454 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6826 0 2457 2456 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6827 2457 2456 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6828 1 2451 2450 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6829 2451 2450 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6830 1 2453 2452 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6831 2453 2452 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6832 1 2455 2454 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6833 2455 2454 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6834 1 2457 2456 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6835 2457 2456 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6836 1 2459 2458 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6837 2459 2458 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6838 1 2461 2460 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6839 2461 2460 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6840 1 2463 2462 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6841 2463 2462 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6842 1 2465 2464 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6843 2465 2464 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6844 0 2459 2458 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6845 2459 2458 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6846 0 2461 2460 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6847 2461 2460 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6848 0 2463 2462 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6849 2463 2462 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6850 0 2465 2464 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6851 2465 2464 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6852 274 524 2458 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6853 275 524 2459 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6854 276 524 2460 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6855 277 524 2461 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6856 278 524 2462 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6857 279 524 2463 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6858 280 524 2464 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6859 281 524 2465 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6860 2466 527 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6861 2467 527 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6862 2468 527 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6863 2469 527 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6864 2470 527 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6865 2471 527 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6866 2472 527 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6867 2473 527 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6868 0 2467 2466 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6869 2467 2466 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6870 0 2469 2468 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6871 2469 2468 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6872 0 2471 2470 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6873 2471 2470 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6874 0 2473 2472 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6875 2473 2472 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6876 1 2467 2466 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6877 2467 2466 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6878 1 2469 2468 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6879 2469 2468 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6880 1 2475 2474 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6881 2475 2474 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6882 1 2477 2476 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6883 2477 2476 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6884 1 2471 2470 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6885 2471 2470 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6886 1 2473 2472 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6887 2473 2472 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6888 1 2479 2478 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6889 2479 2478 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6890 1 2481 2480 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6891 2481 2480 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6892 0 2475 2474 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6893 2475 2474 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6894 0 2477 2476 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6895 2477 2476 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6896 0 2479 2478 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6897 2479 2478 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6898 0 2481 2480 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6899 2481 2480 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6900 274 532 2474 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6901 275 532 2475 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6902 276 532 2476 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6903 277 532 2477 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6904 278 532 2478 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6905 279 532 2479 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6906 280 532 2480 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6907 281 532 2481 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6908 2482 536 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6909 2483 536 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6910 2484 536 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6911 2485 536 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6912 2486 536 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6913 2487 536 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6914 2488 536 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6915 2489 536 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6916 0 2483 2482 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6917 2483 2482 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6918 0 2485 2484 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6919 2485 2484 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6920 0 2487 2486 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6921 2487 2486 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6922 0 2489 2488 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6923 2489 2488 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6924 1 2483 2482 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6925 2483 2482 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6926 1 2485 2484 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6927 2485 2484 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6928 1 2487 2486 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6929 2487 2486 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6930 1 2489 2488 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6931 2489 2488 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6932 1 2491 2490 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6933 2491 2490 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6934 1 2493 2492 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6935 2493 2492 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6936 1 2495 2494 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6937 2495 2494 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6938 1 2497 2496 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6939 2497 2496 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6940 0 2491 2490 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6941 2491 2490 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6942 0 2493 2492 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6943 2493 2492 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6944 0 2495 2494 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6945 2495 2494 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6946 0 2497 2496 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6947 2497 2496 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6948 274 540 2490 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6949 275 540 2491 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6950 276 540 2492 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6951 277 540 2493 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6952 278 540 2494 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m6953 279 540 2495 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6954 280 540 2496 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6955 281 540 2497 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m6956 2498 543 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m6957 2499 543 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6958 2500 543 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6959 2501 543 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6960 2502 543 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m6961 2503 543 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m6962 2504 543 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m6963 2505 543 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m6964 0 2499 2498 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6965 2499 2498 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6966 0 2501 2500 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6967 2501 2500 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6968 0 2503 2502 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6969 2503 2502 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6970 0 2505 2504 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6971 2505 2504 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6972 1 2499 2498 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6973 2499 2498 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6974 1 2501 2500 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6975 2501 2500 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6976 1 2507 2506 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6977 2507 2506 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m6978 1 2509 2508 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6979 2509 2508 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6980 1 2503 2502 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6981 2503 2502 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6982 1 2505 2504 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6983 2505 2504 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6984 1 2511 2510 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m6985 2511 2510 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6986 1 2513 2512 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m6987 2513 2512 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m6988 0 2507 2506 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6989 2507 2506 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6990 0 2509 2508 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m6991 2509 2508 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m6992 0 2511 2510 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6993 2511 2510 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6994 0 2513 2512 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m6995 2513 2512 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m6996 274 548 2506 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m6997 275 548 2507 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m6998 276 548 2508 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m6999 277 548 2509 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7000 278 548 2510 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7001 279 548 2511 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7002 280 548 2512 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7003 281 548 2513 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7004 2514 552 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7005 2515 552 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7006 2516 552 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7007 2517 552 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7008 2518 552 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7009 2519 552 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7010 2520 552 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7011 2521 552 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7012 0 2515 2514 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7013 2515 2514 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7014 0 2517 2516 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7015 2517 2516 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7016 0 2519 2518 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7017 2519 2518 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7018 0 2521 2520 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7019 2521 2520 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7020 1 2515 2514 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7021 2515 2514 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7022 1 2517 2516 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7023 2517 2516 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7024 1 2519 2518 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7025 2519 2518 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7026 1 2521 2520 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7027 2521 2520 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7028 1 2523 2522 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7029 2523 2522 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7030 1 2525 2524 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7031 2525 2524 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7032 1 2527 2526 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7033 2527 2526 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7034 1 2529 2528 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7035 2529 2528 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7036 0 2523 2522 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7037 2523 2522 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7038 0 2525 2524 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7039 2525 2524 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7040 0 2527 2526 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7041 2527 2526 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7042 0 2529 2528 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7043 2529 2528 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7044 274 556 2522 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7045 275 556 2523 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7046 276 556 2524 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7047 277 556 2525 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7048 278 556 2526 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7049 279 556 2527 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7050 280 556 2528 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7051 281 556 2529 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7052 2530 559 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7053 2531 559 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7054 2532 559 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7055 2533 559 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7056 2534 559 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7057 2535 559 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7058 2536 559 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7059 2537 559 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7060 0 2531 2530 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7061 2531 2530 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7062 0 2533 2532 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7063 2533 2532 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7064 0 2535 2534 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7065 2535 2534 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7066 0 2537 2536 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7067 2537 2536 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7068 1 2531 2530 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7069 2531 2530 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7070 1 2533 2532 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7071 2533 2532 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7072 1 2539 2538 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7073 2539 2538 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7074 1 2541 2540 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7075 2541 2540 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7076 1 2535 2534 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7077 2535 2534 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7078 1 2537 2536 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7079 2537 2536 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7080 1 2543 2542 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7081 2543 2542 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7082 1 2545 2544 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7083 2545 2544 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7084 0 2539 2538 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7085 2539 2538 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7086 0 2541 2540 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7087 2541 2540 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7088 0 2543 2542 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7089 2543 2542 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7090 0 2545 2544 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7091 2545 2544 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7092 274 564 2538 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7093 275 564 2539 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7094 276 564 2540 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7095 277 564 2541 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7096 278 564 2542 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7097 279 564 2543 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7098 280 564 2544 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7099 281 564 2545 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7100 2546 568 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7101 2547 568 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7102 2548 568 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7103 2549 568 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7104 2550 568 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7105 2551 568 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7106 2552 568 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7107 2553 568 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7108 0 2547 2546 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7109 2547 2546 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7110 0 2549 2548 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7111 2549 2548 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7112 0 2551 2550 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7113 2551 2550 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7114 0 2553 2552 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7115 2553 2552 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7116 1 2547 2546 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7117 2547 2546 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7118 1 2549 2548 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7119 2549 2548 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7120 1 2551 2550 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7121 2551 2550 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7122 1 2553 2552 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7123 2553 2552 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7124 1 2555 2554 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7125 2555 2554 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7126 1 2557 2556 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7127 2557 2556 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7128 1 2559 2558 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7129 2559 2558 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7130 1 2561 2560 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7131 2561 2560 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7132 0 2555 2554 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7133 2555 2554 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7134 0 2557 2556 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7135 2557 2556 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7136 0 2559 2558 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7137 2559 2558 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7138 0 2561 2560 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7139 2561 2560 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7140 274 572 2554 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7141 275 572 2555 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7142 276 572 2556 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7143 277 572 2557 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7144 278 572 2558 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7145 279 572 2559 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7146 280 572 2560 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7147 281 572 2561 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7148 2562 575 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7149 2563 575 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7150 2564 575 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7151 2565 575 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7152 2566 575 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7153 2567 575 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7154 2568 575 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7155 2569 575 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7156 0 2563 2562 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7157 2563 2562 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7158 0 2565 2564 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7159 2565 2564 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7160 0 2567 2566 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7161 2567 2566 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7162 0 2569 2568 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7163 2569 2568 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7164 1 2563 2562 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7165 2563 2562 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7166 1 2565 2564 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7167 2565 2564 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7168 1 2571 2570 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7169 2571 2570 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7170 1 2573 2572 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7171 2573 2572 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7172 1 2567 2566 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7173 2567 2566 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7174 1 2569 2568 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7175 2569 2568 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7176 1 2575 2574 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7177 2575 2574 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7178 1 2577 2576 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7179 2577 2576 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7180 0 2571 2570 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7181 2571 2570 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7182 0 2573 2572 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7183 2573 2572 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7184 0 2575 2574 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7185 2575 2574 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7186 0 2577 2576 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7187 2577 2576 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7188 274 580 2570 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7189 275 580 2571 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7190 276 580 2572 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7191 277 580 2573 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7192 278 580 2574 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7193 279 580 2575 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7194 280 580 2576 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7195 281 580 2577 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7196 2578 584 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7197 2579 584 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7198 2580 584 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7199 2581 584 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7200 2582 584 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7201 2583 584 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7202 2584 584 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7203 2585 584 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7204 0 2579 2578 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7205 2579 2578 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7206 0 2581 2580 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7207 2581 2580 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7208 0 2583 2582 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7209 2583 2582 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7210 0 2585 2584 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7211 2585 2584 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7212 1 2579 2578 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7213 2579 2578 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7214 1 2581 2580 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7215 2581 2580 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7216 1 2583 2582 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7217 2583 2582 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7218 1 2585 2584 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7219 2585 2584 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7220 1 2587 2586 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7221 2587 2586 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7222 1 2589 2588 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7223 2589 2588 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7224 1 2591 2590 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7225 2591 2590 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7226 1 2593 2592 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7227 2593 2592 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7228 0 2587 2586 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7229 2587 2586 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7230 0 2589 2588 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7231 2589 2588 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7232 0 2591 2590 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7233 2591 2590 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7234 0 2593 2592 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7235 2593 2592 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7236 274 588 2586 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7237 275 588 2587 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7238 276 588 2588 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7239 277 588 2589 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7240 278 588 2590 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7241 279 588 2591 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7242 280 588 2592 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7243 281 588 2593 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7244 2594 591 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7245 2595 591 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7246 2596 591 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7247 2597 591 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7248 2598 591 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7249 2599 591 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7250 2600 591 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7251 2601 591 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7252 0 2595 2594 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7253 2595 2594 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7254 0 2597 2596 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7255 2597 2596 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7256 0 2599 2598 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7257 2599 2598 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7258 0 2601 2600 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7259 2601 2600 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7260 1 2595 2594 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7261 2595 2594 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7262 1 2597 2596 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7263 2597 2596 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7264 1 2603 2602 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7265 2603 2602 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7266 1 2605 2604 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7267 2605 2604 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7268 1 2599 2598 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7269 2599 2598 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7270 1 2601 2600 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7271 2601 2600 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7272 1 2607 2606 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7273 2607 2606 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7274 1 2609 2608 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7275 2609 2608 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7276 0 2603 2602 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7277 2603 2602 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7278 0 2605 2604 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7279 2605 2604 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7280 0 2607 2606 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7281 2607 2606 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7282 0 2609 2608 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7283 2609 2608 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7284 274 596 2602 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7285 275 596 2603 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7286 276 596 2604 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7287 277 596 2605 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7288 278 596 2606 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7289 279 596 2607 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7290 280 596 2608 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7291 281 596 2609 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7292 2610 600 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7293 2611 600 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7294 2612 600 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7295 2613 600 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7296 2614 600 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7297 2615 600 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7298 2616 600 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7299 2617 600 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7300 0 2611 2610 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7301 2611 2610 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7302 0 2613 2612 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7303 2613 2612 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7304 0 2615 2614 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7305 2615 2614 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7306 0 2617 2616 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7307 2617 2616 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7308 1 2611 2610 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7309 2611 2610 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7310 1 2613 2612 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7311 2613 2612 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7312 1 2615 2614 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7313 2615 2614 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7314 1 2617 2616 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7315 2617 2616 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7316 1 2619 2618 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7317 2619 2618 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7318 1 2621 2620 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7319 2621 2620 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7320 1 2623 2622 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7321 2623 2622 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7322 1 2625 2624 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7323 2625 2624 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7324 0 2619 2618 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7325 2619 2618 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7326 0 2621 2620 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7327 2621 2620 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7328 0 2623 2622 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7329 2623 2622 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7330 0 2625 2624 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7331 2625 2624 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7332 274 604 2618 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7333 275 604 2619 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7334 276 604 2620 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7335 277 604 2621 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7336 278 604 2622 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7337 279 604 2623 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7338 280 604 2624 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7339 281 604 2625 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7340 2626 607 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7341 2627 607 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7342 2628 607 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7343 2629 607 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7344 2630 607 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7345 2631 607 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7346 2632 607 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7347 2633 607 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7348 0 2627 2626 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7349 2627 2626 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7350 0 2629 2628 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7351 2629 2628 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7352 0 2631 2630 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7353 2631 2630 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7354 0 2633 2632 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7355 2633 2632 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7356 1 2627 2626 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7357 2627 2626 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7358 1 2629 2628 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7359 2629 2628 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7360 1 2635 2634 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7361 2635 2634 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7362 1 2637 2636 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7363 2637 2636 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7364 1 2631 2630 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7365 2631 2630 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7366 1 2633 2632 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7367 2633 2632 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7368 1 2639 2638 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7369 2639 2638 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7370 1 2641 2640 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7371 2641 2640 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7372 0 2635 2634 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7373 2635 2634 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7374 0 2637 2636 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7375 2637 2636 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7376 0 2639 2638 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7377 2639 2638 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7378 0 2641 2640 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7379 2641 2640 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7380 274 612 2634 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7381 275 612 2635 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7382 276 612 2636 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7383 277 612 2637 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7384 278 612 2638 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7385 279 612 2639 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7386 280 612 2640 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7387 281 612 2641 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7388 2642 616 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7389 2643 616 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7390 2644 616 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7391 2645 616 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7392 2646 616 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7393 2647 616 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7394 2648 616 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7395 2649 616 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7396 0 2643 2642 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7397 2643 2642 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7398 0 2645 2644 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7399 2645 2644 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7400 0 2647 2646 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7401 2647 2646 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7402 0 2649 2648 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7403 2649 2648 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7404 1 2643 2642 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7405 2643 2642 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7406 1 2645 2644 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7407 2645 2644 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7408 1 2647 2646 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7409 2647 2646 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7410 1 2649 2648 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7411 2649 2648 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7412 1 2651 2650 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7413 2651 2650 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7414 1 2653 2652 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7415 2653 2652 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7416 1 2655 2654 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7417 2655 2654 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7418 1 2657 2656 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7419 2657 2656 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7420 0 2651 2650 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7421 2651 2650 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7422 0 2653 2652 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7423 2653 2652 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7424 0 2655 2654 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7425 2655 2654 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7426 0 2657 2656 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7427 2657 2656 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7428 274 620 2650 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7429 275 620 2651 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7430 276 620 2652 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7431 277 620 2653 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7432 278 620 2654 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7433 279 620 2655 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7434 280 620 2656 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7435 281 620 2657 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7436 2658 624 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7437 2659 624 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7438 2660 624 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7439 2661 624 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7440 2662 624 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7441 2663 624 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7442 2664 624 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7443 2665 624 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7444 0 2659 2658 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7445 2659 2658 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7446 0 2661 2660 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7447 2661 2660 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7448 0 2663 2662 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7449 2663 2662 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7450 0 2665 2664 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7451 2665 2664 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7452 1 2659 2658 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7453 2659 2658 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7454 1 2661 2660 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7455 2661 2660 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7456 1 2667 2666 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7457 2667 2666 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7458 1 2669 2668 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7459 2669 2668 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7460 1 2663 2662 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7461 2663 2662 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7462 1 2665 2664 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7463 2665 2664 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7464 1 2671 2670 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7465 2671 2670 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7466 1 2673 2672 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7467 2673 2672 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7468 0 2667 2666 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7469 2667 2666 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7470 0 2669 2668 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7471 2669 2668 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7472 0 2671 2670 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7473 2671 2670 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7474 0 2673 2672 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7475 2673 2672 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7476 274 628 2666 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7477 275 628 2667 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7478 276 628 2668 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7479 277 628 2669 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7480 278 628 2670 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7481 279 628 2671 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7482 280 628 2672 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7483 281 628 2673 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7484 2674 632 274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7485 2675 632 275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7486 2676 632 276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7487 2677 632 277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7488 2678 632 278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7489 2679 632 279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7490 2680 632 280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7491 2681 632 281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7492 0 2675 2674 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7493 2675 2674 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7494 0 2677 2676 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7495 2677 2676 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7496 0 2679 2678 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7497 2679 2678 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7498 0 2681 2680 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7499 2681 2680 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7500 1 2675 2674 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7501 2675 2674 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7502 1 2677 2676 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7503 2677 2676 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7504 1 2679 2678 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7505 2679 2678 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7506 1 2681 2680 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7507 2681 2680 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7508 1 2683 2682 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7509 2683 2682 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7510 1 2685 2684 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7511 2685 2684 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7512 1 2687 2686 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7513 2687 2686 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7514 1 2689 2688 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7515 2689 2688 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7516 0 2683 2682 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7517 2683 2682 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7518 0 2685 2684 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7519 2685 2684 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7520 0 2687 2686 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7521 2687 2686 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7522 0 2689 2688 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7523 2689 2688 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7524 300 380 2682 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7525 301 380 2683 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7526 302 380 2684 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7527 303 380 2685 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7528 304 380 2686 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7529 305 380 2687 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7530 306 380 2688 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7531 307 380 2689 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7532 2690 383 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7533 2691 383 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7534 2692 383 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7535 2693 383 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7536 2694 383 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7537 2695 383 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7538 2696 383 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7539 2697 383 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7540 0 2691 2690 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7541 2691 2690 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7542 0 2693 2692 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7543 2693 2692 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7544 0 2695 2694 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7545 2695 2694 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7546 0 2697 2696 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7547 2697 2696 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7548 1 2691 2690 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7549 2691 2690 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7550 1 2693 2692 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7551 2693 2692 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7552 1 2699 2698 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7553 2699 2698 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7554 1 2701 2700 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7555 2701 2700 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7556 1 2695 2694 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7557 2695 2694 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7558 1 2697 2696 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7559 2697 2696 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7560 1 2703 2702 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7561 2703 2702 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7562 1 2705 2704 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7563 2705 2704 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7564 0 2699 2698 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7565 2699 2698 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7566 0 2701 2700 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7567 2701 2700 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7568 0 2703 2702 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7569 2703 2702 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7570 0 2705 2704 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7571 2705 2704 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7572 300 388 2698 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7573 301 388 2699 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7574 302 388 2700 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7575 303 388 2701 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7576 304 388 2702 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7577 305 388 2703 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7578 306 388 2704 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7579 307 388 2705 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7580 2706 392 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7581 2707 392 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7582 2708 392 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7583 2709 392 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7584 2710 392 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7585 2711 392 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7586 2712 392 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7587 2713 392 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7588 0 2707 2706 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7589 2707 2706 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7590 0 2709 2708 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7591 2709 2708 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7592 0 2711 2710 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7593 2711 2710 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7594 0 2713 2712 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7595 2713 2712 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7596 1 2707 2706 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7597 2707 2706 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7598 1 2709 2708 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7599 2709 2708 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7600 1 2711 2710 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7601 2711 2710 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7602 1 2713 2712 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7603 2713 2712 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7604 1 2715 2714 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7605 2715 2714 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7606 1 2717 2716 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7607 2717 2716 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7608 1 2719 2718 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7609 2719 2718 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7610 1 2721 2720 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7611 2721 2720 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7612 0 2715 2714 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7613 2715 2714 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7614 0 2717 2716 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7615 2717 2716 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7616 0 2719 2718 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7617 2719 2718 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7618 0 2721 2720 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7619 2721 2720 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7620 300 396 2714 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7621 301 396 2715 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7622 302 396 2716 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7623 303 396 2717 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7624 304 396 2718 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7625 305 396 2719 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7626 306 396 2720 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7627 307 396 2721 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7628 2722 399 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7629 2723 399 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7630 2724 399 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7631 2725 399 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7632 2726 399 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7633 2727 399 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7634 2728 399 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7635 2729 399 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7636 0 2723 2722 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7637 2723 2722 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7638 0 2725 2724 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7639 2725 2724 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7640 0 2727 2726 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7641 2727 2726 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7642 0 2729 2728 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7643 2729 2728 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7644 1 2723 2722 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7645 2723 2722 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7646 1 2725 2724 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7647 2725 2724 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7648 1 2731 2730 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7649 2731 2730 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7650 1 2733 2732 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7651 2733 2732 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7652 1 2727 2726 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7653 2727 2726 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7654 1 2729 2728 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7655 2729 2728 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7656 1 2735 2734 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7657 2735 2734 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7658 1 2737 2736 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7659 2737 2736 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7660 0 2731 2730 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7661 2731 2730 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7662 0 2733 2732 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7663 2733 2732 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7664 0 2735 2734 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7665 2735 2734 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7666 0 2737 2736 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7667 2737 2736 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7668 300 404 2730 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7669 301 404 2731 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7670 302 404 2732 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7671 303 404 2733 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7672 304 404 2734 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7673 305 404 2735 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7674 306 404 2736 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7675 307 404 2737 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7676 2738 408 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7677 2739 408 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7678 2740 408 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7679 2741 408 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7680 2742 408 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7681 2743 408 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7682 2744 408 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7683 2745 408 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7684 0 2739 2738 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7685 2739 2738 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7686 0 2741 2740 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7687 2741 2740 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7688 0 2743 2742 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7689 2743 2742 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7690 0 2745 2744 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7691 2745 2744 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7692 1 2739 2738 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7693 2739 2738 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7694 1 2741 2740 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7695 2741 2740 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7696 1 2743 2742 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7697 2743 2742 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7698 1 2745 2744 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7699 2745 2744 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7700 1 2747 2746 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7701 2747 2746 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7702 1 2749 2748 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7703 2749 2748 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7704 1 2751 2750 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7705 2751 2750 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7706 1 2753 2752 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7707 2753 2752 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7708 0 2747 2746 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7709 2747 2746 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7710 0 2749 2748 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7711 2749 2748 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7712 0 2751 2750 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7713 2751 2750 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7714 0 2753 2752 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7715 2753 2752 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7716 300 412 2746 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7717 301 412 2747 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7718 302 412 2748 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7719 303 412 2749 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7720 304 412 2750 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7721 305 412 2751 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7722 306 412 2752 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7723 307 412 2753 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7724 2754 415 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7725 2755 415 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7726 2756 415 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7727 2757 415 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7728 2758 415 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7729 2759 415 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7730 2760 415 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7731 2761 415 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7732 0 2755 2754 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7733 2755 2754 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7734 0 2757 2756 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7735 2757 2756 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7736 0 2759 2758 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7737 2759 2758 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7738 0 2761 2760 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7739 2761 2760 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7740 1 2755 2754 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7741 2755 2754 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7742 1 2757 2756 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7743 2757 2756 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7744 1 2763 2762 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7745 2763 2762 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7746 1 2765 2764 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7747 2765 2764 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7748 1 2759 2758 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7749 2759 2758 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7750 1 2761 2760 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7751 2761 2760 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7752 1 2767 2766 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7753 2767 2766 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7754 1 2769 2768 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7755 2769 2768 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7756 0 2763 2762 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7757 2763 2762 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7758 0 2765 2764 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7759 2765 2764 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7760 0 2767 2766 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7761 2767 2766 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7762 0 2769 2768 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7763 2769 2768 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7764 300 420 2762 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7765 301 420 2763 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7766 302 420 2764 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7767 303 420 2765 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7768 304 420 2766 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7769 305 420 2767 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7770 306 420 2768 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7771 307 420 2769 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7772 2770 424 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7773 2771 424 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7774 2772 424 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7775 2773 424 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7776 2774 424 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7777 2775 424 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7778 2776 424 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7779 2777 424 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7780 0 2771 2770 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7781 2771 2770 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7782 0 2773 2772 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7783 2773 2772 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7784 0 2775 2774 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7785 2775 2774 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7786 0 2777 2776 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7787 2777 2776 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7788 1 2771 2770 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7789 2771 2770 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7790 1 2773 2772 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7791 2773 2772 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7792 1 2775 2774 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7793 2775 2774 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7794 1 2777 2776 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7795 2777 2776 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7796 1 2779 2778 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7797 2779 2778 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7798 1 2781 2780 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7799 2781 2780 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7800 1 2783 2782 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7801 2783 2782 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7802 1 2785 2784 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7803 2785 2784 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7804 0 2779 2778 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7805 2779 2778 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7806 0 2781 2780 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7807 2781 2780 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7808 0 2783 2782 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7809 2783 2782 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7810 0 2785 2784 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7811 2785 2784 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7812 300 428 2778 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7813 301 428 2779 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7814 302 428 2780 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7815 303 428 2781 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7816 304 428 2782 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7817 305 428 2783 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7818 306 428 2784 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7819 307 428 2785 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7820 2786 431 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7821 2787 431 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7822 2788 431 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7823 2789 431 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7824 2790 431 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7825 2791 431 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7826 2792 431 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7827 2793 431 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7828 0 2787 2786 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7829 2787 2786 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7830 0 2789 2788 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7831 2789 2788 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7832 0 2791 2790 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7833 2791 2790 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7834 0 2793 2792 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7835 2793 2792 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7836 1 2787 2786 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7837 2787 2786 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7838 1 2789 2788 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7839 2789 2788 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7840 1 2795 2794 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7841 2795 2794 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7842 1 2797 2796 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7843 2797 2796 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7844 1 2791 2790 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7845 2791 2790 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7846 1 2793 2792 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7847 2793 2792 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7848 1 2799 2798 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7849 2799 2798 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7850 1 2801 2800 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7851 2801 2800 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7852 0 2795 2794 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7853 2795 2794 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7854 0 2797 2796 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7855 2797 2796 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7856 0 2799 2798 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7857 2799 2798 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7858 0 2801 2800 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7859 2801 2800 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7860 300 436 2794 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7861 301 436 2795 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7862 302 436 2796 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7863 303 436 2797 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7864 304 436 2798 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7865 305 436 2799 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7866 306 436 2800 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7867 307 436 2801 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7868 2802 440 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7869 2803 440 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7870 2804 440 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7871 2805 440 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7872 2806 440 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7873 2807 440 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7874 2808 440 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7875 2809 440 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7876 0 2803 2802 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7877 2803 2802 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7878 0 2805 2804 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7879 2805 2804 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7880 0 2807 2806 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7881 2807 2806 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7882 0 2809 2808 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7883 2809 2808 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7884 1 2803 2802 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7885 2803 2802 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7886 1 2805 2804 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7887 2805 2804 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7888 1 2807 2806 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7889 2807 2806 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7890 1 2809 2808 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7891 2809 2808 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7892 1 2811 2810 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7893 2811 2810 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7894 1 2813 2812 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7895 2813 2812 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7896 1 2815 2814 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7897 2815 2814 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7898 1 2817 2816 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7899 2817 2816 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7900 0 2811 2810 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7901 2811 2810 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7902 0 2813 2812 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7903 2813 2812 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7904 0 2815 2814 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7905 2815 2814 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7906 0 2817 2816 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7907 2817 2816 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7908 300 444 2810 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7909 301 444 2811 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7910 302 444 2812 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7911 303 444 2813 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7912 304 444 2814 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7913 305 444 2815 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7914 306 444 2816 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7915 307 444 2817 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7916 2818 447 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7917 2819 447 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7918 2820 447 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7919 2821 447 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7920 2822 447 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7921 2823 447 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7922 2824 447 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7923 2825 447 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7924 0 2819 2818 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7925 2819 2818 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7926 0 2821 2820 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7927 2821 2820 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7928 0 2823 2822 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7929 2823 2822 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7930 0 2825 2824 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7931 2825 2824 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7932 1 2819 2818 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7933 2819 2818 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7934 1 2821 2820 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7935 2821 2820 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7936 1 2827 2826 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7937 2827 2826 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7938 1 2829 2828 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7939 2829 2828 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7940 1 2823 2822 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7941 2823 2822 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7942 1 2825 2824 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7943 2825 2824 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7944 1 2831 2830 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7945 2831 2830 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7946 1 2833 2832 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7947 2833 2832 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7948 0 2827 2826 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7949 2827 2826 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7950 0 2829 2828 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7951 2829 2828 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7952 0 2831 2830 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7953 2831 2830 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7954 0 2833 2832 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7955 2833 2832 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7956 300 452 2826 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m7957 301 452 2827 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7958 302 452 2828 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7959 303 452 2829 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7960 304 452 2830 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m7961 305 452 2831 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m7962 306 452 2832 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m7963 307 452 2833 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m7964 2834 456 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m7965 2835 456 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7966 2836 456 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7967 2837 456 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7968 2838 456 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m7969 2839 456 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m7970 2840 456 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m7971 2841 456 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m7972 0 2835 2834 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7973 2835 2834 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7974 0 2837 2836 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7975 2837 2836 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7976 0 2839 2838 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7977 2839 2838 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7978 0 2841 2840 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m7979 2841 2840 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m7980 1 2835 2834 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7981 2835 2834 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7982 1 2837 2836 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7983 2837 2836 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7984 1 2839 2838 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7985 2839 2838 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7986 1 2841 2840 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7987 2841 2840 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7988 1 2843 2842 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7989 2843 2842 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m7990 1 2845 2844 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7991 2845 2844 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7992 1 2847 2846 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m7993 2847 2846 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7994 1 2849 2848 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m7995 2849 2848 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m7996 0 2843 2842 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7997 2843 2842 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m7998 0 2845 2844 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m7999 2845 2844 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8000 0 2847 2846 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8001 2847 2846 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8002 0 2849 2848 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8003 2849 2848 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8004 300 460 2842 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8005 301 460 2843 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8006 302 460 2844 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8007 303 460 2845 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8008 304 460 2846 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8009 305 460 2847 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8010 306 460 2848 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8011 307 460 2849 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8012 2850 463 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8013 2851 463 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8014 2852 463 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8015 2853 463 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8016 2854 463 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8017 2855 463 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8018 2856 463 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8019 2857 463 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8020 0 2851 2850 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8021 2851 2850 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8022 0 2853 2852 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8023 2853 2852 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8024 0 2855 2854 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8025 2855 2854 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8026 0 2857 2856 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8027 2857 2856 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8028 1 2851 2850 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8029 2851 2850 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8030 1 2853 2852 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8031 2853 2852 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8032 1 2859 2858 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8033 2859 2858 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8034 1 2861 2860 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8035 2861 2860 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8036 1 2855 2854 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8037 2855 2854 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8038 1 2857 2856 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8039 2857 2856 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8040 1 2863 2862 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8041 2863 2862 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8042 1 2865 2864 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8043 2865 2864 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8044 0 2859 2858 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8045 2859 2858 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8046 0 2861 2860 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8047 2861 2860 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8048 0 2863 2862 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8049 2863 2862 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8050 0 2865 2864 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8051 2865 2864 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8052 300 468 2858 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8053 301 468 2859 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8054 302 468 2860 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8055 303 468 2861 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8056 304 468 2862 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8057 305 468 2863 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8058 306 468 2864 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8059 307 468 2865 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8060 2866 472 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8061 2867 472 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8062 2868 472 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8063 2869 472 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8064 2870 472 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8065 2871 472 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8066 2872 472 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8067 2873 472 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8068 0 2867 2866 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8069 2867 2866 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8070 0 2869 2868 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8071 2869 2868 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8072 0 2871 2870 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8073 2871 2870 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8074 0 2873 2872 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8075 2873 2872 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8076 1 2867 2866 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8077 2867 2866 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8078 1 2869 2868 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8079 2869 2868 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8080 1 2871 2870 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8081 2871 2870 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8082 1 2873 2872 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8083 2873 2872 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8084 1 2875 2874 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8085 2875 2874 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8086 1 2877 2876 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8087 2877 2876 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8088 1 2879 2878 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8089 2879 2878 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8090 1 2881 2880 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8091 2881 2880 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8092 0 2875 2874 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8093 2875 2874 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8094 0 2877 2876 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8095 2877 2876 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8096 0 2879 2878 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8097 2879 2878 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8098 0 2881 2880 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8099 2881 2880 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8100 300 476 2874 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8101 301 476 2875 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8102 302 476 2876 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8103 303 476 2877 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8104 304 476 2878 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8105 305 476 2879 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8106 306 476 2880 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8107 307 476 2881 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8108 2882 479 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8109 2883 479 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8110 2884 479 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8111 2885 479 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8112 2886 479 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8113 2887 479 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8114 2888 479 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8115 2889 479 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8116 0 2883 2882 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8117 2883 2882 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8118 0 2885 2884 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8119 2885 2884 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8120 0 2887 2886 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8121 2887 2886 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8122 0 2889 2888 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8123 2889 2888 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8124 1 2883 2882 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8125 2883 2882 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8126 1 2885 2884 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8127 2885 2884 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8128 1 2891 2890 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8129 2891 2890 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8130 1 2893 2892 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8131 2893 2892 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8132 1 2887 2886 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8133 2887 2886 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8134 1 2889 2888 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8135 2889 2888 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8136 1 2895 2894 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8137 2895 2894 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8138 1 2897 2896 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8139 2897 2896 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8140 0 2891 2890 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8141 2891 2890 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8142 0 2893 2892 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8143 2893 2892 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8144 0 2895 2894 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8145 2895 2894 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8146 0 2897 2896 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8147 2897 2896 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8148 300 484 2890 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8149 301 484 2891 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8150 302 484 2892 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8151 303 484 2893 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8152 304 484 2894 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8153 305 484 2895 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8154 306 484 2896 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8155 307 484 2897 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8156 2898 488 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8157 2899 488 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8158 2900 488 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8159 2901 488 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8160 2902 488 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8161 2903 488 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8162 2904 488 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8163 2905 488 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8164 0 2899 2898 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8165 2899 2898 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8166 0 2901 2900 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8167 2901 2900 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8168 0 2903 2902 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8169 2903 2902 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8170 0 2905 2904 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8171 2905 2904 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8172 1 2899 2898 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8173 2899 2898 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8174 1 2901 2900 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8175 2901 2900 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8176 1 2903 2902 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8177 2903 2902 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8178 1 2905 2904 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8179 2905 2904 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8180 1 2907 2906 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8181 2907 2906 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8182 1 2909 2908 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8183 2909 2908 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8184 1 2911 2910 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8185 2911 2910 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8186 1 2913 2912 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8187 2913 2912 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8188 0 2907 2906 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8189 2907 2906 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8190 0 2909 2908 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8191 2909 2908 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8192 0 2911 2910 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8193 2911 2910 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8194 0 2913 2912 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8195 2913 2912 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8196 300 492 2906 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8197 301 492 2907 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8198 302 492 2908 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8199 303 492 2909 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8200 304 492 2910 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8201 305 492 2911 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8202 306 492 2912 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8203 307 492 2913 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8204 2914 495 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8205 2915 495 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8206 2916 495 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8207 2917 495 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8208 2918 495 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8209 2919 495 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8210 2920 495 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8211 2921 495 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8212 0 2915 2914 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8213 2915 2914 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8214 0 2917 2916 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8215 2917 2916 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8216 0 2919 2918 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8217 2919 2918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8218 0 2921 2920 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8219 2921 2920 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8220 1 2915 2914 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8221 2915 2914 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8222 1 2917 2916 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8223 2917 2916 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8224 1 2923 2922 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8225 2923 2922 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8226 1 2925 2924 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8227 2925 2924 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8228 1 2919 2918 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8229 2919 2918 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8230 1 2921 2920 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8231 2921 2920 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8232 1 2927 2926 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8233 2927 2926 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8234 1 2929 2928 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8235 2929 2928 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8236 0 2923 2922 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8237 2923 2922 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8238 0 2925 2924 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8239 2925 2924 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8240 0 2927 2926 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8241 2927 2926 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8242 0 2929 2928 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8243 2929 2928 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8244 300 500 2922 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8245 301 500 2923 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8246 302 500 2924 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8247 303 500 2925 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8248 304 500 2926 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8249 305 500 2927 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8250 306 500 2928 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8251 307 500 2929 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8252 2930 504 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8253 2931 504 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8254 2932 504 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8255 2933 504 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8256 2934 504 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8257 2935 504 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8258 2936 504 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8259 2937 504 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8260 0 2931 2930 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8261 2931 2930 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8262 0 2933 2932 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8263 2933 2932 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8264 0 2935 2934 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8265 2935 2934 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8266 0 2937 2936 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8267 2937 2936 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8268 1 2931 2930 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8269 2931 2930 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8270 1 2933 2932 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8271 2933 2932 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8272 1 2935 2934 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8273 2935 2934 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8274 1 2937 2936 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8275 2937 2936 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8276 1 2939 2938 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8277 2939 2938 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8278 1 2941 2940 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8279 2941 2940 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8280 1 2943 2942 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8281 2943 2942 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8282 1 2945 2944 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8283 2945 2944 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8284 0 2939 2938 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8285 2939 2938 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8286 0 2941 2940 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8287 2941 2940 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8288 0 2943 2942 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8289 2943 2942 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8290 0 2945 2944 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8291 2945 2944 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8292 300 508 2938 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8293 301 508 2939 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8294 302 508 2940 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8295 303 508 2941 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8296 304 508 2942 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8297 305 508 2943 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8298 306 508 2944 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8299 307 508 2945 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8300 2946 511 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8301 2947 511 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8302 2948 511 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8303 2949 511 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8304 2950 511 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8305 2951 511 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8306 2952 511 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8307 2953 511 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8308 0 2947 2946 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8309 2947 2946 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8310 0 2949 2948 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8311 2949 2948 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8312 0 2951 2950 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8313 2951 2950 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8314 0 2953 2952 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8315 2953 2952 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8316 1 2947 2946 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8317 2947 2946 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8318 1 2949 2948 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8319 2949 2948 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8320 1 2955 2954 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8321 2955 2954 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8322 1 2957 2956 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8323 2957 2956 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8324 1 2951 2950 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8325 2951 2950 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8326 1 2953 2952 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8327 2953 2952 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8328 1 2959 2958 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8329 2959 2958 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8330 1 2961 2960 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8331 2961 2960 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8332 0 2955 2954 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8333 2955 2954 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8334 0 2957 2956 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8335 2957 2956 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8336 0 2959 2958 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8337 2959 2958 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8338 0 2961 2960 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8339 2961 2960 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8340 300 516 2954 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8341 301 516 2955 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8342 302 516 2956 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8343 303 516 2957 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8344 304 516 2958 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8345 305 516 2959 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8346 306 516 2960 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8347 307 516 2961 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8348 2962 520 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8349 2963 520 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8350 2964 520 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8351 2965 520 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8352 2966 520 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8353 2967 520 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8354 2968 520 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8355 2969 520 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8356 0 2963 2962 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8357 2963 2962 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8358 0 2965 2964 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8359 2965 2964 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8360 0 2967 2966 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8361 2967 2966 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8362 0 2969 2968 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8363 2969 2968 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8364 1 2963 2962 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8365 2963 2962 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8366 1 2965 2964 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8367 2965 2964 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8368 1 2967 2966 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8369 2967 2966 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8370 1 2969 2968 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8371 2969 2968 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8372 1 2971 2970 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8373 2971 2970 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8374 1 2973 2972 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8375 2973 2972 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8376 1 2975 2974 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8377 2975 2974 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8378 1 2977 2976 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8379 2977 2976 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8380 0 2971 2970 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8381 2971 2970 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8382 0 2973 2972 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8383 2973 2972 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8384 0 2975 2974 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8385 2975 2974 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8386 0 2977 2976 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8387 2977 2976 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8388 300 524 2970 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8389 301 524 2971 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8390 302 524 2972 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8391 303 524 2973 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8392 304 524 2974 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8393 305 524 2975 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8394 306 524 2976 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8395 307 524 2977 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8396 2978 527 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8397 2979 527 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8398 2980 527 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8399 2981 527 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8400 2982 527 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8401 2983 527 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8402 2984 527 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8403 2985 527 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8404 0 2979 2978 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8405 2979 2978 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8406 0 2981 2980 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8407 2981 2980 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8408 0 2983 2982 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8409 2983 2982 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8410 0 2985 2984 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8411 2985 2984 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8412 1 2979 2978 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8413 2979 2978 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8414 1 2981 2980 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8415 2981 2980 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8416 1 2987 2986 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8417 2987 2986 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8418 1 2989 2988 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8419 2989 2988 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8420 1 2983 2982 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8421 2983 2982 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8422 1 2985 2984 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8423 2985 2984 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8424 1 2991 2990 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8425 2991 2990 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8426 1 2993 2992 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8427 2993 2992 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8428 0 2987 2986 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8429 2987 2986 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8430 0 2989 2988 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8431 2989 2988 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8432 0 2991 2990 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8433 2991 2990 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8434 0 2993 2992 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8435 2993 2992 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8436 300 532 2986 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8437 301 532 2987 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8438 302 532 2988 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8439 303 532 2989 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8440 304 532 2990 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8441 305 532 2991 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8442 306 532 2992 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8443 307 532 2993 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8444 2994 536 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8445 2995 536 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8446 2996 536 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8447 2997 536 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8448 2998 536 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8449 2999 536 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8450 3000 536 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8451 3001 536 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8452 0 2995 2994 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8453 2995 2994 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8454 0 2997 2996 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8455 2997 2996 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8456 0 2999 2998 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8457 2999 2998 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8458 0 3001 3000 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8459 3001 3000 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8460 1 2995 2994 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8461 2995 2994 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8462 1 2997 2996 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8463 2997 2996 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8464 1 2999 2998 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8465 2999 2998 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8466 1 3001 3000 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8467 3001 3000 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8468 1 3003 3002 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8469 3003 3002 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8470 1 3005 3004 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8471 3005 3004 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8472 1 3007 3006 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8473 3007 3006 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8474 1 3009 3008 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8475 3009 3008 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8476 0 3003 3002 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8477 3003 3002 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8478 0 3005 3004 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8479 3005 3004 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8480 0 3007 3006 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8481 3007 3006 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8482 0 3009 3008 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8483 3009 3008 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8484 300 540 3002 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8485 301 540 3003 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8486 302 540 3004 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8487 303 540 3005 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8488 304 540 3006 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8489 305 540 3007 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8490 306 540 3008 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8491 307 540 3009 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8492 3010 543 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8493 3011 543 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8494 3012 543 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8495 3013 543 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8496 3014 543 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8497 3015 543 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8498 3016 543 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8499 3017 543 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8500 0 3011 3010 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8501 3011 3010 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8502 0 3013 3012 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8503 3013 3012 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8504 0 3015 3014 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8505 3015 3014 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8506 0 3017 3016 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8507 3017 3016 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8508 1 3011 3010 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8509 3011 3010 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8510 1 3013 3012 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8511 3013 3012 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8512 1 3019 3018 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8513 3019 3018 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8514 1 3021 3020 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8515 3021 3020 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8516 1 3015 3014 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8517 3015 3014 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8518 1 3017 3016 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8519 3017 3016 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8520 1 3023 3022 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8521 3023 3022 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8522 1 3025 3024 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8523 3025 3024 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8524 0 3019 3018 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8525 3019 3018 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8526 0 3021 3020 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8527 3021 3020 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8528 0 3023 3022 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8529 3023 3022 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8530 0 3025 3024 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8531 3025 3024 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8532 300 548 3018 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8533 301 548 3019 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8534 302 548 3020 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8535 303 548 3021 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8536 304 548 3022 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8537 305 548 3023 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8538 306 548 3024 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8539 307 548 3025 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8540 3026 552 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8541 3027 552 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8542 3028 552 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8543 3029 552 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8544 3030 552 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8545 3031 552 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8546 3032 552 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8547 3033 552 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8548 0 3027 3026 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8549 3027 3026 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8550 0 3029 3028 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8551 3029 3028 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8552 0 3031 3030 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8553 3031 3030 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8554 0 3033 3032 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8555 3033 3032 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8556 1 3027 3026 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8557 3027 3026 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8558 1 3029 3028 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8559 3029 3028 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8560 1 3031 3030 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8561 3031 3030 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8562 1 3033 3032 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8563 3033 3032 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8564 1 3035 3034 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8565 3035 3034 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8566 1 3037 3036 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8567 3037 3036 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8568 1 3039 3038 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8569 3039 3038 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8570 1 3041 3040 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8571 3041 3040 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8572 0 3035 3034 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8573 3035 3034 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8574 0 3037 3036 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8575 3037 3036 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8576 0 3039 3038 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8577 3039 3038 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8578 0 3041 3040 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8579 3041 3040 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8580 300 556 3034 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8581 301 556 3035 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8582 302 556 3036 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8583 303 556 3037 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8584 304 556 3038 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8585 305 556 3039 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8586 306 556 3040 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8587 307 556 3041 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8588 3042 559 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8589 3043 559 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8590 3044 559 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8591 3045 559 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8592 3046 559 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8593 3047 559 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8594 3048 559 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8595 3049 559 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8596 0 3043 3042 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8597 3043 3042 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8598 0 3045 3044 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8599 3045 3044 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8600 0 3047 3046 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8601 3047 3046 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8602 0 3049 3048 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8603 3049 3048 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8604 1 3043 3042 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8605 3043 3042 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8606 1 3045 3044 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8607 3045 3044 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8608 1 3051 3050 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8609 3051 3050 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8610 1 3053 3052 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8611 3053 3052 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8612 1 3047 3046 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8613 3047 3046 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8614 1 3049 3048 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8615 3049 3048 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8616 1 3055 3054 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8617 3055 3054 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8618 1 3057 3056 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8619 3057 3056 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8620 0 3051 3050 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8621 3051 3050 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8622 0 3053 3052 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8623 3053 3052 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8624 0 3055 3054 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8625 3055 3054 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8626 0 3057 3056 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8627 3057 3056 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8628 300 564 3050 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8629 301 564 3051 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8630 302 564 3052 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8631 303 564 3053 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8632 304 564 3054 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8633 305 564 3055 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8634 306 564 3056 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8635 307 564 3057 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8636 3058 568 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8637 3059 568 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8638 3060 568 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8639 3061 568 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8640 3062 568 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8641 3063 568 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8642 3064 568 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8643 3065 568 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8644 0 3059 3058 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8645 3059 3058 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8646 0 3061 3060 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8647 3061 3060 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8648 0 3063 3062 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8649 3063 3062 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8650 0 3065 3064 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8651 3065 3064 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8652 1 3059 3058 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8653 3059 3058 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8654 1 3061 3060 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8655 3061 3060 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8656 1 3063 3062 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8657 3063 3062 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8658 1 3065 3064 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8659 3065 3064 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8660 1 3067 3066 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8661 3067 3066 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8662 1 3069 3068 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8663 3069 3068 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8664 1 3071 3070 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8665 3071 3070 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8666 1 3073 3072 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8667 3073 3072 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8668 0 3067 3066 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8669 3067 3066 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8670 0 3069 3068 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8671 3069 3068 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8672 0 3071 3070 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8673 3071 3070 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8674 0 3073 3072 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8675 3073 3072 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8676 300 572 3066 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8677 301 572 3067 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8678 302 572 3068 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8679 303 572 3069 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8680 304 572 3070 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8681 305 572 3071 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8682 306 572 3072 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8683 307 572 3073 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8684 3074 575 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8685 3075 575 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8686 3076 575 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8687 3077 575 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8688 3078 575 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8689 3079 575 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8690 3080 575 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8691 3081 575 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8692 0 3075 3074 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8693 3075 3074 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8694 0 3077 3076 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8695 3077 3076 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8696 0 3079 3078 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8697 3079 3078 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8698 0 3081 3080 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8699 3081 3080 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8700 1 3075 3074 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8701 3075 3074 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8702 1 3077 3076 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8703 3077 3076 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8704 1 3083 3082 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8705 3083 3082 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8706 1 3085 3084 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8707 3085 3084 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8708 1 3079 3078 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8709 3079 3078 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8710 1 3081 3080 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8711 3081 3080 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8712 1 3087 3086 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8713 3087 3086 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8714 1 3089 3088 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8715 3089 3088 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8716 0 3083 3082 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8717 3083 3082 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8718 0 3085 3084 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8719 3085 3084 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8720 0 3087 3086 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8721 3087 3086 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8722 0 3089 3088 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8723 3089 3088 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8724 300 580 3082 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8725 301 580 3083 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8726 302 580 3084 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8727 303 580 3085 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8728 304 580 3086 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8729 305 580 3087 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8730 306 580 3088 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8731 307 580 3089 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8732 3090 584 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8733 3091 584 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8734 3092 584 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8735 3093 584 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8736 3094 584 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8737 3095 584 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8738 3096 584 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8739 3097 584 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8740 0 3091 3090 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8741 3091 3090 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8742 0 3093 3092 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8743 3093 3092 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8744 0 3095 3094 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8745 3095 3094 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8746 0 3097 3096 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8747 3097 3096 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8748 1 3091 3090 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8749 3091 3090 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8750 1 3093 3092 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8751 3093 3092 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8752 1 3095 3094 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8753 3095 3094 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8754 1 3097 3096 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8755 3097 3096 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8756 1 3099 3098 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8757 3099 3098 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8758 1 3101 3100 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8759 3101 3100 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8760 1 3103 3102 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8761 3103 3102 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8762 1 3105 3104 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8763 3105 3104 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8764 0 3099 3098 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8765 3099 3098 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8766 0 3101 3100 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8767 3101 3100 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8768 0 3103 3102 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8769 3103 3102 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8770 0 3105 3104 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8771 3105 3104 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8772 300 588 3098 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8773 301 588 3099 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8774 302 588 3100 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8775 303 588 3101 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8776 304 588 3102 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8777 305 588 3103 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8778 306 588 3104 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8779 307 588 3105 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8780 3106 591 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8781 3107 591 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8782 3108 591 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8783 3109 591 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8784 3110 591 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8785 3111 591 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8786 3112 591 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8787 3113 591 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8788 0 3107 3106 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8789 3107 3106 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8790 0 3109 3108 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8791 3109 3108 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8792 0 3111 3110 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8793 3111 3110 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8794 0 3113 3112 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8795 3113 3112 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8796 1 3107 3106 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8797 3107 3106 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8798 1 3109 3108 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8799 3109 3108 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8800 1 3115 3114 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8801 3115 3114 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8802 1 3117 3116 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8803 3117 3116 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8804 1 3111 3110 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8805 3111 3110 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8806 1 3113 3112 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8807 3113 3112 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8808 1 3119 3118 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8809 3119 3118 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8810 1 3121 3120 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8811 3121 3120 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8812 0 3115 3114 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8813 3115 3114 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8814 0 3117 3116 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8815 3117 3116 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8816 0 3119 3118 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8817 3119 3118 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8818 0 3121 3120 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8819 3121 3120 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8820 300 596 3114 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8821 301 596 3115 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8822 302 596 3116 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8823 303 596 3117 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8824 304 596 3118 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8825 305 596 3119 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8826 306 596 3120 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8827 307 596 3121 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8828 3122 600 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8829 3123 600 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8830 3124 600 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8831 3125 600 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8832 3126 600 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8833 3127 600 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8834 3128 600 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8835 3129 600 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8836 0 3123 3122 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8837 3123 3122 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8838 0 3125 3124 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8839 3125 3124 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8840 0 3127 3126 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8841 3127 3126 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8842 0 3129 3128 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8843 3129 3128 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8844 1 3123 3122 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8845 3123 3122 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8846 1 3125 3124 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8847 3125 3124 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8848 1 3127 3126 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8849 3127 3126 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8850 1 3129 3128 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8851 3129 3128 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8852 1 3131 3130 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8853 3131 3130 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8854 1 3133 3132 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8855 3133 3132 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8856 1 3135 3134 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8857 3135 3134 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8858 1 3137 3136 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8859 3137 3136 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8860 0 3131 3130 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8861 3131 3130 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8862 0 3133 3132 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8863 3133 3132 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8864 0 3135 3134 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8865 3135 3134 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8866 0 3137 3136 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8867 3137 3136 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8868 300 604 3130 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8869 301 604 3131 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8870 302 604 3132 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8871 303 604 3133 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8872 304 604 3134 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8873 305 604 3135 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8874 306 604 3136 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8875 307 604 3137 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8876 3138 607 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8877 3139 607 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8878 3140 607 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8879 3141 607 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8880 3142 607 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8881 3143 607 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8882 3144 607 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8883 3145 607 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8884 0 3139 3138 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8885 3139 3138 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8886 0 3141 3140 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8887 3141 3140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8888 0 3143 3142 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8889 3143 3142 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8890 0 3145 3144 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8891 3145 3144 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8892 1 3139 3138 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8893 3139 3138 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8894 1 3141 3140 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8895 3141 3140 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8896 1 3147 3146 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8897 3147 3146 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8898 1 3149 3148 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8899 3149 3148 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8900 1 3143 3142 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8901 3143 3142 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8902 1 3145 3144 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8903 3145 3144 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8904 1 3151 3150 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8905 3151 3150 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8906 1 3153 3152 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8907 3153 3152 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8908 0 3147 3146 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8909 3147 3146 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8910 0 3149 3148 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8911 3149 3148 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8912 0 3151 3150 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8913 3151 3150 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8914 0 3153 3152 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8915 3153 3152 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8916 300 612 3146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8917 301 612 3147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8918 302 612 3148 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8919 303 612 3149 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8920 304 612 3150 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8921 305 612 3151 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8922 306 612 3152 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8923 307 612 3153 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8924 3154 616 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8925 3155 616 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8926 3156 616 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8927 3157 616 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8928 3158 616 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8929 3159 616 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8930 3160 616 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8931 3161 616 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8932 0 3155 3154 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8933 3155 3154 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8934 0 3157 3156 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8935 3157 3156 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8936 0 3159 3158 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8937 3159 3158 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8938 0 3161 3160 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8939 3161 3160 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8940 1 3155 3154 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8941 3155 3154 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8942 1 3157 3156 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8943 3157 3156 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8944 1 3159 3158 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8945 3159 3158 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8946 1 3161 3160 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8947 3161 3160 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8948 1 3163 3162 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8949 3163 3162 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8950 1 3165 3164 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8951 3165 3164 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8952 1 3167 3166 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8953 3167 3166 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8954 1 3169 3168 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m8955 3169 3168 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8956 0 3163 3162 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8957 3163 3162 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8958 0 3165 3164 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8959 3165 3164 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8960 0 3167 3166 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8961 3167 3166 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8962 0 3169 3168 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8963 3169 3168 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8964 300 620 3162 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m8965 301 620 3163 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8966 302 620 3164 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8967 303 620 3165 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8968 304 620 3166 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m8969 305 620 3167 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m8970 306 620 3168 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m8971 307 620 3169 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m8972 3170 624 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m8973 3171 624 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8974 3172 624 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8975 3173 624 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8976 3174 624 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m8977 3175 624 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m8978 3176 624 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m8979 3177 624 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m8980 0 3171 3170 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8981 3171 3170 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8982 0 3173 3172 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m8983 3173 3172 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m8984 0 3175 3174 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8985 3175 3174 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8986 0 3177 3176 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m8987 3177 3176 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m8988 1 3171 3170 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8989 3171 3170 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8990 1 3173 3172 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8991 3173 3172 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8992 1 3179 3178 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8993 3179 3178 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m8994 1 3181 3180 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8995 3181 3180 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8996 1 3175 3174 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8997 3175 3174 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m8998 1 3177 3176 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m8999 3177 3176 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9000 1 3183 3182 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9001 3183 3182 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9002 1 3185 3184 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9003 3185 3184 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9004 0 3179 3178 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9005 3179 3178 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9006 0 3181 3180 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9007 3181 3180 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9008 0 3183 3182 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9009 3183 3182 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9010 0 3185 3184 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9011 3185 3184 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9012 300 628 3178 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9013 301 628 3179 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9014 302 628 3180 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9015 303 628 3181 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9016 304 628 3182 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9017 305 628 3183 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9018 306 628 3184 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9019 307 628 3185 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9020 3186 632 300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9021 3187 632 301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9022 3188 632 302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9023 3189 632 303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9024 3190 632 304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9025 3191 632 305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9026 3192 632 306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9027 3193 632 307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9028 0 3187 3186 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9029 3187 3186 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9030 0 3189 3188 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9031 3189 3188 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9032 0 3191 3190 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9033 3191 3190 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9034 0 3193 3192 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9035 3193 3192 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9036 1 3187 3186 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9037 3187 3186 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9038 1 3189 3188 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9039 3189 3188 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9040 1 3191 3190 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9041 3191 3190 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9042 1 3193 3192 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9043 3193 3192 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9044 1 3195 3194 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9045 3195 3194 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9046 1 3197 3196 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9047 3197 3196 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9048 1 3199 3198 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9049 3199 3198 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9050 1 3201 3200 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9051 3201 3200 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9052 0 3195 3194 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9053 3195 3194 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9054 0 3197 3196 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9055 3197 3196 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9056 0 3199 3198 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9057 3199 3198 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9058 0 3201 3200 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9059 3201 3200 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9060 326 380 3194 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9061 327 380 3195 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9062 328 380 3196 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9063 329 380 3197 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9064 330 380 3198 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9065 331 380 3199 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9066 332 380 3200 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9067 333 380 3201 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9068 3202 383 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9069 3203 383 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9070 3204 383 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9071 3205 383 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9072 3206 383 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9073 3207 383 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9074 3208 383 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9075 3209 383 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9076 0 3203 3202 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9077 3203 3202 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9078 0 3205 3204 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9079 3205 3204 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9080 0 3207 3206 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9081 3207 3206 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9082 0 3209 3208 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9083 3209 3208 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9084 1 3203 3202 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9085 3203 3202 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9086 1 3205 3204 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9087 3205 3204 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9088 1 3211 3210 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9089 3211 3210 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9090 1 3213 3212 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9091 3213 3212 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9092 1 3207 3206 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9093 3207 3206 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9094 1 3209 3208 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9095 3209 3208 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9096 1 3215 3214 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9097 3215 3214 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9098 1 3217 3216 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9099 3217 3216 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9100 0 3211 3210 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9101 3211 3210 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9102 0 3213 3212 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9103 3213 3212 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9104 0 3215 3214 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9105 3215 3214 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9106 0 3217 3216 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9107 3217 3216 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9108 326 388 3210 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9109 327 388 3211 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9110 328 388 3212 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9111 329 388 3213 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9112 330 388 3214 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9113 331 388 3215 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9114 332 388 3216 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9115 333 388 3217 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9116 3218 392 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9117 3219 392 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9118 3220 392 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9119 3221 392 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9120 3222 392 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9121 3223 392 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9122 3224 392 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9123 3225 392 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9124 0 3219 3218 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9125 3219 3218 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9126 0 3221 3220 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9127 3221 3220 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9128 0 3223 3222 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9129 3223 3222 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9130 0 3225 3224 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9131 3225 3224 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9132 1 3219 3218 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9133 3219 3218 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9134 1 3221 3220 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9135 3221 3220 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9136 1 3223 3222 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9137 3223 3222 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9138 1 3225 3224 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9139 3225 3224 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9140 1 3227 3226 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9141 3227 3226 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9142 1 3229 3228 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9143 3229 3228 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9144 1 3231 3230 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9145 3231 3230 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9146 1 3233 3232 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9147 3233 3232 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9148 0 3227 3226 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9149 3227 3226 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9150 0 3229 3228 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9151 3229 3228 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9152 0 3231 3230 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9153 3231 3230 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9154 0 3233 3232 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9155 3233 3232 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9156 326 396 3226 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9157 327 396 3227 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9158 328 396 3228 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9159 329 396 3229 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9160 330 396 3230 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9161 331 396 3231 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9162 332 396 3232 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9163 333 396 3233 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9164 3234 399 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9165 3235 399 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9166 3236 399 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9167 3237 399 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9168 3238 399 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9169 3239 399 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9170 3240 399 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9171 3241 399 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9172 0 3235 3234 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9173 3235 3234 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9174 0 3237 3236 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9175 3237 3236 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9176 0 3239 3238 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9177 3239 3238 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9178 0 3241 3240 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9179 3241 3240 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9180 1 3235 3234 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9181 3235 3234 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9182 1 3237 3236 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9183 3237 3236 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9184 1 3243 3242 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9185 3243 3242 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9186 1 3245 3244 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9187 3245 3244 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9188 1 3239 3238 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9189 3239 3238 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9190 1 3241 3240 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9191 3241 3240 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9192 1 3247 3246 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9193 3247 3246 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9194 1 3249 3248 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9195 3249 3248 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9196 0 3243 3242 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9197 3243 3242 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9198 0 3245 3244 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9199 3245 3244 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9200 0 3247 3246 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9201 3247 3246 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9202 0 3249 3248 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9203 3249 3248 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9204 326 404 3242 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9205 327 404 3243 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9206 328 404 3244 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9207 329 404 3245 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9208 330 404 3246 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9209 331 404 3247 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9210 332 404 3248 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9211 333 404 3249 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9212 3250 408 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9213 3251 408 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9214 3252 408 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9215 3253 408 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9216 3254 408 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9217 3255 408 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9218 3256 408 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9219 3257 408 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9220 0 3251 3250 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9221 3251 3250 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9222 0 3253 3252 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9223 3253 3252 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9224 0 3255 3254 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9225 3255 3254 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9226 0 3257 3256 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9227 3257 3256 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9228 1 3251 3250 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9229 3251 3250 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9230 1 3253 3252 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9231 3253 3252 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9232 1 3255 3254 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9233 3255 3254 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9234 1 3257 3256 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9235 3257 3256 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9236 1 3259 3258 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9237 3259 3258 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9238 1 3261 3260 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9239 3261 3260 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9240 1 3263 3262 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9241 3263 3262 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9242 1 3265 3264 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9243 3265 3264 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9244 0 3259 3258 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9245 3259 3258 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9246 0 3261 3260 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9247 3261 3260 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9248 0 3263 3262 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9249 3263 3262 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9250 0 3265 3264 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9251 3265 3264 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9252 326 412 3258 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9253 327 412 3259 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9254 328 412 3260 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9255 329 412 3261 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9256 330 412 3262 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9257 331 412 3263 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9258 332 412 3264 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9259 333 412 3265 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9260 3266 415 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9261 3267 415 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9262 3268 415 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9263 3269 415 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9264 3270 415 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9265 3271 415 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9266 3272 415 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9267 3273 415 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9268 0 3267 3266 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9269 3267 3266 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9270 0 3269 3268 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9271 3269 3268 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9272 0 3271 3270 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9273 3271 3270 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9274 0 3273 3272 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9275 3273 3272 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9276 1 3267 3266 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9277 3267 3266 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9278 1 3269 3268 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9279 3269 3268 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9280 1 3275 3274 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9281 3275 3274 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9282 1 3277 3276 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9283 3277 3276 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9284 1 3271 3270 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9285 3271 3270 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9286 1 3273 3272 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9287 3273 3272 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9288 1 3279 3278 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9289 3279 3278 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9290 1 3281 3280 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9291 3281 3280 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9292 0 3275 3274 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9293 3275 3274 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9294 0 3277 3276 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9295 3277 3276 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9296 0 3279 3278 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9297 3279 3278 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9298 0 3281 3280 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9299 3281 3280 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9300 326 420 3274 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9301 327 420 3275 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9302 328 420 3276 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9303 329 420 3277 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9304 330 420 3278 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9305 331 420 3279 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9306 332 420 3280 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9307 333 420 3281 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9308 3282 424 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9309 3283 424 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9310 3284 424 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9311 3285 424 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9312 3286 424 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9313 3287 424 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9314 3288 424 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9315 3289 424 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9316 0 3283 3282 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9317 3283 3282 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9318 0 3285 3284 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9319 3285 3284 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9320 0 3287 3286 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9321 3287 3286 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9322 0 3289 3288 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9323 3289 3288 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9324 1 3283 3282 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9325 3283 3282 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9326 1 3285 3284 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9327 3285 3284 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9328 1 3287 3286 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9329 3287 3286 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9330 1 3289 3288 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9331 3289 3288 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9332 1 3291 3290 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9333 3291 3290 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9334 1 3293 3292 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9335 3293 3292 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9336 1 3295 3294 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9337 3295 3294 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9338 1 3297 3296 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9339 3297 3296 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9340 0 3291 3290 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9341 3291 3290 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9342 0 3293 3292 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9343 3293 3292 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9344 0 3295 3294 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9345 3295 3294 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9346 0 3297 3296 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9347 3297 3296 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9348 326 428 3290 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9349 327 428 3291 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9350 328 428 3292 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9351 329 428 3293 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9352 330 428 3294 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9353 331 428 3295 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9354 332 428 3296 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9355 333 428 3297 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9356 3298 431 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9357 3299 431 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9358 3300 431 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9359 3301 431 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9360 3302 431 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9361 3303 431 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9362 3304 431 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9363 3305 431 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9364 0 3299 3298 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9365 3299 3298 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9366 0 3301 3300 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9367 3301 3300 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9368 0 3303 3302 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9369 3303 3302 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9370 0 3305 3304 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9371 3305 3304 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9372 1 3299 3298 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9373 3299 3298 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9374 1 3301 3300 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9375 3301 3300 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9376 1 3307 3306 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9377 3307 3306 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9378 1 3309 3308 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9379 3309 3308 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9380 1 3303 3302 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9381 3303 3302 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9382 1 3305 3304 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9383 3305 3304 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9384 1 3311 3310 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9385 3311 3310 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9386 1 3313 3312 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9387 3313 3312 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9388 0 3307 3306 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9389 3307 3306 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9390 0 3309 3308 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9391 3309 3308 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9392 0 3311 3310 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9393 3311 3310 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9394 0 3313 3312 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9395 3313 3312 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9396 326 436 3306 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9397 327 436 3307 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9398 328 436 3308 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9399 329 436 3309 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9400 330 436 3310 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9401 331 436 3311 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9402 332 436 3312 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9403 333 436 3313 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9404 3314 440 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9405 3315 440 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9406 3316 440 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9407 3317 440 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9408 3318 440 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9409 3319 440 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9410 3320 440 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9411 3321 440 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9412 0 3315 3314 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9413 3315 3314 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9414 0 3317 3316 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9415 3317 3316 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9416 0 3319 3318 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9417 3319 3318 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9418 0 3321 3320 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9419 3321 3320 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9420 1 3315 3314 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9421 3315 3314 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9422 1 3317 3316 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9423 3317 3316 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9424 1 3319 3318 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9425 3319 3318 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9426 1 3321 3320 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9427 3321 3320 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9428 1 3323 3322 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9429 3323 3322 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9430 1 3325 3324 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9431 3325 3324 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9432 1 3327 3326 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9433 3327 3326 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9434 1 3329 3328 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9435 3329 3328 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9436 0 3323 3322 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9437 3323 3322 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9438 0 3325 3324 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9439 3325 3324 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9440 0 3327 3326 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9441 3327 3326 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9442 0 3329 3328 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9443 3329 3328 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9444 326 444 3322 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9445 327 444 3323 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9446 328 444 3324 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9447 329 444 3325 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9448 330 444 3326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9449 331 444 3327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9450 332 444 3328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9451 333 444 3329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9452 3330 447 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9453 3331 447 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9454 3332 447 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9455 3333 447 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9456 3334 447 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9457 3335 447 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9458 3336 447 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9459 3337 447 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9460 0 3331 3330 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9461 3331 3330 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9462 0 3333 3332 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9463 3333 3332 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9464 0 3335 3334 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9465 3335 3334 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9466 0 3337 3336 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9467 3337 3336 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9468 1 3331 3330 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9469 3331 3330 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9470 1 3333 3332 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9471 3333 3332 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9472 1 3339 3338 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9473 3339 3338 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9474 1 3341 3340 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9475 3341 3340 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9476 1 3335 3334 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9477 3335 3334 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9478 1 3337 3336 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9479 3337 3336 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9480 1 3343 3342 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9481 3343 3342 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9482 1 3345 3344 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9483 3345 3344 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9484 0 3339 3338 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9485 3339 3338 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9486 0 3341 3340 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9487 3341 3340 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9488 0 3343 3342 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9489 3343 3342 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9490 0 3345 3344 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9491 3345 3344 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9492 326 452 3338 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9493 327 452 3339 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9494 328 452 3340 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9495 329 452 3341 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9496 330 452 3342 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9497 331 452 3343 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9498 332 452 3344 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9499 333 452 3345 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9500 3346 456 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9501 3347 456 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9502 3348 456 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9503 3349 456 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9504 3350 456 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9505 3351 456 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9506 3352 456 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9507 3353 456 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9508 0 3347 3346 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9509 3347 3346 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9510 0 3349 3348 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9511 3349 3348 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9512 0 3351 3350 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9513 3351 3350 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9514 0 3353 3352 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9515 3353 3352 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9516 1 3347 3346 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9517 3347 3346 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9518 1 3349 3348 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9519 3349 3348 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9520 1 3351 3350 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9521 3351 3350 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9522 1 3353 3352 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9523 3353 3352 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9524 1 3355 3354 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9525 3355 3354 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9526 1 3357 3356 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9527 3357 3356 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9528 1 3359 3358 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9529 3359 3358 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9530 1 3361 3360 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9531 3361 3360 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9532 0 3355 3354 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9533 3355 3354 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9534 0 3357 3356 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9535 3357 3356 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9536 0 3359 3358 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9537 3359 3358 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9538 0 3361 3360 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9539 3361 3360 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9540 326 460 3354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9541 327 460 3355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9542 328 460 3356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9543 329 460 3357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9544 330 460 3358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9545 331 460 3359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9546 332 460 3360 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9547 333 460 3361 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9548 3362 463 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9549 3363 463 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9550 3364 463 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9551 3365 463 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9552 3366 463 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9553 3367 463 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9554 3368 463 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9555 3369 463 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9556 0 3363 3362 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9557 3363 3362 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9558 0 3365 3364 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9559 3365 3364 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9560 0 3367 3366 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9561 3367 3366 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9562 0 3369 3368 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9563 3369 3368 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9564 1 3363 3362 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9565 3363 3362 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9566 1 3365 3364 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9567 3365 3364 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9568 1 3371 3370 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9569 3371 3370 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9570 1 3373 3372 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9571 3373 3372 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9572 1 3367 3366 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9573 3367 3366 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9574 1 3369 3368 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9575 3369 3368 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9576 1 3375 3374 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9577 3375 3374 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9578 1 3377 3376 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9579 3377 3376 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9580 0 3371 3370 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9581 3371 3370 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9582 0 3373 3372 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9583 3373 3372 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9584 0 3375 3374 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9585 3375 3374 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9586 0 3377 3376 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9587 3377 3376 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9588 326 468 3370 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9589 327 468 3371 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9590 328 468 3372 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9591 329 468 3373 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9592 330 468 3374 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9593 331 468 3375 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9594 332 468 3376 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9595 333 468 3377 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9596 3378 472 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9597 3379 472 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9598 3380 472 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9599 3381 472 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9600 3382 472 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9601 3383 472 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9602 3384 472 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9603 3385 472 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9604 0 3379 3378 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9605 3379 3378 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9606 0 3381 3380 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9607 3381 3380 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9608 0 3383 3382 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9609 3383 3382 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9610 0 3385 3384 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9611 3385 3384 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9612 1 3379 3378 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9613 3379 3378 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9614 1 3381 3380 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9615 3381 3380 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9616 1 3383 3382 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9617 3383 3382 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9618 1 3385 3384 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9619 3385 3384 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9620 1 3387 3386 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9621 3387 3386 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9622 1 3389 3388 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9623 3389 3388 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9624 1 3391 3390 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9625 3391 3390 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9626 1 3393 3392 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9627 3393 3392 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9628 0 3387 3386 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9629 3387 3386 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9630 0 3389 3388 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9631 3389 3388 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9632 0 3391 3390 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9633 3391 3390 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9634 0 3393 3392 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9635 3393 3392 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9636 326 476 3386 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9637 327 476 3387 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9638 328 476 3388 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9639 329 476 3389 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9640 330 476 3390 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9641 331 476 3391 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9642 332 476 3392 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9643 333 476 3393 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9644 3394 479 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9645 3395 479 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9646 3396 479 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9647 3397 479 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9648 3398 479 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9649 3399 479 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9650 3400 479 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9651 3401 479 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9652 0 3395 3394 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9653 3395 3394 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9654 0 3397 3396 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9655 3397 3396 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9656 0 3399 3398 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9657 3399 3398 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9658 0 3401 3400 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9659 3401 3400 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9660 1 3395 3394 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9661 3395 3394 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9662 1 3397 3396 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9663 3397 3396 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9664 1 3403 3402 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9665 3403 3402 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9666 1 3405 3404 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9667 3405 3404 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9668 1 3399 3398 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9669 3399 3398 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9670 1 3401 3400 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9671 3401 3400 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9672 1 3407 3406 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9673 3407 3406 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9674 1 3409 3408 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9675 3409 3408 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9676 0 3403 3402 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9677 3403 3402 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9678 0 3405 3404 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9679 3405 3404 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9680 0 3407 3406 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9681 3407 3406 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9682 0 3409 3408 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9683 3409 3408 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9684 326 484 3402 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9685 327 484 3403 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9686 328 484 3404 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9687 329 484 3405 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9688 330 484 3406 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9689 331 484 3407 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9690 332 484 3408 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9691 333 484 3409 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9692 3410 488 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9693 3411 488 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9694 3412 488 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9695 3413 488 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9696 3414 488 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9697 3415 488 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9698 3416 488 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9699 3417 488 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9700 0 3411 3410 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9701 3411 3410 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9702 0 3413 3412 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9703 3413 3412 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9704 0 3415 3414 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9705 3415 3414 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9706 0 3417 3416 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9707 3417 3416 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9708 1 3411 3410 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9709 3411 3410 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9710 1 3413 3412 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9711 3413 3412 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9712 1 3415 3414 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9713 3415 3414 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9714 1 3417 3416 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9715 3417 3416 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9716 1 3419 3418 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9717 3419 3418 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9718 1 3421 3420 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9719 3421 3420 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9720 1 3423 3422 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9721 3423 3422 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9722 1 3425 3424 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9723 3425 3424 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9724 0 3419 3418 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9725 3419 3418 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9726 0 3421 3420 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9727 3421 3420 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9728 0 3423 3422 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9729 3423 3422 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9730 0 3425 3424 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9731 3425 3424 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9732 326 492 3418 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9733 327 492 3419 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9734 328 492 3420 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9735 329 492 3421 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9736 330 492 3422 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9737 331 492 3423 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9738 332 492 3424 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9739 333 492 3425 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9740 3426 495 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9741 3427 495 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9742 3428 495 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9743 3429 495 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9744 3430 495 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9745 3431 495 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9746 3432 495 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9747 3433 495 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9748 0 3427 3426 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9749 3427 3426 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9750 0 3429 3428 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9751 3429 3428 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9752 0 3431 3430 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9753 3431 3430 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9754 0 3433 3432 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9755 3433 3432 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9756 1 3427 3426 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9757 3427 3426 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9758 1 3429 3428 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9759 3429 3428 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9760 1 3435 3434 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9761 3435 3434 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9762 1 3437 3436 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9763 3437 3436 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9764 1 3431 3430 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9765 3431 3430 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9766 1 3433 3432 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9767 3433 3432 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9768 1 3439 3438 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9769 3439 3438 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9770 1 3441 3440 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9771 3441 3440 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9772 0 3435 3434 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9773 3435 3434 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9774 0 3437 3436 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9775 3437 3436 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9776 0 3439 3438 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9777 3439 3438 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9778 0 3441 3440 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9779 3441 3440 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9780 326 500 3434 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9781 327 500 3435 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9782 328 500 3436 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9783 329 500 3437 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9784 330 500 3438 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9785 331 500 3439 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9786 332 500 3440 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9787 333 500 3441 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9788 3442 504 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9789 3443 504 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9790 3444 504 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9791 3445 504 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9792 3446 504 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9793 3447 504 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9794 3448 504 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9795 3449 504 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9796 0 3443 3442 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9797 3443 3442 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9798 0 3445 3444 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9799 3445 3444 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9800 0 3447 3446 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9801 3447 3446 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9802 0 3449 3448 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9803 3449 3448 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9804 1 3443 3442 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9805 3443 3442 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9806 1 3445 3444 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9807 3445 3444 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9808 1 3447 3446 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9809 3447 3446 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9810 1 3449 3448 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9811 3449 3448 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9812 1 3451 3450 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9813 3451 3450 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9814 1 3453 3452 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9815 3453 3452 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9816 1 3455 3454 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9817 3455 3454 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9818 1 3457 3456 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9819 3457 3456 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9820 0 3451 3450 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9821 3451 3450 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9822 0 3453 3452 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9823 3453 3452 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9824 0 3455 3454 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9825 3455 3454 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9826 0 3457 3456 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9827 3457 3456 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9828 326 508 3450 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9829 327 508 3451 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9830 328 508 3452 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9831 329 508 3453 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9832 330 508 3454 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9833 331 508 3455 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9834 332 508 3456 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9835 333 508 3457 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9836 3458 511 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9837 3459 511 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9838 3460 511 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9839 3461 511 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9840 3462 511 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9841 3463 511 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9842 3464 511 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9843 3465 511 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9844 0 3459 3458 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9845 3459 3458 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9846 0 3461 3460 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9847 3461 3460 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9848 0 3463 3462 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9849 3463 3462 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9850 0 3465 3464 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9851 3465 3464 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9852 1 3459 3458 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9853 3459 3458 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9854 1 3461 3460 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9855 3461 3460 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9856 1 3467 3466 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9857 3467 3466 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9858 1 3469 3468 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9859 3469 3468 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9860 1 3463 3462 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9861 3463 3462 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9862 1 3465 3464 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9863 3465 3464 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9864 1 3471 3470 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9865 3471 3470 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9866 1 3473 3472 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9867 3473 3472 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9868 0 3467 3466 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9869 3467 3466 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9870 0 3469 3468 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9871 3469 3468 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9872 0 3471 3470 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9873 3471 3470 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9874 0 3473 3472 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9875 3473 3472 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9876 326 516 3466 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9877 327 516 3467 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9878 328 516 3468 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9879 329 516 3469 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9880 330 516 3470 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9881 331 516 3471 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9882 332 516 3472 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9883 333 516 3473 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9884 3474 520 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9885 3475 520 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9886 3476 520 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9887 3477 520 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9888 3478 520 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9889 3479 520 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9890 3480 520 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9891 3481 520 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9892 0 3475 3474 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9893 3475 3474 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9894 0 3477 3476 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9895 3477 3476 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9896 0 3479 3478 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9897 3479 3478 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9898 0 3481 3480 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9899 3481 3480 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9900 1 3475 3474 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9901 3475 3474 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9902 1 3477 3476 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9903 3477 3476 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9904 1 3479 3478 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9905 3479 3478 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9906 1 3481 3480 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9907 3481 3480 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9908 1 3483 3482 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9909 3483 3482 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9910 1 3485 3484 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9911 3485 3484 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9912 1 3487 3486 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9913 3487 3486 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9914 1 3489 3488 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9915 3489 3488 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9916 0 3483 3482 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9917 3483 3482 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9918 0 3485 3484 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9919 3485 3484 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9920 0 3487 3486 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9921 3487 3486 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9922 0 3489 3488 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9923 3489 3488 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9924 326 524 3482 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9925 327 524 3483 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9926 328 524 3484 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9927 329 524 3485 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9928 330 524 3486 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9929 331 524 3487 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9930 332 524 3488 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9931 333 524 3489 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9932 3490 527 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9933 3491 527 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9934 3492 527 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9935 3493 527 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9936 3494 527 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9937 3495 527 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9938 3496 527 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9939 3497 527 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9940 0 3491 3490 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9941 3491 3490 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9942 0 3493 3492 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9943 3493 3492 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9944 0 3495 3494 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9945 3495 3494 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9946 0 3497 3496 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9947 3497 3496 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9948 1 3491 3490 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9949 3491 3490 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9950 1 3493 3492 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9951 3493 3492 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9952 1 3499 3498 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9953 3499 3498 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m9954 1 3501 3500 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9955 3501 3500 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9956 1 3495 3494 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9957 3495 3494 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9958 1 3497 3496 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9959 3497 3496 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9960 1 3503 3502 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9961 3503 3502 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9962 1 3505 3504 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m9963 3505 3504 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9964 0 3499 3498 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9965 3499 3498 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9966 0 3501 3500 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9967 3501 3500 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9968 0 3503 3502 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9969 3503 3502 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9970 0 3505 3504 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9971 3505 3504 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9972 326 532 3498 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m9973 327 532 3499 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9974 328 532 3500 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9975 329 532 3501 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9976 330 532 3502 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m9977 331 532 3503 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m9978 332 532 3504 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m9979 333 532 3505 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m9980 3506 536 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m9981 3507 536 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9982 3508 536 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9983 3509 536 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9984 3510 536 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m9985 3511 536 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m9986 3512 536 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m9987 3513 536 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m9988 0 3507 3506 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9989 3507 3506 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9990 0 3509 3508 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m9991 3509 3508 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m9992 0 3511 3510 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9993 3511 3510 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9994 0 3513 3512 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m9995 3513 3512 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m9996 1 3507 3506 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9997 3507 3506 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m9998 1 3509 3508 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m9999 3509 3508 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10000 1 3511 3510 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10001 3511 3510 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10002 1 3513 3512 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10003 3513 3512 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10004 1 3515 3514 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10005 3515 3514 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10006 1 3517 3516 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10007 3517 3516 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10008 1 3519 3518 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10009 3519 3518 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10010 1 3521 3520 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10011 3521 3520 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10012 0 3515 3514 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10013 3515 3514 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10014 0 3517 3516 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10015 3517 3516 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10016 0 3519 3518 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10017 3519 3518 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10018 0 3521 3520 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10019 3521 3520 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10020 326 540 3514 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10021 327 540 3515 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10022 328 540 3516 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10023 329 540 3517 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10024 330 540 3518 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10025 331 540 3519 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10026 332 540 3520 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10027 333 540 3521 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10028 3522 543 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10029 3523 543 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10030 3524 543 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10031 3525 543 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10032 3526 543 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10033 3527 543 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10034 3528 543 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10035 3529 543 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10036 0 3523 3522 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10037 3523 3522 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10038 0 3525 3524 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10039 3525 3524 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10040 0 3527 3526 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10041 3527 3526 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10042 0 3529 3528 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10043 3529 3528 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10044 1 3523 3522 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10045 3523 3522 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10046 1 3525 3524 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10047 3525 3524 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10048 1 3531 3530 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10049 3531 3530 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10050 1 3533 3532 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10051 3533 3532 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10052 1 3527 3526 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10053 3527 3526 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10054 1 3529 3528 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10055 3529 3528 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10056 1 3535 3534 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10057 3535 3534 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10058 1 3537 3536 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10059 3537 3536 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10060 0 3531 3530 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10061 3531 3530 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10062 0 3533 3532 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10063 3533 3532 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10064 0 3535 3534 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10065 3535 3534 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10066 0 3537 3536 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10067 3537 3536 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10068 326 548 3530 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10069 327 548 3531 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10070 328 548 3532 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10071 329 548 3533 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10072 330 548 3534 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10073 331 548 3535 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10074 332 548 3536 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10075 333 548 3537 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10076 3538 552 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10077 3539 552 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10078 3540 552 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10079 3541 552 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10080 3542 552 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10081 3543 552 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10082 3544 552 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10083 3545 552 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10084 0 3539 3538 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10085 3539 3538 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10086 0 3541 3540 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10087 3541 3540 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10088 0 3543 3542 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10089 3543 3542 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10090 0 3545 3544 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10091 3545 3544 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10092 1 3539 3538 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10093 3539 3538 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10094 1 3541 3540 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10095 3541 3540 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10096 1 3543 3542 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10097 3543 3542 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10098 1 3545 3544 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10099 3545 3544 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10100 1 3547 3546 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10101 3547 3546 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10102 1 3549 3548 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10103 3549 3548 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10104 1 3551 3550 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10105 3551 3550 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10106 1 3553 3552 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10107 3553 3552 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10108 0 3547 3546 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10109 3547 3546 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10110 0 3549 3548 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10111 3549 3548 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10112 0 3551 3550 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10113 3551 3550 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10114 0 3553 3552 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10115 3553 3552 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10116 326 556 3546 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10117 327 556 3547 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10118 328 556 3548 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10119 329 556 3549 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10120 330 556 3550 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10121 331 556 3551 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10122 332 556 3552 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10123 333 556 3553 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10124 3554 559 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10125 3555 559 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10126 3556 559 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10127 3557 559 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10128 3558 559 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10129 3559 559 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10130 3560 559 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10131 3561 559 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10132 0 3555 3554 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10133 3555 3554 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10134 0 3557 3556 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10135 3557 3556 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10136 0 3559 3558 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10137 3559 3558 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10138 0 3561 3560 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10139 3561 3560 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10140 1 3555 3554 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10141 3555 3554 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10142 1 3557 3556 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10143 3557 3556 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10144 1 3563 3562 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10145 3563 3562 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10146 1 3565 3564 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10147 3565 3564 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10148 1 3559 3558 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10149 3559 3558 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10150 1 3561 3560 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10151 3561 3560 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10152 1 3567 3566 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10153 3567 3566 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10154 1 3569 3568 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10155 3569 3568 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10156 0 3563 3562 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10157 3563 3562 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10158 0 3565 3564 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10159 3565 3564 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10160 0 3567 3566 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10161 3567 3566 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10162 0 3569 3568 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10163 3569 3568 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10164 326 564 3562 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10165 327 564 3563 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10166 328 564 3564 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10167 329 564 3565 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10168 330 564 3566 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10169 331 564 3567 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10170 332 564 3568 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10171 333 564 3569 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10172 3570 568 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10173 3571 568 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10174 3572 568 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10175 3573 568 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10176 3574 568 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10177 3575 568 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10178 3576 568 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10179 3577 568 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10180 0 3571 3570 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10181 3571 3570 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10182 0 3573 3572 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10183 3573 3572 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10184 0 3575 3574 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10185 3575 3574 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10186 0 3577 3576 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10187 3577 3576 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10188 1 3571 3570 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10189 3571 3570 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10190 1 3573 3572 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10191 3573 3572 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10192 1 3575 3574 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10193 3575 3574 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10194 1 3577 3576 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10195 3577 3576 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10196 1 3579 3578 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10197 3579 3578 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10198 1 3581 3580 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10199 3581 3580 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10200 1 3583 3582 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10201 3583 3582 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10202 1 3585 3584 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10203 3585 3584 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10204 0 3579 3578 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10205 3579 3578 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10206 0 3581 3580 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10207 3581 3580 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10208 0 3583 3582 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10209 3583 3582 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10210 0 3585 3584 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10211 3585 3584 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10212 326 572 3578 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10213 327 572 3579 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10214 328 572 3580 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10215 329 572 3581 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10216 330 572 3582 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10217 331 572 3583 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10218 332 572 3584 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10219 333 572 3585 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10220 3586 575 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10221 3587 575 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10222 3588 575 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10223 3589 575 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10224 3590 575 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10225 3591 575 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10226 3592 575 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10227 3593 575 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10228 0 3587 3586 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10229 3587 3586 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10230 0 3589 3588 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10231 3589 3588 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10232 0 3591 3590 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10233 3591 3590 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10234 0 3593 3592 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10235 3593 3592 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10236 1 3587 3586 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10237 3587 3586 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10238 1 3589 3588 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10239 3589 3588 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10240 1 3595 3594 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10241 3595 3594 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10242 1 3597 3596 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10243 3597 3596 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10244 1 3591 3590 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10245 3591 3590 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10246 1 3593 3592 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10247 3593 3592 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10248 1 3599 3598 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10249 3599 3598 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10250 1 3601 3600 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10251 3601 3600 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10252 0 3595 3594 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10253 3595 3594 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10254 0 3597 3596 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10255 3597 3596 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10256 0 3599 3598 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10257 3599 3598 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10258 0 3601 3600 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10259 3601 3600 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10260 326 580 3594 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10261 327 580 3595 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10262 328 580 3596 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10263 329 580 3597 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10264 330 580 3598 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10265 331 580 3599 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10266 332 580 3600 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10267 333 580 3601 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10268 3602 584 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10269 3603 584 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10270 3604 584 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10271 3605 584 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10272 3606 584 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10273 3607 584 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10274 3608 584 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10275 3609 584 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10276 0 3603 3602 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10277 3603 3602 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10278 0 3605 3604 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10279 3605 3604 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10280 0 3607 3606 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10281 3607 3606 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10282 0 3609 3608 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10283 3609 3608 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10284 1 3603 3602 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10285 3603 3602 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10286 1 3605 3604 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10287 3605 3604 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10288 1 3607 3606 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10289 3607 3606 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10290 1 3609 3608 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10291 3609 3608 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10292 1 3611 3610 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10293 3611 3610 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10294 1 3613 3612 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10295 3613 3612 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10296 1 3615 3614 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10297 3615 3614 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10298 1 3617 3616 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10299 3617 3616 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10300 0 3611 3610 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10301 3611 3610 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10302 0 3613 3612 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10303 3613 3612 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10304 0 3615 3614 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10305 3615 3614 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10306 0 3617 3616 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10307 3617 3616 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10308 326 588 3610 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10309 327 588 3611 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10310 328 588 3612 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10311 329 588 3613 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10312 330 588 3614 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10313 331 588 3615 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10314 332 588 3616 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10315 333 588 3617 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10316 3618 591 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10317 3619 591 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10318 3620 591 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10319 3621 591 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10320 3622 591 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10321 3623 591 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10322 3624 591 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10323 3625 591 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10324 0 3619 3618 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10325 3619 3618 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10326 0 3621 3620 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10327 3621 3620 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10328 0 3623 3622 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10329 3623 3622 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10330 0 3625 3624 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10331 3625 3624 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10332 1 3619 3618 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10333 3619 3618 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10334 1 3621 3620 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10335 3621 3620 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10336 1 3627 3626 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10337 3627 3626 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10338 1 3629 3628 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10339 3629 3628 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10340 1 3623 3622 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10341 3623 3622 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10342 1 3625 3624 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10343 3625 3624 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10344 1 3631 3630 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10345 3631 3630 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10346 1 3633 3632 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10347 3633 3632 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10348 0 3627 3626 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10349 3627 3626 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10350 0 3629 3628 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10351 3629 3628 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10352 0 3631 3630 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10353 3631 3630 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10354 0 3633 3632 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10355 3633 3632 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10356 326 596 3626 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10357 327 596 3627 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10358 328 596 3628 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10359 329 596 3629 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10360 330 596 3630 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10361 331 596 3631 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10362 332 596 3632 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10363 333 596 3633 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10364 3634 600 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10365 3635 600 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10366 3636 600 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10367 3637 600 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10368 3638 600 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10369 3639 600 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10370 3640 600 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10371 3641 600 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10372 0 3635 3634 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10373 3635 3634 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10374 0 3637 3636 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10375 3637 3636 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10376 0 3639 3638 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10377 3639 3638 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10378 0 3641 3640 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10379 3641 3640 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10380 1 3635 3634 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10381 3635 3634 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10382 1 3637 3636 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10383 3637 3636 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10384 1 3639 3638 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10385 3639 3638 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10386 1 3641 3640 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10387 3641 3640 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10388 1 3643 3642 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10389 3643 3642 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10390 1 3645 3644 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10391 3645 3644 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10392 1 3647 3646 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10393 3647 3646 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10394 1 3649 3648 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10395 3649 3648 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10396 0 3643 3642 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10397 3643 3642 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10398 0 3645 3644 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10399 3645 3644 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10400 0 3647 3646 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10401 3647 3646 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10402 0 3649 3648 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10403 3649 3648 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10404 326 604 3642 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10405 327 604 3643 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10406 328 604 3644 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10407 329 604 3645 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10408 330 604 3646 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10409 331 604 3647 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10410 332 604 3648 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10411 333 604 3649 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10412 3650 607 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10413 3651 607 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10414 3652 607 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10415 3653 607 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10416 3654 607 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10417 3655 607 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10418 3656 607 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10419 3657 607 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10420 0 3651 3650 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10421 3651 3650 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10422 0 3653 3652 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10423 3653 3652 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10424 0 3655 3654 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10425 3655 3654 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10426 0 3657 3656 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10427 3657 3656 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10428 1 3651 3650 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10429 3651 3650 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10430 1 3653 3652 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10431 3653 3652 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10432 1 3659 3658 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10433 3659 3658 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10434 1 3661 3660 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10435 3661 3660 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10436 1 3655 3654 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10437 3655 3654 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10438 1 3657 3656 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10439 3657 3656 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10440 1 3663 3662 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10441 3663 3662 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10442 1 3665 3664 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10443 3665 3664 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10444 0 3659 3658 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10445 3659 3658 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10446 0 3661 3660 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10447 3661 3660 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10448 0 3663 3662 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10449 3663 3662 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10450 0 3665 3664 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10451 3665 3664 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10452 326 612 3658 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10453 327 612 3659 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10454 328 612 3660 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10455 329 612 3661 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10456 330 612 3662 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10457 331 612 3663 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10458 332 612 3664 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10459 333 612 3665 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10460 3666 616 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10461 3667 616 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10462 3668 616 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10463 3669 616 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10464 3670 616 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10465 3671 616 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10466 3672 616 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10467 3673 616 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10468 0 3667 3666 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10469 3667 3666 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10470 0 3669 3668 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10471 3669 3668 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10472 0 3671 3670 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10473 3671 3670 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10474 0 3673 3672 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10475 3673 3672 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10476 1 3667 3666 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10477 3667 3666 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10478 1 3669 3668 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10479 3669 3668 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10480 1 3671 3670 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10481 3671 3670 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10482 1 3673 3672 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10483 3673 3672 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10484 1 3675 3674 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10485 3675 3674 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10486 1 3677 3676 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10487 3677 3676 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10488 1 3679 3678 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10489 3679 3678 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10490 1 3681 3680 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10491 3681 3680 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10492 0 3675 3674 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10493 3675 3674 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10494 0 3677 3676 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10495 3677 3676 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10496 0 3679 3678 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10497 3679 3678 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10498 0 3681 3680 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10499 3681 3680 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10500 326 620 3674 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10501 327 620 3675 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10502 328 620 3676 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10503 329 620 3677 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10504 330 620 3678 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10505 331 620 3679 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10506 332 620 3680 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10507 333 620 3681 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10508 3682 624 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10509 3683 624 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10510 3684 624 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10511 3685 624 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10512 3686 624 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10513 3687 624 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10514 3688 624 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10515 3689 624 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10516 0 3683 3682 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10517 3683 3682 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10518 0 3685 3684 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10519 3685 3684 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10520 0 3687 3686 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10521 3687 3686 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10522 0 3689 3688 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10523 3689 3688 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10524 1 3683 3682 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10525 3683 3682 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10526 1 3685 3684 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10527 3685 3684 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10528 1 3691 3690 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10529 3691 3690 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10530 1 3693 3692 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10531 3693 3692 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10532 1 3687 3686 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10533 3687 3686 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10534 1 3689 3688 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10535 3689 3688 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10536 1 3695 3694 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10537 3695 3694 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10538 1 3697 3696 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10539 3697 3696 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10540 0 3691 3690 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10541 3691 3690 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10542 0 3693 3692 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10543 3693 3692 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10544 0 3695 3694 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10545 3695 3694 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10546 0 3697 3696 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10547 3697 3696 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10548 326 628 3690 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10549 327 628 3691 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10550 328 628 3692 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10551 329 628 3693 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10552 330 628 3694 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10553 331 628 3695 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10554 332 628 3696 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10555 333 628 3697 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10556 3698 632 326 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10557 3699 632 327 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10558 3700 632 328 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10559 3701 632 329 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10560 3702 632 330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10561 3703 632 331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10562 3704 632 332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10563 3705 632 333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10564 0 3699 3698 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10565 3699 3698 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10566 0 3701 3700 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10567 3701 3700 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10568 0 3703 3702 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10569 3703 3702 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10570 0 3705 3704 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10571 3705 3704 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10572 1 3699 3698 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10573 3699 3698 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10574 1 3701 3700 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10575 3701 3700 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10576 1 3703 3702 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10577 3703 3702 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10578 1 3705 3704 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10579 3705 3704 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10580 1 3707 3706 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10581 3707 3706 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10582 1 3709 3708 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10583 3709 3708 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10584 1 3711 3710 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10585 3711 3710 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10586 1 3713 3712 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10587 3713 3712 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10588 0 3707 3706 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10589 3707 3706 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10590 0 3709 3708 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10591 3709 3708 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10592 0 3711 3710 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10593 3711 3710 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10594 0 3713 3712 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10595 3713 3712 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10596 352 380 3706 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10597 353 380 3707 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10598 354 380 3708 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10599 355 380 3709 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10600 356 380 3710 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10601 357 380 3711 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10602 358 380 3712 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10603 359 380 3713 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10604 3714 383 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10605 3715 383 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10606 3716 383 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10607 3717 383 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10608 3718 383 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10609 3719 383 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10610 3720 383 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10611 3721 383 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10612 0 3715 3714 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10613 3715 3714 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10614 0 3717 3716 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10615 3717 3716 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10616 0 3719 3718 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10617 3719 3718 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10618 0 3721 3720 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10619 3721 3720 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10620 1 3715 3714 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10621 3715 3714 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10622 1 3717 3716 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10623 3717 3716 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10624 1 3723 3722 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10625 3723 3722 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10626 1 3725 3724 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10627 3725 3724 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10628 1 3719 3718 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10629 3719 3718 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10630 1 3721 3720 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10631 3721 3720 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10632 1 3727 3726 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10633 3727 3726 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10634 1 3729 3728 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10635 3729 3728 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10636 0 3723 3722 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10637 3723 3722 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10638 0 3725 3724 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10639 3725 3724 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10640 0 3727 3726 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10641 3727 3726 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10642 0 3729 3728 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10643 3729 3728 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10644 352 388 3722 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10645 353 388 3723 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10646 354 388 3724 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10647 355 388 3725 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10648 356 388 3726 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10649 357 388 3727 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10650 358 388 3728 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10651 359 388 3729 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10652 3730 392 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10653 3731 392 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10654 3732 392 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10655 3733 392 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10656 3734 392 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10657 3735 392 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10658 3736 392 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10659 3737 392 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10660 0 3731 3730 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10661 3731 3730 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10662 0 3733 3732 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10663 3733 3732 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10664 0 3735 3734 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10665 3735 3734 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10666 0 3737 3736 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10667 3737 3736 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10668 1 3731 3730 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10669 3731 3730 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10670 1 3733 3732 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10671 3733 3732 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10672 1 3735 3734 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10673 3735 3734 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10674 1 3737 3736 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10675 3737 3736 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10676 1 3739 3738 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10677 3739 3738 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10678 1 3741 3740 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10679 3741 3740 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10680 1 3743 3742 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10681 3743 3742 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10682 1 3745 3744 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10683 3745 3744 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10684 0 3739 3738 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10685 3739 3738 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10686 0 3741 3740 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10687 3741 3740 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10688 0 3743 3742 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10689 3743 3742 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10690 0 3745 3744 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10691 3745 3744 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10692 352 396 3738 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10693 353 396 3739 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10694 354 396 3740 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10695 355 396 3741 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10696 356 396 3742 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10697 357 396 3743 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10698 358 396 3744 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10699 359 396 3745 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10700 3746 399 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10701 3747 399 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10702 3748 399 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10703 3749 399 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10704 3750 399 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10705 3751 399 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10706 3752 399 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10707 3753 399 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10708 0 3747 3746 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10709 3747 3746 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10710 0 3749 3748 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10711 3749 3748 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10712 0 3751 3750 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10713 3751 3750 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10714 0 3753 3752 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10715 3753 3752 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10716 1 3747 3746 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10717 3747 3746 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10718 1 3749 3748 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10719 3749 3748 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10720 1 3755 3754 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10721 3755 3754 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10722 1 3757 3756 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10723 3757 3756 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10724 1 3751 3750 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10725 3751 3750 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10726 1 3753 3752 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10727 3753 3752 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10728 1 3759 3758 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10729 3759 3758 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10730 1 3761 3760 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10731 3761 3760 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10732 0 3755 3754 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10733 3755 3754 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10734 0 3757 3756 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10735 3757 3756 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10736 0 3759 3758 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10737 3759 3758 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10738 0 3761 3760 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10739 3761 3760 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10740 352 404 3754 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10741 353 404 3755 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10742 354 404 3756 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10743 355 404 3757 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10744 356 404 3758 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10745 357 404 3759 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10746 358 404 3760 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10747 359 404 3761 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10748 3762 408 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10749 3763 408 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10750 3764 408 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10751 3765 408 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10752 3766 408 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10753 3767 408 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10754 3768 408 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10755 3769 408 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10756 0 3763 3762 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10757 3763 3762 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10758 0 3765 3764 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10759 3765 3764 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10760 0 3767 3766 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10761 3767 3766 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10762 0 3769 3768 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10763 3769 3768 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10764 1 3763 3762 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10765 3763 3762 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10766 1 3765 3764 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10767 3765 3764 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10768 1 3767 3766 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10769 3767 3766 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10770 1 3769 3768 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10771 3769 3768 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10772 1 3771 3770 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10773 3771 3770 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10774 1 3773 3772 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10775 3773 3772 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10776 1 3775 3774 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10777 3775 3774 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10778 1 3777 3776 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10779 3777 3776 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10780 0 3771 3770 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10781 3771 3770 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10782 0 3773 3772 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10783 3773 3772 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10784 0 3775 3774 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10785 3775 3774 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10786 0 3777 3776 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10787 3777 3776 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10788 352 412 3770 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10789 353 412 3771 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10790 354 412 3772 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10791 355 412 3773 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10792 356 412 3774 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10793 357 412 3775 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10794 358 412 3776 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10795 359 412 3777 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10796 3778 415 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10797 3779 415 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10798 3780 415 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10799 3781 415 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10800 3782 415 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10801 3783 415 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10802 3784 415 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10803 3785 415 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10804 0 3779 3778 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10805 3779 3778 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10806 0 3781 3780 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10807 3781 3780 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10808 0 3783 3782 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10809 3783 3782 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10810 0 3785 3784 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10811 3785 3784 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10812 1 3779 3778 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10813 3779 3778 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10814 1 3781 3780 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10815 3781 3780 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10816 1 3787 3786 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10817 3787 3786 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10818 1 3789 3788 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10819 3789 3788 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10820 1 3783 3782 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10821 3783 3782 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10822 1 3785 3784 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10823 3785 3784 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10824 1 3791 3790 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10825 3791 3790 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10826 1 3793 3792 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10827 3793 3792 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10828 0 3787 3786 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10829 3787 3786 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10830 0 3789 3788 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10831 3789 3788 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10832 0 3791 3790 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10833 3791 3790 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10834 0 3793 3792 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10835 3793 3792 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10836 352 420 3786 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10837 353 420 3787 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10838 354 420 3788 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10839 355 420 3789 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10840 356 420 3790 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10841 357 420 3791 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10842 358 420 3792 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10843 359 420 3793 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10844 3794 424 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10845 3795 424 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10846 3796 424 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10847 3797 424 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10848 3798 424 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10849 3799 424 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10850 3800 424 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10851 3801 424 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10852 0 3795 3794 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10853 3795 3794 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10854 0 3797 3796 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10855 3797 3796 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10856 0 3799 3798 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10857 3799 3798 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10858 0 3801 3800 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10859 3801 3800 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10860 1 3795 3794 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10861 3795 3794 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10862 1 3797 3796 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10863 3797 3796 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10864 1 3799 3798 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10865 3799 3798 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10866 1 3801 3800 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10867 3801 3800 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10868 1 3803 3802 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10869 3803 3802 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10870 1 3805 3804 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10871 3805 3804 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10872 1 3807 3806 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10873 3807 3806 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10874 1 3809 3808 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10875 3809 3808 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10876 0 3803 3802 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10877 3803 3802 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10878 0 3805 3804 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10879 3805 3804 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10880 0 3807 3806 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10881 3807 3806 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10882 0 3809 3808 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10883 3809 3808 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10884 352 428 3802 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10885 353 428 3803 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10886 354 428 3804 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10887 355 428 3805 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10888 356 428 3806 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10889 357 428 3807 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10890 358 428 3808 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10891 359 428 3809 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10892 3810 431 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10893 3811 431 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10894 3812 431 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10895 3813 431 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10896 3814 431 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10897 3815 431 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10898 3816 431 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10899 3817 431 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10900 0 3811 3810 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10901 3811 3810 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10902 0 3813 3812 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10903 3813 3812 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10904 0 3815 3814 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10905 3815 3814 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10906 0 3817 3816 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10907 3817 3816 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10908 1 3811 3810 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10909 3811 3810 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10910 1 3813 3812 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10911 3813 3812 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10912 1 3819 3818 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10913 3819 3818 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10914 1 3821 3820 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10915 3821 3820 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10916 1 3815 3814 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10917 3815 3814 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10918 1 3817 3816 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10919 3817 3816 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10920 1 3823 3822 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10921 3823 3822 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10922 1 3825 3824 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10923 3825 3824 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10924 0 3819 3818 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10925 3819 3818 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10926 0 3821 3820 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10927 3821 3820 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10928 0 3823 3822 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10929 3823 3822 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10930 0 3825 3824 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10931 3825 3824 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10932 352 436 3818 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10933 353 436 3819 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10934 354 436 3820 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10935 355 436 3821 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10936 356 436 3822 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10937 357 436 3823 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10938 358 436 3824 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10939 359 436 3825 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10940 3826 440 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10941 3827 440 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10942 3828 440 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10943 3829 440 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10944 3830 440 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10945 3831 440 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10946 3832 440 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10947 3833 440 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10948 0 3827 3826 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10949 3827 3826 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10950 0 3829 3828 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10951 3829 3828 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10952 0 3831 3830 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10953 3831 3830 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10954 0 3833 3832 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10955 3833 3832 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10956 1 3827 3826 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10957 3827 3826 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10958 1 3829 3828 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10959 3829 3828 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10960 1 3831 3830 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10961 3831 3830 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10962 1 3833 3832 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10963 3833 3832 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10964 1 3835 3834 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10965 3835 3834 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m10966 1 3837 3836 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10967 3837 3836 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10968 1 3839 3838 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m10969 3839 3838 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10970 1 3841 3840 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m10971 3841 3840 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m10972 0 3835 3834 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10973 3835 3834 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10974 0 3837 3836 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10975 3837 3836 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10976 0 3839 3838 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10977 3839 3838 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10978 0 3841 3840 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m10979 3841 3840 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m10980 352 444 3834 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m10981 353 444 3835 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10982 354 444 3836 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10983 355 444 3837 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10984 356 444 3838 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m10985 357 444 3839 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m10986 358 444 3840 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m10987 359 444 3841 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m10988 3842 447 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m10989 3843 447 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10990 3844 447 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10991 3845 447 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10992 3846 447 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m10993 3847 447 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m10994 3848 447 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m10995 3849 447 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m10996 0 3843 3842 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10997 3843 3842 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m10998 0 3845 3844 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m10999 3845 3844 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11000 0 3847 3846 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11001 3847 3846 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11002 0 3849 3848 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11003 3849 3848 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11004 1 3843 3842 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11005 3843 3842 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11006 1 3845 3844 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11007 3845 3844 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11008 1 3851 3850 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11009 3851 3850 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11010 1 3853 3852 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11011 3853 3852 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11012 1 3847 3846 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11013 3847 3846 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11014 1 3849 3848 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11015 3849 3848 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11016 1 3855 3854 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11017 3855 3854 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11018 1 3857 3856 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11019 3857 3856 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11020 0 3851 3850 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11021 3851 3850 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11022 0 3853 3852 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11023 3853 3852 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11024 0 3855 3854 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11025 3855 3854 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11026 0 3857 3856 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11027 3857 3856 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11028 352 452 3850 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11029 353 452 3851 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11030 354 452 3852 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11031 355 452 3853 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11032 356 452 3854 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11033 357 452 3855 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11034 358 452 3856 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11035 359 452 3857 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11036 3858 456 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11037 3859 456 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11038 3860 456 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11039 3861 456 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11040 3862 456 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11041 3863 456 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11042 3864 456 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11043 3865 456 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11044 0 3859 3858 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11045 3859 3858 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11046 0 3861 3860 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11047 3861 3860 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11048 0 3863 3862 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11049 3863 3862 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11050 0 3865 3864 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11051 3865 3864 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11052 1 3859 3858 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11053 3859 3858 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11054 1 3861 3860 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11055 3861 3860 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11056 1 3863 3862 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11057 3863 3862 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11058 1 3865 3864 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11059 3865 3864 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11060 1 3867 3866 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11061 3867 3866 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11062 1 3869 3868 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11063 3869 3868 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11064 1 3871 3870 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11065 3871 3870 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11066 1 3873 3872 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11067 3873 3872 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11068 0 3867 3866 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11069 3867 3866 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11070 0 3869 3868 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11071 3869 3868 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11072 0 3871 3870 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11073 3871 3870 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11074 0 3873 3872 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11075 3873 3872 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11076 352 460 3866 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11077 353 460 3867 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11078 354 460 3868 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11079 355 460 3869 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11080 356 460 3870 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11081 357 460 3871 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11082 358 460 3872 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11083 359 460 3873 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11084 3874 463 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11085 3875 463 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11086 3876 463 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11087 3877 463 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11088 3878 463 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11089 3879 463 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11090 3880 463 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11091 3881 463 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11092 0 3875 3874 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11093 3875 3874 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11094 0 3877 3876 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11095 3877 3876 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11096 0 3879 3878 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11097 3879 3878 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11098 0 3881 3880 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11099 3881 3880 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11100 1 3875 3874 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11101 3875 3874 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11102 1 3877 3876 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11103 3877 3876 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11104 1 3883 3882 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11105 3883 3882 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11106 1 3885 3884 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11107 3885 3884 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11108 1 3879 3878 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11109 3879 3878 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11110 1 3881 3880 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11111 3881 3880 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11112 1 3887 3886 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11113 3887 3886 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11114 1 3889 3888 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11115 3889 3888 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11116 0 3883 3882 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11117 3883 3882 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11118 0 3885 3884 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11119 3885 3884 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11120 0 3887 3886 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11121 3887 3886 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11122 0 3889 3888 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11123 3889 3888 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11124 352 468 3882 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11125 353 468 3883 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11126 354 468 3884 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11127 355 468 3885 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11128 356 468 3886 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11129 357 468 3887 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11130 358 468 3888 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11131 359 468 3889 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11132 3890 472 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11133 3891 472 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11134 3892 472 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11135 3893 472 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11136 3894 472 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11137 3895 472 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11138 3896 472 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11139 3897 472 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11140 0 3891 3890 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11141 3891 3890 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11142 0 3893 3892 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11143 3893 3892 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11144 0 3895 3894 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11145 3895 3894 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11146 0 3897 3896 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11147 3897 3896 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11148 1 3891 3890 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11149 3891 3890 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11150 1 3893 3892 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11151 3893 3892 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11152 1 3895 3894 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11153 3895 3894 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11154 1 3897 3896 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11155 3897 3896 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11156 1 3899 3898 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11157 3899 3898 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11158 1 3901 3900 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11159 3901 3900 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11160 1 3903 3902 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11161 3903 3902 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11162 1 3905 3904 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11163 3905 3904 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11164 0 3899 3898 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11165 3899 3898 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11166 0 3901 3900 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11167 3901 3900 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11168 0 3903 3902 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11169 3903 3902 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11170 0 3905 3904 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11171 3905 3904 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11172 352 476 3898 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11173 353 476 3899 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11174 354 476 3900 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11175 355 476 3901 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11176 356 476 3902 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11177 357 476 3903 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11178 358 476 3904 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11179 359 476 3905 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11180 3906 479 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11181 3907 479 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11182 3908 479 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11183 3909 479 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11184 3910 479 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11185 3911 479 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11186 3912 479 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11187 3913 479 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11188 0 3907 3906 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11189 3907 3906 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11190 0 3909 3908 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11191 3909 3908 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11192 0 3911 3910 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11193 3911 3910 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11194 0 3913 3912 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11195 3913 3912 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11196 1 3907 3906 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11197 3907 3906 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11198 1 3909 3908 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11199 3909 3908 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11200 1 3915 3914 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11201 3915 3914 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11202 1 3917 3916 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11203 3917 3916 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11204 1 3911 3910 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11205 3911 3910 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11206 1 3913 3912 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11207 3913 3912 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11208 1 3919 3918 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11209 3919 3918 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11210 1 3921 3920 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11211 3921 3920 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11212 0 3915 3914 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11213 3915 3914 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11214 0 3917 3916 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11215 3917 3916 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11216 0 3919 3918 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11217 3919 3918 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11218 0 3921 3920 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11219 3921 3920 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11220 352 484 3914 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11221 353 484 3915 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11222 354 484 3916 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11223 355 484 3917 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11224 356 484 3918 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11225 357 484 3919 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11226 358 484 3920 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11227 359 484 3921 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11228 3922 488 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11229 3923 488 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11230 3924 488 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11231 3925 488 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11232 3926 488 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11233 3927 488 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11234 3928 488 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11235 3929 488 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11236 0 3923 3922 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11237 3923 3922 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11238 0 3925 3924 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11239 3925 3924 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11240 0 3927 3926 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11241 3927 3926 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11242 0 3929 3928 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11243 3929 3928 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11244 1 3923 3922 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11245 3923 3922 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11246 1 3925 3924 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11247 3925 3924 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11248 1 3927 3926 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11249 3927 3926 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11250 1 3929 3928 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11251 3929 3928 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11252 1 3931 3930 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11253 3931 3930 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11254 1 3933 3932 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11255 3933 3932 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11256 1 3935 3934 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11257 3935 3934 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11258 1 3937 3936 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11259 3937 3936 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11260 0 3931 3930 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11261 3931 3930 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11262 0 3933 3932 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11263 3933 3932 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11264 0 3935 3934 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11265 3935 3934 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11266 0 3937 3936 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11267 3937 3936 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11268 352 492 3930 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11269 353 492 3931 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11270 354 492 3932 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11271 355 492 3933 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11272 356 492 3934 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11273 357 492 3935 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11274 358 492 3936 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11275 359 492 3937 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11276 3938 495 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11277 3939 495 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11278 3940 495 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11279 3941 495 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11280 3942 495 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11281 3943 495 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11282 3944 495 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11283 3945 495 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11284 0 3939 3938 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11285 3939 3938 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11286 0 3941 3940 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11287 3941 3940 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11288 0 3943 3942 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11289 3943 3942 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11290 0 3945 3944 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11291 3945 3944 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11292 1 3939 3938 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11293 3939 3938 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11294 1 3941 3940 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11295 3941 3940 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11296 1 3947 3946 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11297 3947 3946 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11298 1 3949 3948 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11299 3949 3948 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11300 1 3943 3942 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11301 3943 3942 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11302 1 3945 3944 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11303 3945 3944 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11304 1 3951 3950 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11305 3951 3950 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11306 1 3953 3952 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11307 3953 3952 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11308 0 3947 3946 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11309 3947 3946 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11310 0 3949 3948 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11311 3949 3948 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11312 0 3951 3950 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11313 3951 3950 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11314 0 3953 3952 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11315 3953 3952 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11316 352 500 3946 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11317 353 500 3947 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11318 354 500 3948 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11319 355 500 3949 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11320 356 500 3950 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11321 357 500 3951 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11322 358 500 3952 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11323 359 500 3953 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11324 3954 504 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11325 3955 504 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11326 3956 504 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11327 3957 504 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11328 3958 504 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11329 3959 504 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11330 3960 504 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11331 3961 504 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11332 0 3955 3954 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11333 3955 3954 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11334 0 3957 3956 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11335 3957 3956 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11336 0 3959 3958 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11337 3959 3958 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11338 0 3961 3960 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11339 3961 3960 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11340 1 3955 3954 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11341 3955 3954 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11342 1 3957 3956 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11343 3957 3956 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11344 1 3959 3958 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11345 3959 3958 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11346 1 3961 3960 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11347 3961 3960 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11348 1 3963 3962 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11349 3963 3962 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11350 1 3965 3964 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11351 3965 3964 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11352 1 3967 3966 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11353 3967 3966 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11354 1 3969 3968 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11355 3969 3968 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11356 0 3963 3962 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11357 3963 3962 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11358 0 3965 3964 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11359 3965 3964 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11360 0 3967 3966 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11361 3967 3966 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11362 0 3969 3968 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11363 3969 3968 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11364 352 508 3962 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11365 353 508 3963 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11366 354 508 3964 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11367 355 508 3965 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11368 356 508 3966 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11369 357 508 3967 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11370 358 508 3968 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11371 359 508 3969 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11372 3970 511 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11373 3971 511 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11374 3972 511 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11375 3973 511 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11376 3974 511 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11377 3975 511 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11378 3976 511 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11379 3977 511 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11380 0 3971 3970 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11381 3971 3970 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11382 0 3973 3972 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11383 3973 3972 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11384 0 3975 3974 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11385 3975 3974 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11386 0 3977 3976 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11387 3977 3976 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11388 1 3971 3970 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11389 3971 3970 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11390 1 3973 3972 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11391 3973 3972 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11392 1 3979 3978 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11393 3979 3978 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11394 1 3981 3980 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11395 3981 3980 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11396 1 3975 3974 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11397 3975 3974 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11398 1 3977 3976 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11399 3977 3976 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11400 1 3983 3982 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11401 3983 3982 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11402 1 3985 3984 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11403 3985 3984 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11404 0 3979 3978 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11405 3979 3978 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11406 0 3981 3980 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11407 3981 3980 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11408 0 3983 3982 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11409 3983 3982 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11410 0 3985 3984 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11411 3985 3984 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11412 352 516 3978 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11413 353 516 3979 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11414 354 516 3980 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11415 355 516 3981 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11416 356 516 3982 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11417 357 516 3983 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11418 358 516 3984 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11419 359 516 3985 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11420 3986 520 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11421 3987 520 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11422 3988 520 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11423 3989 520 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11424 3990 520 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11425 3991 520 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11426 3992 520 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11427 3993 520 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11428 0 3987 3986 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11429 3987 3986 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11430 0 3989 3988 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11431 3989 3988 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11432 0 3991 3990 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11433 3991 3990 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11434 0 3993 3992 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11435 3993 3992 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11436 1 3987 3986 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11437 3987 3986 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11438 1 3989 3988 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11439 3989 3988 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11440 1 3991 3990 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11441 3991 3990 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11442 1 3993 3992 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11443 3993 3992 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11444 1 3995 3994 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11445 3995 3994 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11446 1 3997 3996 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11447 3997 3996 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11448 1 3999 3998 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11449 3999 3998 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11450 1 4001 4000 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11451 4001 4000 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11452 0 3995 3994 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11453 3995 3994 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11454 0 3997 3996 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11455 3997 3996 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11456 0 3999 3998 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11457 3999 3998 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11458 0 4001 4000 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11459 4001 4000 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11460 352 524 3994 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11461 353 524 3995 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11462 354 524 3996 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11463 355 524 3997 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11464 356 524 3998 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11465 357 524 3999 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11466 358 524 4000 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11467 359 524 4001 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11468 4002 527 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11469 4003 527 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11470 4004 527 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11471 4005 527 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11472 4006 527 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11473 4007 527 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11474 4008 527 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11475 4009 527 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11476 0 4003 4002 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11477 4003 4002 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11478 0 4005 4004 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11479 4005 4004 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11480 0 4007 4006 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11481 4007 4006 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11482 0 4009 4008 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11483 4009 4008 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11484 1 4003 4002 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11485 4003 4002 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11486 1 4005 4004 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11487 4005 4004 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11488 1 4011 4010 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11489 4011 4010 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11490 1 4013 4012 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11491 4013 4012 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11492 1 4007 4006 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11493 4007 4006 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11494 1 4009 4008 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11495 4009 4008 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11496 1 4015 4014 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11497 4015 4014 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11498 1 4017 4016 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11499 4017 4016 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11500 0 4011 4010 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11501 4011 4010 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11502 0 4013 4012 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11503 4013 4012 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11504 0 4015 4014 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11505 4015 4014 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11506 0 4017 4016 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11507 4017 4016 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11508 352 532 4010 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11509 353 532 4011 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11510 354 532 4012 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11511 355 532 4013 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11512 356 532 4014 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11513 357 532 4015 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11514 358 532 4016 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11515 359 532 4017 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11516 4018 536 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11517 4019 536 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11518 4020 536 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11519 4021 536 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11520 4022 536 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11521 4023 536 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11522 4024 536 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11523 4025 536 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11524 0 4019 4018 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11525 4019 4018 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11526 0 4021 4020 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11527 4021 4020 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11528 0 4023 4022 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11529 4023 4022 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11530 0 4025 4024 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11531 4025 4024 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11532 1 4019 4018 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11533 4019 4018 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11534 1 4021 4020 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11535 4021 4020 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11536 1 4023 4022 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11537 4023 4022 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11538 1 4025 4024 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11539 4025 4024 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11540 1 4027 4026 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11541 4027 4026 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11542 1 4029 4028 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11543 4029 4028 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11544 1 4031 4030 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11545 4031 4030 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11546 1 4033 4032 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11547 4033 4032 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11548 0 4027 4026 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11549 4027 4026 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11550 0 4029 4028 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11551 4029 4028 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11552 0 4031 4030 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11553 4031 4030 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11554 0 4033 4032 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11555 4033 4032 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11556 352 540 4026 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11557 353 540 4027 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11558 354 540 4028 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11559 355 540 4029 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11560 356 540 4030 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11561 357 540 4031 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11562 358 540 4032 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11563 359 540 4033 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11564 4034 543 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11565 4035 543 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11566 4036 543 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11567 4037 543 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11568 4038 543 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11569 4039 543 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11570 4040 543 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11571 4041 543 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11572 0 4035 4034 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11573 4035 4034 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11574 0 4037 4036 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11575 4037 4036 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11576 0 4039 4038 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11577 4039 4038 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11578 0 4041 4040 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11579 4041 4040 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11580 1 4035 4034 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11581 4035 4034 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11582 1 4037 4036 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11583 4037 4036 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11584 1 4043 4042 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11585 4043 4042 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11586 1 4045 4044 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11587 4045 4044 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11588 1 4039 4038 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11589 4039 4038 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11590 1 4041 4040 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11591 4041 4040 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11592 1 4047 4046 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11593 4047 4046 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11594 1 4049 4048 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11595 4049 4048 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11596 0 4043 4042 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11597 4043 4042 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11598 0 4045 4044 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11599 4045 4044 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11600 0 4047 4046 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11601 4047 4046 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11602 0 4049 4048 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11603 4049 4048 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11604 352 548 4042 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11605 353 548 4043 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11606 354 548 4044 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11607 355 548 4045 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11608 356 548 4046 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11609 357 548 4047 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11610 358 548 4048 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11611 359 548 4049 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11612 4050 552 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11613 4051 552 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11614 4052 552 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11615 4053 552 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11616 4054 552 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11617 4055 552 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11618 4056 552 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11619 4057 552 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11620 0 4051 4050 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11621 4051 4050 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11622 0 4053 4052 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11623 4053 4052 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11624 0 4055 4054 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11625 4055 4054 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11626 0 4057 4056 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11627 4057 4056 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11628 1 4051 4050 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11629 4051 4050 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11630 1 4053 4052 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11631 4053 4052 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11632 1 4055 4054 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11633 4055 4054 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11634 1 4057 4056 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11635 4057 4056 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11636 1 4059 4058 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11637 4059 4058 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11638 1 4061 4060 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11639 4061 4060 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11640 1 4063 4062 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11641 4063 4062 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11642 1 4065 4064 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11643 4065 4064 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11644 0 4059 4058 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11645 4059 4058 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11646 0 4061 4060 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11647 4061 4060 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11648 0 4063 4062 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11649 4063 4062 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11650 0 4065 4064 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11651 4065 4064 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11652 352 556 4058 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11653 353 556 4059 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11654 354 556 4060 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11655 355 556 4061 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11656 356 556 4062 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11657 357 556 4063 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11658 358 556 4064 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11659 359 556 4065 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11660 4066 559 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11661 4067 559 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11662 4068 559 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11663 4069 559 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11664 4070 559 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11665 4071 559 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11666 4072 559 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11667 4073 559 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11668 0 4067 4066 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11669 4067 4066 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11670 0 4069 4068 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11671 4069 4068 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11672 0 4071 4070 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11673 4071 4070 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11674 0 4073 4072 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11675 4073 4072 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11676 1 4067 4066 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11677 4067 4066 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11678 1 4069 4068 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11679 4069 4068 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11680 1 4075 4074 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11681 4075 4074 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11682 1 4077 4076 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11683 4077 4076 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11684 1 4071 4070 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11685 4071 4070 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11686 1 4073 4072 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11687 4073 4072 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11688 1 4079 4078 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11689 4079 4078 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11690 1 4081 4080 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11691 4081 4080 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11692 0 4075 4074 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11693 4075 4074 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11694 0 4077 4076 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11695 4077 4076 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11696 0 4079 4078 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11697 4079 4078 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11698 0 4081 4080 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11699 4081 4080 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11700 352 564 4074 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11701 353 564 4075 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11702 354 564 4076 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11703 355 564 4077 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11704 356 564 4078 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11705 357 564 4079 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11706 358 564 4080 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11707 359 564 4081 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11708 4082 568 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11709 4083 568 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11710 4084 568 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11711 4085 568 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11712 4086 568 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11713 4087 568 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11714 4088 568 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11715 4089 568 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11716 0 4083 4082 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11717 4083 4082 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11718 0 4085 4084 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11719 4085 4084 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11720 0 4087 4086 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11721 4087 4086 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11722 0 4089 4088 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11723 4089 4088 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11724 1 4083 4082 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11725 4083 4082 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11726 1 4085 4084 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11727 4085 4084 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11728 1 4087 4086 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11729 4087 4086 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11730 1 4089 4088 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11731 4089 4088 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11732 1 4091 4090 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11733 4091 4090 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11734 1 4093 4092 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11735 4093 4092 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11736 1 4095 4094 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11737 4095 4094 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11738 1 4097 4096 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11739 4097 4096 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11740 0 4091 4090 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11741 4091 4090 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11742 0 4093 4092 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11743 4093 4092 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11744 0 4095 4094 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11745 4095 4094 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11746 0 4097 4096 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11747 4097 4096 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11748 352 572 4090 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11749 353 572 4091 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11750 354 572 4092 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11751 355 572 4093 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11752 356 572 4094 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11753 357 572 4095 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11754 358 572 4096 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11755 359 572 4097 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11756 4098 575 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11757 4099 575 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11758 4100 575 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11759 4101 575 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11760 4102 575 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11761 4103 575 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11762 4104 575 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11763 4105 575 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11764 0 4099 4098 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11765 4099 4098 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11766 0 4101 4100 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11767 4101 4100 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11768 0 4103 4102 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11769 4103 4102 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11770 0 4105 4104 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11771 4105 4104 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11772 1 4099 4098 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11773 4099 4098 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11774 1 4101 4100 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11775 4101 4100 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11776 1 4107 4106 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11777 4107 4106 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11778 1 4109 4108 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11779 4109 4108 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11780 1 4103 4102 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11781 4103 4102 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11782 1 4105 4104 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11783 4105 4104 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11784 1 4111 4110 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11785 4111 4110 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11786 1 4113 4112 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11787 4113 4112 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11788 0 4107 4106 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11789 4107 4106 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11790 0 4109 4108 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11791 4109 4108 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11792 0 4111 4110 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11793 4111 4110 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11794 0 4113 4112 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11795 4113 4112 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11796 352 580 4106 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11797 353 580 4107 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11798 354 580 4108 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11799 355 580 4109 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11800 356 580 4110 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11801 357 580 4111 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11802 358 580 4112 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11803 359 580 4113 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11804 4114 584 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11805 4115 584 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11806 4116 584 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11807 4117 584 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11808 4118 584 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11809 4119 584 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11810 4120 584 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11811 4121 584 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11812 0 4115 4114 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11813 4115 4114 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11814 0 4117 4116 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11815 4117 4116 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11816 0 4119 4118 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11817 4119 4118 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11818 0 4121 4120 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11819 4121 4120 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11820 1 4115 4114 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11821 4115 4114 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11822 1 4117 4116 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11823 4117 4116 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11824 1 4119 4118 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11825 4119 4118 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11826 1 4121 4120 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11827 4121 4120 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11828 1 4123 4122 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11829 4123 4122 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11830 1 4125 4124 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11831 4125 4124 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11832 1 4127 4126 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11833 4127 4126 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11834 1 4129 4128 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11835 4129 4128 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11836 0 4123 4122 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11837 4123 4122 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11838 0 4125 4124 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11839 4125 4124 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11840 0 4127 4126 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11841 4127 4126 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11842 0 4129 4128 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11843 4129 4128 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11844 352 588 4122 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11845 353 588 4123 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11846 354 588 4124 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11847 355 588 4125 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11848 356 588 4126 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11849 357 588 4127 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11850 358 588 4128 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11851 359 588 4129 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11852 4130 591 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11853 4131 591 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11854 4132 591 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11855 4133 591 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11856 4134 591 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11857 4135 591 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11858 4136 591 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11859 4137 591 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11860 0 4131 4130 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11861 4131 4130 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11862 0 4133 4132 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11863 4133 4132 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11864 0 4135 4134 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11865 4135 4134 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11866 0 4137 4136 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11867 4137 4136 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11868 1 4131 4130 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11869 4131 4130 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11870 1 4133 4132 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11871 4133 4132 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11872 1 4139 4138 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11873 4139 4138 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11874 1 4141 4140 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11875 4141 4140 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11876 1 4135 4134 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11877 4135 4134 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11878 1 4137 4136 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11879 4137 4136 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11880 1 4143 4142 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11881 4143 4142 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11882 1 4145 4144 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11883 4145 4144 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11884 0 4139 4138 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11885 4139 4138 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11886 0 4141 4140 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11887 4141 4140 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11888 0 4143 4142 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11889 4143 4142 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11890 0 4145 4144 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11891 4145 4144 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11892 352 596 4138 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11893 353 596 4139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11894 354 596 4140 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11895 355 596 4141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11896 356 596 4142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11897 357 596 4143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11898 358 596 4144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11899 359 596 4145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11900 4146 600 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11901 4147 600 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11902 4148 600 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11903 4149 600 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11904 4150 600 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11905 4151 600 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11906 4152 600 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11907 4153 600 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11908 0 4147 4146 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11909 4147 4146 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11910 0 4149 4148 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11911 4149 4148 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11912 0 4151 4150 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11913 4151 4150 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11914 0 4153 4152 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11915 4153 4152 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11916 1 4147 4146 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11917 4147 4146 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11918 1 4149 4148 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11919 4149 4148 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11920 1 4151 4150 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11921 4151 4150 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11922 1 4153 4152 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11923 4153 4152 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11924 1 4155 4154 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11925 4155 4154 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11926 1 4157 4156 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11927 4157 4156 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11928 1 4159 4158 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11929 4159 4158 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11930 1 4161 4160 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11931 4161 4160 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11932 0 4155 4154 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11933 4155 4154 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11934 0 4157 4156 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11935 4157 4156 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11936 0 4159 4158 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11937 4159 4158 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11938 0 4161 4160 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11939 4161 4160 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11940 352 604 4154 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11941 353 604 4155 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11942 354 604 4156 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11943 355 604 4157 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11944 356 604 4158 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11945 357 604 4159 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11946 358 604 4160 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11947 359 604 4161 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11948 4162 607 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11949 4163 607 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11950 4164 607 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11951 4165 607 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11952 4166 607 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m11953 4167 607 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11954 4168 607 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11955 4169 607 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m11956 0 4163 4162 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11957 4163 4162 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11958 0 4165 4164 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11959 4165 4164 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11960 0 4167 4166 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11961 4167 4166 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11962 0 4169 4168 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11963 4169 4168 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11964 1 4163 4162 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11965 4163 4162 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11966 1 4165 4164 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11967 4165 4164 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11968 1 4171 4170 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11969 4171 4170 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m11970 1 4173 4172 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11971 4173 4172 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11972 1 4167 4166 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11973 4167 4166 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11974 1 4169 4168 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11975 4169 4168 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11976 1 4175 4174 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m11977 4175 4174 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11978 1 4177 4176 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m11979 4177 4176 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m11980 0 4171 4170 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11981 4171 4170 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11982 0 4173 4172 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m11983 4173 4172 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m11984 0 4175 4174 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11985 4175 4174 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11986 0 4177 4176 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m11987 4177 4176 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m11988 352 612 4170 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m11989 353 612 4171 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11990 354 612 4172 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11991 355 612 4173 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11992 356 612 4174 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m11993 357 612 4175 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m11994 358 612 4176 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m11995 359 612 4177 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m11996 4178 616 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m11997 4179 616 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m11998 4180 616 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m11999 4181 616 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12000 4182 616 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12001 4183 616 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12002 4184 616 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12003 4185 616 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12004 0 4179 4178 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12005 4179 4178 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12006 0 4181 4180 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12007 4181 4180 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12008 0 4183 4182 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12009 4183 4182 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12010 0 4185 4184 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12011 4185 4184 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12012 1 4179 4178 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12013 4179 4178 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12014 1 4181 4180 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12015 4181 4180 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12016 1 4183 4182 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12017 4183 4182 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12018 1 4185 4184 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12019 4185 4184 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12020 1 4187 4186 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12021 4187 4186 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12022 1 4189 4188 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12023 4189 4188 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12024 1 4191 4190 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12025 4191 4190 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12026 1 4193 4192 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12027 4193 4192 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12028 0 4187 4186 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12029 4187 4186 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12030 0 4189 4188 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12031 4189 4188 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12032 0 4191 4190 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12033 4191 4190 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12034 0 4193 4192 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12035 4193 4192 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12036 352 620 4186 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12037 353 620 4187 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12038 354 620 4188 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12039 355 620 4189 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12040 356 620 4190 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12041 357 620 4191 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12042 358 620 4192 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12043 359 620 4193 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12044 4194 624 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12045 4195 624 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12046 4196 624 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12047 4197 624 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12048 4198 624 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12049 4199 624 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12050 4200 624 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12051 4201 624 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12052 0 4195 4194 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12053 4195 4194 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12054 0 4197 4196 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12055 4197 4196 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12056 0 4199 4198 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12057 4199 4198 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12058 0 4201 4200 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12059 4201 4200 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12060 1 4195 4194 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12061 4195 4194 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12062 1 4197 4196 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12063 4197 4196 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12064 1 4203 4202 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12065 4203 4202 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12066 1 4205 4204 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12067 4205 4204 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12068 1 4199 4198 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12069 4199 4198 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12070 1 4201 4200 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12071 4201 4200 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12072 1 4207 4206 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12073 4207 4206 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12074 1 4209 4208 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12075 4209 4208 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12076 0 4203 4202 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12077 4203 4202 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12078 0 4205 4204 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12079 4205 4204 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12080 0 4207 4206 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12081 4207 4206 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12082 0 4209 4208 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12083 4209 4208 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12084 352 628 4202 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12085 353 628 4203 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12086 354 628 4204 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12087 355 628 4205 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12088 356 628 4206 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12089 357 628 4207 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12090 358 628 4208 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12091 359 628 4209 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12092 4210 632 352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12093 4211 632 353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12094 4212 632 354 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12095 4213 632 355 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12096 4214 632 356 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12097 4215 632 357 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12098 4216 632 358 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12099 4217 632 359 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12100 0 4211 4210 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12101 4211 4210 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12102 0 4213 4212 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12103 4213 4212 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12104 0 4215 4214 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12105 4215 4214 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12106 0 4217 4216 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12107 4217 4216 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12108 1 4211 4210 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12109 4211 4210 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12110 1 4213 4212 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12111 4213 4212 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12112 1 4215 4214 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12113 4215 4214 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12114 1 4217 4216 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12115 4217 4216 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12116 1 4219 4218 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12117 4219 4218 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12118 1 4221 4220 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12119 4221 4220 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12120 1 4223 4222 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12121 4223 4222 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12122 1 4225 4224 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12123 4225 4224 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12124 0 4219 4218 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12125 4219 4218 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12126 0 4221 4220 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12127 4221 4220 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12128 0 4223 4222 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12129 4223 4222 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12130 0 4225 4224 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12131 4225 4224 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12132 139 380 4218 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12133 141 380 4219 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12134 142 380 4220 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12135 143 380 4221 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12136 144 380 4222 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12137 145 380 4223 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12138 146 380 4224 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12139 147 380 4225 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12140 4226 383 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12141 4227 383 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12142 4228 383 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12143 4229 383 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12144 4230 383 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12145 4231 383 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12146 4232 383 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12147 4233 383 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12148 0 4227 4226 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12149 4227 4226 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12150 0 4229 4228 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12151 4229 4228 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12152 0 4231 4230 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12153 4231 4230 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12154 0 4233 4232 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12155 4233 4232 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12156 1 4227 4226 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12157 4227 4226 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12158 1 4229 4228 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12159 4229 4228 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12160 1 4235 4234 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12161 4235 4234 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12162 1 4237 4236 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12163 4237 4236 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12164 1 4231 4230 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12165 4231 4230 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12166 1 4233 4232 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12167 4233 4232 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12168 1 4239 4238 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12169 4239 4238 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12170 1 4241 4240 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12171 4241 4240 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12172 0 4235 4234 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12173 4235 4234 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12174 0 4237 4236 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12175 4237 4236 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12176 0 4239 4238 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12177 4239 4238 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12178 0 4241 4240 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12179 4241 4240 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12180 139 388 4234 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12181 141 388 4235 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12182 142 388 4236 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12183 143 388 4237 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12184 144 388 4238 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12185 145 388 4239 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12186 146 388 4240 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12187 147 388 4241 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12188 4242 392 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12189 4243 392 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12190 4244 392 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12191 4245 392 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12192 4246 392 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12193 4247 392 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12194 4248 392 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12195 4249 392 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12196 0 4243 4242 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12197 4243 4242 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12198 0 4245 4244 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12199 4245 4244 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12200 0 4247 4246 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12201 4247 4246 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12202 0 4249 4248 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12203 4249 4248 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12204 1 4243 4242 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12205 4243 4242 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12206 1 4245 4244 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12207 4245 4244 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12208 1 4247 4246 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12209 4247 4246 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12210 1 4249 4248 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12211 4249 4248 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12212 1 4251 4250 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12213 4251 4250 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12214 1 4253 4252 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12215 4253 4252 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12216 1 4255 4254 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12217 4255 4254 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12218 1 4257 4256 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12219 4257 4256 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12220 0 4251 4250 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12221 4251 4250 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12222 0 4253 4252 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12223 4253 4252 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12224 0 4255 4254 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12225 4255 4254 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12226 0 4257 4256 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12227 4257 4256 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12228 139 396 4250 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12229 141 396 4251 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12230 142 396 4252 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12231 143 396 4253 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12232 144 396 4254 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12233 145 396 4255 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12234 146 396 4256 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12235 147 396 4257 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12236 4258 399 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12237 4259 399 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12238 4260 399 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12239 4261 399 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12240 4262 399 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12241 4263 399 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12242 4264 399 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12243 4265 399 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12244 0 4259 4258 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12245 4259 4258 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12246 0 4261 4260 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12247 4261 4260 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12248 0 4263 4262 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12249 4263 4262 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12250 0 4265 4264 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12251 4265 4264 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12252 1 4259 4258 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12253 4259 4258 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12254 1 4261 4260 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12255 4261 4260 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12256 1 4267 4266 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12257 4267 4266 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12258 1 4269 4268 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12259 4269 4268 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12260 1 4263 4262 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12261 4263 4262 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12262 1 4265 4264 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12263 4265 4264 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12264 1 4271 4270 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12265 4271 4270 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12266 1 4273 4272 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12267 4273 4272 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12268 0 4267 4266 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12269 4267 4266 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12270 0 4269 4268 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12271 4269 4268 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12272 0 4271 4270 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12273 4271 4270 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12274 0 4273 4272 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12275 4273 4272 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12276 139 404 4266 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12277 141 404 4267 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12278 142 404 4268 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12279 143 404 4269 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12280 144 404 4270 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12281 145 404 4271 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12282 146 404 4272 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12283 147 404 4273 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12284 4274 408 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12285 4275 408 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12286 4276 408 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12287 4277 408 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12288 4278 408 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12289 4279 408 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12290 4280 408 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12291 4281 408 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12292 0 4275 4274 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12293 4275 4274 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12294 0 4277 4276 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12295 4277 4276 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12296 0 4279 4278 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12297 4279 4278 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12298 0 4281 4280 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12299 4281 4280 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12300 1 4275 4274 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12301 4275 4274 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12302 1 4277 4276 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12303 4277 4276 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12304 1 4279 4278 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12305 4279 4278 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12306 1 4281 4280 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12307 4281 4280 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12308 1 4283 4282 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12309 4283 4282 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12310 1 4285 4284 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12311 4285 4284 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12312 1 4287 4286 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12313 4287 4286 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12314 1 4289 4288 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12315 4289 4288 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12316 0 4283 4282 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12317 4283 4282 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12318 0 4285 4284 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12319 4285 4284 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12320 0 4287 4286 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12321 4287 4286 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12322 0 4289 4288 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12323 4289 4288 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12324 139 412 4282 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12325 141 412 4283 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12326 142 412 4284 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12327 143 412 4285 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12328 144 412 4286 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12329 145 412 4287 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12330 146 412 4288 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12331 147 412 4289 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12332 4290 415 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12333 4291 415 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12334 4292 415 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12335 4293 415 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12336 4294 415 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12337 4295 415 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12338 4296 415 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12339 4297 415 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12340 0 4291 4290 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12341 4291 4290 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12342 0 4293 4292 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12343 4293 4292 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12344 0 4295 4294 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12345 4295 4294 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12346 0 4297 4296 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12347 4297 4296 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12348 1 4291 4290 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12349 4291 4290 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12350 1 4293 4292 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12351 4293 4292 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12352 1 4299 4298 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12353 4299 4298 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12354 1 4301 4300 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12355 4301 4300 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12356 1 4295 4294 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12357 4295 4294 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12358 1 4297 4296 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12359 4297 4296 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12360 1 4303 4302 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12361 4303 4302 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12362 1 4305 4304 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12363 4305 4304 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12364 0 4299 4298 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12365 4299 4298 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12366 0 4301 4300 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12367 4301 4300 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12368 0 4303 4302 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12369 4303 4302 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12370 0 4305 4304 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12371 4305 4304 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12372 139 420 4298 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12373 141 420 4299 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12374 142 420 4300 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12375 143 420 4301 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12376 144 420 4302 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12377 145 420 4303 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12378 146 420 4304 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12379 147 420 4305 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12380 4306 424 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12381 4307 424 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12382 4308 424 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12383 4309 424 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12384 4310 424 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12385 4311 424 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12386 4312 424 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12387 4313 424 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12388 0 4307 4306 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12389 4307 4306 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12390 0 4309 4308 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12391 4309 4308 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12392 0 4311 4310 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12393 4311 4310 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12394 0 4313 4312 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12395 4313 4312 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12396 1 4307 4306 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12397 4307 4306 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12398 1 4309 4308 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12399 4309 4308 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12400 1 4311 4310 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12401 4311 4310 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12402 1 4313 4312 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12403 4313 4312 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12404 1 4315 4314 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12405 4315 4314 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12406 1 4317 4316 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12407 4317 4316 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12408 1 4319 4318 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12409 4319 4318 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12410 1 4321 4320 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12411 4321 4320 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12412 0 4315 4314 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12413 4315 4314 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12414 0 4317 4316 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12415 4317 4316 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12416 0 4319 4318 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12417 4319 4318 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12418 0 4321 4320 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12419 4321 4320 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12420 139 428 4314 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12421 141 428 4315 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12422 142 428 4316 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12423 143 428 4317 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12424 144 428 4318 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12425 145 428 4319 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12426 146 428 4320 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12427 147 428 4321 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12428 4322 431 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12429 4323 431 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12430 4324 431 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12431 4325 431 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12432 4326 431 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12433 4327 431 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12434 4328 431 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12435 4329 431 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12436 0 4323 4322 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12437 4323 4322 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12438 0 4325 4324 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12439 4325 4324 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12440 0 4327 4326 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12441 4327 4326 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12442 0 4329 4328 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12443 4329 4328 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12444 1 4323 4322 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12445 4323 4322 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12446 1 4325 4324 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12447 4325 4324 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12448 1 4331 4330 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12449 4331 4330 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12450 1 4333 4332 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12451 4333 4332 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12452 1 4327 4326 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12453 4327 4326 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12454 1 4329 4328 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12455 4329 4328 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12456 1 4335 4334 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12457 4335 4334 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12458 1 4337 4336 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12459 4337 4336 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12460 0 4331 4330 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12461 4331 4330 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12462 0 4333 4332 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12463 4333 4332 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12464 0 4335 4334 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12465 4335 4334 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12466 0 4337 4336 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12467 4337 4336 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12468 139 436 4330 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12469 141 436 4331 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12470 142 436 4332 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12471 143 436 4333 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12472 144 436 4334 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12473 145 436 4335 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12474 146 436 4336 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12475 147 436 4337 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12476 4338 440 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12477 4339 440 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12478 4340 440 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12479 4341 440 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12480 4342 440 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12481 4343 440 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12482 4344 440 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12483 4345 440 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12484 0 4339 4338 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12485 4339 4338 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12486 0 4341 4340 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12487 4341 4340 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12488 0 4343 4342 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12489 4343 4342 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12490 0 4345 4344 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12491 4345 4344 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12492 1 4339 4338 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12493 4339 4338 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12494 1 4341 4340 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12495 4341 4340 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12496 1 4343 4342 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12497 4343 4342 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12498 1 4345 4344 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12499 4345 4344 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12500 1 4347 4346 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12501 4347 4346 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12502 1 4349 4348 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12503 4349 4348 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12504 1 4351 4350 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12505 4351 4350 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12506 1 4353 4352 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12507 4353 4352 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12508 0 4347 4346 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12509 4347 4346 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12510 0 4349 4348 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12511 4349 4348 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12512 0 4351 4350 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12513 4351 4350 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12514 0 4353 4352 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12515 4353 4352 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12516 139 444 4346 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12517 141 444 4347 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12518 142 444 4348 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12519 143 444 4349 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12520 144 444 4350 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12521 145 444 4351 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12522 146 444 4352 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12523 147 444 4353 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12524 4354 447 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12525 4355 447 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12526 4356 447 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12527 4357 447 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12528 4358 447 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12529 4359 447 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12530 4360 447 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12531 4361 447 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12532 0 4355 4354 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12533 4355 4354 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12534 0 4357 4356 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12535 4357 4356 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12536 0 4359 4358 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12537 4359 4358 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12538 0 4361 4360 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12539 4361 4360 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12540 1 4355 4354 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12541 4355 4354 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12542 1 4357 4356 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12543 4357 4356 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12544 1 4363 4362 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12545 4363 4362 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12546 1 4365 4364 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12547 4365 4364 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12548 1 4359 4358 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12549 4359 4358 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12550 1 4361 4360 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12551 4361 4360 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12552 1 4367 4366 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12553 4367 4366 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12554 1 4369 4368 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12555 4369 4368 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12556 0 4363 4362 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12557 4363 4362 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12558 0 4365 4364 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12559 4365 4364 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12560 0 4367 4366 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12561 4367 4366 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12562 0 4369 4368 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12563 4369 4368 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12564 139 452 4362 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12565 141 452 4363 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12566 142 452 4364 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12567 143 452 4365 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12568 144 452 4366 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12569 145 452 4367 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12570 146 452 4368 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12571 147 452 4369 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12572 4370 456 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12573 4371 456 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12574 4372 456 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12575 4373 456 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12576 4374 456 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12577 4375 456 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12578 4376 456 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12579 4377 456 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12580 0 4371 4370 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12581 4371 4370 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12582 0 4373 4372 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12583 4373 4372 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12584 0 4375 4374 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12585 4375 4374 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12586 0 4377 4376 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12587 4377 4376 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12588 1 4371 4370 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12589 4371 4370 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12590 1 4373 4372 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12591 4373 4372 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12592 1 4375 4374 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12593 4375 4374 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12594 1 4377 4376 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12595 4377 4376 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12596 1 4379 4378 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12597 4379 4378 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12598 1 4381 4380 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12599 4381 4380 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12600 1 4383 4382 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12601 4383 4382 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12602 1 4385 4384 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12603 4385 4384 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12604 0 4379 4378 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12605 4379 4378 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12606 0 4381 4380 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12607 4381 4380 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12608 0 4383 4382 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12609 4383 4382 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12610 0 4385 4384 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12611 4385 4384 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12612 139 460 4378 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12613 141 460 4379 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12614 142 460 4380 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12615 143 460 4381 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12616 144 460 4382 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12617 145 460 4383 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12618 146 460 4384 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12619 147 460 4385 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12620 4386 463 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12621 4387 463 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12622 4388 463 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12623 4389 463 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12624 4390 463 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12625 4391 463 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12626 4392 463 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12627 4393 463 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12628 0 4387 4386 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12629 4387 4386 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12630 0 4389 4388 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12631 4389 4388 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12632 0 4391 4390 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12633 4391 4390 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12634 0 4393 4392 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12635 4393 4392 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12636 1 4387 4386 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12637 4387 4386 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12638 1 4389 4388 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12639 4389 4388 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12640 1 4395 4394 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12641 4395 4394 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12642 1 4397 4396 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12643 4397 4396 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12644 1 4391 4390 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12645 4391 4390 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12646 1 4393 4392 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12647 4393 4392 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12648 1 4399 4398 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12649 4399 4398 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12650 1 4401 4400 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12651 4401 4400 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12652 0 4395 4394 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12653 4395 4394 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12654 0 4397 4396 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12655 4397 4396 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12656 0 4399 4398 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12657 4399 4398 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12658 0 4401 4400 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12659 4401 4400 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12660 139 468 4394 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12661 141 468 4395 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12662 142 468 4396 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12663 143 468 4397 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12664 144 468 4398 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12665 145 468 4399 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12666 146 468 4400 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12667 147 468 4401 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12668 4402 472 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12669 4403 472 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12670 4404 472 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12671 4405 472 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12672 4406 472 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12673 4407 472 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12674 4408 472 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12675 4409 472 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12676 0 4403 4402 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12677 4403 4402 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12678 0 4405 4404 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12679 4405 4404 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12680 0 4407 4406 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12681 4407 4406 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12682 0 4409 4408 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12683 4409 4408 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12684 1 4403 4402 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12685 4403 4402 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12686 1 4405 4404 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12687 4405 4404 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12688 1 4407 4406 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12689 4407 4406 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12690 1 4409 4408 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12691 4409 4408 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12692 1 4411 4410 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12693 4411 4410 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12694 1 4413 4412 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12695 4413 4412 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12696 1 4415 4414 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12697 4415 4414 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12698 1 4417 4416 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12699 4417 4416 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12700 0 4411 4410 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12701 4411 4410 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12702 0 4413 4412 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12703 4413 4412 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12704 0 4415 4414 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12705 4415 4414 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12706 0 4417 4416 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12707 4417 4416 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12708 139 476 4410 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12709 141 476 4411 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12710 142 476 4412 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12711 143 476 4413 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12712 144 476 4414 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12713 145 476 4415 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12714 146 476 4416 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12715 147 476 4417 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12716 4418 479 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12717 4419 479 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12718 4420 479 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12719 4421 479 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12720 4422 479 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12721 4423 479 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12722 4424 479 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12723 4425 479 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12724 0 4419 4418 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12725 4419 4418 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12726 0 4421 4420 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12727 4421 4420 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12728 0 4423 4422 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12729 4423 4422 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12730 0 4425 4424 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12731 4425 4424 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12732 1 4419 4418 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12733 4419 4418 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12734 1 4421 4420 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12735 4421 4420 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12736 1 4427 4426 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12737 4427 4426 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12738 1 4429 4428 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12739 4429 4428 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12740 1 4423 4422 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12741 4423 4422 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12742 1 4425 4424 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12743 4425 4424 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12744 1 4431 4430 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12745 4431 4430 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12746 1 4433 4432 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12747 4433 4432 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12748 0 4427 4426 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12749 4427 4426 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12750 0 4429 4428 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12751 4429 4428 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12752 0 4431 4430 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12753 4431 4430 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12754 0 4433 4432 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12755 4433 4432 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12756 139 484 4426 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12757 141 484 4427 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12758 142 484 4428 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12759 143 484 4429 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12760 144 484 4430 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12761 145 484 4431 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12762 146 484 4432 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12763 147 484 4433 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12764 4434 488 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12765 4435 488 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12766 4436 488 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12767 4437 488 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12768 4438 488 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12769 4439 488 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12770 4440 488 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12771 4441 488 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12772 0 4435 4434 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12773 4435 4434 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12774 0 4437 4436 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12775 4437 4436 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12776 0 4439 4438 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12777 4439 4438 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12778 0 4441 4440 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12779 4441 4440 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12780 1 4435 4434 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12781 4435 4434 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12782 1 4437 4436 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12783 4437 4436 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12784 1 4439 4438 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12785 4439 4438 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12786 1 4441 4440 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12787 4441 4440 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12788 1 4443 4442 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12789 4443 4442 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12790 1 4445 4444 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12791 4445 4444 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12792 1 4447 4446 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12793 4447 4446 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12794 1 4449 4448 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12795 4449 4448 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12796 0 4443 4442 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12797 4443 4442 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12798 0 4445 4444 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12799 4445 4444 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12800 0 4447 4446 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12801 4447 4446 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12802 0 4449 4448 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12803 4449 4448 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12804 139 492 4442 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12805 141 492 4443 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12806 142 492 4444 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12807 143 492 4445 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12808 144 492 4446 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12809 145 492 4447 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12810 146 492 4448 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12811 147 492 4449 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12812 4450 495 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12813 4451 495 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12814 4452 495 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12815 4453 495 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12816 4454 495 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12817 4455 495 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12818 4456 495 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12819 4457 495 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12820 0 4451 4450 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12821 4451 4450 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12822 0 4453 4452 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12823 4453 4452 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12824 0 4455 4454 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12825 4455 4454 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12826 0 4457 4456 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12827 4457 4456 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12828 1 4451 4450 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12829 4451 4450 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12830 1 4453 4452 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12831 4453 4452 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12832 1 4459 4458 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12833 4459 4458 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12834 1 4461 4460 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12835 4461 4460 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12836 1 4455 4454 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12837 4455 4454 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12838 1 4457 4456 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12839 4457 4456 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12840 1 4463 4462 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12841 4463 4462 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12842 1 4465 4464 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12843 4465 4464 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12844 0 4459 4458 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12845 4459 4458 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12846 0 4461 4460 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12847 4461 4460 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12848 0 4463 4462 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12849 4463 4462 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12850 0 4465 4464 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12851 4465 4464 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12852 139 500 4458 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12853 141 500 4459 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12854 142 500 4460 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12855 143 500 4461 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12856 144 500 4462 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12857 145 500 4463 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12858 146 500 4464 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12859 147 500 4465 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12860 4466 504 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12861 4467 504 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12862 4468 504 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12863 4469 504 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12864 4470 504 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12865 4471 504 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12866 4472 504 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12867 4473 504 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12868 0 4467 4466 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12869 4467 4466 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12870 0 4469 4468 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12871 4469 4468 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12872 0 4471 4470 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12873 4471 4470 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12874 0 4473 4472 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12875 4473 4472 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12876 1 4467 4466 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12877 4467 4466 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12878 1 4469 4468 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12879 4469 4468 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12880 1 4471 4470 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12881 4471 4470 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12882 1 4473 4472 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12883 4473 4472 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12884 1 4475 4474 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12885 4475 4474 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12886 1 4477 4476 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12887 4477 4476 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12888 1 4479 4478 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12889 4479 4478 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12890 1 4481 4480 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12891 4481 4480 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12892 0 4475 4474 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12893 4475 4474 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12894 0 4477 4476 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12895 4477 4476 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12896 0 4479 4478 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12897 4479 4478 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12898 0 4481 4480 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12899 4481 4480 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12900 139 508 4474 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12901 141 508 4475 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12902 142 508 4476 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12903 143 508 4477 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12904 144 508 4478 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12905 145 508 4479 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12906 146 508 4480 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12907 147 508 4481 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12908 4482 511 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12909 4483 511 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12910 4484 511 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12911 4485 511 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12912 4486 511 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12913 4487 511 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12914 4488 511 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12915 4489 511 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12916 0 4483 4482 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12917 4483 4482 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12918 0 4485 4484 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12919 4485 4484 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12920 0 4487 4486 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12921 4487 4486 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12922 0 4489 4488 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12923 4489 4488 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12924 1 4483 4482 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12925 4483 4482 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12926 1 4485 4484 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12927 4485 4484 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12928 1 4491 4490 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12929 4491 4490 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12930 1 4493 4492 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12931 4493 4492 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12932 1 4487 4486 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12933 4487 4486 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12934 1 4489 4488 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12935 4489 4488 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12936 1 4495 4494 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12937 4495 4494 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12938 1 4497 4496 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12939 4497 4496 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12940 0 4491 4490 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12941 4491 4490 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12942 0 4493 4492 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12943 4493 4492 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12944 0 4495 4494 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12945 4495 4494 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12946 0 4497 4496 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12947 4497 4496 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12948 139 516 4490 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12949 141 516 4491 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12950 142 516 4492 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12951 143 516 4493 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12952 144 516 4494 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m12953 145 516 4495 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12954 146 516 4496 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12955 147 516 4497 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m12956 4498 520 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m12957 4499 520 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12958 4500 520 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12959 4501 520 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12960 4502 520 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m12961 4503 520 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m12962 4504 520 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m12963 4505 520 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m12964 0 4499 4498 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12965 4499 4498 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12966 0 4501 4500 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12967 4501 4500 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12968 0 4503 4502 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12969 4503 4502 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12970 0 4505 4504 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12971 4505 4504 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12972 1 4499 4498 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12973 4499 4498 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12974 1 4501 4500 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12975 4501 4500 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12976 1 4503 4502 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12977 4503 4502 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12978 1 4505 4504 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12979 4505 4504 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12980 1 4507 4506 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12981 4507 4506 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m12982 1 4509 4508 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12983 4509 4508 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12984 1 4511 4510 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m12985 4511 4510 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12986 1 4513 4512 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m12987 4513 4512 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m12988 0 4507 4506 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12989 4507 4506 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12990 0 4509 4508 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m12991 4509 4508 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m12992 0 4511 4510 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12993 4511 4510 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12994 0 4513 4512 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m12995 4513 4512 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m12996 139 524 4506 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m12997 141 524 4507 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m12998 142 524 4508 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m12999 143 524 4509 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13000 144 524 4510 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13001 145 524 4511 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13002 146 524 4512 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13003 147 524 4513 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m13004 4514 527 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m13005 4515 527 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13006 4516 527 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13007 4517 527 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13008 4518 527 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13009 4519 527 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13010 4520 527 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13011 4521 527 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m13012 0 4515 4514 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13013 4515 4514 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13014 0 4517 4516 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13015 4517 4516 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13016 0 4519 4518 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13017 4519 4518 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13018 0 4521 4520 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13019 4521 4520 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13020 1 4515 4514 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13021 4515 4514 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13022 1 4517 4516 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13023 4517 4516 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13024 1 4523 4522 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13025 4523 4522 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m13026 1 4525 4524 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13027 4525 4524 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13028 1 4519 4518 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13029 4519 4518 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13030 1 4521 4520 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13031 4521 4520 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13032 1 4527 4526 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13033 4527 4526 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13034 1 4529 4528 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m13035 4529 4528 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13036 0 4523 4522 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13037 4523 4522 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13038 0 4525 4524 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13039 4525 4524 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13040 0 4527 4526 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13041 4527 4526 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13042 0 4529 4528 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13043 4529 4528 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13044 139 532 4522 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m13045 141 532 4523 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13046 142 532 4524 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13047 143 532 4525 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13048 144 532 4526 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13049 145 532 4527 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13050 146 532 4528 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13051 147 532 4529 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m13052 4530 536 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m13053 4531 536 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13054 4532 536 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13055 4533 536 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13056 4534 536 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13057 4535 536 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13058 4536 536 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13059 4537 536 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m13060 0 4531 4530 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13061 4531 4530 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13062 0 4533 4532 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13063 4533 4532 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13064 0 4535 4534 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13065 4535 4534 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13066 0 4537 4536 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13067 4537 4536 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13068 1 4531 4530 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13069 4531 4530 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13070 1 4533 4532 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13071 4533 4532 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13072 1 4535 4534 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13073 4535 4534 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13074 1 4537 4536 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13075 4537 4536 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13076 1 4539 4538 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13077 4539 4538 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m13078 1 4541 4540 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13079 4541 4540 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13080 1 4543 4542 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13081 4543 4542 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13082 1 4545 4544 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m13083 4545 4544 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13084 0 4539 4538 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13085 4539 4538 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13086 0 4541 4540 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13087 4541 4540 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13088 0 4543 4542 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13089 4543 4542 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13090 0 4545 4544 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13091 4545 4544 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13092 139 540 4538 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m13093 141 540 4539 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13094 142 540 4540 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13095 143 540 4541 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13096 144 540 4542 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13097 145 540 4543 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13098 146 540 4544 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13099 147 540 4545 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m13100 4546 543 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m13101 4547 543 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13102 4548 543 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13103 4549 543 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13104 4550 543 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13105 4551 543 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13106 4552 543 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13107 4553 543 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m13108 0 4547 4546 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13109 4547 4546 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13110 0 4549 4548 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13111 4549 4548 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13112 0 4551 4550 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13113 4551 4550 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13114 0 4553 4552 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13115 4553 4552 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13116 1 4547 4546 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13117 4547 4546 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13118 1 4549 4548 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13119 4549 4548 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13120 1 4555 4554 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13121 4555 4554 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m13122 1 4557 4556 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13123 4557 4556 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13124 1 4551 4550 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13125 4551 4550 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13126 1 4553 4552 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13127 4553 4552 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13128 1 4559 4558 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13129 4559 4558 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13130 1 4561 4560 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m13131 4561 4560 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13132 0 4555 4554 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13133 4555 4554 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13134 0 4557 4556 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13135 4557 4556 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13136 0 4559 4558 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13137 4559 4558 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13138 0 4561 4560 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13139 4561 4560 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13140 139 548 4554 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m13141 141 548 4555 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13142 142 548 4556 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13143 143 548 4557 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13144 144 548 4558 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13145 145 548 4559 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13146 146 548 4560 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13147 147 548 4561 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m13148 4562 552 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m13149 4563 552 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13150 4564 552 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13151 4565 552 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13152 4566 552 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13153 4567 552 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13154 4568 552 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13155 4569 552 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m13156 0 4563 4562 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13157 4563 4562 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13158 0 4565 4564 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13159 4565 4564 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13160 0 4567 4566 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13161 4567 4566 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13162 0 4569 4568 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13163 4569 4568 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13164 1 4563 4562 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13165 4563 4562 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13166 1 4565 4564 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13167 4565 4564 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13168 1 4567 4566 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13169 4567 4566 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13170 1 4569 4568 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13171 4569 4568 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13172 1 4571 4570 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13173 4571 4570 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m13174 1 4573 4572 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13175 4573 4572 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13176 1 4575 4574 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13177 4575 4574 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13178 1 4577 4576 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m13179 4577 4576 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13180 0 4571 4570 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13181 4571 4570 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13182 0 4573 4572 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13183 4573 4572 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13184 0 4575 4574 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13185 4575 4574 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13186 0 4577 4576 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13187 4577 4576 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13188 139 556 4570 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m13189 141 556 4571 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13190 142 556 4572 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13191 143 556 4573 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13192 144 556 4574 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13193 145 556 4575 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13194 146 556 4576 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13195 147 556 4577 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m13196 4578 559 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m13197 4579 559 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13198 4580 559 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13199 4581 559 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13200 4582 559 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13201 4583 559 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13202 4584 559 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13203 4585 559 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m13204 0 4579 4578 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13205 4579 4578 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13206 0 4581 4580 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13207 4581 4580 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13208 0 4583 4582 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13209 4583 4582 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13210 0 4585 4584 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13211 4585 4584 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13212 1 4579 4578 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13213 4579 4578 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13214 1 4581 4580 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13215 4581 4580 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13216 1 4587 4586 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13217 4587 4586 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m13218 1 4589 4588 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13219 4589 4588 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13220 1 4583 4582 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13221 4583 4582 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13222 1 4585 4584 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13223 4585 4584 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13224 1 4591 4590 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13225 4591 4590 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13226 1 4593 4592 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m13227 4593 4592 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13228 0 4587 4586 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13229 4587 4586 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13230 0 4589 4588 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13231 4589 4588 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13232 0 4591 4590 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13233 4591 4590 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13234 0 4593 4592 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13235 4593 4592 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13236 139 564 4586 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m13237 141 564 4587 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13238 142 564 4588 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13239 143 564 4589 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13240 144 564 4590 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13241 145 564 4591 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13242 146 564 4592 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13243 147 564 4593 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m13244 4594 568 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m13245 4595 568 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13246 4596 568 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13247 4597 568 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13248 4598 568 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13249 4599 568 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13250 4600 568 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13251 4601 568 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m13252 0 4595 4594 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13253 4595 4594 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13254 0 4597 4596 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13255 4597 4596 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13256 0 4599 4598 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13257 4599 4598 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13258 0 4601 4600 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13259 4601 4600 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13260 1 4595 4594 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13261 4595 4594 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13262 1 4597 4596 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13263 4597 4596 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13264 1 4599 4598 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13265 4599 4598 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13266 1 4601 4600 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13267 4601 4600 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13268 1 4603 4602 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13269 4603 4602 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m13270 1 4605 4604 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13271 4605 4604 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13272 1 4607 4606 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13273 4607 4606 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13274 1 4609 4608 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m13275 4609 4608 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13276 0 4603 4602 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13277 4603 4602 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13278 0 4605 4604 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13279 4605 4604 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13280 0 4607 4606 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13281 4607 4606 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13282 0 4609 4608 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13283 4609 4608 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13284 139 572 4602 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m13285 141 572 4603 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13286 142 572 4604 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13287 143 572 4605 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13288 144 572 4606 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13289 145 572 4607 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13290 146 572 4608 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13291 147 572 4609 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m13292 4610 575 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m13293 4611 575 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13294 4612 575 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13295 4613 575 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13296 4614 575 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13297 4615 575 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13298 4616 575 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13299 4617 575 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m13300 0 4611 4610 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13301 4611 4610 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13302 0 4613 4612 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13303 4613 4612 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13304 0 4615 4614 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13305 4615 4614 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13306 0 4617 4616 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13307 4617 4616 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13308 1 4611 4610 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13309 4611 4610 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13310 1 4613 4612 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13311 4613 4612 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13312 1 4619 4618 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13313 4619 4618 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m13314 1 4621 4620 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13315 4621 4620 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13316 1 4615 4614 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13317 4615 4614 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13318 1 4617 4616 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13319 4617 4616 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13320 1 4623 4622 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13321 4623 4622 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13322 1 4625 4624 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m13323 4625 4624 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13324 0 4619 4618 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13325 4619 4618 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13326 0 4621 4620 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13327 4621 4620 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13328 0 4623 4622 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13329 4623 4622 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13330 0 4625 4624 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13331 4625 4624 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13332 139 580 4618 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m13333 141 580 4619 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13334 142 580 4620 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13335 143 580 4621 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13336 144 580 4622 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13337 145 580 4623 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13338 146 580 4624 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13339 147 580 4625 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m13340 4626 584 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m13341 4627 584 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13342 4628 584 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13343 4629 584 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13344 4630 584 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13345 4631 584 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13346 4632 584 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13347 4633 584 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m13348 0 4627 4626 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13349 4627 4626 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13350 0 4629 4628 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13351 4629 4628 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13352 0 4631 4630 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13353 4631 4630 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13354 0 4633 4632 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13355 4633 4632 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13356 1 4627 4626 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13357 4627 4626 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13358 1 4629 4628 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13359 4629 4628 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13360 1 4631 4630 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13361 4631 4630 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13362 1 4633 4632 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13363 4633 4632 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13364 1 4635 4634 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13365 4635 4634 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m13366 1 4637 4636 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13367 4637 4636 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13368 1 4639 4638 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13369 4639 4638 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13370 1 4641 4640 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m13371 4641 4640 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13372 0 4635 4634 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13373 4635 4634 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13374 0 4637 4636 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13375 4637 4636 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13376 0 4639 4638 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13377 4639 4638 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13378 0 4641 4640 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13379 4641 4640 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13380 139 588 4634 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m13381 141 588 4635 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13382 142 588 4636 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13383 143 588 4637 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13384 144 588 4638 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13385 145 588 4639 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13386 146 588 4640 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13387 147 588 4641 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m13388 4642 591 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m13389 4643 591 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13390 4644 591 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13391 4645 591 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13392 4646 591 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13393 4647 591 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13394 4648 591 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13395 4649 591 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m13396 0 4643 4642 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13397 4643 4642 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13398 0 4645 4644 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13399 4645 4644 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13400 0 4647 4646 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13401 4647 4646 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13402 0 4649 4648 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13403 4649 4648 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13404 1 4643 4642 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13405 4643 4642 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13406 1 4645 4644 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13407 4645 4644 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13408 1 4651 4650 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13409 4651 4650 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m13410 1 4653 4652 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13411 4653 4652 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13412 1 4647 4646 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13413 4647 4646 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13414 1 4649 4648 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13415 4649 4648 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13416 1 4655 4654 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13417 4655 4654 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13418 1 4657 4656 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m13419 4657 4656 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13420 0 4651 4650 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13421 4651 4650 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13422 0 4653 4652 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13423 4653 4652 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13424 0 4655 4654 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13425 4655 4654 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13426 0 4657 4656 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13427 4657 4656 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13428 139 596 4650 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m13429 141 596 4651 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13430 142 596 4652 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13431 143 596 4653 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13432 144 596 4654 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13433 145 596 4655 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13434 146 596 4656 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13435 147 596 4657 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m13436 4658 600 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m13437 4659 600 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13438 4660 600 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13439 4661 600 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13440 4662 600 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13441 4663 600 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13442 4664 600 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13443 4665 600 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m13444 0 4659 4658 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13445 4659 4658 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13446 0 4661 4660 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13447 4661 4660 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13448 0 4663 4662 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13449 4663 4662 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13450 0 4665 4664 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13451 4665 4664 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13452 1 4659 4658 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13453 4659 4658 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13454 1 4661 4660 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13455 4661 4660 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13456 1 4663 4662 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13457 4663 4662 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13458 1 4665 4664 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13459 4665 4664 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13460 1 4667 4666 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13461 4667 4666 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m13462 1 4669 4668 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13463 4669 4668 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13464 1 4671 4670 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13465 4671 4670 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13466 1 4673 4672 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m13467 4673 4672 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13468 0 4667 4666 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13469 4667 4666 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13470 0 4669 4668 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13471 4669 4668 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13472 0 4671 4670 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13473 4671 4670 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13474 0 4673 4672 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13475 4673 4672 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13476 139 604 4666 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m13477 141 604 4667 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13478 142 604 4668 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13479 143 604 4669 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13480 144 604 4670 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13481 145 604 4671 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13482 146 604 4672 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13483 147 604 4673 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m13484 4674 607 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m13485 4675 607 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13486 4676 607 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13487 4677 607 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13488 4678 607 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13489 4679 607 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13490 4680 607 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13491 4681 607 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m13492 0 4675 4674 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13493 4675 4674 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13494 0 4677 4676 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13495 4677 4676 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13496 0 4679 4678 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13497 4679 4678 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13498 0 4681 4680 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13499 4681 4680 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13500 1 4675 4674 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13501 4675 4674 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13502 1 4677 4676 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13503 4677 4676 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13504 1 4683 4682 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13505 4683 4682 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m13506 1 4685 4684 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13507 4685 4684 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13508 1 4679 4678 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13509 4679 4678 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13510 1 4681 4680 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13511 4681 4680 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13512 1 4687 4686 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13513 4687 4686 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13514 1 4689 4688 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m13515 4689 4688 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13516 0 4683 4682 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13517 4683 4682 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13518 0 4685 4684 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13519 4685 4684 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13520 0 4687 4686 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13521 4687 4686 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13522 0 4689 4688 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13523 4689 4688 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13524 139 612 4682 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m13525 141 612 4683 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13526 142 612 4684 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13527 143 612 4685 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13528 144 612 4686 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13529 145 612 4687 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13530 146 612 4688 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13531 147 612 4689 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m13532 4690 616 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m13533 4691 616 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13534 4692 616 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13535 4693 616 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13536 4694 616 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13537 4695 616 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13538 4696 616 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13539 4697 616 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m13540 0 4691 4690 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13541 4691 4690 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13542 0 4693 4692 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13543 4693 4692 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13544 0 4695 4694 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13545 4695 4694 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13546 0 4697 4696 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13547 4697 4696 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13548 1 4691 4690 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13549 4691 4690 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13550 1 4693 4692 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13551 4693 4692 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13552 1 4695 4694 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13553 4695 4694 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13554 1 4697 4696 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13555 4697 4696 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13556 1 4699 4698 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13557 4699 4698 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m13558 1 4701 4700 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13559 4701 4700 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13560 1 4703 4702 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13561 4703 4702 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13562 1 4705 4704 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m13563 4705 4704 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13564 0 4699 4698 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13565 4699 4698 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13566 0 4701 4700 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13567 4701 4700 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13568 0 4703 4702 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13569 4703 4702 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13570 0 4705 4704 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13571 4705 4704 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13572 139 620 4698 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m13573 141 620 4699 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13574 142 620 4700 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13575 143 620 4701 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13576 144 620 4702 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13577 145 620 4703 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13578 146 620 4704 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13579 147 620 4705 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m13580 4706 624 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m13581 4707 624 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13582 4708 624 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13583 4709 624 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13584 4710 624 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13585 4711 624 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13586 4712 624 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13587 4713 624 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m13588 0 4707 4706 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13589 4707 4706 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13590 0 4709 4708 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13591 4709 4708 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13592 0 4711 4710 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13593 4711 4710 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13594 0 4713 4712 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13595 4713 4712 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13596 1 4707 4706 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13597 4707 4706 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13598 1 4709 4708 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13599 4709 4708 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13600 1 4715 4714 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13601 4715 4714 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=4.41e-12 ad=8.39e-12 ps=8.4e-06 pd=8.67e-06 
+ nrs=1 nrd=1.9 
m13602 1 4717 4716 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13603 4717 4716 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13604 1 4711 4710 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13605 4711 4710 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13606 1 4713 4712 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13607 4713 4712 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13608 1 4719 4718 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13609 4719 4718 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13610 1 4721 4720 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=4.41e-12 ps=8.67e-06 pd=8.4e-06 
+ nrs=1.9 nrd=1 
m13611 4721 4720 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13612 0 4715 4714 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13613 4715 4714 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13614 0 4717 4716 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13615 4717 4716 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13616 0 4719 4718 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13617 4719 4718 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13618 0 4721 4720 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13619 4721 4720 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13620 139 628 4714 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.229e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.79 nrd=1.52 
m13621 141 628 4715 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13622 142 628 4716 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13623 143 628 4717 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13624 144 628 4718 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.088e-11 ad=6.09e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.47 nrd=1.38 
m13625 145 628 4719 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.72e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.52 
m13626 146 628 4720 0 nenh l=1.1e-06 w=2.1e-06 
+ as=9.47e-12 ad=6.09e-12 ps=1.43e-05 pd=9e-06 
+ nrs=2.15 nrd=1.38 
m13627 147 628 4721 0 nenh l=1.1e-06 w=2.1e-06 
+ as=1.158e-11 ad=6.72e-12 ps=1.497e-05 pd=9e-06 
+ nrs=2.63 nrd=1.52 
m13628 4722 632 139 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.229e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.79 
m13629 4723 632 141 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13630 4724 632 142 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13631 4725 632 143 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13632 4726 632 144 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=1.088e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.38 nrd=2.47 
m13633 4727 632 145 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.52 nrd=2.15 
m13634 4728 632 146 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.09e-12 ad=9.47e-12 ps=9e-06 pd=1.43e-05 
+ nrs=1.38 nrd=2.15 
m13635 4729 632 147 0 nenh l=1.1e-06 w=2.1e-06 
+ as=6.72e-12 ad=1.158e-11 ps=9e-06 pd=1.497e-05 
+ nrs=1.52 nrd=2.63 
m13636 0 4723 4722 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13637 4723 4722 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13638 0 4725 4724 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.96e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.14 
m13639 4725 4724 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.12e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.04 nrd=1.06 
m13640 0 4727 4726 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13641 4727 4726 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13642 0 4729 4728 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.33e-12 ad=8.12e-12 ps=8.76e-06 pd=1.2e-05 
+ nrs=1.06 nrd=1.04 
m13643 4729 4728 0 0 nenh l=1.1e-06 w=2.8e-06 
+ as=8.96e-12 ad=8.33e-12 ps=1.2e-05 pd=8.76e-06 
+ nrs=1.14 nrd=1.06 
m13644 1 4723 4722 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13645 4723 4722 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13646 1 4725 4724 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13647 4725 4724 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13648 1 4727 4726 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13649 4727 4726 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13650 1 4729 4728 1 penh l=1.1e-06 w=2.1e-06 
+ as=8.39e-12 ad=2.94e-12 ps=8.67e-06 pd=7e-06 
+ nrs=1.9 nrd=0.67 
m13651 4729 4728 1 1 penh l=1.1e-06 w=2.1e-06 
+ as=2.94e-12 ad=8.39e-12 ps=7e-06 pd=8.67e-06 
+ nrs=0.67 nrd=1.9 
m13652 4730 4732 4731 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13653 4733 4734 4730 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13654 4730 4736 4735 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13655 4737 4738 4730 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13656 4739 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13657 4741 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13658 4739 196 4742 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13659 4731 197 4739 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13660 4743 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13661 4744 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13662 4741 198 4745 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13663 4733 199 4741 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13664 4743 200 4746 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13665 4735 201 4743 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13666 4744 202 4747 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13667 4737 203 4744 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13668 1 4742 4742 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13669 4731 4742 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13670 1 4745 4745 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13671 4733 4745 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13672 1 4746 4746 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13673 4735 4746 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13674 1 4747 4747 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13675 4737 4747 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13676 4748 4732 4749 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13677 4750 4734 4748 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13678 4748 4736 4751 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13679 4752 4738 4748 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13680 4753 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13681 4754 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13682 4753 222 4755 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13683 4749 223 4753 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13684 4756 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13685 4757 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13686 4754 224 4758 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13687 4750 225 4754 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13688 4756 226 4759 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13689 4751 227 4756 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13690 4757 228 4760 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13691 4752 229 4757 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13692 1 4755 4755 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13693 4749 4755 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13694 1 4758 4758 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13695 4750 4758 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13696 1 4759 4759 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13697 4751 4759 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13698 1 4760 4760 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13699 4752 4760 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13700 4761 4732 4762 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13701 4763 4734 4761 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13702 4761 4736 4764 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13703 4765 4738 4761 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13704 4766 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13705 4767 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13706 4766 248 4768 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13707 4762 249 4766 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13708 4769 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13709 4770 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13710 4767 250 4771 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13711 4763 251 4767 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13712 4769 252 4772 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13713 4764 253 4769 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13714 4770 254 4773 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13715 4765 255 4770 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13716 1 4768 4768 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13717 4762 4768 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13718 1 4771 4771 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13719 4763 4771 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13720 1 4772 4772 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13721 4764 4772 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13722 1 4773 4773 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13723 4765 4773 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13724 4774 4732 4775 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13725 4776 4734 4774 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13726 4774 4736 4777 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13727 4778 4738 4774 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13728 4779 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13729 4780 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13730 4779 274 4781 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13731 4775 275 4779 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13732 4782 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13733 4783 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13734 4780 276 4784 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13735 4776 277 4780 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13736 4782 278 4785 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13737 4777 279 4782 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13738 4783 280 4786 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13739 4778 281 4783 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13740 1 4781 4781 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13741 4775 4781 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13742 1 4784 4784 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13743 4776 4784 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13744 1 4785 4785 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13745 4777 4785 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13746 1 4786 4786 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13747 4778 4786 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13748 4787 4732 4788 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13749 4789 4734 4787 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13750 4787 4736 4790 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13751 4791 4738 4787 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13752 4792 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13753 4793 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13754 4792 300 4794 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13755 4788 301 4792 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13756 4795 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13757 4796 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13758 4793 302 4797 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13759 4789 303 4793 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13760 4795 304 4798 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13761 4790 305 4795 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13762 4796 306 4799 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13763 4791 307 4796 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13764 1 4794 4794 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13765 4788 4794 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13766 1 4797 4797 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13767 4789 4797 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13768 1 4798 4798 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13769 4790 4798 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13770 1 4799 4799 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13771 4791 4799 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13772 4800 4732 4801 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13773 4802 4734 4800 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13774 4800 4736 4803 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13775 4804 4738 4800 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13776 4805 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13777 4806 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13778 4805 326 4807 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13779 4801 327 4805 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13780 4808 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13781 4809 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13782 4806 328 4810 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13783 4802 329 4806 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13784 4808 330 4811 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13785 4803 331 4808 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13786 4809 332 4812 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13787 4804 333 4809 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13788 1 4807 4807 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13789 4801 4807 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13790 1 4810 4810 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13791 4802 4810 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13792 1 4811 4811 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13793 4803 4811 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13794 1 4812 4812 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13795 4804 4812 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13796 4813 4732 4814 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13797 4815 4734 4813 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13798 4813 4736 4816 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13799 4817 4738 4813 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13800 4818 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13801 4819 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13802 4818 352 4820 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13803 4814 353 4818 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13804 4821 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13805 4822 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13806 4819 354 4823 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13807 4815 355 4819 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13808 4821 356 4824 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13809 4816 357 4821 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13810 4822 358 4825 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13811 4817 359 4822 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13812 1 4820 4820 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13813 4814 4820 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13814 1 4823 4823 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13815 4815 4823 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13816 1 4824 4824 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13817 4816 4824 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13818 1 4825 4825 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13819 4817 4825 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13820 4826 4827 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m13821 4828 167 0 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=2.917e-11 ps=2.1e-05 pd=3.068e-05 
+ nrs=0.07 nrd=0.3 
m13822 4828 167 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m13823 4732 4826 0 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=2.917e-11 ps=2.1e-05 pd=3.068e-05 
+ nrs=0.07 nrd=0.3 
m13824 4732 4826 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m13825 4829 4827 0 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=2.917e-11 ps=1.12e-05 pd=3.068e-05 
+ nrs=0.07 nrd=0.3 
m13826 4826 4828 4829 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=6.86e-12 ps=2.1e-05 pd=1.12e-05 
+ nrs=0.07 nrd=0.07 
m13827 1 4828 4826 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m13828 4830 4828 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m13829 4831 4828 4830 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=6.86e-12 ps=1.12e-05 pd=2.1e-05 
+ nrs=0.07 nrd=0.07 
m13830 0 187 4831 0 nenh l=1.1e-06 w=9.8e-06 
+ as=2.917e-11 ad=6.86e-12 ps=3.068e-05 pd=1.12e-05 
+ nrs=0.3 nrd=0.07 
m13831 1 4830 4736 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m13832 0 4830 4736 0 nenh l=1.1e-06 w=9.8e-06 
+ as=2.917e-11 ad=6.86e-12 ps=3.068e-05 pd=2.1e-05 
+ nrs=0.3 nrd=0.07 
m13833 1 187 4830 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m13834 4832 4732 4833 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13835 4834 4734 4832 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13836 4832 4736 4835 0 nenh l=1.1e-06 w=2.8e-06 
+ as=1.96e-12 ad=2.8e-12 ps=7e-06 pd=8e-06 
+ nrs=0.25 nrd=0.36 
m13837 4836 4738 4832 0 nenh l=1.1e-06 w=2.8e-06 
+ as=2.8e-12 ad=1.96e-12 ps=8e-06 pd=7e-06 
+ nrs=0.36 nrd=0.25 
m13838 0 4837 4738 0 nenh l=1.1e-06 w=9.8e-06 
+ as=2.917e-11 ad=6.86e-12 ps=3.068e-05 pd=2.1e-05 
+ nrs=0.3 nrd=0.07 
m13839 1 4837 4738 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m13840 0 4838 4734 0 nenh l=1.1e-06 w=9.8e-06 
+ as=2.917e-11 ad=6.86e-12 ps=3.068e-05 pd=2.1e-05 
+ nrs=0.3 nrd=0.07 
m13841 4838 167 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m13842 4839 167 4838 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=6.86e-12 ps=1.12e-05 pd=2.1e-05 
+ nrs=0.07 nrd=0.07 
m13843 1 4838 4734 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m13844 0 4827 4839 0 nenh l=1.1e-06 w=9.8e-06 
+ as=2.917e-11 ad=6.86e-12 ps=3.068e-05 pd=1.12e-05 
+ nrs=0.3 nrd=0.07 
m13845 1 4827 4838 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m13846 4840 167 4837 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=6.86e-12 ps=1.12e-05 pd=2.1e-05 
+ nrs=0.07 nrd=0.07 
m13847 4837 167 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m13848 0 187 4840 0 nenh l=1.1e-06 w=9.8e-06 
+ as=2.917e-11 ad=6.86e-12 ps=3.068e-05 pd=1.12e-05 
+ nrs=0.3 nrd=0.07 
m13849 4841 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13850 4842 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13851 4841 139 4843 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13852 4833 141 4841 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13853 4844 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13854 4845 4740 0 0 nenh l=1.1e-06 w=4.9e-06 
+ as=2.005e-11 ad=1.458e-11 ps=1.432e-05 pd=1.534e-05 
+ nrs=0.84 nrd=0.61 
m13855 4842 142 4846 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13856 4834 143 4842 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13857 4844 144 4847 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13858 4835 145 4844 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13859 1 187 4837 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m13860 4845 146 4848 0 nenh l=1.1e-06 w=2.1e-06 
+ as=8.59e-12 ad=2.94e-12 ps=6.14e-06 pd=7e-06 
+ nrs=1.95 nrd=0.67 
m13861 4836 147 4845 0 nenh l=1.1e-06 w=2.1e-06 
+ as=2.1e-12 ad=8.59e-12 ps=6e-06 pd=6.14e-06 
+ nrs=0.48 nrd=1.95 
m13862 4827 187 0 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=2.917e-11 ps=2.1e-05 pd=3.068e-05 
+ nrs=0.07 nrd=0.3 
m13863 4827 187 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m13864 4740 4849 0 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=2.917e-11 ps=2.1e-05 pd=3.068e-05 
+ nrs=0.07 nrd=0.3 
m13865 4849 169 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=7.35e-12 ad=4.194e-11 ps=2.24e-05 pd=4.335e-05 
+ nrs=0.07 nrd=0.38 
m13866 4740 4849 1 1 penh l=1.1e-06 w=1.05e-05 
+ as=8.33e-12 ad=4.194e-11 ps=2.45e-05 pd=4.335e-05 
+ nrs=0.08 nrd=0.38 
m13867 0 4849 4740 0 nenh l=1.1e-06 w=9.8e-06 
+ as=2.917e-11 ad=6.86e-12 ps=3.068e-05 pd=2.1e-05 
+ nrs=0.3 nrd=0.07 
m13868 4850 169 4849 0 nenh l=1.1e-06 w=9.8e-06 
+ as=6.86e-12 ad=6.86e-12 ps=1.12e-05 pd=2.1e-05 
+ nrs=0.07 nrd=0.07 
m13869 1 185 4849 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=7.35e-12 ps=4.335e-05 pd=2.24e-05 
+ nrs=0.38 nrd=0.07 
m13870 0 185 4850 0 nenh l=1.1e-06 w=9.8e-06 
+ as=2.917e-11 ad=6.86e-12 ps=3.068e-05 pd=1.12e-05 
+ nrs=0.3 nrd=0.07 
m13871 1 4849 4740 1 penh l=1.1e-06 w=1.05e-05 
+ as=4.194e-11 ad=8.33e-12 ps=4.335e-05 pd=2.45e-05 
+ nrs=0.38 nrd=0.08 
m13872 1 4843 4843 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13873 4833 4843 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13874 1 4846 4846 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13875 4834 4846 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
m13876 1 4847 4847 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.568e-11 ps=2.89e-05 pd=2.24e-05 
+ nrs=0.57 nrd=0.32 
m13877 4835 4847 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.274e-11 ad=2.796e-11 ps=1.96e-05 pd=2.89e-05 
+ nrs=0.26 nrd=0.57 
m13878 1 4848 4848 1 penh l=1.1e-06 w=7e-06 
+ as=2.796e-11 ad=1.274e-11 ps=2.89e-05 pd=1.96e-05 
+ nrs=0.57 nrd=0.26 
m13879 4836 4848 1 1 penh l=1.1e-06 w=7e-06 
+ as=1.568e-11 ad=2.796e-11 ps=2.24e-05 pd=2.89e-05 
+ nrs=0.32 nrd=0.57 
c0 185 0 4.35e-13
c1 4740 0 2.16e-13
c2 147 0 3.29e-13
c3 146 0 3.45e-13
c4 145 0 3.46e-13
c5 144 0 3.31e-13
c6 143 0 3.29e-13
c7 142 0 3.46e-13
c8 141 0 3.46e-13
c9 139 0 3.31e-13
c10 4734 0 1.92e-13
c11 4738 0 2.09e-13
c12 4736 0 2e-13
c13 4732 0 1.92e-13
c14 359 0 3.29e-13
c15 358 0 3.45e-13
c16 357 0 3.46e-13
c17 356 0 3.31e-13
c18 355 0 3.29e-13
c19 354 0 3.46e-13
c20 353 0 3.46e-13
c21 352 0 3.3e-13
c22 333 0 3.29e-13
c23 332 0 3.45e-13
c24 331 0 3.46e-13
c25 330 0 3.31e-13
c26 329 0 3.29e-13
c27 328 0 3.46e-13
c28 327 0 3.46e-13
c29 326 0 3.3e-13
c30 307 0 3.29e-13
c31 306 0 3.45e-13
c32 305 0 3.46e-13
c33 304 0 3.31e-13
c34 303 0 3.29e-13
c35 302 0 3.46e-13
c36 301 0 3.46e-13
c37 300 0 3.3e-13
c38 281 0 3.29e-13
c39 280 0 3.45e-13
c40 279 0 3.46e-13
c41 278 0 3.31e-13
c42 277 0 3.29e-13
c43 276 0 3.46e-13
c44 275 0 3.46e-13
c45 274 0 3.3e-13
c46 255 0 3.29e-13
c47 254 0 3.45e-13
c48 253 0 3.46e-13
c49 252 0 3.31e-13
c50 251 0 3.29e-13
c51 250 0 3.46e-13
c52 249 0 3.46e-13
c53 248 0 3.3e-13
c54 229 0 3.29e-13
c55 228 0 3.45e-13
c56 227 0 3.46e-13
c57 226 0 3.31e-13
c58 225 0 3.29e-13
c59 224 0 3.46e-13
c60 223 0 3.46e-13
c61 222 0 3.3e-13
c62 203 0 3.29e-13
c63 202 0 3.45e-13
c64 201 0 3.46e-13
c65 200 0 3.31e-13
c66 199 0 3.29e-13
c67 198 0 3.46e-13
c68 197 0 3.46e-13
c69 196 0 3.3e-13
c70 632 0 2.32e-13
c71 628 0 2.32e-13
c72 624 0 2.32e-13
c73 620 0 2.32e-13
c74 616 0 2.31e-13
c75 612 0 2.31e-13
c76 607 0 2.31e-13
c77 604 0 2.31e-13
c78 600 0 2.31e-13
c79 596 0 2.31e-13
c80 591 0 2.31e-13
c81 588 0 2.31e-13
c82 584 0 2.31e-13
c83 580 0 2.31e-13
c84 575 0 2.31e-13
c85 572 0 2.31e-13
c86 568 0 2.31e-13
c87 564 0 2.31e-13
c88 559 0 2.31e-13
c89 556 0 2.31e-13
c90 552 0 2.31e-13
c91 548 0 2.31e-13
c92 543 0 2.31e-13
c93 540 0 2.31e-13
c94 536 0 2.31e-13
c95 532 0 2.31e-13
c96 527 0 2.31e-13
c97 524 0 2.31e-13
c98 520 0 2.31e-13
c99 516 0 2.31e-13
c100 511 0 2.31e-13
c101 508 0 2.31e-13
c102 504 0 2.31e-13
c103 500 0 2.31e-13
c104 495 0 2.31e-13
c105 492 0 2.31e-13
c106 488 0 2.31e-13
c107 484 0 2.31e-13
c108 479 0 2.31e-13
c109 476 0 2.31e-13
c110 472 0 2.31e-13
c111 468 0 2.31e-13
c112 463 0 2.31e-13
c113 460 0 2.31e-13
c114 456 0 2.31e-13
c115 452 0 2.31e-13
c116 447 0 2.31e-13
c117 444 0 2.31e-13
c118 440 0 2.31e-13
c119 436 0 2.31e-13
c120 431 0 2.31e-13
c121 428 0 2.31e-13
c122 424 0 2.31e-13
c123 420 0 2.31e-13
c124 415 0 2.31e-13
c125 412 0 2.31e-13
c126 408 0 2.31e-13
c127 404 0 2.31e-13
c128 399 0 2.31e-13
c129 396 0 2.31e-13
c130 392 0 2.31e-13
c131 388 0 2.31e-13
c132 383 0 2.31e-13
c133 380 0 2.31e-13
c134 140 0 1.728e-12
c135 150 0 3.87e-13
c136 148 0 3.87e-13
c137 151 0 3.94e-13
c138 149 0 3.95e-13
c139 182 0 1.96e-13
c140 185 0 1.97e-13
c141 183 0 2.21e-13
c142 172 0 2.11e-13
c143 162 0 2.43e-13
c144 159 0 2.74e-13
c145 156 0 2.5e-13
c146 153 0 2.53e-13
c147 43 0 4.79e-13
c148 26 0 4.88e-13
c149 17 0 4.87e-13
c150 5 0 4.75e-13
c151 8 0 5.2e-13
c152 7 0 4.88e-13
c153 6 0 4.62e-13
c154 76 0 4.91e-13
c155 1 0 1.1018e-11
Vid2 245 0 0 
Vid3 271 0 0 
Vid4 297 0 0 
Vid5 323 0 0 
Vid6 349 0 0 
Vid7 375 0 0 
Vresetbar 182 0 0 
Vphi1H 172 0 pwl (0 3 2e-08 3 2.1e-08 0 5e-08 0 
+ 5.1e-08 3 7e-08 3 7.1e-08 0 1e-07 0 
+ 1.01e-07 3 1.2e-07 3 1.21e-07 0 1.5e-07 0 
+ 1.51e-07 3 1.7e-07 3 1.71e-07 0 2e-07 0 
+ 2.01e-07 3 2.2e-07 3 2.21e-07 0 2.5e-07 0 
+ 2.51e-07 3 2.7e-07 3 2.71e-07 0 3e-07 0 
+ 3.01e-07 3 3.2e-07 3 3.21e-07 0 3.5e-07 0 
+ 3.51e-07 3 3.7e-07 3 3.71e-07 0 4e-07 0 
+ 4.01e-07 3 4.2e-07 3 4.21e-07 0 4.5e-07 0 
+ 4.51e-07 3 4.7e-07 3 4.71e-07 0 5e-07 0 
+ 5.01e-07 3 5.2e-07 3 5.21e-07 0 5.5e-07 0 
+ 5.51e-07 3 5.7e-07 3 5.71e-07 0 6e-07 0 
+ 6.01e-07 3 )
Vphi2H 185 0 pwl (0 0 2.5e-08 0 2.6e-08 3 4.5e-08 3 
+ 4.6e-08 0 5e-08 0 7.5e-08 0 7.6e-08 3 
+ 9.5e-08 3 9.6e-08 0 1e-07 0 1.25e-07 0 
+ 1.26e-07 3 1.45e-07 3 1.46e-07 0 1.5e-07 0 
+ 1.75e-07 0 1.76e-07 3 1.95e-07 3 1.96e-07 0 
+ 2e-07 0 2.25e-07 0 2.26e-07 3 2.45e-07 3 
+ 2.46e-07 0 2.5e-07 0 2.75e-07 0 2.76e-07 3 
+ 2.95e-07 3 2.96e-07 0 3e-07 0 3.25e-07 0 
+ 3.26e-07 3 3.45e-07 3 3.46e-07 0 3.5e-07 0 
+ 3.75e-07 0 3.76e-07 3 3.95e-07 3 3.96e-07 0 
+ 4e-07 0 4.25e-07 0 4.26e-07 3 4.45e-07 3 
+ 4.46e-07 0 4.5e-07 0 4.75e-07 0 4.76e-07 3 
+ 4.95e-07 3 4.96e-07 0 5e-07 0 5.25e-07 0 
+ 5.26e-07 3 5.45e-07 3 5.46e-07 0 5.5e-07 0 
+ 5.75e-07 0 5.76e-07 3 5.95e-07 3 5.96e-07 0 
+ 6e-07 0 )
Vphi1L 140 0 pwl (0 0 2e-08 0 2.1e-08 3 5e-08 3 
+ 5.1e-08 0 7e-08 0 7.1e-08 3 1e-07 3 
+ 1.01e-07 0 1.2e-07 0 1.21e-07 3 1.5e-07 3 
+ 1.51e-07 0 1.7e-07 0 1.71e-07 3 2e-07 3 
+ 2.01e-07 0 2.2e-07 0 2.21e-07 3 2.5e-07 3 
+ 2.51e-07 0 2.7e-07 0 2.71e-07 3 3e-07 3 
+ 3.01e-07 0 3.2e-07 0 3.21e-07 3 3.5e-07 3 
+ 3.51e-07 0 3.7e-07 0 3.71e-07 3 4e-07 3 
+ 4.01e-07 0 4.2e-07 0 4.21e-07 3 4.5e-07 3 
+ 4.51e-07 0 4.7e-07 0 4.71e-07 3 5e-07 3 
+ 5.01e-07 0 5.2e-07 0 5.21e-07 3 5.5e-07 3 
+ 5.51e-07 0 5.7e-07 0 5.71e-07 3 6e-07 3 
+ 6.01e-07 0 )
Vphi2L 183 0 pwl (0 3 2.5e-08 3 2.6e-08 0 4.5e-08 0 
+ 4.6e-08 3 5e-08 3 7.5e-08 3 7.6e-08 0 
+ 9.5e-08 0 9.6e-08 3 1e-07 3 1.25e-07 3 
+ 1.26e-07 0 1.45e-07 0 1.46e-07 3 1.5e-07 3 
+ 1.75e-07 3 1.76e-07 0 1.95e-07 0 1.96e-07 3 
+ 2e-07 3 2.25e-07 3 2.26e-07 0 2.45e-07 0 
+ 2.46e-07 3 2.5e-07 3 2.75e-07 3 2.76e-07 0 
+ 2.95e-07 0 2.96e-07 3 3e-07 3 3.25e-07 3 
+ 3.26e-07 0 3.45e-07 0 3.46e-07 3 3.5e-07 3 
+ 3.75e-07 3 3.76e-07 0 3.95e-07 0 3.96e-07 3 
+ 4e-07 3 4.25e-07 3 4.26e-07 0 4.45e-07 0 
+ 4.46e-07 3 4.5e-07 3 4.75e-07 3 4.76e-07 0 
+ 4.95e-07 0 4.96e-07 3 5e-07 3 5.25e-07 3 
+ 5.26e-07 0 5.45e-07 0 5.46e-07 3 5.5e-07 3 
+ 5.75e-07 3 5.76e-07 0 5.95e-07 0 5.96e-07 3 
+ 6e-07 3 )
Vid1 219 0 pwl (0 0 1e-07 0 1.01e-07 3 1.5e-07 3 
+ 1.51e-07 0 2e-07 0 2.01e-07 3 2.5e-07 3 
+ 2.51e-07 0 3.5e-07 0 3.51e-07 3 4e-07 3 
+ 4.01e-07 0 4.5e-07 0 4.51e-07 3 5.5e-07 3 
+ 5.51e-07 0 6e-07 0 6.01e-07 3 6.5e-07 3 
+ 6.51e-07 0 7.5e-07 0 7.51e-07 3 8e-07 3 
+ 8.01e-07 0 8.5e-07 0 8.51e-07 3 9.5e-07 3 
+ 9.51e-07 0 1e-06 0 1.001e-06 3 1.05e-06 3 
+ 1.051e-06 0 1.15e-06 0 1.151e-06 3 1.2e-06 3 
+ 1.201e-06 0 1.25e-06 0 1.251e-06 3 1.35e-06 3 
+ 1.351e-06 0 1.4e-06 0 1.401e-06 3 1.45e-06 3 
+ 1.451e-06 0 1.55e-06 0 1.551e-06 3 1.6e-06 3 
+ 1.601e-06 0 1.65e-06 0 1.651e-06 3 1.75e-06 3 
+ 1.751e-06 0 1.8e-06 0 1.801e-06 3 1.85e-06 3 
+ 1.851e-06 0 1.95e-06 0 1.951e-06 3 2e-06 3 
+ 2.001e-06 0 2.05e-06 0 2.051e-06 3 2.15e-06 3 
+ 2.151e-06 0 2.2e-06 0 2.201e-06 3 2.25e-06 3 
+ 2.251e-06 0 2.35e-06 0 2.351e-06 3 2.4e-06 3 
+ 2.401e-06 0 2.45e-06 0 2.451e-06 3 2.55e-06 3 
+ 2.551e-06 0 2.6e-06 0 2.601e-06 3 2.65e-06 3 
+ 2.651e-06 0 2.75e-06 0 2.751e-06 3 2.8e-06 3 
+ 2.801e-06 0 2.85e-06 0 2.851e-06 3 2.95e-06 3 
+ 2.951e-06 0 3e-06 0 3.001e-06 3 3.05e-06 3 
+ 3.051e-06 0 3.15e-06 0 3.151e-06 3 3.2e-06 3 
+ 3.201e-06 0 3.25e-06 0 3.251e-06 3 3.3e-06 3 
+ 3.301e-06 0 )
Vid8 184 0 pwl (0 0 1e-07 0 1.01e-07 3 1.5e-07 3 
+ 1.51e-07 0 2e-07 0 2.01e-07 3 2.5e-07 3 
+ 2.51e-07 0 3.5e-07 0 3.51e-07 3 4e-07 3 
+ 4.01e-07 0 4.5e-07 0 4.51e-07 3 5.5e-07 3 
+ 5.51e-07 0 6e-07 0 6.01e-07 3 6.5e-07 3 
+ 6.51e-07 0 7.5e-07 0 7.51e-07 3 8e-07 3 
+ 8.01e-07 0 8.5e-07 0 8.51e-07 3 9.5e-07 3 
+ 9.51e-07 0 1e-06 0 1.001e-06 3 1.05e-06 3 
+ 1.051e-06 0 1.15e-06 0 1.151e-06 3 1.2e-06 3 
+ 1.201e-06 0 1.25e-06 0 1.251e-06 3 1.35e-06 3 
+ 1.351e-06 0 1.4e-06 0 1.401e-06 3 1.45e-06 3 
+ 1.451e-06 0 1.55e-06 0 1.551e-06 3 1.6e-06 3 
+ 1.601e-06 0 1.65e-06 0 1.651e-06 3 1.75e-06 3 
+ 1.751e-06 0 1.8e-06 0 1.801e-06 3 1.85e-06 3 
+ 1.851e-06 0 1.95e-06 0 1.951e-06 3 2e-06 3 
+ 2.001e-06 0 2.05e-06 0 2.051e-06 3 2.15e-06 3 
+ 2.151e-06 0 2.2e-06 0 2.201e-06 3 2.25e-06 3 
+ 2.251e-06 0 2.35e-06 0 2.351e-06 3 2.4e-06 3 
+ 2.401e-06 0 2.45e-06 0 2.451e-06 3 2.55e-06 3 
+ 2.551e-06 0 2.6e-06 0 2.601e-06 3 2.65e-06 3 
+ 2.651e-06 0 2.75e-06 0 2.751e-06 3 2.8e-06 3 
+ 2.801e-06 0 2.85e-06 0 2.851e-06 3 2.95e-06 3 
+ 2.951e-06 0 3e-06 0 3.001e-06 3 3.05e-06 3 
+ 3.051e-06 0 3.15e-06 0 3.151e-06 3 3.2e-06 3 
+ 3.201e-06 0 3.25e-06 0 3.251e-06 3 3.3e-06 3 
+ 3.301e-06 0 )
Vrw 169 0 pwl (0 0 5e-07 0 5.01e-07 3 9e-07 3 
+ 9.01e-07 0 1.3e-06 0 1.301e-06 3 1.7e-06 3 
+ 1.701e-06 0 2.1e-06 0 2.101e-06 3 2.5e-06 3 
+ 2.501e-06 0 2.9e-06 0 2.901e-06 3 3.3e-06 3 
+ 3.301e-06 0 )
Vadr7 5 0 pwl (0 0 3.3e-06 0 )
Vadr6 6 0 pwl (0 0 3.3e-06 0 )
Vadr5 7 0 pwl (0 0 3.3e-06 0 )
Vadr4 8 0 pwl (0 0 3.3e-06 0 )
Vadr3 149 0 pwl (0 0 2e-07 0 2.01e-07 3 3e-07 3 
+ 3.01e-07 0 4e-07 0 4.01e-07 3 5e-07 3 
+ 5.01e-07 0 6e-07 0 6.01e-07 3 7e-07 3 
+ 7.01e-07 0 8e-07 0 8.01e-07 3 9e-07 3 
+ 9.01e-07 0 1e-06 0 1.001e-06 3 1.1e-06 3 
+ 1.101e-06 0 1.2e-06 0 1.201e-06 3 1.3e-06 3 
+ 1.301e-06 0 1.4e-06 0 1.401e-06 3 1.5e-06 3 
+ 1.501e-06 0 1.6e-06 0 1.601e-06 3 1.7e-06 3 
+ 1.701e-06 0 1.8e-06 0 1.801e-06 3 1.9e-06 3 
+ 1.901e-06 0 2e-06 0 2.001e-06 3 2.1e-06 3 
+ 2.101e-06 0 2.2e-06 0 2.201e-06 3 2.3e-06 3 
+ 2.301e-06 0 2.4e-06 0 2.401e-06 3 2.5e-06 3 
+ 2.501e-06 0 2.6e-06 0 2.601e-06 3 2.7e-06 3 
+ 2.701e-06 0 2.8e-06 0 2.801e-06 3 2.9e-06 3 
+ 2.901e-06 0 3e-06 0 3.001e-06 3 3.1e-06 3 
+ 3.101e-06 0 3.2e-06 0 3.201e-06 3 3.3e-06 3 
+ 3.301e-06 0 )
Vadr2 151 0 pwl (0 0 1.5e-07 0 1.51e-07 3 2e-07 3 
+ 2.01e-07 0 2.5e-07 0 2.51e-07 3 3e-07 3 
+ 3.01e-07 0 3.5e-07 0 3.51e-07 3 4e-07 3 
+ 4.01e-07 0 4.5e-07 0 4.51e-07 3 5e-07 3 
+ 5.01e-07 0 5.5e-07 0 5.51e-07 3 6e-07 3 
+ 6.01e-07 0 6.5e-07 0 6.51e-07 3 7e-07 3 
+ 7.01e-07 0 7.5e-07 0 7.51e-07 3 8e-07 3 
+ 8.01e-07 0 8.5e-07 0 8.51e-07 3 9e-07 3 
+ 9.01e-07 0 9.5e-07 0 9.51e-07 3 1e-06 3 
+ 1.001e-06 0 1.05e-06 0 1.051e-06 3 1.1e-06 3 
+ 1.101e-06 0 1.15e-06 0 1.151e-06 3 1.2e-06 3 
+ 1.201e-06 0 1.25e-06 0 1.251e-06 3 1.3e-06 3 
+ 1.301e-06 0 1.35e-06 0 1.351e-06 3 1.4e-06 3 
+ 1.401e-06 0 1.45e-06 0 1.451e-06 3 1.5e-06 3 
+ 1.501e-06 0 1.55e-06 0 1.551e-06 3 1.6e-06 3 
+ 1.601e-06 0 1.65e-06 0 1.651e-06 3 1.7e-06 3 
+ 1.701e-06 0 1.75e-06 0 1.751e-06 3 1.8e-06 3 
+ 1.801e-06 0 1.85e-06 0 1.851e-06 3 1.9e-06 3 
+ 1.901e-06 0 1.95e-06 0 1.951e-06 3 2e-06 3 
+ 2.001e-06 0 2.05e-06 0 2.051e-06 3 2.1e-06 3 
+ 2.101e-06 0 2.15e-06 0 2.151e-06 3 2.2e-06 3 
+ 2.201e-06 0 2.25e-06 0 2.251e-06 3 2.3e-06 3 
+ 2.301e-06 0 2.35e-06 0 2.351e-06 3 2.4e-06 3 
+ 2.401e-06 0 2.45e-06 0 2.451e-06 3 2.5e-06 3 
+ 2.501e-06 0 2.55e-06 0 2.551e-06 3 2.6e-06 3 
+ 2.601e-06 0 2.65e-06 0 2.651e-06 3 2.7e-06 3 
+ 2.701e-06 0 2.75e-06 0 2.751e-06 3 2.8e-06 3 
+ 2.801e-06 0 2.85e-06 0 2.851e-06 3 2.9e-06 3 
+ 2.901e-06 0 2.95e-06 0 2.951e-06 3 3e-06 3 
+ 3.001e-06 0 3.05e-06 0 3.051e-06 3 3.1e-06 3 
+ 3.101e-06 0 3.15e-06 0 3.151e-06 3 3.2e-06 3 
+ 3.201e-06 0 3.25e-06 0 3.251e-06 3 3.3e-06 3 
+ 3.301e-06 0 )
Vadr1 167 0 pwl (0 0 3e-07 0 3.01e-07 3 5e-07 3 
+ 5.01e-07 0 7e-07 0 7.01e-07 3 9e-07 3 
+ 9.01e-07 0 1.1e-06 0 1.101e-06 3 1.3e-06 3 
+ 1.301e-06 0 1.5e-06 0 1.501e-06 3 1.7e-06 3 
+ 1.701e-06 0 1.9e-06 0 1.901e-06 3 2.1e-06 3 
+ 2.101e-06 0 2.3e-06 0 2.301e-06 3 2.5e-06 3 
+ 2.501e-06 0 2.7e-06 0 2.701e-06 3 2.9e-06 3 
+ 2.901e-06 0 3.1e-06 0 3.101e-06 3 3.3e-06 3 
+ 3.301e-06 0 )
Vadr0 187 0 pwl (0 0 9e-07 0 9.01e-07 3 1.7e-06 3 
+ 1.701e-06 0 2.5e-06 0 2.501e-06 3 3.3e-06 3 
+ 3.301e-06 0 )
VVdd 1 0 3 
.options device temp=70 
.print TRAN v(140) v(169) v(153) v(156) v(620) v(624) 
+v(628) v(632) v(213) v(165) v(196) v(197) 
+v(198) v(199) v(139) v(141) v(142) v(143) 
+v(4740) v(4732) v(4734) v(4730) v(4832) 
*.options limpts=50000 itl5=50000
.options timeint abstol=1.0e-5 nlnearconv=1
.TRAN 1e-09 6e-07
.end
