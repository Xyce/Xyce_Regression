* This netlist is equivalent to Step 1 for the
* DotStep_fftAccurateOne.cir netlist.  It has VS1:VA=600.
***********************************************************

.TRAN 0 1
.OPTIONS FFT FFT_ACCURATE=1 FFTOUT=1

V1 1 0 SIN(0 600 1)
V3 3 0 SIN(0 200 2)
R1 1 2 1
R2 2 0 1
R3 3 2 1

.FFT V(2) NP=16 WINDOW=HANN FORMAT=UNORM
.PRINT TRAN V(1) V(2) V(3)

.END
