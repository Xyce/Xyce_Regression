* https://en.wikipedia.org/wiki/Lotka%E2%80%93Volterra_equations
*
* Also see chapter 2, example 2.10 of this book:
*
*  https://www.springer.com/us/book/9781461404774
*
* " Stochastic Approaches for Systems Biology"
*  Authors: Ullah, Mukhtar, Wolkenhauer, Olaf 
*-------------------------------------------------------------------------
VBASE BAS 0 0.5V
VEMIT  GND 0 0.0V
YRXN r1  BAS  GND  rxn1
+ transport=false  
+ scalerxn=false
+ dirichletbc=false
+ tecplotlevel=0
*-------------------------------------------------------------------------

.MODEL rxn1 rxn (LEVEL=1
+ REACTION_FILE=lotkaVolterraRxn
+ NUMBER_REGIONS=1
+ )

.options timeint debuglevel=-10   reltol=1.0e-5 

.TRAN 3.0E-8 30.0

.PRINT TRAN delimiter=tab N(yrxn!r1_000_conc_xspec) N(yrxn!r1_000_conc_yspec)

.END

