********************************************************
* Test .PRINT PCE ES for .DC for FORMAT = STD,
* CSV and NOINDEX.  Also output all of the samples
* for the quadrature points.
*
* See SON Bug 1231 for more details.
********************************************************

.global_param R1value={1000.0}
.global_param R2value={1000.0}

R2 1 0 {R2value}
R1 1 2 {R1value}
Von 2 0 5

.dc Von 5 5 1

.print dc v(1)
.PRINT PCE PRECISION=6 outputAllSamples=true
.PRINT PCE PRECISION=6 FORMAT=CSV FILE=pce-dc-prn.cir.PCE.csv
+ outputAllSamples=true
.PRINT PCE PRECISION=6 FORMAT=NOINDEX FILE=pce-dc-prn.cir.PCE.noindex.prn
+ outputAllSamples=true

.PCE
+ param=R1value
+ type=normal
+ means=1000.0
+ std_deviations=200.0

.options PCES
+ order=2
+ outputs={v(2)},{v(1)}

.options nonlin nox=0

.end
