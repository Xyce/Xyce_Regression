*********************************************************************
* This tests the error messages, from remeasure, that should occur
* if a TRAN mode measure is included in a netlist that is doing a 
* .DC analysis.  
* 
* See SON Bug 889 for more details.
*
*
*********************************************************************

vsrc1   1a 0 1
rload1a 1a 1b 0.1
rload1b 1b 0 1

.DC vsrc1 1 5 1
.print dc vsrc1:DCV0 v(1a) v(1b)

* Test what happens when a TRAN measure is requested in a .DC netlist 
* during remeasure
.MEASURE TRAN tranmax max v(1a)


.END


