****************************************************
* Test .PRINT AC SP() YP() ZP() output in radians.
*
* See SON Bug 1208 for more details.
****************************************************

* RC ladder circuit
* Note that all ports (P devices) must use a common
* Reference Node, which is 0 here.
P1 1  0  port=1  z0=50
P2 12 0  port=2  z0=50

C1 2 0 1e-2
Rgs 1 2 0.02

.subckt RCBlock IN OUT GND
R1 IN OUT 20
C1 IN OUT 1p
Cg1 OUT GND 1p
.ends

X1 2 3 0 RCBlock
X2 3 4 0 RCBlock
X3 4 5 0 RCBlock
X4 5 6 0 RCBlock
X5 6 7 0 RCBlock
X6 7 8 0 RCBlock
X7 8 9 0 RCBlock
X8 9 10 0 RCBlock
X9 10 11 0 RCBlock
X10 11 12 0 RCBlock

.AC DEC 10 10  1e5

.LIN DATAFORMAT=MA LINTYPE=S
*.LIN DATAFORMAT=MA LINTYPE=Y FILE=sparams-phase-in-degrees.yparams.s2p
*.LIN DATAFORMAT=MA LINTYPE=Z FILE=sparams-phase-in-degrees.zparams.s2p

.PRINT AC SP(1,1) SP(1,2) SP(2,1) SP(2,2)
+ YP(1,1) YP(1,2) YP(2,1) YP(2,2)
+ ZP(1,1) ZP(1,2) ZP(2,1) ZP(2,2)

.OPTIONS OUTPUT PHASE_OUTPUT_RADIANS=true

.END
