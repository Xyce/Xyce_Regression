test multiplier

Vin 1 0 1.0
Rin 1 2 1.0

Xtest1 2 3 test 
Xtest2 3 0 test 

.global_param Mval=2

.subckt test A B 
Xtest A B test2 M={Mval}
.ends

.global_param Mval2=2.5

.subckt test2 A B 
R1 A B 0.5 M={Mval2}
.ends

.DC Vin 1 1 1
.PRINT DC V(1) V(2) V(3) I(Vin) 

