* Lead Current test for inductors for a .NOISE analysis

* NOISE ANALYSIS: RESISTOR DIVIDER, AMP, AND HP FILTER
*
* RESISTOR DIVIDER
V1  1 0 DC 5.0 AC  1.0
R1  1 2 100K
R2  2 0 100K
*
* AMP AND HP FILTER
EAMP  3 0 2 0 1
RLP1  3 4 100
LLP1  4 4b 1m
VMON  4b 0 0

.OP
.NOISE  V(4)  V1  DEC  5 100 1e5
.PRINT NOISE VM(4) I(LLP1) I(VMON)

.END

