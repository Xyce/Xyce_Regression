* Transient sensitivity example, pulse source "dummy" file to provide variable 
* list to xyce_verify.  This file is not run as part of the test, just parsed.
.param cap=0.1u
.param res=1K

c1 1 0 cap
c2 2 0 cap
R1 1 3 res
R2 1 2 res

Vin 3 0 PULSE(0V 1V 0S 10US 10US 100US 220US)

* Transient commands
.tran 0 1.5ms 
.options timeint reltol=1e-6 abstol=1e-6

*comp V(2) offset=0.1
*comp V(2)_V1 offset=0.1
*comp V(2)_V2  offset=0.1
*comp V(2)_TD offset=10000.0
*comp V(2)_TR  offset=1500.0
*comp V(2)_TF offset=-1.0
*comp V(2)_PW   offset=1.0
*comp V(2)_PER  offset=100000.0

.print tran v(2) 
+ V(2)_V1
+V(2)_V2
+V(2)_TD
+V(2)_TR
+V(2)_TF
+V(2)_PW
+V(2)_PER

.end

