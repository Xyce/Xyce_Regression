* DC simulation for xyce
.options device temp=27
.subckt mysub c_x b_x e_x s_x
e_c c_v 0 c_x 0 -1
v_c c_v c 0
f_c c_x 0 v_c   1
e_b b_v 0 b_x 0 -1
v_b b_v b 0
f_b b_x 0 v_b   1
e_e e_v 0 e_x 0 -1
v_e e_v e 0
f_e e_x 0 v_e   1
e_s s_v 0 s_x 0 -1
v_s s_v s 0
f_s s_x 0 v_s   1
q1 c b e s mymodel
.model mymodel pnp level=12
+ IS=4.70047e-25
+ NF=1.09575
+ NR=1.020
+ IBEI=1.484e-23
+ NEI=1.302
+ IBEN=6.096e-18
+ NEN=2.081
+ IBCI=5.618e-24
+ NCI=1.110
+ IBCN=3.297e-14
+ NCN=2.000
+ RCX=10.26
+ RCI=0.001
+ RBX=122.23
+ RBI=0.001
+ RE=17.61
+ RS=1
+ RBP=1
+ VEF=800
+ VER=700
+ CJE=7e-15
+ CJC=11e-15
+ CJCP=3e-15
+ TF=2.3e-12
+ RTH=159.177
+ EA=1.1095
+ EAIE=1.489271313
+ EANE=1.489271313
+ EAIC=1.489271313
+ EANC=1.489271313
+ XRE=2
+ XRBX=2
+ XRBI=2
+ XRCX=2
+ XRCI=2
+ XRS=2
+ GMIN=0.0
.ends
v_c c c_b 0
e_c c_b 0 b 0 1
v_b b 0 0.49
v_e e 0 0
v_s s 0 0
x1 c b e s mysub
.dc v_b 0.50 2.00 0.01
.print dc V(b)
+ i(v_c)
+ i(v_b)
.end
