Netlist to Test the Xyce Voltage-Controlled Voltage Source Model
******************************************************************************
* Tier No.:	1                                                             
* Description:	Test of Xyce voltage controlled voltage source
*		model using a voltage amplifier circuit.  A transient ramped
*		analysis is performed to obtain the transfer
*		function characteristics of the circuit (i.e., Rin, 
*		Rout, and voltage gain, Vout/Vin) and node voltages.
* Input:	0-10V Ramped Source, V
* Output:	V(2), V(3), V(4), Rin, Rout, V(4)/VIN
* Circuit Elements: resistors (4), VCVS
* Analysis:
*		The VCVS, E, is controlled by the independent source, VIN,
*		in the circuit. The VCVS has a factor k*VIN=2*VIN, which gives
*			E = V(3) = 2 * VIN
*		The voltages at nodes 2 and 4 are
*			V(2) = VIN * R2/(R1+R2) = VIN * 0.9975
*			V(4) = V(3) * R4/(R3+R4) = VIN * 1.9231V
*		Additionally, Rin, Rout and the voltage gain are
*			Rin  = R1 + R2 = 100K + 250 =			100.25K
*			Rout = R3||R4 = 40||1K =			38.46 Ohms
*			V(4)/VIN = 					1.923 		
****************************************************************************** 
VIN 1 0 0V PWL(0.0 0.0 1.0 10.0)
E 3 0 1 0 2V
R1 1 2 250
R2 2 0 100K
R3 3 4 40
R4 4 0 1K
.TRAN 0.0 1.0
.PRINT TRAN V(1) V(2) V(3) V(4)
.END
