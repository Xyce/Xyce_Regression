*Test of bug fix for bug 864 (SON)
* Prior to the fix, Xyce would hang while parsing the expression in the
* parameter definition of "foo".  After the fix it exits with an error
* saying "Unable to resolve parameter FOO found in .PARAM statement."
*
vd d 0 dc 1.8
vg g 0 dc 0
xM1 d g 0 0 mymos w=0.4u l=3.57u
.dc vg 0 1.8 0.01
.print dc i(vd)
.subckt mymos 1 2 3 4 w=0 l=0
.param foo = '(meh != 1)'
r1 1 3 1k
r2 2 3 4k
r3 4 3 100
.ends mymos
.end
