* test of coupled inductor parameters on the .PRINT line
V1 1 0 SIN(0 1 1KHz)
R1 1 0 2
R2 2 0 2

* mutual inductor definition (nonlnear level=1)
L1 1 0 100
L2 2 0 100
K1 L1 L2 1.00 nlcore

* perturbation circuit
* test of coupled inductor parameters on the .PRINT line
V1b 1b 0 SIN(0 1 1KHz)
R1b 1b 0 2
R2b 2b 0 2

* mutual inductor definition (nonlnear level=1)
L1b 1b 0 {100+1e-5}
L2b 2b 0 100
K1b L1b L2b 1.00 nlcore

.model nlcore core level=2 c=0.001

.TRAN 0 0.3ms 
.PRINT TRAN V(2) {((V(2b)-V(2))/1.0e-5)}

.options timeint reltol=1e-6 abstol=1e-6 method=gear

.END 

