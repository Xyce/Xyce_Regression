Test for OCT capability in DC sweeps with expressions
*
VT1 4 0 0V
R1  4 5 10
R2  5 0 5

.param start=0.125
.param end=66
.param segs=3

.DC OCT VT1   {start} {end} {segs}
.print DC V(4) V(5)

.END

