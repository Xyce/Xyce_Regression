***********************************************************************
* Netlist to test that .SENS output in RAW format defaults to
* STD format (.prn file with an Index column)
*
* It uses a level=1 diode circuit
***********************************************************************
R1 1 2 0.0001
V2 2 0 0.21
V1 3 0 0.0
D2 1 3 DA

.MODEL DA D (RS=6.5e-05 IS=1.0e-09 N=1.037)

.SENS objfunc={I(V1)} param=DA:RS,DA:IS
.options SENSITIVITY adjoint=1 direct=0  STDOUTPUT=0
.DC V2 0.1 2.0 0.1
.print DC format=RAW v(2) I(V1)  
.print SENS format=raw v(2) I(V1)
.END

