Transmission Line Test Circuit
*
.OPTIONS TIMEINT ABSTOL=1e-04 RELTOL=1e-02 
.options PARALLEL partitioner=0

* Slow pulse to drive 10K lump dual microstrip or simple transfer load
VSLOW 1 22 DC 0 EXP(0v 10v 3ms 10ms 200ms 10ms)
RS 1 11 50

* Enable xtstcir for 10K lump dual microstrip transmission line
* Or enable RT, RB, & RG for simple transfer load
xtstcir 11 22 33 44 microstrip
* RT 11 33 50
* RB 22 44 50
* RG 22 0 1u

* Terminator
RL 33 44 10K

**************************************************************
.subckt microstrip 1 2 3 4 
xcouple1 1 2 3 4 l3dsub1
.ends microstrip
***********************************
*** subcircuit: l3dsc1
*** Parasitic Model: microstrip
*** Only one segment
***
.subckt l3dsc1 1 3 2 4 
C01 1 0 4.540e-12
RG01 1 0 7.816e+03
L1 1 5 3.718e-08
R1 5 2 4.300e-01
C1 2 0 4.540e-12
RG1 2 0 7.816e+03
C02 3 0 4.540e-12
RG02 3 0 7.816e+03
L2 3 6 3.668e-08
R2 6 4 4.184e-01
C2 4 0 4.540e-12
RG2 4 0 7.816e+03
CM012 1 3 5.288e-13
KM12 L1 L2 2.229e-01
CM12 2 4 5.288e-13
.ends l3dsc1
***********************************
*** subcircuit: l3dsub1
*** Parasitic Model: microstrip
*** All segments
***
.subckt l3dsub1 1 2 2001 2002 
X1 1 2 3 4 l3dsc1
X2 3 4 5 6 l3dsc1
X3 5 6 7 8 l3dsc1
X4 7 8 9 10 l3dsc1
X5 9 10 11 12 l3dsc1
X6 11 12 13 14 l3dsc1
X7 13 14 15 16 l3dsc1
X8 15 16 17 18 l3dsc1
X9 17 18 19 20 l3dsc1
X10 19 20 21 22 l3dsc1
X11 21 22 23 24 l3dsc1
X12 23 24 25 26 l3dsc1
X13 25 26 27 28 l3dsc1
X14 27 28 29 30 l3dsc1
X15 29 30 31 32 l3dsc1
X16 31 32 33 34 l3dsc1
X17 33 34 35 36 l3dsc1
X18 35 36 37 38 l3dsc1
X19 37 38 39 40 l3dsc1
X20 39 40 41 42 l3dsc1
X21 41 42 43 44 l3dsc1
X22 43 44 45 46 l3dsc1
X23 45 46 47 48 l3dsc1
X24 47 48 49 50 l3dsc1
X25 49 50 51 52 l3dsc1
X26 51 52 53 54 l3dsc1
X27 53 54 55 56 l3dsc1
X28 55 56 57 58 l3dsc1
X29 57 58 59 60 l3dsc1
X30 59 60 61 62 l3dsc1
X31 61 62 63 64 l3dsc1
X32 63 64 65 66 l3dsc1
X33 65 66 67 68 l3dsc1
X34 67 68 69 70 l3dsc1
X35 69 70 71 72 l3dsc1
X36 71 72 73 74 l3dsc1
X37 73 74 75 76 l3dsc1
X38 75 76 77 78 l3dsc1
X39 77 78 79 80 l3dsc1
X40 79 80 81 82 l3dsc1
X41 81 82 83 84 l3dsc1
X42 83 84 85 86 l3dsc1
X43 85 86 87 88 l3dsc1
X44 87 88 89 90 l3dsc1
X45 89 90 91 92 l3dsc1
X46 91 92 93 94 l3dsc1
X47 93 94 95 96 l3dsc1
X48 95 96 97 98 l3dsc1
X49 97 98 99 100 l3dsc1
X50 99 100 101 102 l3dsc1
X51 101 102 103 104 l3dsc1
X52 103 104 105 106 l3dsc1
X53 105 106 107 108 l3dsc1
X54 107 108 109 110 l3dsc1
X55 109 110 111 112 l3dsc1
X56 111 112 113 114 l3dsc1
X57 113 114 115 116 l3dsc1
X58 115 116 117 118 l3dsc1
X59 117 118 119 120 l3dsc1
X60 119 120 121 122 l3dsc1
X61 121 122 123 124 l3dsc1
X62 123 124 125 126 l3dsc1
X63 125 126 127 128 l3dsc1
X64 127 128 129 130 l3dsc1
X65 129 130 131 132 l3dsc1
X66 131 132 133 134 l3dsc1
X67 133 134 135 136 l3dsc1
X68 135 136 137 138 l3dsc1
X69 137 138 139 140 l3dsc1
X70 139 140 141 142 l3dsc1
X71 141 142 143 144 l3dsc1
X72 143 144 145 146 l3dsc1
X73 145 146 147 148 l3dsc1
X74 147 148 149 150 l3dsc1
X75 149 150 151 152 l3dsc1
X76 151 152 153 154 l3dsc1
X77 153 154 155 156 l3dsc1
X78 155 156 157 158 l3dsc1
X79 157 158 159 160 l3dsc1
X80 159 160 161 162 l3dsc1
X81 161 162 163 164 l3dsc1
X82 163 164 165 166 l3dsc1
X83 165 166 167 168 l3dsc1
X84 167 168 169 170 l3dsc1
X85 169 170 171 172 l3dsc1
X86 171 172 173 174 l3dsc1
X87 173 174 175 176 l3dsc1
X88 175 176 177 178 l3dsc1
X89 177 178 179 180 l3dsc1
X90 179 180 181 182 l3dsc1
X91 181 182 183 184 l3dsc1
X92 183 184 185 186 l3dsc1
X93 185 186 187 188 l3dsc1
X94 187 188 189 190 l3dsc1
X95 189 190 191 192 l3dsc1
X96 191 192 193 194 l3dsc1
X97 193 194 195 196 l3dsc1
X98 195 196 197 198 l3dsc1
X99 197 198 199 200 l3dsc1
X100 199 200 201 202 l3dsc1
X101 201 202 203 204 l3dsc1
X102 203 204 205 206 l3dsc1
X103 205 206 207 208 l3dsc1
X104 207 208 209 210 l3dsc1
X105 209 210 211 212 l3dsc1
X106 211 212 213 214 l3dsc1
X107 213 214 215 216 l3dsc1
X108 215 216 217 218 l3dsc1
X109 217 218 219 220 l3dsc1
X110 219 220 221 222 l3dsc1
X111 221 222 223 224 l3dsc1
X112 223 224 225 226 l3dsc1
X113 225 226 227 228 l3dsc1
X114 227 228 229 230 l3dsc1
X115 229 230 231 232 l3dsc1
X116 231 232 233 234 l3dsc1
X117 233 234 235 236 l3dsc1
X118 235 236 237 238 l3dsc1
X119 237 238 239 240 l3dsc1
X120 239 240 241 242 l3dsc1
X121 241 242 243 244 l3dsc1
X122 243 244 245 246 l3dsc1
X123 245 246 247 248 l3dsc1
X124 247 248 249 250 l3dsc1
X125 249 250 251 252 l3dsc1
X126 251 252 253 254 l3dsc1
X127 253 254 255 256 l3dsc1
X128 255 256 257 258 l3dsc1
X129 257 258 259 260 l3dsc1
X130 259 260 261 262 l3dsc1
X131 261 262 263 264 l3dsc1
X132 263 264 265 266 l3dsc1
X133 265 266 267 268 l3dsc1
X134 267 268 269 270 l3dsc1
X135 269 270 271 272 l3dsc1
X136 271 272 273 274 l3dsc1
X137 273 274 275 276 l3dsc1
X138 275 276 277 278 l3dsc1
X139 277 278 279 280 l3dsc1
X140 279 280 281 282 l3dsc1
X141 281 282 283 284 l3dsc1
X142 283 284 285 286 l3dsc1
X143 285 286 287 288 l3dsc1
X144 287 288 289 290 l3dsc1
X145 289 290 291 292 l3dsc1
X146 291 292 293 294 l3dsc1
X147 293 294 295 296 l3dsc1
X148 295 296 297 298 l3dsc1
X149 297 298 299 300 l3dsc1
X150 299 300 301 302 l3dsc1
X151 301 302 303 304 l3dsc1
X152 303 304 305 306 l3dsc1
X153 305 306 307 308 l3dsc1
X154 307 308 309 310 l3dsc1
X155 309 310 311 312 l3dsc1
X156 311 312 313 314 l3dsc1
X157 313 314 315 316 l3dsc1
X158 315 316 317 318 l3dsc1
X159 317 318 319 320 l3dsc1
X160 319 320 321 322 l3dsc1
X161 321 322 323 324 l3dsc1
X162 323 324 325 326 l3dsc1
X163 325 326 327 328 l3dsc1
X164 327 328 329 330 l3dsc1
X165 329 330 331 332 l3dsc1
X166 331 332 333 334 l3dsc1
X167 333 334 335 336 l3dsc1
X168 335 336 337 338 l3dsc1
X169 337 338 339 340 l3dsc1
X170 339 340 341 342 l3dsc1
X171 341 342 343 344 l3dsc1
X172 343 344 345 346 l3dsc1
X173 345 346 347 348 l3dsc1
X174 347 348 349 350 l3dsc1
X175 349 350 351 352 l3dsc1
X176 351 352 353 354 l3dsc1
X177 353 354 355 356 l3dsc1
X178 355 356 357 358 l3dsc1
X179 357 358 359 360 l3dsc1
X180 359 360 361 362 l3dsc1
X181 361 362 363 364 l3dsc1
X182 363 364 365 366 l3dsc1
X183 365 366 367 368 l3dsc1
X184 367 368 369 370 l3dsc1
X185 369 370 371 372 l3dsc1
X186 371 372 373 374 l3dsc1
X187 373 374 375 376 l3dsc1
X188 375 376 377 378 l3dsc1
X189 377 378 379 380 l3dsc1
X190 379 380 381 382 l3dsc1
X191 381 382 383 384 l3dsc1
X192 383 384 385 386 l3dsc1
X193 385 386 387 388 l3dsc1
X194 387 388 389 390 l3dsc1
X195 389 390 391 392 l3dsc1
X196 391 392 393 394 l3dsc1
X197 393 394 395 396 l3dsc1
X198 395 396 397 398 l3dsc1
X199 397 398 399 400 l3dsc1
X200 399 400 401 402 l3dsc1
X201 401 402 403 404 l3dsc1
X202 403 404 405 406 l3dsc1
X203 405 406 407 408 l3dsc1
X204 407 408 409 410 l3dsc1
X205 409 410 411 412 l3dsc1
X206 411 412 413 414 l3dsc1
X207 413 414 415 416 l3dsc1
X208 415 416 417 418 l3dsc1
X209 417 418 419 420 l3dsc1
X210 419 420 421 422 l3dsc1
X211 421 422 423 424 l3dsc1
X212 423 424 425 426 l3dsc1
X213 425 426 427 428 l3dsc1
X214 427 428 429 430 l3dsc1
X215 429 430 431 432 l3dsc1
X216 431 432 433 434 l3dsc1
X217 433 434 435 436 l3dsc1
X218 435 436 437 438 l3dsc1
X219 437 438 439 440 l3dsc1
X220 439 440 441 442 l3dsc1
X221 441 442 443 444 l3dsc1
X222 443 444 445 446 l3dsc1
X223 445 446 447 448 l3dsc1
X224 447 448 449 450 l3dsc1
X225 449 450 451 452 l3dsc1
X226 451 452 453 454 l3dsc1
X227 453 454 455 456 l3dsc1
X228 455 456 457 458 l3dsc1
X229 457 458 459 460 l3dsc1
X230 459 460 461 462 l3dsc1
X231 461 462 463 464 l3dsc1
X232 463 464 465 466 l3dsc1
X233 465 466 467 468 l3dsc1
X234 467 468 469 470 l3dsc1
X235 469 470 471 472 l3dsc1
X236 471 472 473 474 l3dsc1
X237 473 474 475 476 l3dsc1
X238 475 476 477 478 l3dsc1
X239 477 478 479 480 l3dsc1
X240 479 480 481 482 l3dsc1
X241 481 482 483 484 l3dsc1
X242 483 484 485 486 l3dsc1
X243 485 486 487 488 l3dsc1
X244 487 488 489 490 l3dsc1
X245 489 490 491 492 l3dsc1
X246 491 492 493 494 l3dsc1
X247 493 494 495 496 l3dsc1
X248 495 496 497 498 l3dsc1
X249 497 498 499 500 l3dsc1
X250 499 500 501 502 l3dsc1
X251 501 502 503 504 l3dsc1
X252 503 504 505 506 l3dsc1
X253 505 506 507 508 l3dsc1
X254 507 508 509 510 l3dsc1
X255 509 510 511 512 l3dsc1
X256 511 512 513 514 l3dsc1
X257 513 514 515 516 l3dsc1
X258 515 516 517 518 l3dsc1
X259 517 518 519 520 l3dsc1
X260 519 520 521 522 l3dsc1
X261 521 522 523 524 l3dsc1
X262 523 524 525 526 l3dsc1
X263 525 526 527 528 l3dsc1
X264 527 528 529 530 l3dsc1
X265 529 530 531 532 l3dsc1
X266 531 532 533 534 l3dsc1
X267 533 534 535 536 l3dsc1
X268 535 536 537 538 l3dsc1
X269 537 538 539 540 l3dsc1
X270 539 540 541 542 l3dsc1
X271 541 542 543 544 l3dsc1
X272 543 544 545 546 l3dsc1
X273 545 546 547 548 l3dsc1
X274 547 548 549 550 l3dsc1
X275 549 550 551 552 l3dsc1
X276 551 552 553 554 l3dsc1
X277 553 554 555 556 l3dsc1
X278 555 556 557 558 l3dsc1
X279 557 558 559 560 l3dsc1
X280 559 560 561 562 l3dsc1
X281 561 562 563 564 l3dsc1
X282 563 564 565 566 l3dsc1
X283 565 566 567 568 l3dsc1
X284 567 568 569 570 l3dsc1
X285 569 570 571 572 l3dsc1
X286 571 572 573 574 l3dsc1
X287 573 574 575 576 l3dsc1
X288 575 576 577 578 l3dsc1
X289 577 578 579 580 l3dsc1
X290 579 580 581 582 l3dsc1
X291 581 582 583 584 l3dsc1
X292 583 584 585 586 l3dsc1
X293 585 586 587 588 l3dsc1
X294 587 588 589 590 l3dsc1
X295 589 590 591 592 l3dsc1
X296 591 592 593 594 l3dsc1
X297 593 594 595 596 l3dsc1
X298 595 596 597 598 l3dsc1
X299 597 598 599 600 l3dsc1
X300 599 600 601 602 l3dsc1
X301 601 602 603 604 l3dsc1
X302 603 604 605 606 l3dsc1
X303 605 606 607 608 l3dsc1
X304 607 608 609 610 l3dsc1
X305 609 610 611 612 l3dsc1
X306 611 612 613 614 l3dsc1
X307 613 614 615 616 l3dsc1
X308 615 616 617 618 l3dsc1
X309 617 618 619 620 l3dsc1
X310 619 620 621 622 l3dsc1
X311 621 622 623 624 l3dsc1
X312 623 624 625 626 l3dsc1
X313 625 626 627 628 l3dsc1
X314 627 628 629 630 l3dsc1
X315 629 630 631 632 l3dsc1
X316 631 632 633 634 l3dsc1
X317 633 634 635 636 l3dsc1
X318 635 636 637 638 l3dsc1
X319 637 638 639 640 l3dsc1
X320 639 640 641 642 l3dsc1
X321 641 642 643 644 l3dsc1
X322 643 644 645 646 l3dsc1
X323 645 646 647 648 l3dsc1
X324 647 648 649 650 l3dsc1
X325 649 650 651 652 l3dsc1
X326 651 652 653 654 l3dsc1
X327 653 654 655 656 l3dsc1
X328 655 656 657 658 l3dsc1
X329 657 658 659 660 l3dsc1
X330 659 660 661 662 l3dsc1
X331 661 662 663 664 l3dsc1
X332 663 664 665 666 l3dsc1
X333 665 666 667 668 l3dsc1
X334 667 668 669 670 l3dsc1
X335 669 670 671 672 l3dsc1
X336 671 672 673 674 l3dsc1
X337 673 674 675 676 l3dsc1
X338 675 676 677 678 l3dsc1
X339 677 678 679 680 l3dsc1
X340 679 680 681 682 l3dsc1
X341 681 682 683 684 l3dsc1
X342 683 684 685 686 l3dsc1
X343 685 686 687 688 l3dsc1
X344 687 688 689 690 l3dsc1
X345 689 690 691 692 l3dsc1
X346 691 692 693 694 l3dsc1
X347 693 694 695 696 l3dsc1
X348 695 696 697 698 l3dsc1
X349 697 698 699 700 l3dsc1
X350 699 700 701 702 l3dsc1
X351 701 702 703 704 l3dsc1
X352 703 704 705 706 l3dsc1
X353 705 706 707 708 l3dsc1
X354 707 708 709 710 l3dsc1
X355 709 710 711 712 l3dsc1
X356 711 712 713 714 l3dsc1
X357 713 714 715 716 l3dsc1
X358 715 716 717 718 l3dsc1
X359 717 718 719 720 l3dsc1
X360 719 720 721 722 l3dsc1
X361 721 722 723 724 l3dsc1
X362 723 724 725 726 l3dsc1
X363 725 726 727 728 l3dsc1
X364 727 728 729 730 l3dsc1
X365 729 730 731 732 l3dsc1
X366 731 732 733 734 l3dsc1
X367 733 734 735 736 l3dsc1
X368 735 736 737 738 l3dsc1
X369 737 738 739 740 l3dsc1
X370 739 740 741 742 l3dsc1
X371 741 742 743 744 l3dsc1
X372 743 744 745 746 l3dsc1
X373 745 746 747 748 l3dsc1
X374 747 748 749 750 l3dsc1
X375 749 750 751 752 l3dsc1
X376 751 752 753 754 l3dsc1
X377 753 754 755 756 l3dsc1
X378 755 756 757 758 l3dsc1
X379 757 758 759 760 l3dsc1
X380 759 760 761 762 l3dsc1
X381 761 762 763 764 l3dsc1
X382 763 764 765 766 l3dsc1
X383 765 766 767 768 l3dsc1
X384 767 768 769 770 l3dsc1
X385 769 770 771 772 l3dsc1
X386 771 772 773 774 l3dsc1
X387 773 774 775 776 l3dsc1
X388 775 776 777 778 l3dsc1
X389 777 778 779 780 l3dsc1
X390 779 780 781 782 l3dsc1
X391 781 782 783 784 l3dsc1
X392 783 784 785 786 l3dsc1
X393 785 786 787 788 l3dsc1
X394 787 788 789 790 l3dsc1
X395 789 790 791 792 l3dsc1
X396 791 792 793 794 l3dsc1
X397 793 794 795 796 l3dsc1
X398 795 796 797 798 l3dsc1
X399 797 798 799 800 l3dsc1
X400 799 800 801 802 l3dsc1
X401 801 802 803 804 l3dsc1
X402 803 804 805 806 l3dsc1
X403 805 806 807 808 l3dsc1
X404 807 808 809 810 l3dsc1
X405 809 810 811 812 l3dsc1
X406 811 812 813 814 l3dsc1
X407 813 814 815 816 l3dsc1
X408 815 816 817 818 l3dsc1
X409 817 818 819 820 l3dsc1
X410 819 820 821 822 l3dsc1
X411 821 822 823 824 l3dsc1
X412 823 824 825 826 l3dsc1
X413 825 826 827 828 l3dsc1
X414 827 828 829 830 l3dsc1
X415 829 830 831 832 l3dsc1
X416 831 832 833 834 l3dsc1
X417 833 834 835 836 l3dsc1
X418 835 836 837 838 l3dsc1
X419 837 838 839 840 l3dsc1
X420 839 840 841 842 l3dsc1
X421 841 842 843 844 l3dsc1
X422 843 844 845 846 l3dsc1
X423 845 846 847 848 l3dsc1
X424 847 848 849 850 l3dsc1
X425 849 850 851 852 l3dsc1
X426 851 852 853 854 l3dsc1
X427 853 854 855 856 l3dsc1
X428 855 856 857 858 l3dsc1
X429 857 858 859 860 l3dsc1
X430 859 860 861 862 l3dsc1
X431 861 862 863 864 l3dsc1
X432 863 864 865 866 l3dsc1
X433 865 866 867 868 l3dsc1
X434 867 868 869 870 l3dsc1
X435 869 870 871 872 l3dsc1
X436 871 872 873 874 l3dsc1
X437 873 874 875 876 l3dsc1
X438 875 876 877 878 l3dsc1
X439 877 878 879 880 l3dsc1
X440 879 880 881 882 l3dsc1
X441 881 882 883 884 l3dsc1
X442 883 884 885 886 l3dsc1
X443 885 886 887 888 l3dsc1
X444 887 888 889 890 l3dsc1
X445 889 890 891 892 l3dsc1
X446 891 892 893 894 l3dsc1
X447 893 894 895 896 l3dsc1
X448 895 896 897 898 l3dsc1
X449 897 898 899 900 l3dsc1
X450 899 900 901 902 l3dsc1
X451 901 902 903 904 l3dsc1
X452 903 904 905 906 l3dsc1
X453 905 906 907 908 l3dsc1
X454 907 908 909 910 l3dsc1
X455 909 910 911 912 l3dsc1
X456 911 912 913 914 l3dsc1
X457 913 914 915 916 l3dsc1
X458 915 916 917 918 l3dsc1
X459 917 918 919 920 l3dsc1
X460 919 920 921 922 l3dsc1
X461 921 922 923 924 l3dsc1
X462 923 924 925 926 l3dsc1
X463 925 926 927 928 l3dsc1
X464 927 928 929 930 l3dsc1
X465 929 930 931 932 l3dsc1
X466 931 932 933 934 l3dsc1
X467 933 934 935 936 l3dsc1
X468 935 936 937 938 l3dsc1
X469 937 938 939 940 l3dsc1
X470 939 940 941 942 l3dsc1
X471 941 942 943 944 l3dsc1
X472 943 944 945 946 l3dsc1
X473 945 946 947 948 l3dsc1
X474 947 948 949 950 l3dsc1
X475 949 950 951 952 l3dsc1
X476 951 952 953 954 l3dsc1
X477 953 954 955 956 l3dsc1
X478 955 956 957 958 l3dsc1
X479 957 958 959 960 l3dsc1
X480 959 960 961 962 l3dsc1
X481 961 962 963 964 l3dsc1
X482 963 964 965 966 l3dsc1
X483 965 966 967 968 l3dsc1
X484 967 968 969 970 l3dsc1
X485 969 970 971 972 l3dsc1
X486 971 972 973 974 l3dsc1
X487 973 974 975 976 l3dsc1
X488 975 976 977 978 l3dsc1
X489 977 978 979 980 l3dsc1
X490 979 980 981 982 l3dsc1
X491 981 982 983 984 l3dsc1
X492 983 984 985 986 l3dsc1
X493 985 986 987 988 l3dsc1
X494 987 988 989 990 l3dsc1
X495 989 990 991 992 l3dsc1
X496 991 992 993 994 l3dsc1
X497 993 994 995 996 l3dsc1
X498 995 996 997 998 l3dsc1
X499 997 998 999 1000 l3dsc1
X500 999 1000 1001 1002 l3dsc1
X501 1001 1002 1003 1004 l3dsc1
X502 1003 1004 1005 1006 l3dsc1
X503 1005 1006 1007 1008 l3dsc1
X504 1007 1008 1009 1010 l3dsc1
X505 1009 1010 1011 1012 l3dsc1
X506 1011 1012 1013 1014 l3dsc1
X507 1013 1014 1015 1016 l3dsc1
X508 1015 1016 1017 1018 l3dsc1
X509 1017 1018 1019 1020 l3dsc1
X510 1019 1020 1021 1022 l3dsc1
X511 1021 1022 1023 1024 l3dsc1
X512 1023 1024 1025 1026 l3dsc1
X513 1025 1026 1027 1028 l3dsc1
X514 1027 1028 1029 1030 l3dsc1
X515 1029 1030 1031 1032 l3dsc1
X516 1031 1032 1033 1034 l3dsc1
X517 1033 1034 1035 1036 l3dsc1
X518 1035 1036 1037 1038 l3dsc1
X519 1037 1038 1039 1040 l3dsc1
X520 1039 1040 1041 1042 l3dsc1
X521 1041 1042 1043 1044 l3dsc1
X522 1043 1044 1045 1046 l3dsc1
X523 1045 1046 1047 1048 l3dsc1
X524 1047 1048 1049 1050 l3dsc1
X525 1049 1050 1051 1052 l3dsc1
X526 1051 1052 1053 1054 l3dsc1
X527 1053 1054 1055 1056 l3dsc1
X528 1055 1056 1057 1058 l3dsc1
X529 1057 1058 1059 1060 l3dsc1
X530 1059 1060 1061 1062 l3dsc1
X531 1061 1062 1063 1064 l3dsc1
X532 1063 1064 1065 1066 l3dsc1
X533 1065 1066 1067 1068 l3dsc1
X534 1067 1068 1069 1070 l3dsc1
X535 1069 1070 1071 1072 l3dsc1
X536 1071 1072 1073 1074 l3dsc1
X537 1073 1074 1075 1076 l3dsc1
X538 1075 1076 1077 1078 l3dsc1
X539 1077 1078 1079 1080 l3dsc1
X540 1079 1080 1081 1082 l3dsc1
X541 1081 1082 1083 1084 l3dsc1
X542 1083 1084 1085 1086 l3dsc1
X543 1085 1086 1087 1088 l3dsc1
X544 1087 1088 1089 1090 l3dsc1
X545 1089 1090 1091 1092 l3dsc1
X546 1091 1092 1093 1094 l3dsc1
X547 1093 1094 1095 1096 l3dsc1
X548 1095 1096 1097 1098 l3dsc1
X549 1097 1098 1099 1100 l3dsc1
X550 1099 1100 1101 1102 l3dsc1
X551 1101 1102 1103 1104 l3dsc1
X552 1103 1104 1105 1106 l3dsc1
X553 1105 1106 1107 1108 l3dsc1
X554 1107 1108 1109 1110 l3dsc1
X555 1109 1110 1111 1112 l3dsc1
X556 1111 1112 1113 1114 l3dsc1
X557 1113 1114 1115 1116 l3dsc1
X558 1115 1116 1117 1118 l3dsc1
X559 1117 1118 1119 1120 l3dsc1
X560 1119 1120 1121 1122 l3dsc1
X561 1121 1122 1123 1124 l3dsc1
X562 1123 1124 1125 1126 l3dsc1
X563 1125 1126 1127 1128 l3dsc1
X564 1127 1128 1129 1130 l3dsc1
X565 1129 1130 1131 1132 l3dsc1
X566 1131 1132 1133 1134 l3dsc1
X567 1133 1134 1135 1136 l3dsc1
X568 1135 1136 1137 1138 l3dsc1
X569 1137 1138 1139 1140 l3dsc1
X570 1139 1140 1141 1142 l3dsc1
X571 1141 1142 1143 1144 l3dsc1
X572 1143 1144 1145 1146 l3dsc1
X573 1145 1146 1147 1148 l3dsc1
X574 1147 1148 1149 1150 l3dsc1
X575 1149 1150 1151 1152 l3dsc1
X576 1151 1152 1153 1154 l3dsc1
X577 1153 1154 1155 1156 l3dsc1
X578 1155 1156 1157 1158 l3dsc1
X579 1157 1158 1159 1160 l3dsc1
X580 1159 1160 1161 1162 l3dsc1
X581 1161 1162 1163 1164 l3dsc1
X582 1163 1164 1165 1166 l3dsc1
X583 1165 1166 1167 1168 l3dsc1
X584 1167 1168 1169 1170 l3dsc1
X585 1169 1170 1171 1172 l3dsc1
X586 1171 1172 1173 1174 l3dsc1
X587 1173 1174 1175 1176 l3dsc1
X588 1175 1176 1177 1178 l3dsc1
X589 1177 1178 1179 1180 l3dsc1
X590 1179 1180 1181 1182 l3dsc1
X591 1181 1182 1183 1184 l3dsc1
X592 1183 1184 1185 1186 l3dsc1
X593 1185 1186 1187 1188 l3dsc1
X594 1187 1188 1189 1190 l3dsc1
X595 1189 1190 1191 1192 l3dsc1
X596 1191 1192 1193 1194 l3dsc1
X597 1193 1194 1195 1196 l3dsc1
X598 1195 1196 1197 1198 l3dsc1
X599 1197 1198 1199 1200 l3dsc1
X600 1199 1200 1201 1202 l3dsc1
X601 1201 1202 1203 1204 l3dsc1
X602 1203 1204 1205 1206 l3dsc1
X603 1205 1206 1207 1208 l3dsc1
X604 1207 1208 1209 1210 l3dsc1
X605 1209 1210 1211 1212 l3dsc1
X606 1211 1212 1213 1214 l3dsc1
X607 1213 1214 1215 1216 l3dsc1
X608 1215 1216 1217 1218 l3dsc1
X609 1217 1218 1219 1220 l3dsc1
X610 1219 1220 1221 1222 l3dsc1
X611 1221 1222 1223 1224 l3dsc1
X612 1223 1224 1225 1226 l3dsc1
X613 1225 1226 1227 1228 l3dsc1
X614 1227 1228 1229 1230 l3dsc1
X615 1229 1230 1231 1232 l3dsc1
X616 1231 1232 1233 1234 l3dsc1
X617 1233 1234 1235 1236 l3dsc1
X618 1235 1236 1237 1238 l3dsc1
X619 1237 1238 1239 1240 l3dsc1
X620 1239 1240 1241 1242 l3dsc1
X621 1241 1242 1243 1244 l3dsc1
X622 1243 1244 1245 1246 l3dsc1
X623 1245 1246 1247 1248 l3dsc1
X624 1247 1248 1249 1250 l3dsc1
X625 1249 1250 1251 1252 l3dsc1
X626 1251 1252 1253 1254 l3dsc1
X627 1253 1254 1255 1256 l3dsc1
X628 1255 1256 1257 1258 l3dsc1
X629 1257 1258 1259 1260 l3dsc1
X630 1259 1260 1261 1262 l3dsc1
X631 1261 1262 1263 1264 l3dsc1
X632 1263 1264 1265 1266 l3dsc1
X633 1265 1266 1267 1268 l3dsc1
X634 1267 1268 1269 1270 l3dsc1
X635 1269 1270 1271 1272 l3dsc1
X636 1271 1272 1273 1274 l3dsc1
X637 1273 1274 1275 1276 l3dsc1
X638 1275 1276 1277 1278 l3dsc1
X639 1277 1278 1279 1280 l3dsc1
X640 1279 1280 1281 1282 l3dsc1
X641 1281 1282 1283 1284 l3dsc1
X642 1283 1284 1285 1286 l3dsc1
X643 1285 1286 1287 1288 l3dsc1
X644 1287 1288 1289 1290 l3dsc1
X645 1289 1290 1291 1292 l3dsc1
X646 1291 1292 1293 1294 l3dsc1
X647 1293 1294 1295 1296 l3dsc1
X648 1295 1296 1297 1298 l3dsc1
X649 1297 1298 1299 1300 l3dsc1
X650 1299 1300 1301 1302 l3dsc1
X651 1301 1302 1303 1304 l3dsc1
X652 1303 1304 1305 1306 l3dsc1
X653 1305 1306 1307 1308 l3dsc1
X654 1307 1308 1309 1310 l3dsc1
X655 1309 1310 1311 1312 l3dsc1
X656 1311 1312 1313 1314 l3dsc1
X657 1313 1314 1315 1316 l3dsc1
X658 1315 1316 1317 1318 l3dsc1
X659 1317 1318 1319 1320 l3dsc1
X660 1319 1320 1321 1322 l3dsc1
X661 1321 1322 1323 1324 l3dsc1
X662 1323 1324 1325 1326 l3dsc1
X663 1325 1326 1327 1328 l3dsc1
X664 1327 1328 1329 1330 l3dsc1
X665 1329 1330 1331 1332 l3dsc1
X666 1331 1332 1333 1334 l3dsc1
X667 1333 1334 1335 1336 l3dsc1
X668 1335 1336 1337 1338 l3dsc1
X669 1337 1338 1339 1340 l3dsc1
X670 1339 1340 1341 1342 l3dsc1
X671 1341 1342 1343 1344 l3dsc1
X672 1343 1344 1345 1346 l3dsc1
X673 1345 1346 1347 1348 l3dsc1
X674 1347 1348 1349 1350 l3dsc1
X675 1349 1350 1351 1352 l3dsc1
X676 1351 1352 1353 1354 l3dsc1
X677 1353 1354 1355 1356 l3dsc1
X678 1355 1356 1357 1358 l3dsc1
X679 1357 1358 1359 1360 l3dsc1
X680 1359 1360 1361 1362 l3dsc1
X681 1361 1362 1363 1364 l3dsc1
X682 1363 1364 1365 1366 l3dsc1
X683 1365 1366 1367 1368 l3dsc1
X684 1367 1368 1369 1370 l3dsc1
X685 1369 1370 1371 1372 l3dsc1
X686 1371 1372 1373 1374 l3dsc1
X687 1373 1374 1375 1376 l3dsc1
X688 1375 1376 1377 1378 l3dsc1
X689 1377 1378 1379 1380 l3dsc1
X690 1379 1380 1381 1382 l3dsc1
X691 1381 1382 1383 1384 l3dsc1
X692 1383 1384 1385 1386 l3dsc1
X693 1385 1386 1387 1388 l3dsc1
X694 1387 1388 1389 1390 l3dsc1
X695 1389 1390 1391 1392 l3dsc1
X696 1391 1392 1393 1394 l3dsc1
X697 1393 1394 1395 1396 l3dsc1
X698 1395 1396 1397 1398 l3dsc1
X699 1397 1398 1399 1400 l3dsc1
X700 1399 1400 1401 1402 l3dsc1
X701 1401 1402 1403 1404 l3dsc1
X702 1403 1404 1405 1406 l3dsc1
X703 1405 1406 1407 1408 l3dsc1
X704 1407 1408 1409 1410 l3dsc1
X705 1409 1410 1411 1412 l3dsc1
X706 1411 1412 1413 1414 l3dsc1
X707 1413 1414 1415 1416 l3dsc1
X708 1415 1416 1417 1418 l3dsc1
X709 1417 1418 1419 1420 l3dsc1
X710 1419 1420 1421 1422 l3dsc1
X711 1421 1422 1423 1424 l3dsc1
X712 1423 1424 1425 1426 l3dsc1
X713 1425 1426 1427 1428 l3dsc1
X714 1427 1428 1429 1430 l3dsc1
X715 1429 1430 1431 1432 l3dsc1
X716 1431 1432 1433 1434 l3dsc1
X717 1433 1434 1435 1436 l3dsc1
X718 1435 1436 1437 1438 l3dsc1
X719 1437 1438 1439 1440 l3dsc1
X720 1439 1440 1441 1442 l3dsc1
X721 1441 1442 1443 1444 l3dsc1
X722 1443 1444 1445 1446 l3dsc1
X723 1445 1446 1447 1448 l3dsc1
X724 1447 1448 1449 1450 l3dsc1
X725 1449 1450 1451 1452 l3dsc1
X726 1451 1452 1453 1454 l3dsc1
X727 1453 1454 1455 1456 l3dsc1
X728 1455 1456 1457 1458 l3dsc1
X729 1457 1458 1459 1460 l3dsc1
X730 1459 1460 1461 1462 l3dsc1
X731 1461 1462 1463 1464 l3dsc1
X732 1463 1464 1465 1466 l3dsc1
X733 1465 1466 1467 1468 l3dsc1
X734 1467 1468 1469 1470 l3dsc1
X735 1469 1470 1471 1472 l3dsc1
X736 1471 1472 1473 1474 l3dsc1
X737 1473 1474 1475 1476 l3dsc1
X738 1475 1476 1477 1478 l3dsc1
X739 1477 1478 1479 1480 l3dsc1
X740 1479 1480 1481 1482 l3dsc1
X741 1481 1482 1483 1484 l3dsc1
X742 1483 1484 1485 1486 l3dsc1
X743 1485 1486 1487 1488 l3dsc1
X744 1487 1488 1489 1490 l3dsc1
X745 1489 1490 1491 1492 l3dsc1
X746 1491 1492 1493 1494 l3dsc1
X747 1493 1494 1495 1496 l3dsc1
X748 1495 1496 1497 1498 l3dsc1
X749 1497 1498 1499 1500 l3dsc1
X750 1499 1500 1501 1502 l3dsc1
X751 1501 1502 1503 1504 l3dsc1
X752 1503 1504 1505 1506 l3dsc1
X753 1505 1506 1507 1508 l3dsc1
X754 1507 1508 1509 1510 l3dsc1
X755 1509 1510 1511 1512 l3dsc1
X756 1511 1512 1513 1514 l3dsc1
X757 1513 1514 1515 1516 l3dsc1
X758 1515 1516 1517 1518 l3dsc1
X759 1517 1518 1519 1520 l3dsc1
X760 1519 1520 1521 1522 l3dsc1
X761 1521 1522 1523 1524 l3dsc1
X762 1523 1524 1525 1526 l3dsc1
X763 1525 1526 1527 1528 l3dsc1
X764 1527 1528 1529 1530 l3dsc1
X765 1529 1530 1531 1532 l3dsc1
X766 1531 1532 1533 1534 l3dsc1
X767 1533 1534 1535 1536 l3dsc1
X768 1535 1536 1537 1538 l3dsc1
X769 1537 1538 1539 1540 l3dsc1
X770 1539 1540 1541 1542 l3dsc1
X771 1541 1542 1543 1544 l3dsc1
X772 1543 1544 1545 1546 l3dsc1
X773 1545 1546 1547 1548 l3dsc1
X774 1547 1548 1549 1550 l3dsc1
X775 1549 1550 1551 1552 l3dsc1
X776 1551 1552 1553 1554 l3dsc1
X777 1553 1554 1555 1556 l3dsc1
X778 1555 1556 1557 1558 l3dsc1
X779 1557 1558 1559 1560 l3dsc1
X780 1559 1560 1561 1562 l3dsc1
X781 1561 1562 1563 1564 l3dsc1
X782 1563 1564 1565 1566 l3dsc1
X783 1565 1566 1567 1568 l3dsc1
X784 1567 1568 1569 1570 l3dsc1
X785 1569 1570 1571 1572 l3dsc1
X786 1571 1572 1573 1574 l3dsc1
X787 1573 1574 1575 1576 l3dsc1
X788 1575 1576 1577 1578 l3dsc1
X789 1577 1578 1579 1580 l3dsc1
X790 1579 1580 1581 1582 l3dsc1
X791 1581 1582 1583 1584 l3dsc1
X792 1583 1584 1585 1586 l3dsc1
X793 1585 1586 1587 1588 l3dsc1
X794 1587 1588 1589 1590 l3dsc1
X795 1589 1590 1591 1592 l3dsc1
X796 1591 1592 1593 1594 l3dsc1
X797 1593 1594 1595 1596 l3dsc1
X798 1595 1596 1597 1598 l3dsc1
X799 1597 1598 1599 1600 l3dsc1
X800 1599 1600 1601 1602 l3dsc1
X801 1601 1602 1603 1604 l3dsc1
X802 1603 1604 1605 1606 l3dsc1
X803 1605 1606 1607 1608 l3dsc1
X804 1607 1608 1609 1610 l3dsc1
X805 1609 1610 1611 1612 l3dsc1
X806 1611 1612 1613 1614 l3dsc1
X807 1613 1614 1615 1616 l3dsc1
X808 1615 1616 1617 1618 l3dsc1
X809 1617 1618 1619 1620 l3dsc1
X810 1619 1620 1621 1622 l3dsc1
X811 1621 1622 1623 1624 l3dsc1
X812 1623 1624 1625 1626 l3dsc1
X813 1625 1626 1627 1628 l3dsc1
X814 1627 1628 1629 1630 l3dsc1
X815 1629 1630 1631 1632 l3dsc1
X816 1631 1632 1633 1634 l3dsc1
X817 1633 1634 1635 1636 l3dsc1
X818 1635 1636 1637 1638 l3dsc1
X819 1637 1638 1639 1640 l3dsc1
X820 1639 1640 1641 1642 l3dsc1
X821 1641 1642 1643 1644 l3dsc1
X822 1643 1644 1645 1646 l3dsc1
X823 1645 1646 1647 1648 l3dsc1
X824 1647 1648 1649 1650 l3dsc1
X825 1649 1650 1651 1652 l3dsc1
X826 1651 1652 1653 1654 l3dsc1
X827 1653 1654 1655 1656 l3dsc1
X828 1655 1656 1657 1658 l3dsc1
X829 1657 1658 1659 1660 l3dsc1
X830 1659 1660 1661 1662 l3dsc1
X831 1661 1662 1663 1664 l3dsc1
X832 1663 1664 1665 1666 l3dsc1
X833 1665 1666 1667 1668 l3dsc1
X834 1667 1668 1669 1670 l3dsc1
X835 1669 1670 1671 1672 l3dsc1
X836 1671 1672 1673 1674 l3dsc1
X837 1673 1674 1675 1676 l3dsc1
X838 1675 1676 1677 1678 l3dsc1
X839 1677 1678 1679 1680 l3dsc1
X840 1679 1680 1681 1682 l3dsc1
X841 1681 1682 1683 1684 l3dsc1
X842 1683 1684 1685 1686 l3dsc1
X843 1685 1686 1687 1688 l3dsc1
X844 1687 1688 1689 1690 l3dsc1
X845 1689 1690 1691 1692 l3dsc1
X846 1691 1692 1693 1694 l3dsc1
X847 1693 1694 1695 1696 l3dsc1
X848 1695 1696 1697 1698 l3dsc1
X849 1697 1698 1699 1700 l3dsc1
X850 1699 1700 1701 1702 l3dsc1
X851 1701 1702 1703 1704 l3dsc1
X852 1703 1704 1705 1706 l3dsc1
X853 1705 1706 1707 1708 l3dsc1
X854 1707 1708 1709 1710 l3dsc1
X855 1709 1710 1711 1712 l3dsc1
X856 1711 1712 1713 1714 l3dsc1
X857 1713 1714 1715 1716 l3dsc1
X858 1715 1716 1717 1718 l3dsc1
X859 1717 1718 1719 1720 l3dsc1
X860 1719 1720 1721 1722 l3dsc1
X861 1721 1722 1723 1724 l3dsc1
X862 1723 1724 1725 1726 l3dsc1
X863 1725 1726 1727 1728 l3dsc1
X864 1727 1728 1729 1730 l3dsc1
X865 1729 1730 1731 1732 l3dsc1
X866 1731 1732 1733 1734 l3dsc1
X867 1733 1734 1735 1736 l3dsc1
X868 1735 1736 1737 1738 l3dsc1
X869 1737 1738 1739 1740 l3dsc1
X870 1739 1740 1741 1742 l3dsc1
X871 1741 1742 1743 1744 l3dsc1
X872 1743 1744 1745 1746 l3dsc1
X873 1745 1746 1747 1748 l3dsc1
X874 1747 1748 1749 1750 l3dsc1
X875 1749 1750 1751 1752 l3dsc1
X876 1751 1752 1753 1754 l3dsc1
X877 1753 1754 1755 1756 l3dsc1
X878 1755 1756 1757 1758 l3dsc1
X879 1757 1758 1759 1760 l3dsc1
X880 1759 1760 1761 1762 l3dsc1
X881 1761 1762 1763 1764 l3dsc1
X882 1763 1764 1765 1766 l3dsc1
X883 1765 1766 1767 1768 l3dsc1
X884 1767 1768 1769 1770 l3dsc1
X885 1769 1770 1771 1772 l3dsc1
X886 1771 1772 1773 1774 l3dsc1
X887 1773 1774 1775 1776 l3dsc1
X888 1775 1776 1777 1778 l3dsc1
X889 1777 1778 1779 1780 l3dsc1
X890 1779 1780 1781 1782 l3dsc1
X891 1781 1782 1783 1784 l3dsc1
X892 1783 1784 1785 1786 l3dsc1
X893 1785 1786 1787 1788 l3dsc1
X894 1787 1788 1789 1790 l3dsc1
X895 1789 1790 1791 1792 l3dsc1
X896 1791 1792 1793 1794 l3dsc1
X897 1793 1794 1795 1796 l3dsc1
X898 1795 1796 1797 1798 l3dsc1
X899 1797 1798 1799 1800 l3dsc1
X900 1799 1800 1801 1802 l3dsc1
X901 1801 1802 1803 1804 l3dsc1
X902 1803 1804 1805 1806 l3dsc1
X903 1805 1806 1807 1808 l3dsc1
X904 1807 1808 1809 1810 l3dsc1
X905 1809 1810 1811 1812 l3dsc1
X906 1811 1812 1813 1814 l3dsc1
X907 1813 1814 1815 1816 l3dsc1
X908 1815 1816 1817 1818 l3dsc1
X909 1817 1818 1819 1820 l3dsc1
X910 1819 1820 1821 1822 l3dsc1
X911 1821 1822 1823 1824 l3dsc1
X912 1823 1824 1825 1826 l3dsc1
X913 1825 1826 1827 1828 l3dsc1
X914 1827 1828 1829 1830 l3dsc1
X915 1829 1830 1831 1832 l3dsc1
X916 1831 1832 1833 1834 l3dsc1
X917 1833 1834 1835 1836 l3dsc1
X918 1835 1836 1837 1838 l3dsc1
X919 1837 1838 1839 1840 l3dsc1
X920 1839 1840 1841 1842 l3dsc1
X921 1841 1842 1843 1844 l3dsc1
X922 1843 1844 1845 1846 l3dsc1
X923 1845 1846 1847 1848 l3dsc1
X924 1847 1848 1849 1850 l3dsc1
X925 1849 1850 1851 1852 l3dsc1
X926 1851 1852 1853 1854 l3dsc1
X927 1853 1854 1855 1856 l3dsc1
X928 1855 1856 1857 1858 l3dsc1
X929 1857 1858 1859 1860 l3dsc1
X930 1859 1860 1861 1862 l3dsc1
X931 1861 1862 1863 1864 l3dsc1
X932 1863 1864 1865 1866 l3dsc1
X933 1865 1866 1867 1868 l3dsc1
X934 1867 1868 1869 1870 l3dsc1
X935 1869 1870 1871 1872 l3dsc1
X936 1871 1872 1873 1874 l3dsc1
X937 1873 1874 1875 1876 l3dsc1
X938 1875 1876 1877 1878 l3dsc1
X939 1877 1878 1879 1880 l3dsc1
X940 1879 1880 1881 1882 l3dsc1
X941 1881 1882 1883 1884 l3dsc1
X942 1883 1884 1885 1886 l3dsc1
X943 1885 1886 1887 1888 l3dsc1
X944 1887 1888 1889 1890 l3dsc1
X945 1889 1890 1891 1892 l3dsc1
X946 1891 1892 1893 1894 l3dsc1
X947 1893 1894 1895 1896 l3dsc1
X948 1895 1896 1897 1898 l3dsc1
X949 1897 1898 1899 1900 l3dsc1
X950 1899 1900 1901 1902 l3dsc1
X951 1901 1902 1903 1904 l3dsc1
X952 1903 1904 1905 1906 l3dsc1
X953 1905 1906 1907 1908 l3dsc1
X954 1907 1908 1909 1910 l3dsc1
X955 1909 1910 1911 1912 l3dsc1
X956 1911 1912 1913 1914 l3dsc1
X957 1913 1914 1915 1916 l3dsc1
X958 1915 1916 1917 1918 l3dsc1
X959 1917 1918 1919 1920 l3dsc1
X960 1919 1920 1921 1922 l3dsc1
X961 1921 1922 1923 1924 l3dsc1
X962 1923 1924 1925 1926 l3dsc1
X963 1925 1926 1927 1928 l3dsc1
X964 1927 1928 1929 1930 l3dsc1
X965 1929 1930 1931 1932 l3dsc1
X966 1931 1932 1933 1934 l3dsc1
X967 1933 1934 1935 1936 l3dsc1
X968 1935 1936 1937 1938 l3dsc1
X969 1937 1938 1939 1940 l3dsc1
X970 1939 1940 1941 1942 l3dsc1
X971 1941 1942 1943 1944 l3dsc1
X972 1943 1944 1945 1946 l3dsc1
X973 1945 1946 1947 1948 l3dsc1
X974 1947 1948 1949 1950 l3dsc1
X975 1949 1950 1951 1952 l3dsc1
X976 1951 1952 1953 1954 l3dsc1
X977 1953 1954 1955 1956 l3dsc1
X978 1955 1956 1957 1958 l3dsc1
X979 1957 1958 1959 1960 l3dsc1
X980 1959 1960 1961 1962 l3dsc1
X981 1961 1962 1963 1964 l3dsc1
X982 1963 1964 1965 1966 l3dsc1
X983 1965 1966 1967 1968 l3dsc1
X984 1967 1968 1969 1970 l3dsc1
X985 1969 1970 1971 1972 l3dsc1
X986 1971 1972 1973 1974 l3dsc1
X987 1973 1974 1975 1976 l3dsc1
X988 1975 1976 1977 1978 l3dsc1
X989 1977 1978 1979 1980 l3dsc1
X990 1979 1980 1981 1982 l3dsc1
X991 1981 1982 1983 1984 l3dsc1
X992 1983 1984 1985 1986 l3dsc1
X993 1985 1986 1987 1988 l3dsc1
X994 1987 1988 1989 1990 l3dsc1
X995 1989 1990 1991 1992 l3dsc1
X996 1991 1992 1993 1994 l3dsc1
X997 1993 1994 1995 1996 l3dsc1
X998 1995 1996 1997 1998 l3dsc1
X999 1997 1998 1999 2000 l3dsc1
X1000 1999 2000 2001 2002 l3dsc1
.ends l3dsub1

* Isolated High Speed Circuit
*
* High Speed source
* VFAST 8 0 DC 0 SIN(5v 10v 400MEGhz 1ms) NO CHANCE, Too expensive
*VFAST 8 0 DC 0 SIN(5v 10v 400Khz 1ms 0)
*VFAST 8 0 DC 0 SIN(5v 10v 4Khz 1ms 0)
*RFSS 8 9 0.5

* High Speed RLC load
*LFS  8 9 3n
*RFSP 9 0 1K
*CFS  9 0 680p

.tran 100us 300ms 

*COMP v(1) reltol=0.02 abstol=2e-6
*COMP v(11) reltol=0.02 abstol=1e-6
*COMP v(22) reltol=0.02 abstol=1e-6
*COMP v(33) reltol=0.02 abstol=1e-6
*COMP v(44) reltol=0.02 abstol=1e-6
.print  tran v(1) v(11) v(22) v(33) v(44)

.END
