Bug 668 output format test. (format=tecplot)

R1 1 0 10
V1 1 0 sin (0 10 10MEG 0 0)
R2 2 0 10
V2 2 0 sin (0 10 5MEG 0 0)
R3 3 0 10
V3 3 0 sin (0 10 10MEG 0 0)
R4 4 0 10
V4 4 0 sin (0 10 5MEG 0 0)
R5 5 0 10
V5 5 0 sin (0 10 10MEG 0 0)
R6 6 0 10
V6 6 0 sin (0 10 5MEG 0 0)
R7 7 0 10
V7 7 0 sin (0 10 10MEG 0 0)
R8 8 0 10
V8 8 0 sin (0 10 5MEG 0 0)
R9 9 0 10
V9 9 0 sin (0 10 10MEG 0 0)

.print tran format=tecplot v(1) v(2) v(3) v(4) v(5) v(6) v(7) v(8) v(9) I(v1) I(v2) I(v3) I(v4) I(v5) I(v6) I(v7) I(v8) I(v9) 

.tran 1ns 1us

.end
