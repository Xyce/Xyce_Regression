* test of coupled inductor parameters on the .PRINT line, when inside subcircuit
V1 1 0 SIN(0 1 1KHz)
R1 1 0 2
R2 2 0 2

X1 1 2 foo

.subckt foo a b
* mutual inductor definition (nonlnear level=2)
L1 a 0 100
L2 b 0 100
K1 L1 L2 1.00 nlcore
.ends

.model nlcore core level=2 c=0.001

.TRAN 0 1ms 
.PRINT TRAN V(1) V(2) X1:L1:L {X1:L1:L} {2.0*X1:L1:L} {X1:L1:L**2} {(X1:L1:L)*R1:R}
.END 

