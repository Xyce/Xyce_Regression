*******************************************************************************
* This netlist is equivalent to Step 3 for the MaxTest.cir netlist.
* It has VS1:VA=2 and VS3:V0=-0.5
*
*******************************************************************************
*
* a few sources of different types
VS1  1  0  SIN(0 2 1KHz 0 0)
VP   2  0  PULSE( 0 100 0.2ms 0.2ms 0.2ms 1ms 2ms )
VS3  3  0  SIN(-0.5 1.0 1KHZ 0 500)
VS4  4  0  SIN(0.5 -1.0 1KHZ 0 500)

R1  1  0  100
R2  2  0  100
R3  3  0  100
R4  4  0  100

.TRAN 0  3ms
.PRINT TRAN FORMAT=NOINDEX V(1) V(2) V(3) V(4)

* plain test
.measure tran maxSine max V(1)
.measure tran max2 MAX v(2)

* add TO-FROM modifiers
.measure tran maxHalfSine max V(1) from=0 to=0.5e-3

* mix in TDs before and after FROM value.
.measure tran sine60 max V(1) FROM=0.5e-3 TO=0.75e-3 TD=0.6e-3
.measure tran sine70 max V(1) FROM=0.7e-3 TO=0.75e-3 TD=0.6e-3

* these tests should return -1 and -100
.measure tran returnNegOne max V(1) FROM=0.2e-3 TO=0.25e-3 TD=0.5e-3
.measure tran returnNeg100 max V(1) FROM=0.2e-3 TO=0.25e-3 TD=0.5e-3 default_val=-100

* add tests for rise/fall/cross.  VS2 and VS3 have a DC offset
* and are damped sinusoids
.measure tran maxv3fall2 max v(3) fall=2
.measure tran maxv4rise1 max v(4) rise=1
.measure tran maxv3cross3 max v(3) cross=3

* test LAST for rise/fall/cross
.measure tran maxv3falllast max v(3) fall=last
.measure tran maxv4riselast max v(4) rise=last
.measure tran maxv3crosslast max v(3) cross=last
.measure tran maxv4crosslast max v(4) cross=last

* test RFC_LEVEL keyword
.measure tran maxv1Rise1RFClevel50 max V(1) RFC_LEVEL=0.5 RISE=1
.measure tran maxv1Fall1RFClevel50 max V(1) RFC_LEVEL=0.5 FALL=1
.measure tran maxv1Cross1RFClevel50 max V(1) RFC_LEVEL=0.5 CROSS=1 

*test Failed measures for rise/fall/cross
.measure tran maxv3fallfail max v(3) fall=10
.measure tran maxv4risefail max v(4) rise=10
.measure tran maxv3crossfail max v(3) cross=10

.END

