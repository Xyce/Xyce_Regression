RAW File Output test for the N-Channel MESFET.
************************************************************
* This test has two purposes:
*   1) Verify that the variable type (e.g., "voltage") and 
*      variable name is correct for the MESFET. This test
*      just has a non-zero source and drain conductivity.  
*      So, both drainprime and sourceprime properly show 
*      up as an internal voltage nodes.  
*
*   2) Verify that the data is actually correct for all of
*      the time-steps in the .RAW file output 
*
* The "gold" .RAW file output was generated by manually
* comparing that "gold" file with a .PRN file.  It was 
* generated for a limited set of fixed time-steps, so that
* a file comparison could be used to verify the test output's
* .RAW file against that "gold" .RAW file.
*
************************************************************
*
VDS 2 0 2V
VGS 3 0 pulse (-1 1 1ns 1ns 1ns 1us 2us)
VSS 4 0 0
Z1 2 3 4 MESMOD AREA=1.4
.MODEL MESMOD NMF
+ LEVEL=1 BETA=1.4E-3
+ RD=46 RS=46 VTO=-1.3 LAMBDA=0.03 ALPHA=3 CGS=1uf CGD=1uf

.options timeint method=gear
.options nonlin-tran rhstol=1.0e-7
.options output initial_interval=0.5us
.tran 1ns 10us

* .PRINT statement is not actually used for .RAW output.
* It was included in the netslit so that the "gold" .RAW 
* file output could manually verified against a .PRN file
* during test development
.print tran v(2) v(3) v(4) I(VDS) I(VGS) I(VSS)
+ N(z1_drainprime) N(z1_sourceprime)
 
.end

