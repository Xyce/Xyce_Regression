* Test of duplicate measure names in Xyce.  The first
* M1 and M2 definitions should be ignored and produce
* warning messages.  The EQN measures should produce
* the values given by the second M1 and M2 definitions.
*
* See SON Bug 1300 for more details.
******************************************************
.TRAN 0 1
.PRINT TRAN V(1) V(2)

V1 1 0 PWL 0 0 0.5 1 1 0
R1 1 0 1

V2 2 0 PWL 0 1 0.5 0 1 1
R2 2 0 1

.MEASURE TRAN M1 MIN V(1)
.MEASURE TRAN M1 MAX V(1)
.MEASURE TRAN EQNM1 EQN M1

.MEASURE TRAN EQNM2 EQN M2
.MEASURE TRAN M2 MAX V(2)
.MEASURE TRAN M2 MIN V(2)

.END
