Test of ABM power function
**********************************************************
* This circuit tests the that the minus sign in the 
* argument is handled correctly in the floating 
* point exponent (not integer) case.
* Passing this test certifies bug #8 (joseki bugzilla).
**********************************************************
VS  1  0  -2.5
R1  1  0  1.0
B5  5  0  V = { (V(1))**2.1 }
R5  5  0  1
B6  6  0  V = { (-V(1))**3.1 }
R6  6  0  1
*
.DC VS -2.5 2.5 0.2
.PRINT DC V(1) V(5) V(6)
.END
