* Test NOISE mode support for the NOISE_CONT version of
* FIND-AT, FIND-WHEN and WHEN measures.
*
* See SON Bugs 1274 and 1313 for more details.
********************************************************************

* Used to adjust reference frequency from 1Hz to 1KHz
.PARAM scaleFactor=1e3

* RESISTOR DIVIDER
V1  1 0 DC 5.0 AC  1.0
R1  1 2 100K
R2  2 0 100K
*
* AMP AND LP FILTER
EAMP   3 0 2 0 2
* 7th order Chebychev LPF with 2dB of passband ripple.
* This is not a realistic passbad ripple level, but is
* useful for this test.
RS 3 b 1
C1 b 0 {2.865/scaleFactor}
L2 b c {0.912/scaleFactor}
C3 c 0 {3.8774/scaleFactor}
L4 c d {0.9537/scaleFactor}
C5 d 0 {3.8774/scaleFactor}
L6 d e {0.912/scaleFactor}
C7 e 0 {2.8650/scaleFactor}
RL e 0 1.0

.NOISE  V(E)  V1  DEC  20 1 1000
.STEP RL 1 1.5 0.5
.PRINT NOISE VM(3) vm(b) vm(c) vm(d) vm(e)

* The non-continuous version should return the first crossing.
* The continuous version should return all crossings.
.MEASURE NOISE whenCrossTest1 WHEN vm(e)=0.45
.MEASURE NOISE_CONT whenCrossContTest1 WHEN vm(e)=0.45

* Non-continuous version should return first crossing.
* Continuous version should return all crossings, starting
* with the first one.
.MEASURE NOISE whenCrossTest2 WHEN VM(e)=0.45 CROSS=1
.MEASURE NOISE_CONT whenCrossContTest2 WHEN VM(e)=0.45 CROSS=1

* Non-continuous version should return second crossing.
* Continuous version should return all crossings, starting
* with the second one.
.MEASURE NOISE whenCrossTest3 WHEN VM(e)=0.45 CROSS=2
.MEASURE NOISE_CONT whenCrossContTest3 WHEN VM(e)=0.45 CROSS=2

* These should both return the last crossing
.MEASURE NOISE whenCrossTest4 WHEN VM(e)=0.45 CROSS=LAST
.MEASURE NOISE_CONT whenCrossContTest4 WHEN VM(e)=0.45 CROSS=LAST

* FIND-AT measures
* These should give the same answer
.MEASURE NOISE atTest FIND VM(e) AT=20
.MEASURE NOISE_CONT atContTest FIND VM(e) AT=20

******************************************************
* Repeat WHEN tests as FIND-WHEN measures
.MEASURE NOISE findCrossTest1 FIND VM(d) WHEN VM(e)=0.45
.MEASURE NOISE_CONT findCrossContTest1 FIND VM(d) WHEN VM(e)=0.45

.MEASURE NOISE findCrossTest2 FIND VM(d) WHEN VM(e)=0.45 CROSS=1
.MEASURE NOISE_CONT findCrossContTest2 FIND VM(d) WHEN VM(e)=0.45 CROSS=1

.MEASURE NOISE findCrossTest3 FIND VM(d) WHEN VM(e)=0.45 CROSS=2
.MEASURE NOISE_CONT findCrossContTest3 FIND VM(d) WHEN VM(e)=0.45 CROSS=2

.MEASURE NOISE findCrossTest4 FIND VM(d) WHEN VM(e)=0.45 CROSS=LAST
.MEASURE NOISE_CONT findCrossContTest4 FIND VM(d) WHEN VM(e)=0.45 CROSS=LAST

*****************************************************
* test RISE and FAll qualifiers for WHEN and FIND-WHEN
.MEASURE NOISE_CONT whenRiseContTest1 WHEN VM(e)=0.45 RISE=1
.MEASURE NOISE_CONT whenRiseContTest2 WHEN VM(e)=0.45 RISE=2
.MEASURE NOISE_CONT whenRiseContTest3 WHEN VM(e)=0.45 RISE=LAST

.MEASURE NOISE_CONT whenFallContTest1 WHEN VM(e)=0.45 FALL=1
.MEASURE NOISE_CONT whenFallContTest2 WHEN VM(e)=0.45 FALL=2
.MEASURE NOISE_CONT whenFallContTest3 WHEN VM(e)=0.45 FALL=LAST

.MEASURE NOISE_CONT findRiseContTest1 FIND VM(b) WHEN VM(e)=0.45 RISE=1
.MEASURE NOISE_CONT findRiseContTest2 FIND VM(b) WHEN VM(e)=0.45 RISE=2
.MEASURE NOISE_CONT findRiseContTest3 FIND VM(b) WHEN VM(e)=0.45 RISE=LAST

.MEASURE NOISE_CONT findFallContTest1 FIND VM(b) WHEN VM(e)=0.45 FALL=1
.MEASURE NOISE_CONT findFallContTest2 FIND VM(b) WHEN VM(e)=0.45 FALL=2
.MEASURE NOISE_CONT findFallContTest3 FIND VM(b) WHEN VM(e)=0.45 FALL=LAST

*********************************************************
* Test negative values
.MEASURE NOISE_CONT whenCrossContNeg1 WHEN VM(e)=0.45 CROSS=-1
.MEASURE NOISE_CONT whenCrossContNeg2 WHEN VM(e)=0.45 CROSS=-2
.MEASURE NOISE_CONT whenCrossContNeg3 WHEN VM(e)=0.45 CROSS=-3
.MEASURE NOISE_CONT whenCrossContNeg6 WHEN VM(e)=0.45 CROSS=-6

.MEASURE NOISE_CONT whenRiseContNeg1 WHEN VM(e)=0.45 RISE=-1
.MEASURE NOISE_CONT whenRiseContNeg2 WHEN VM(e)=0.45 RISE=-2
.MEASURE NOISE_CONT whenRiseContNeg3 WHEN VM(e)=0.45 RISE=-3

.MEASURE NOISE_CONT whenFallContNeg1 WHEN VM(e)=0.45 FALL=-1
.MEASURE NOISE_CONT whenFallContNeg2 WHEN VM(e)=0.45 FALL=-2
.MEASURE NOISE_CONT whenFallContNeg3 WHEN VM(e)=0.45 FALL=-4

*************************************************
* test failed measures
.MEASURE NOISE_CONT whenCrossContFail1 WHEN VM(e)=1
.MEASURE NOISE_CONT atContFail FIND VM(e) at=2000
.MEASURE NOISE_CONT whenCrossContFail2 WHEN VM(e)=0.45 CROSS=6
.MEASURE NOISE_CONT whenRiseContFail WHEN VM(e)=0.45 RISE=4
.MEASURE NOISE_CONT whenFallContFail WHEN VM(e)=0.45 FALL=4

* Signifies end of test. .sh file looks for a measure named lastMeasure.
* This is needed for compatibility for testing with a verbose build, which
* is often used by the Xyce developers.
.measure NOISE lastMeasure max VM(e)

.END

