power test for BJT 
*
*
vie1 0 Emitter1 0
vic1 0 Collector1 5
vib1 0 Base1 pulse(0 1 1ns 1ns 1ns 1us) 
q1 Collector1 Base1 Emitter1 0 qjunk1 

vie2 0 Emitter2 0
vic2 0 Collector2 5
vib2 0 Base2 pulse(0 1 1ns 1ns 1ns 1us) 
q2 Collector2 Base2 Emitter2 0 qjunk2 

.model qjunk1 npn
+ level=12
+ RCX=10 RCI=10 RBX=1 RBI=10 RE=1 RBP=10 RS=10
+ IBEN=1.0e-13 RTH=100

.model qjunk2 pnp
+ level=12
+ RCX=10 RCI=10 RBX=1 RBI=10 RE=1 RBP=10 RS=10
+ IBEN=1.0e-13 RTH=100

.options timeint method=gear
.options nonlin-tran rhstol=1.0e-8
.tran 1ns 20us

.PRINT TRAN  v(Collector1) V(Base1) v(Emitter1) i(vic1) i(vib1)
+ {abs(i(vic1)*(v(Collector1)-v(Emitter1)))+abs(i(vib1)*(V(Base1)-v(Emitter1)))} p(q1) w(q1)
+ v(Collector2) v(Base2) v(Emitter2) i(vic2) i(vib2)
+ {abs(i(vic2)*(v(Collector2)-v(Emitter2)))+abs(i(vib2)*(v(Base2)-v(Emitter2)))} p(q2) w(q2)

.END
