**********************************************************************
* Purpose of circuit is to test:
*
*   1) whether xdm query mode can "ignore" .MEASURE statements.  
*    
*   2) the 'D' option for query mode (-q D)
* 
* This circuit was used as a test-example during xdm development,
* and is a likely example-case for a Query Mode section of the eventual 
* xdm Users Guide.
*
* Note: the -q D output for this netlist ends up in the file
* diodeClipperMeasure.cir.xdm.D.gs.out.
***********************************************************************

* Voltage Sources
VCC 1 0 5V
VIN 3 0 SIN(0V 10V 1kHz)
* Analysis Command
.TRAN 2ns 2ms
* Output and .MEASURE statements
.PRINT TRAN V(3) V(2) V(4)
.MEASURE TRAN MAXV3 MAX V(3) FROM=0 TO=1e-3
.MEASURE TRAN MAXV4 MAX V(4) FROM=0 TO=1e-3
.MEASURE TRAN MAXV3minusV4 MAX {V(3) - V(4)} FROM=0 TO=1e-3
.MEASURE TRAN MINV3 MIN V(3) FROM=0 TO=1e-3
.MEASURE TRAN MINV4 MIN V(4) FROM=0 TO=1e-3
.MEASURE TRAN MAXABSV3minusV4 MAX {abs(V(3) - V(4))} FROM=0 TO=1e-3

* Diodes
D1 2 1 D1N3940
D2 0 2 D1N3940
* Resistors
R1 2 3 1K
R2 1 2 3.3K
R3 2 0 3.3K
R4 4 0 5.6K
* Capacitor
C1 2 4 0.47u
*
* GENERIC FUNCTIONAL EQUIVALENT = 1N3940
* TYPE: DIODE
* SUBTYPE: RECTIFIER
.MODEL D1N3940 D(
+ IS = 4E-10
+ RS = .105
+ N = 1.48
+ TT = 8E-7
+ CJO = 1.95E-11
+ VJ = .4
+ M = .38
+ EG = 1.36
+ XTI = -8
+ KF = 0
+ AF = 1
+ FC = .9
+ BV = 600
+ IBV = 1E-4)
*
.END


