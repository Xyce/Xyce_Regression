* Sensitivity of collector current to amplifier component
* This circuit was found  on page 298 of the book,
* "PSPICE and MATLAB for Electronics: An Integrated Approach" by John Okyere Attia.
*
* The relevant pages are excerpted in google books, and includes a printout of the
* PSPICE output.
*
.global_param VCCvalue=10V

VCC 4 0 DC {VCCvalue}
RB1 4 1 40k
RB2 1 0 10k
RE 2 0 1K
RC 5 3 6K
VM 4 5 DC 0; monitor collector current
Q1 3 1 2 0 0 mymodel

.DC VCCvalue 1 10 0.4

.print dc v(4) I(VM)
.print sens v(4)


.SENS param=
+ mymodel:ibes,
+ mymodel:rci0,
+ mymodel:tnom
+objfunc={I(VM)}

.options SENSITIVITY direct=1 adjoint=0  forcedevicefd=1  debuglevel=2

.model mymodel npn level=230
+ mcf= 1 
+ rbi0= 4.444 
+ rbx= 2.568 
+ fgeo= 0.7409 
+ re= 1.511 
+ rcx= 2.483 
+ itss= 0 
+ msf= 1 
+ iscs= 0 
+ msc= 1 
+ cjci0= 3.58e-015 
+ vdci= 0.8201 
+ zci= 0.2857 
+ vptci= 1.79 
+ cjcx0= 6.299e-015 
+ vdcx= 0.8201 
+ zcx= 0.2863 
+ vptcx= 1.977 
+ cjs0= 2.6e-014 
+ vds= 0.9997 
+ zs= 0.4295 
+ vpts= 100 
+ t0= 2.089e-013 
+ dt0h= 8e-014 
+ tbvl= 8.25e-014 
+ tef0= 3.271e-013 
+ thcs= 5.001e-012 
+ ahc= 0.05 
+ rci0= 9.523 
+ vlim= 0.6999 
+ vces= 0.01 
+ vpt= 2 
+ tr= 0 
+ cbepar= 2.609e-014 
+ cbcpar= 1.64512e-014 
+ alqf= 0.166667 
+ alit= 0.333333 
+ flnqs= 0 
+ kf= 0 
+ af= 2 
+ vgb= 0.91 
+ alt0= 0.004 
+ kt0= 6.588e-005 
+ zetaci= 0.58 
+ alvs= 0.001 
+ alces= -0.2286 
+ zetarbi= 0.3002 
+ zetarbx= 0.06011 
+ zetarcx= -0.02768 
+ zetare= -0.9605 
+ vge= 1.17 
+ vgc= 1.17 
+ vgs= 1.17 
+ f1vg= -0.000102377 
+ f2vg= 0.00043215 
+ zetact= 5 
+ zetabet= 4.892 
+ flsh= 1 
+ rth= 1113.4 
+ cth= 6.841e-012 
+ zetarth= 0 
+ tnom= 26.85 
+ zetavgbe= 0.7 
