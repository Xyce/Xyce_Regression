Polynomial Source Netlist for a single input, fourth order polynomial
***********************************************************************
*		B = V(3) = 3 + 2*V(2) + V(2)^2 + 3*V(2)^3 + 4*V(2)^4
***********************************************************************
.param C0=3.0
.param C1=2.0
.param C2=1.0
.param C3=3.0
.param C4=4.0

* POLY function
.func polyVersion(x1) {POLY(1) x1 C0 C1 C2 C3 C4}

* POLY version:
VINPUT 1 0 1.0
B 3 0 V ={3.0*(polyVersion(V(2)))}
R1 1 2 1K
R2 2 0 1K
R3 3 4 2K
R4 4 0 2K

* expression style function,  implementing the same polynomial:
.func exprVersion(x1) { (C0 + C1*x1+ C2*pow(x1,2.0) + C3*pow(x1,3.0) + C4*pow(x1,4.0)  ) } 

Ba 3a 0 V ={3.0*(exprVersion(V(2a)))}
R1a 1 2a 1K
R2a 2a 0 1K
R3a 3a 4a 2K
R4a 4a 0 2K

.DC VINPUT -4 4 1
.PRINT DC V(1) {100.0-abs(V(3)-V(3a))}

.END
