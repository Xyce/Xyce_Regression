*Sample netlist for BSIM-MG 
*Drain current symmetry for nmos

*.options nonlin abstol=1e-6 reltol=1e-6 
.options device temp=25 

.include "modelcard.nmos_xyce"

* --- Voltage Sources ---
vdrain drain 0 dc 0
esource source 0 drain 0 -1
vgate gate  0 dc 1.0
vbulk bulk 0 dc 0.0


* --- single Transistor ---
Vdamm drain drainsingle 0
Vgamm gate gatesingle 0
Vsamm source sourcesingle 0
Vbamm bulk bulksingle 0
M1 drainsingle gatesingle sourcesingle bulksingle nmos1 TFIN=15n L=30n NFIN=10 NRS=1 NRD=1

* --- multiple Transistor ---
Vdamm2 drain drainmultiple 0
Vgamm2 gate gatemultiple 0
Vsamm2 source sourcemultiple 0
Vbamm2 bulk bulkmultiple 0
M2 drainmultiple gatemultiple sourcemultiple bulkmultiple nmos1 M=10 TFIN=15n L=30n NFIN=10 NRS=1 NRD=1

* --- DC Analysis ---
.dc vdrain -0.1 0.1 0.001 vgate 0.0 1.0 0.2
.print dc v(drain) v(gate) {-I(Vdamm)} {-I(Vgamm)} {-I(Vsamm)} {-I(Vbamm)} {-I(Vdamm2)} {-I(Vgamm2)} {-I(Vsamm2)} {-I(Vbamm2)}

.end
