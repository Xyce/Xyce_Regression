Diode clipper circuit with transient analysis statement
* This is from Figure 3.5 of the Users Guide
*
* Voltage Sources
VCC 1 0 10V
VIN 3 0 SIN(0V 10V 1kHz) AC 1
* Analysis Command
.noise V(4) VIN DEC 5 100 100MEG
* Output
.PRINT noise {log(inoise)} {log(onoise)} {log(DNI(D1))} {log(DNO(D2))} {log(DNI(D2))} {log(DNO(D2))} {log(DNO(D1,flicker_a_aik_flicker))} {log(DNO(D1,white_aik_k_thermal))} {log(DNO(D1,white_a_aik_shot))}
* Diodes
D1 2 1 D1mod
D2 0 2 D1mod
* Resistors
R1 2 3 1K
R2 1 2 3.3K
R3 2 0 3.3K
R4 4 0 5.6K
* Capacitor
C1 2 4 0.47u
.MODEL D1mod D(level=2002)

.END
