*********************************************************
* This netlist tests SON Bug 1033, using the level 1
* resistor device.  It tests that bug for both instance
* and model parameters that depend on TEMP and VT.  This 
* test is also related to SON Bugs 606 and 654.  
*******************************************************

V1 1 0 1
R1 1 0 {TEMP}

V2 2 0 1
R2 2 0 {Vt}

V3 3 0 1
R3 3 0 RMOD1 1

V4 4 0 1
R4 4 0 RMOD2 1

.MODEL RMOD1 R R={TEMP}
.MODEL RMOD2 R R={VT}

.DC V1 1 1 1
.STEP TEMP 27 37 10
.PRINT DC V(1) TEMP {1/TEMP} VT {1/VT}
+ R1:R I(R1) R2:R I(R2) 
+ R3:R I(R3) R4:R I(R4)
.END

