AC test of print output format with .OP and .STEP
*
* Trivial resistor circuit, just do a AC sweep and watch the output
*

R1 1 0 10
V1 1 0 DC 0V

.print AC v(1) I(v1)
.ac dec 10 100Hz 1000MegHz
.step temp -10 10 10
.op

.end
