*A Simple MOSFET Gain Stage. AC Analysis.

*M1 3 2 0 0 nmos w=4u l=1u 
*Rsource 1 2 100k
Rload 3 vdd 25k

Vdd1 vdd 0 5 
*Vin 1 0 1.44 ac .1
Iin 1 0 1.44e-5 ac 0.1e-5 sin(0 1 1e+5 0 0) 
Rsource 1 0  100k
M1 3 1 0 0 nmos w=4u l=1u

*.options noacct
.ac dec 10 100 1000Meg 
.print ac v(3)

.model nmos nmos level=9

.end

