********************************************************
* Test error messsage when .DATA line has an freq
* entry that is not > 0
*
* See SON Bug 1042 for more details.
********************************************************

.global_param mag=1
.global_param phase=0.1

v1  1 0 dc 5.0 ac  {mag} {phase}
r1  1 2 100k
r2  2 0 100k
*
* amp and lp filter
eamp  3 0 2 0 1
rlp1  3 4 100
clp1  4 0 1.59nf
*
.noise  v(4)  v1  data=table

.print noise V(4) {log(onoise)} {log(inoise)}
+ {log(dno(rlp1))} {log(dno(r2))} {log(dno(r1))}
+ {log(dni(rlp1))} {log(dni(r2))} {log(dni(r1))}

.DATA table
+  mag  phase   freq
+  1.0   0.1   1.0e0
+  2.0   0.2   1.0e1
+  3.0   0.3   1.0e2
+  4.0   0.4   1.0e3
+  5.0   0.5   1.0e4
+  6.0   0.6   1.0e5
+  1.0   0.1   0.0e0
.enddata

.end
