* Reference circuit for bug4_issue694.  This circuit is equivalent, but the sensitivities are computed via a crude finite difference.

.model nfet_model nmos level = 54 

.options device temp=25 

* --- Voltage Sources ---
vdd   supply  0 dc 1.8
VIN1 vi 0 PWL(0S 0V  100ps 0V 300ps 1.8V )

* using option scale:
.option scale=1.0e-6
.param Wparam=650000u
.param Lparam=150000u

* Not using option scale:
*.param Wparam=0.65u
*.param Lparam=0.15u

m_nfet 0 vi vo 0 nfet_model l = {Lparam} w = {Wparam}

* --- Transient Analysis ---
.tran 2ps 1ns

.print tran v(*)


.end
