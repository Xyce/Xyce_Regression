Inverter example circuit
*
* This example is used only to look for correct warnings about unsupported
* versions or parameters.

* This circuit does NOT use model binning, intentionally.  
.model nch.1 nmos ( version=4.5 level=54 lmin=0.1u lmax=20u wmin=0.1u wmax=10u   TEMPEOT=300.15)
.model nch.2 nmos ( version=4.65 level=54 lmin=0.1u lmax=20u wmin=10u  wmax=100u  TEMPEOT=300.15)
.model pch.1 pmos ( version=4.7 level=54 lmin=0.1u lmax=20u wmin=0.1u wmax=10u   TEMPEOT=300.15)
.model pch.2 pmos ( version=4.8 level=54 lmin=0.1u lmax=20u wmin=10u  wmax=100u  TEMPEOT=300.15)
*
* parameters
.param vp     = 1.0v

.param drise  = 400ps
.param dfall  = 100ps
.param trise  = 100ps
.param tfall  = 100ps
.param period = 1ns
.param skew_meas = 'vp/2'
*
* parameterized subckt
.subckt inv in out vdd gnd 
mp out in vdd vdd pch.2 w=60 l=0.10
mn out in gnd gnd nch.2 w=20 l=0.10
.ends

.subckt inv2 in out vdd gnd 
mp out in vdd vdd pch.1 w=60 l=0.10
mn out in gnd gnd nch.1 w=20 l=0.10
.ends

v0 vdd 0 'vp'

* vsrc with repeat
v1 in 0 pwl
+ 0ns                       'vp'
+ 'dfall-0.8*tfall'         'vp'
+ 'dfall-0.4*tfall'         '0.9*vp'
+ 'dfall+0.4*tfall'         '0.1*vp'
+ 'dfall+0.8*tfall'         0v
+ 'drise-0.8*trise'         0v
+ 'drise-0.4*trise'         '0.1*vp'
+ 'drise+0.4*trise'         '0.9*vp'
+ 'drise+0.8*trise'         'vp'
+ 'period+dfall-0.8*tfall'  'vp'
+ r='dfall-0.8*tfall'

x1 in out vdd 0 inv pw=60 nw=20
c1 out 0 220fF

x2 in out2 vdd 0 inv2 pw=60 nw=20
c2 out2 0 220fF

.tran 1ps 4ns
.print tran v(vdd) v(in) v(out) v(out2)

.options parser scale=1.0e-6

.end
