Diode Circuit Netlist
VIN 1 0 1
VMON 1 2 0
D1 2 0 DMOD PJ=0.5
.MODEL DMOD D (IS=1e-15 CJO=1e-15 RS=1 JSW=1e-15 CJSW=1e-15 nbv=0.3 bv=15)
.DC VIN -25 1 .5

.PRINT DC V(1) I(VMON) N(D1:Cd)
*
.END
