Simple RC circuit, baseline version
* 
* Eric Keiter, SNL
*
Isrc 1 0 AC 1 0 
R1 1 0 1e3
C1 1 0 2e-6

.print ac v(1)
.AC DEC 1 1 1e8

.END
