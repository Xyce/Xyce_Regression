* Test AC mode support for AVG measures.
* To be conservative, there are subtests for each
* valid operator (V, VR, VI, VP, VM and VDB) for
* each measure type. Expressions are also tested.
*
* See SON Bug 1267 for more details
*****************************************************

* Trivial high-pass filter (V-C-R) circuit
R1 b 0 2
C1 a b 1u
V1 a 0 DC 0V AC 1

.print AC vr(b) vi(b) vm(b) vp(b) vdb(b)
.ac dec 5 100Hz 1e6
.STEP R1 0.5 2 1.5

* MAX
.MEASURE AC avgvb avg v(b)
.MEASURE AC avgvmb avg vm(b)
.MEASURE AC avgvrb avg vr(b)
.MEASURE AC avgvib avg vi(b)
.MEASURE AC avgvpb avg vp(b)
.MEASURE AC avgvdbb avg vdb(b)

* Use expression
.MEASURE AC avgvrbExp avg {1+vr(b)}

* add FROM-TO
*.MEASURE AC avgvmbFromTo avg vm(b) FROM=1e3 TO=1e5

* Tests should return -1 or -100, since the FROM-T0 window
* has various problems.
.measure ac avgReturnNegOne avg v(b) FROM=1e7 TO=1e8
.measure ac avgReturnNeg100 avg vr(b) FROM=1e6 TO=1e2 DEFAULT_VAL=-100

* Signifies end of test. .sh file looks for a measure named lastMeasure.
* This is needed for compatibility for testing with a verbose build, which
* is often used by the Xyce developers.
.measure ac lastMeasure avg vm(b)

.end
