First test of .func/.param resolution, per bug 224
*
* This test doesn't use functions in subcircuits, they are defined outside

.param coef1=1
.param coef2=2
.Func F1(X) {coef1*X*X}
.Func F2(X) {coef2*X*X}
.Param resistance1=10k
.param resistance2=5k

.DC V1 0 5 .1
.print DC v(1) v(2) v(3) v(4) v(5)

*Stupid little circuit to generate a voltage  feed into B source
V1 1 0 5V
R0 1 0 1K
X1 2 3 1 FooCkt
X2 4 5 1 FooCkt2

.subckt FooCkt A B CTL
* Voltage divider, fed by B source
B1 A 0 V={F1(V(CTL))}
R1 A B {resistance1}
R2 B 0 {resistance2}
.ends

.subckt FooCkt2 A B CTL
* Voltage divider, fed by B source
B1 A 0 V={F2(V(CTL))}
R1 A B {resistance1}
R2 B 0 {resistance2}
.ends

.end
