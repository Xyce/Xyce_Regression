*A Simple MOSFET Gain Stage. AC Analysis.

M1 3 2 0 0 nmos w=4u l=1u 
*pd=5e-6 ps=5e-6 
Rsource 1 2 100k
Rload 3 vdd 25k

Vdd1 vdd 0 5 
Vin 1 0 1.44 ac .1 sin(0 1 1e+5 0 0) 

*.options noacct
.op 
.ac dec 10 100 1000Meg 
.print ac v(3)

.include nmos_3_2.mod  
*.model nmos nmos level=10 cgdo=0  cgso=0 k2=-0.0186 k1=0.53 xj=1e-7 xrcrg1=12 xrcrg2=1

.end

