COMPARATOR - BSIM3 Transient Analysis
* Will comment netlist at a later time.  Regina 6/11/01
*
*One Bit Comparator. Takes Two Inputs (A and B), and returns Two Ouputs -
*node 8 - (high when two signalsare equal) and node 9 (high when A is Larger Then B).
* Transient Analysis

*circuit description

.param dtempParam=-37

M1 Anot A E1 E1  PMOS w=3.6u l=1.2u   dtemp={dtempParam}
M2 Anot A 0 0 NMOS w=1.8u l=1.2u  dtemp={dtempParam}
M3 Bnot B E1 E1  PMOS w=3.6u l=1.2u  dtemp={dtempParam}
M4 Bnot B 0 0 NMOS w=1.8u l=1.2u  dtemp={dtempParam}
M5 AorBnot 0 E1 E1 PMOS w=1.8u l=3.6u  dtemp={dtempParam}
M6 AorBnot B 1 0 NMOS w=1.8u l=1.2u  dtemp={dtempParam}
M7 1 Anot 0 0 NMOS w=1.8u l=1.2u  dtemp={dtempParam}
M8 Lnot 0 E1 E1 PMOS w=1.8u l=3.6u  dtemp={dtempParam}
M9 Lnot Bnot 2 0 NMOS w=1.8u l=1.2u  dtemp={dtempParam}
M10 2 A 0 0 NMOS w=1.8u l=1.2u  dtemp={dtempParam}
M11 Qnot 0 E1 E1  PMOS w=3.6u l=3.6u  dtemp={dtempParam}
M12 Qnot AorBnot 3 0 NMOS w=1.8u l=1.2u  dtemp={dtempParam}
M13 3 Lnot 0 0 NMOS w=1.8u l=1.2u  dtemp={dtempParam}
MQLO 8 Qnot E1 E1  PMOS w=3.6u l=1.2u  dtemp={dtempParam}
MQL1 8 Qnot 0 0 NMOS w=1.8u l=1.2u  dtemp={dtempParam}
MLTO 9 Lnot E1 E1  PMOS w=3.6u l=1.2u  dtemp={dtempParam}
MLT1 9 Lnot 0 0 NMOS w=1.8u l=1.2u  dtemp={dtempParam}
CQ Qnot 0 30f  dtemp={dtempParam}
CL Lnot 0 10f  dtemp={dtempParam}

Vdd E1 0 5
Va A 0  pulse(0 5 0ns .1ns .1ns 15ns 30ns)
Vb B 0 0

.model nmos nmos (level=9)
.model pmos pmos (level=9)

* transient analysis
.step vdd 7 5 -1
*.step temp -10 10 10
.step dtempParam -37 -17 10

*.tran 1ns 60ns
.tran 1ns 1ns

.options timeint reltol=1e-4
.print tran precision=12 width=21 {v(9)+0.2} 


.END

