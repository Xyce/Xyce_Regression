********************************************************
* Test FORMAT=GNUPLOT with .STEP.  This should produce 
* the same .NOISE.prn file as FORMAT=STD, but with two 
* blank lines before steps 1,2, ... N-1.  Note that
* first step is "step 0".  In this netlist, N is 4. 
*
********************************************************

V1  1 0 DC 5.0 AC  1.0   
R1  1 2 100K
R2  2 0 100K
*
* AMP AND LP FILTER
EAMP  3 0 2 0 1
RLP1  3 3a 100
RLP2  3a 4 100
CLP1  4 0 1.59NF

* step over two variables
.STEP RLP1 1e2 1e3 9e2
.STEP RLP2 5e2 15e2 10e2

.NOISE  V(4)  V1  DEC  5 100 100MEG 1
.PRINT NOISE FORMAT=GNUPLOT RLP1:R RLP2:R INOISE ONOISE

.END
