Netlist to Test the bsrc with multipliers, subcircuit implicit multiplier, nested subckt
****************************************************************************** 
VIN 1 0 DC 12V
Xtest 3 0 2 0 gsrcSub1 m=5

.subckt gsrcSub1 A B C D M=1
Xtest A B C D gsrcSub2 m=2
.ends

.subckt gsrcSub2 A B C D M=1
B1 A B I='v(C,D)*0.02'
.ends

R1 1 2 300
R2 2 0 900
R3 3 0 200
R4 3 0 200
.DC VIN 1 12 1
.PRINT DC V(1) V(2) V(3) 
* NOTE: XYCE DOES NOT CURRENTLY SUPPORT TRANSFER FUNCTION ANALYSIS 
* THIS PORTION HAS BEEN COMMENTED OUT UNTIL TF IS SUPPORTED
*.TF V(3) V
.END
