*Sample netlist for BSIM-MG 
*Drain current symmetry for nmos

*.options nonlin abstol=1e-6 reltol=1e-6 
.options device temp=25 

.include "modelcard111.nmos_binned"

* --- Voltage Sources ---
vdrain drain 0 dc 0
esource source 0 drain 0 -1
vgate gate  0 dc 1.0
vbulk bulk 0 dc 0.0


* --- Transistor ---
M1 drain gate source bulk nmos1 TFIN=15n L=30n NFIN=10 NRS=1 NRD=1

* --- DC Analysis ---
.dc vdrain -0.1 0.1 0.001 vgate 0.0 1.0 0.2
.print dc v(drain) v(gate) {-I(vdrain)}
.end
