*Testing Gummel-Poon BJT Model TEMP setting
*
* As part of BUG 647 (SON) fix, the instance TEMP should be getting set
* in processParams, not the instance constructor.  Test this by
* doing a .step over the instance TEMP and comparing to a .step over the
* global temp, to make sure things are getting set properly.

V1 1 0 DC 0 PWL (0 0 1 1) 
Q1 1 1 0 Qmod  TEMP=30
.model Qmod NPN level=1 ISE=1e-12 IS=1e-10 NE=1 IKF=1 CJE=10n
.tran 1u .8
.print tran V(1) I(V1) Q1:TEMP
.step lin Q1:TEMP 30 35 1
.end
