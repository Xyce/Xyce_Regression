Basic voltage divider circuit test of subcircuit usage
* Should produce results identical to Double_Resist_Control.
* Tests use of expressions in params of subcircuit *and* context issues 
* regarding those params.

.param R0=10k
XR1 1 2 Rsub R={R0}
XR2 2 0 Rsub R={R0*0.5}
V1 1 0 DC 5V

.subckt Rsub 1 2 R=1K
R1 1 2 {R}
.ends

.dc V1 0 5 1
.print DC v(1) v(2) I(v1)
.end
