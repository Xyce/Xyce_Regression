* DC simulation for xyce
.options device temp=27
.subckt mysub d_x g_x s_x b_x
e_d d_v 0 d_x 0 1
v_d d_v d 0
f_d d_x 0 v_d   -1
e_g g_v 0 g_x 0 1
v_g g_v g 0
f_g g_x 0 v_g   -1
e_s s_v 0 s_x 0 1
v_s s_v s 0
f_s s_x 0 v_s   -1
e_b b_v 0 b_x 0 1
v_b b_v b 0
f_b b_x 0 v_b   -1
m1 d g s b mymodel
+ W=10.0e-6
+ L=0.1e-6
+ AS=5e-12
+ AD=5e-12
+ PS=21e-6
+ PD=21e-6
.model mymodel nmos level=102
+ LEVEL=102.0
+ TR=27.0
+ DTA=0
+ QMC=1.0
+ LVARO=-10.0E-9
+ LVARL=0
+ LVARW=0
+ LAP=10.0E-9
+ WVARO=10.0E-9
+ WVARL=0
+ WVARW=0
+ WOT=0
+ DLQ=0
+ DWQ=0
+ VFBO=-1.1
+ VFBL=0
+ VFBW=0
+ VFBLW=0
+ STVFBO=5.0E-4
+ STVFBL=0
+ STVFBW=0
+ STVFBLW=0
+ TOXO=1.5E-9
+ EPSROXO=3.9
+ NSUBO=3.0E+23
+ NSUBW=0
+ WSEG=1.5E-10
+ NPCK=1.0E+24
+ NPCKW=0
+ WSEGP=0.9E-8
+ LPCK=5.5E-8
+ LPCKW=0
+ FOL1=2.0E-2
+ FOL2=5.0E-6
+ VNSUBO=0
+ NSLPO=0.05
+ DNSUBO=0
+ DPHIBO=0
+ DPHIBL=0
+ DPHIBLEXP=1.0
+ DPHIBW=0
+ DPHIBLW=0
+ NPO=1.5E+26
+ NPL=10.0E-18
+ CTO=5.0E-15
+ CTL=4.0E-2
+ CTLEXP=0.6
+ CTW=0
+ CTLW=0
+ TOXOVO=1.5E-9
+ TOXOVDO=2.0E-9
+ LOV=10.0E-9
+ LOVD=0
+ NOVO=7.5E+25
+ NOVDO=5.0e+25
+ CFL=3.0E-4
+ CFLEXP=2.0
+ CFW=5.0E-3
+ CFBO=0.3
+ UO=3.5E-2
+ FBET1=-0.3
+ FBET1W=0.15
+ LP1=1.5E-7
+ LP1W=-2.5E-2
+ FBET2=50.0
+ LP2=8.5E-10
+ BETW1=5.0E-2
+ BETW2=-2.0E-2
+ WBET=5.0E-10
+ STBETO=1.75
+ STBETL=-2.0E-2
+ STBETW=-2.0E-3
+ STBETLW=-3.0E-3
+ MUEO=0.6
+ MUEW=-1.2E-2
+ STMUEO=0.5
+ THEMUO=2.75
+ STTHEMUO=-0.1
+ CSO=1.0E-2
+ CSL=0
+ CSLEXP=1
+ CSW=0
+ CSLW=0
+ STCSO=-5.0
+ XCORO=0.15
+ XCORL=2.0E-3
+ XCORW=-3.0E-2
+ XCORLW=-3.5E-3
+ STXCORO=1.25
+ FETAO=1
+ RSW1=50
+ RSW2=5.0E-2
+ STRSO=-2.0
+ RSBO=0
+ RSGO=0
+ THESATO=1.0E-6
+ THESATL=0.6
+ THESATLEXP=0.75
+ THESATW=-1.0E-2
+ THESATLW=0
+ STTHESATO=1.5
+ STTHESATL=-2.5E-2
+ STTHESATW=-2.0E-2
+ STTHESATLW=-5.0E-3
+ THESATBO=0.15
+ THESATGO=0.75
+ AXO=20
+ AXL=0.2
+ ALPL=7.0E-3
+ ALPLEXP=0.6
+ ALPW=5.0E-2
+ ALP1L1=2.5E-2
+ ALP1LEXP=0.4
+ ALP1L2=0.1
+ ALP1W=8.5E-3
+ ALP2L1=0.5
+ ALP2LEXP=0
+ ALP2L2=0.5
+ ALP2W=-0.2
+ VPO=0.25
+ A1O=1.0
+ A1L=0
+ A1W=0
+ A2O=10.0
+ STA2O=-0.5
+ A3O=1.0
+ A3L=0
+ A3W=0
+ A4O=0
+ A4L=0
+ A4W=0
+ GCOO=5.0
+ IGINVLW=50.0
+ IGOVW=10.0
+ IGOVDW=0
+ STIGO=1.5
+ GC2O=1.0
+ GC3O=-1.0
+ CHIBO=3.1
+ AGIDLW=50.0
+ AGIDLDW=0
+ BGIDLO=35.0
+ BGIDLDO=41
+ STBGIDLO=-5.0E-4
+ STBGIDLDO=0
+ CGIDLO=0.15
+ CGIDLDO=0
+ CGBOVL=0
+ CFRW=5.0E-17
+ CFRDW=0
+ FNTO=1
+ NFALW=8.0E+22
+ NFBLW=3.0E7
+ NFCLW=0
+ RGO=0
+ RINT=0
+ RVPOLY=0
+ RSHG=0
+ DLSIL=0
+ RBULKO=0
+ RWELLO=0
+ RJUNDO=0
+ RJUNSO=0
+ TRJ=27.0
+ IMAX=1.0E3
+ VJUNREF=2.5
+ FJUNQ=0.03
+ CJORBOT=1.0E-3
+ CJORSTI=1.0E-9
+ CJORGAT=0.5E-9
+ VBIRBOT=0.75
+ VBIRSTI=1.0
+ VBIRGAT=0.75
+ PBOT=0.35
+ PSTI=0.35
+ PGAT=0.6
+ PHIGBOT=1.16
+ PHIGSTI=1.16
+ PHIGGAT=1.16
+ IDSATRBOT=5.0E-9
+ IDSATRSTI=1.0E-18
+ IDSATRGAT=1.0E-18
+ CSRHBOT=5.0E2
+ CSRHSTI=0
+ CSRHGAT=1.0E3
+ XJUNSTI=1.0E-8
+ XJUNGAT=1.0E-9
+ CTATBOT=5.0E2
+ CTATSTI=0
+ CTATGAT=1.0E3
+ MEFFTATBOT=0.25
+ MEFFTATSTI=0.25
+ MEFFTATGAT=0.25
+ CBBTBOT=1.0E-12
+ CBBTSTI=1.0E-18
+ CBBTGAT=1.0E-18
+ FBBTRBOT=1.0E9
+ FBBTRSTI=1.0E9
+ FBBTRGAT=1.0E9
+ STFBBTBOT=-1.0E-3
+ STFBBTSTI=-1.0E-3
+ STFBBTGAT=-1.0E-2
+ VBRBOT=10.0
+ VBRSTI=10.0
+ VBRGAT=10.0
+ PBRBOT=3
+ PBRSTI=4
+ PBRGAT=3
+ VJUNREFD=2.5
+ FJUNQD=0.03
+ CJORBOTD=1.0E-3
+ CJORSTID=1.0E-9
+ CJORGATD=1.0E-9
+ VBIRBOTD=1.0
+ VBIRSTID=1.0
+ VBIRGATD=1.0
+ PBOTD=0.5
+ PSTID=0.5
+ PGATD=0.5
+ PHIGBOTD=1.16
+ PHIGSTID=1.16
+ PHIGGATD=1.16
+ IDSATRBOTD=1.0E-12
+ IDSATRSTID=1.0E-18
+ IDSATRGATD=1.0E-18
+ CSRHBOTD=1.0E+2
+ CSRHSTID=1.0E-4
+ CSRHGATD=1.0E-4
+ XJUNSTID=1.0E-7
+ XJUNGATD=1.0E-7
+ CTATBOTD=1.0E+2
+ CTATSTID=1.0E-4
+ CTATGATD=1.0E-4
+ MEFFTATBOTD=0.25
+ MEFFTATSTID=0.25
+ MEFFTATGATD=0.25
+ CBBTBOTD=1.0E-12
+ CBBTSTID=1.0E-18
+ CBBTGATD=1.0E-18
+ FBBTRBOTD=1.0E9
+ FBBTRSTID=1.0E9
+ FBBTRGATD=1.0E9
+ STFBBTBOTD=-1.0E-3
+ STFBBTSTID=-1.0E-3
+ STFBBTGATD=-1.0E-3
+ VBRBOTD=10.0
+ VBRSTID=10.0
+ VBRGATD=10.0
+ PBRBOTD=4
+ PBRSTID=4
+ PBRGATD=4
+ SWIGATE=1
+ SWIMPACT=1
+ SWGIDL=1
+ SWJUNCAP=3
+ SWJUNASYM=0
.ends
v_d d 0 1.0
v_g g 0 -1.01
v_s s 0 0
v_b b 0 0
x1 d g s b mysub

*Second transistor for finite differencing
Bdrain d2 0 V={V(d)}
Bgate g2 0  V={V(g)+((V(g)==0)?.00000001:(1e-8*abs(v(g))))}
Bsource s2 0 V={V(s)}
Bbulk b2 0 V={V(b)}

x2 d2 g2 s2 b2 mysub

.dc v_g -1.0 1.2 0.01
*COMP {N(X1:M1:gm)-{((N(X2:M1:ids)+N(X2:M1:idb)-N(X2:M1:igd))-(N(X1:M1:ids)+N(X1:M1:idb)-N(X1:M1:igd)))/(V(g2)-V(g))}} abstol=1e-8 offset=3.2e-5
*COMP {((N(X2:M1:ids)+N(X2:M1:idb)-N(X2:M1:igd))-(N(X1:M1:ids)+N(X1:M1:idb)-N(X1:M1:igd)))/(V(g2)-V(g))} abstol=1e-8 offset=2.7e-5
*COMP {N(X1:M1:gm)} abstol=1e-8 reltol=2e-2 offset=5e-6
* PSP "Ids" is only one term of the thing gm differentiates.
.print dc v(g) v(d) {N(X1:M1:ids)+N(X1:M1:idb)-N(X1:M1:igd)}
+ {((N(X2:M1:ids)+N(X2:M1:idb)-N(X2:M1:igd))-(N(X1:M1:ids)+N(X1:M1:idb)-N(X1:M1:igd)))/(V(g2)-V(g))}
+ N(X1:M1:gm)
+ {N(X1:M1:gm)-{((N(X2:M1:ids)+N(X2:M1:idb)-N(X2:M1:igd))-(N(X1:M1:ids)+N(X1:M1:idb)-N(X1:M1:igd)))/(V(g2)-V(g))}}  N(X1:M1:Vth) N(X1:M1:Vds) N(X1:M1:Vsb) N(X1:M1:Vgs) N(X1:M1:Vdss)

.end
