* Test all three documented HSPICE syntaxes for an .INC line

.INC incFile1
.INCL incFile2
.INCLUDE incFile3

V1 1 0 1

.DC V1 1 2 1
.PRINT DC V(1) V(2) V(3)

.END
