********************************************************
* * Test -o command line option for .PRINT PCE.  The
* parameters FORMAT=CSV and FILE=pceFoo on the .PRINT PCE
* line should be ignored.  Also, no output should occur
* from the .PRINT DC line.
*
* See SON Bug 1231 for more details.
********************************************************

.global_param R1value={1000.0}
.global_param R2value={1000.0}

R2 1 0 {R2value}
R1 1 2 {R1value}
Von 2 0 5

.dc Von 5 5 1

.print dc v(1)
.PRINT PCE PRECISION=6 FORMAT=CSV FILE=pceFoo

.PCE
+ param=R1value
+ type=normal
+ means=1000.0
+ std_deviations=200.0

.options PCES
+ order=2
+ outputs={v(1)}

.options nonlin nox=0

.end
