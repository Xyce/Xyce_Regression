Transient sensitivity example, sine source, analytical sensitivity, device-level specification
*****************************************************************************
.param v0=0.3
.param va=1
.param f=500hz
.param td=0
.param phase=500
.param theta=0

* original
isin 0 1 sin({v0} {va} {f} {td} {phase} {theta})
r1   1 0 1

.tran 0.06ms 6ms
.print tran i(isin)

* Sensitivity commands
.print sens 
.sens objfunc={v(1)} sensdevicename=isin
.options sensitivity direct=1 adjoint=0 forceanalytic=true
.end
