******************************************************************
* For testing -o (SON Bug 911), the key point is that the .sh 
* file will try to overwrite the netlist (nooverwrite.cir) and 
* also to send the output to another "netlist file" (noover.cir).
* It both cases, .prn will be appended to the requested -o file.
******************************************************************

V1 1 0 PWL 0 0 1 1
R1 1 2 1
R2 2 0 1

.TRAN 0 1
.PRINT TRAN FORMAT=CSV V(1) 
.PRINT TRAN FILE=nooverwriteFoo V(2)
.OPTIONS OUTPUT INITIAL_INTERVAL=0.2 

.END


