Simple test of .RESULT capability
*

R1 a b 10.0
R2 b c 2.0
R3 c d 3.0
R4 d e 4.0
R5 e f 5.0
R6 f g 6.0
R7 g h 7.0
R8 h 0 8.0

*            V0  VA FREQ TD THETA
Va a 0  sin ( 5.0  {v_amplitude} 0.05 0.0 0.0)

* transient analysis
* Note:  For this test to work, this needs to be a format=tecplot file!
* This is because the perl script needs to determine the value of R1, 
* and that isn't output in a standard format *prn file.  It is, however, 
* in the AUXDATA that is output for tecplot.
.tran 0.5s 60s
.print tran format=tecplot v(a) v(b) {(abs(v(a)))-10.0} {((v(b)+2.0)**2.0)*1.0e3}

.global_param v_amplitude=2.0

.step R1 10.0 15.0 1 
.step v_amplitude 1.0 3.0 1.0

.result {v(a)}
.result {v(b)}
.result {(abs(v(a)))-10.0 }
.result {((v(b)+2.0)**2.0)*1.0e3}

.END
