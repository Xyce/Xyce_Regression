Test Circuit for the Hyperbolic Tangent and Hyperbolic Arctangent Functions
*******************************************************************************
* Tier No.:     1
* Directory/Circuit Name: ABM_ATANH_TANH/atanh_tanh.cir
* Description:  Test of the Xyce analog behavioral modeling hyperbolic tangent
* and hyperbolic arctangent functions.
* Input: VS
* Output: V(1), V(2), V(3)
* Analysis:
*	A sinusoidal source voltage, VS or V(1),  with a 100V amplitude and
* 	1KHZ freq. is the input to the circuit.  Two nonlinear dependent
*  	voltage sources are used to define the functions as follows:
*		V(2)=B2=TANH(V(1)) = tanh of input sine function = V(2)
*		V(3)=B3=ATANH(V(2)) = inverse tanh of B2 (or TANH(VS))=V(1)
*		        = value of the input source VS
*	A transient analysis is performed and the output recorded is the node
* 	voltages defined by the input source, V(1), the hyperbolic tangent,
*  	V(2),  and inverse hyperbolic tangent, V(3), functions.
*
*	This table is a set of hand calculations for the TANH and ATANH
* 	functions:
*	 	X		TANH(X)		ATANH(TANH(X))
*		-1.00		-0.76159416	-1.00
*		 0.00		 0.00		 0.00
*		 1.00		 0.76159416 	 1.00
*
*******************************************************************************
VS  1  0  SIN(0 100 1KHZ 0 0)
R1  1  0  1
B2  2  0  V={TANH(V(1))}
R2  2  0  1
B3  3  0  V={ATANH(V(2))}
R3  3  0  1
.TRAN 0.1MS 2MS

*COMP V(1) OFFSET=1
*COMP V(2) OFFSET=1
*COMP V(3) OFFSET=1
.PRINT TRAN V(1) V(2) V(3)
.options nonlin-tran searchmethod=1


.options  timeint method=7 erroption=1 delmax=2e-5
.END
