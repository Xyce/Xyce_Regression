RAW File Output test for B, E and F Sources.
************************************************************
* This test has two purposes:
*   1) Verify that the variable type (e.g., "current") and 
*      variable names for all the B, E and F controlled 
*      sources in the header info in the .RAW file output
*
*   2) Verify that the data is actually correct for all of
*      the time-steps in the .RAW file output 
*
* The "gold" .RAW file output was generated by manually
* comparing that "gold" file with a .PRN file.  It was 
* generated for a limited set of fixed time-steps, so that
* a file comparison could be used to verify the test output's
* .RAW file against that "gold" .RAW file.
************************************************************  

* Test linear, POLY, VALUE and TABLE formats
ELIN  3 0 1 0 1
R3    3 4 1K
R4    0 4 100

EPOLY 5 0 POLY(2) 3 0 4 0 0 .5 .5
R5    5 6 1K
R6    0 6 100

EVALUE 7 0 VALUE = 5V*SQRT(V(1,0))
R7     7 8 1K
R8     0 8 100

ETABLE  9 0 TABLE V(1,0) = (0,1) (1,2)
R9      9 10 1K
R10     0 10 100

* Test both linear and POLY formats
FLIN   11  0 B1 1
R11    11 12 1K
R12     0 12 100

FPOLY  13  0 POLY(1) B1 0 1
R13    13 14 1K
R14     0 14 100

B1   1 0 V={2.0*sin(2*pi*TIME) }
R1   1 2 1K
R2   0 2 100

* Add a V source for good measure
V15 15 0 1
R15 15 0 1

.options output initial_interval=0.05
.TRAN 0 1.0

* .PRINT statement is not actually used for .RAW output.
* It was included in the netslit so that the "gold" .RAW 
* file output could manually verified against a .PRN file
* during test development
.PRINT TRAN v(1) v(10) v(11) v(12) v(13) v(14) 
+ v(15) v(2) v(3) v(4) v(5) v(6) v(7) v(8) v(9)
+ I(B1) I(ELIN) I(EPOLY) I(ETABLE) I(EVALUE) I(V15)

.END
