*******************************************************************************
* This netlist is equivalent to Step 3 for the IntegralTest.cir netlist.
* It has VS1:VA=2 and VS3:V0=-0.5
*
*******************************************************************************
*
* a few sources of different types
VS1  1  0  SIN(0 2 50Hz 0 0)
VP  2  0  PULSE( 0 100 0.2ms 0.2ms 0.2ms 1ms 2ms )
VS3  3  0  SIN(-0.5 1.0 250HZ 0 500)
VS4  4  0  SIN(0.5 -1.0 250HZ 0 500)

R1  1  0  100
R2  2  0  100
R3  3  0  100
R4  4  0  100

* Use MEASFAIL to test the reset of the default calculation value
.OPTIONS MEASURE MEASFAIL=0

.TRAN 0  10ms
.PRINT TRAN FORMAT=NOINDEX V(1) V(2) V(3) V(4)

.measure tran intAll INTEGRAL v(1)
.measure tran intTop INTEG v(2)

* add TO-FROM modifiers
.measure tran sineHalfInterval Integ V(1) from=0 to=0.001

* mix in TDs before and after FROM value.
.measure tran sineTDbetween integ V(1) FROM=0 TO=0.005 TD=0.001
.measure tran sineTDbefore integ V(1) FROM=0.002 TO=0.005 TD=0.001

* these tests should return -1 and -100
.measure tran returnNegOne integ V(1) FROM=0.2e-3 TO=0.25e-3 TD=0.5e-3 default_val=-1
.measure tran returnNeg100 integ V(1) FROM=0.2e-3 TO=0.25e-3 TD=0.5e-3 default_val=-100

.END

