Regression test for simple normal distribution sampling

R2 1 0 {agauss(2k,0.2k,1)}
R1 1 2 {agauss(3k,0.1k,1)}
v1 2 0 10V

.dc v1 10 10 1

.print dc format=tecplot v(1)

.SAMPLING 
+ useExpr=true

.options SAMPLES numsamples=50
+ projection_pce=true
*+ regression_pce=true
+ output_pce_coeffs=true
+ order=3
+ outputs={v(1)}
+ sample_type=lhs
+ stdoutput=true

.end

