cable simulation - rallpack 1 with 1000 level 1 neurons


.tran 0 0.25  
.options output initial_interval=5.0e-5
.options timeint method=7 newlte=1 newbpstepping=1 reltol=1e-3
.options linsol type=klu

* rallpack 1 calls for a steady current input.  But we need to use PULSE so
* that the current will be off during dcop calculation
Iin 0 in0 PULSE( 0 1.0e-10 1.0e-12 0.0 0.0 1.0e10 1.0e10)

* cable is 1mm long and 1 micron in diameter
* 1000 segments, each 1 micron long and 1 micron in diameter
.param nSeg = 1000
.param segLength = 1.0e-4     ; [cm]
.param segDiameter = 1.0e-4   ; [cm]
.param segSurfaceArea = { 3.14159 * segDiameter * segLength }

* specific membrane capacitance 1uF/cm^2 
.param memC = { 1.0e-6 * segSurfaceArea } ; [F]

* leak current has membrane resistivity of 40,000 ohm cm^2, with reversal potential of -65mV
.param rm = { 4.0e4 / segSurfaceArea }    ; [ohm]
.param memG = { 1 / rm }                  ; [1/ohm]
.param revE = -0.065                      ; [V]

* no active conductances, so set g values to 0; E values don't matter
.param gks  = 0.0
.param gnas = 0.0

* neuron model
.model segParams neuron level=1 cMem={memC}  gMem={memG} eLeak={revE}  gNa={gnas}  gK={gks} vRest={revE}

* segments are connected by a resistor; axial resistance is 4*Ra*l/(pi*d^2); Ra for rallpack 1 is 100 ohm cm
* if segments were different, we'd want two resistors between each pair of segments to handle the differences, but here it doesnt' matter
.param Ra = 100.0
.param rInterSeg = { 4 * Ra * segLength / ( 3.14159 * segDiameter * segDiameter ) }

* here is how we define one neuron
* yneuron neuron1 in1 0 segParams

* loop below creates a resistor between each pair of neuron devices, which means one less resistor than compartments
* add a resistor with resistivity for half a compartment at each end of the cable
* this is the first one
R01 in0 in1 {rInterSeg/2.0} 
 
  
yneuron neuron1 in1 0 segParams
R12 in1 in2 {rInterSeg}
yneuron neuron2 in2 0 segParams
R23 in2 in3 {rInterSeg}
yneuron neuron3 in3 0 segParams
R34 in3 in4 {rInterSeg}
yneuron neuron4 in4 0 segParams
R45 in4 in5 {rInterSeg}
yneuron neuron5 in5 0 segParams
R56 in5 in6 {rInterSeg}
yneuron neuron6 in6 0 segParams
R67 in6 in7 {rInterSeg}
yneuron neuron7 in7 0 segParams
R78 in7 in8 {rInterSeg}
yneuron neuron8 in8 0 segParams
R89 in8 in9 {rInterSeg}
yneuron neuron9 in9 0 segParams
R910 in9 in10 {rInterSeg}
yneuron neuron10 in10 0 segParams
R1011 in10 in11 {rInterSeg}
yneuron neuron11 in11 0 segParams
R1112 in11 in12 {rInterSeg}
yneuron neuron12 in12 0 segParams
R1213 in12 in13 {rInterSeg}
yneuron neuron13 in13 0 segParams
R1314 in13 in14 {rInterSeg}
yneuron neuron14 in14 0 segParams
R1415 in14 in15 {rInterSeg}
yneuron neuron15 in15 0 segParams
R1516 in15 in16 {rInterSeg}
yneuron neuron16 in16 0 segParams
R1617 in16 in17 {rInterSeg}
yneuron neuron17 in17 0 segParams
R1718 in17 in18 {rInterSeg}
yneuron neuron18 in18 0 segParams
R1819 in18 in19 {rInterSeg}
yneuron neuron19 in19 0 segParams
R1920 in19 in20 {rInterSeg}
yneuron neuron20 in20 0 segParams
R2021 in20 in21 {rInterSeg}
yneuron neuron21 in21 0 segParams
R2122 in21 in22 {rInterSeg}
yneuron neuron22 in22 0 segParams
R2223 in22 in23 {rInterSeg}
yneuron neuron23 in23 0 segParams
R2324 in23 in24 {rInterSeg}
yneuron neuron24 in24 0 segParams
R2425 in24 in25 {rInterSeg}
yneuron neuron25 in25 0 segParams
R2526 in25 in26 {rInterSeg}
yneuron neuron26 in26 0 segParams
R2627 in26 in27 {rInterSeg}
yneuron neuron27 in27 0 segParams
R2728 in27 in28 {rInterSeg}
yneuron neuron28 in28 0 segParams
R2829 in28 in29 {rInterSeg}
yneuron neuron29 in29 0 segParams
R2930 in29 in30 {rInterSeg}
yneuron neuron30 in30 0 segParams
R3031 in30 in31 {rInterSeg}
yneuron neuron31 in31 0 segParams
R3132 in31 in32 {rInterSeg}
yneuron neuron32 in32 0 segParams
R3233 in32 in33 {rInterSeg}
yneuron neuron33 in33 0 segParams
R3334 in33 in34 {rInterSeg}
yneuron neuron34 in34 0 segParams
R3435 in34 in35 {rInterSeg}
yneuron neuron35 in35 0 segParams
R3536 in35 in36 {rInterSeg}
yneuron neuron36 in36 0 segParams
R3637 in36 in37 {rInterSeg}
yneuron neuron37 in37 0 segParams
R3738 in37 in38 {rInterSeg}
yneuron neuron38 in38 0 segParams
R3839 in38 in39 {rInterSeg}
yneuron neuron39 in39 0 segParams
R3940 in39 in40 {rInterSeg}
yneuron neuron40 in40 0 segParams
R4041 in40 in41 {rInterSeg}
yneuron neuron41 in41 0 segParams
R4142 in41 in42 {rInterSeg}
yneuron neuron42 in42 0 segParams
R4243 in42 in43 {rInterSeg}
yneuron neuron43 in43 0 segParams
R4344 in43 in44 {rInterSeg}
yneuron neuron44 in44 0 segParams
R4445 in44 in45 {rInterSeg}
yneuron neuron45 in45 0 segParams
R4546 in45 in46 {rInterSeg}
yneuron neuron46 in46 0 segParams
R4647 in46 in47 {rInterSeg}
yneuron neuron47 in47 0 segParams
R4748 in47 in48 {rInterSeg}
yneuron neuron48 in48 0 segParams
R4849 in48 in49 {rInterSeg}
yneuron neuron49 in49 0 segParams
R4950 in49 in50 {rInterSeg}
yneuron neuron50 in50 0 segParams
R5051 in50 in51 {rInterSeg}
yneuron neuron51 in51 0 segParams
R5152 in51 in52 {rInterSeg}
yneuron neuron52 in52 0 segParams
R5253 in52 in53 {rInterSeg}
yneuron neuron53 in53 0 segParams
R5354 in53 in54 {rInterSeg}
yneuron neuron54 in54 0 segParams
R5455 in54 in55 {rInterSeg}
yneuron neuron55 in55 0 segParams
R5556 in55 in56 {rInterSeg}
yneuron neuron56 in56 0 segParams
R5657 in56 in57 {rInterSeg}
yneuron neuron57 in57 0 segParams
R5758 in57 in58 {rInterSeg}
yneuron neuron58 in58 0 segParams
R5859 in58 in59 {rInterSeg}
yneuron neuron59 in59 0 segParams
R5960 in59 in60 {rInterSeg}
yneuron neuron60 in60 0 segParams
R6061 in60 in61 {rInterSeg}
yneuron neuron61 in61 0 segParams
R6162 in61 in62 {rInterSeg}
yneuron neuron62 in62 0 segParams
R6263 in62 in63 {rInterSeg}
yneuron neuron63 in63 0 segParams
R6364 in63 in64 {rInterSeg}
yneuron neuron64 in64 0 segParams
R6465 in64 in65 {rInterSeg}
yneuron neuron65 in65 0 segParams
R6566 in65 in66 {rInterSeg}
yneuron neuron66 in66 0 segParams
R6667 in66 in67 {rInterSeg}
yneuron neuron67 in67 0 segParams
R6768 in67 in68 {rInterSeg}
yneuron neuron68 in68 0 segParams
R6869 in68 in69 {rInterSeg}
yneuron neuron69 in69 0 segParams
R6970 in69 in70 {rInterSeg}
yneuron neuron70 in70 0 segParams
R7071 in70 in71 {rInterSeg}
yneuron neuron71 in71 0 segParams
R7172 in71 in72 {rInterSeg}
yneuron neuron72 in72 0 segParams
R7273 in72 in73 {rInterSeg}
yneuron neuron73 in73 0 segParams
R7374 in73 in74 {rInterSeg}
yneuron neuron74 in74 0 segParams
R7475 in74 in75 {rInterSeg}
yneuron neuron75 in75 0 segParams
R7576 in75 in76 {rInterSeg}
yneuron neuron76 in76 0 segParams
R7677 in76 in77 {rInterSeg}
yneuron neuron77 in77 0 segParams
R7778 in77 in78 {rInterSeg}
yneuron neuron78 in78 0 segParams
R7879 in78 in79 {rInterSeg}
yneuron neuron79 in79 0 segParams
R7980 in79 in80 {rInterSeg}
yneuron neuron80 in80 0 segParams
R8081 in80 in81 {rInterSeg}
yneuron neuron81 in81 0 segParams
R8182 in81 in82 {rInterSeg}
yneuron neuron82 in82 0 segParams
R8283 in82 in83 {rInterSeg}
yneuron neuron83 in83 0 segParams
R8384 in83 in84 {rInterSeg}
yneuron neuron84 in84 0 segParams
R8485 in84 in85 {rInterSeg}
yneuron neuron85 in85 0 segParams
R8586 in85 in86 {rInterSeg}
yneuron neuron86 in86 0 segParams
R8687 in86 in87 {rInterSeg}
yneuron neuron87 in87 0 segParams
R8788 in87 in88 {rInterSeg}
yneuron neuron88 in88 0 segParams
R8889 in88 in89 {rInterSeg}
yneuron neuron89 in89 0 segParams
R8990 in89 in90 {rInterSeg}
yneuron neuron90 in90 0 segParams
R9091 in90 in91 {rInterSeg}
yneuron neuron91 in91 0 segParams
R9192 in91 in92 {rInterSeg}
yneuron neuron92 in92 0 segParams
R9293 in92 in93 {rInterSeg}
yneuron neuron93 in93 0 segParams
R9394 in93 in94 {rInterSeg}
yneuron neuron94 in94 0 segParams
R9495 in94 in95 {rInterSeg}
yneuron neuron95 in95 0 segParams
R9596 in95 in96 {rInterSeg}
yneuron neuron96 in96 0 segParams
R9697 in96 in97 {rInterSeg}
yneuron neuron97 in97 0 segParams
R9798 in97 in98 {rInterSeg}
yneuron neuron98 in98 0 segParams
R9899 in98 in99 {rInterSeg}
yneuron neuron99 in99 0 segParams
R99100 in99 in100 {rInterSeg}
yneuron neuron100 in100 0 segParams
R100101 in100 in101 {rInterSeg}
yneuron neuron101 in101 0 segParams
R101102 in101 in102 {rInterSeg}
yneuron neuron102 in102 0 segParams
R102103 in102 in103 {rInterSeg}
yneuron neuron103 in103 0 segParams
R103104 in103 in104 {rInterSeg}
yneuron neuron104 in104 0 segParams
R104105 in104 in105 {rInterSeg}
yneuron neuron105 in105 0 segParams
R105106 in105 in106 {rInterSeg}
yneuron neuron106 in106 0 segParams
R106107 in106 in107 {rInterSeg}
yneuron neuron107 in107 0 segParams
R107108 in107 in108 {rInterSeg}
yneuron neuron108 in108 0 segParams
R108109 in108 in109 {rInterSeg}
yneuron neuron109 in109 0 segParams
R109110 in109 in110 {rInterSeg}
yneuron neuron110 in110 0 segParams
R110111 in110 in111 {rInterSeg}
yneuron neuron111 in111 0 segParams
R111112 in111 in112 {rInterSeg}
yneuron neuron112 in112 0 segParams
R112113 in112 in113 {rInterSeg}
yneuron neuron113 in113 0 segParams
R113114 in113 in114 {rInterSeg}
yneuron neuron114 in114 0 segParams
R114115 in114 in115 {rInterSeg}
yneuron neuron115 in115 0 segParams
R115116 in115 in116 {rInterSeg}
yneuron neuron116 in116 0 segParams
R116117 in116 in117 {rInterSeg}
yneuron neuron117 in117 0 segParams
R117118 in117 in118 {rInterSeg}
yneuron neuron118 in118 0 segParams
R118119 in118 in119 {rInterSeg}
yneuron neuron119 in119 0 segParams
R119120 in119 in120 {rInterSeg}
yneuron neuron120 in120 0 segParams
R120121 in120 in121 {rInterSeg}
yneuron neuron121 in121 0 segParams
R121122 in121 in122 {rInterSeg}
yneuron neuron122 in122 0 segParams
R122123 in122 in123 {rInterSeg}
yneuron neuron123 in123 0 segParams
R123124 in123 in124 {rInterSeg}
yneuron neuron124 in124 0 segParams
R124125 in124 in125 {rInterSeg}
yneuron neuron125 in125 0 segParams
R125126 in125 in126 {rInterSeg}
yneuron neuron126 in126 0 segParams
R126127 in126 in127 {rInterSeg}
yneuron neuron127 in127 0 segParams
R127128 in127 in128 {rInterSeg}
yneuron neuron128 in128 0 segParams
R128129 in128 in129 {rInterSeg}
yneuron neuron129 in129 0 segParams
R129130 in129 in130 {rInterSeg}
yneuron neuron130 in130 0 segParams
R130131 in130 in131 {rInterSeg}
yneuron neuron131 in131 0 segParams
R131132 in131 in132 {rInterSeg}
yneuron neuron132 in132 0 segParams
R132133 in132 in133 {rInterSeg}
yneuron neuron133 in133 0 segParams
R133134 in133 in134 {rInterSeg}
yneuron neuron134 in134 0 segParams
R134135 in134 in135 {rInterSeg}
yneuron neuron135 in135 0 segParams
R135136 in135 in136 {rInterSeg}
yneuron neuron136 in136 0 segParams
R136137 in136 in137 {rInterSeg}
yneuron neuron137 in137 0 segParams
R137138 in137 in138 {rInterSeg}
yneuron neuron138 in138 0 segParams
R138139 in138 in139 {rInterSeg}
yneuron neuron139 in139 0 segParams
R139140 in139 in140 {rInterSeg}
yneuron neuron140 in140 0 segParams
R140141 in140 in141 {rInterSeg}
yneuron neuron141 in141 0 segParams
R141142 in141 in142 {rInterSeg}
yneuron neuron142 in142 0 segParams
R142143 in142 in143 {rInterSeg}
yneuron neuron143 in143 0 segParams
R143144 in143 in144 {rInterSeg}
yneuron neuron144 in144 0 segParams
R144145 in144 in145 {rInterSeg}
yneuron neuron145 in145 0 segParams
R145146 in145 in146 {rInterSeg}
yneuron neuron146 in146 0 segParams
R146147 in146 in147 {rInterSeg}
yneuron neuron147 in147 0 segParams
R147148 in147 in148 {rInterSeg}
yneuron neuron148 in148 0 segParams
R148149 in148 in149 {rInterSeg}
yneuron neuron149 in149 0 segParams
R149150 in149 in150 {rInterSeg}
yneuron neuron150 in150 0 segParams
R150151 in150 in151 {rInterSeg}
yneuron neuron151 in151 0 segParams
R151152 in151 in152 {rInterSeg}
yneuron neuron152 in152 0 segParams
R152153 in152 in153 {rInterSeg}
yneuron neuron153 in153 0 segParams
R153154 in153 in154 {rInterSeg}
yneuron neuron154 in154 0 segParams
R154155 in154 in155 {rInterSeg}
yneuron neuron155 in155 0 segParams
R155156 in155 in156 {rInterSeg}
yneuron neuron156 in156 0 segParams
R156157 in156 in157 {rInterSeg}
yneuron neuron157 in157 0 segParams
R157158 in157 in158 {rInterSeg}
yneuron neuron158 in158 0 segParams
R158159 in158 in159 {rInterSeg}
yneuron neuron159 in159 0 segParams
R159160 in159 in160 {rInterSeg}
yneuron neuron160 in160 0 segParams
R160161 in160 in161 {rInterSeg}
yneuron neuron161 in161 0 segParams
R161162 in161 in162 {rInterSeg}
yneuron neuron162 in162 0 segParams
R162163 in162 in163 {rInterSeg}
yneuron neuron163 in163 0 segParams
R163164 in163 in164 {rInterSeg}
yneuron neuron164 in164 0 segParams
R164165 in164 in165 {rInterSeg}
yneuron neuron165 in165 0 segParams
R165166 in165 in166 {rInterSeg}
yneuron neuron166 in166 0 segParams
R166167 in166 in167 {rInterSeg}
yneuron neuron167 in167 0 segParams
R167168 in167 in168 {rInterSeg}
yneuron neuron168 in168 0 segParams
R168169 in168 in169 {rInterSeg}
yneuron neuron169 in169 0 segParams
R169170 in169 in170 {rInterSeg}
yneuron neuron170 in170 0 segParams
R170171 in170 in171 {rInterSeg}
yneuron neuron171 in171 0 segParams
R171172 in171 in172 {rInterSeg}
yneuron neuron172 in172 0 segParams
R172173 in172 in173 {rInterSeg}
yneuron neuron173 in173 0 segParams
R173174 in173 in174 {rInterSeg}
yneuron neuron174 in174 0 segParams
R174175 in174 in175 {rInterSeg}
yneuron neuron175 in175 0 segParams
R175176 in175 in176 {rInterSeg}
yneuron neuron176 in176 0 segParams
R176177 in176 in177 {rInterSeg}
yneuron neuron177 in177 0 segParams
R177178 in177 in178 {rInterSeg}
yneuron neuron178 in178 0 segParams
R178179 in178 in179 {rInterSeg}
yneuron neuron179 in179 0 segParams
R179180 in179 in180 {rInterSeg}
yneuron neuron180 in180 0 segParams
R180181 in180 in181 {rInterSeg}
yneuron neuron181 in181 0 segParams
R181182 in181 in182 {rInterSeg}
yneuron neuron182 in182 0 segParams
R182183 in182 in183 {rInterSeg}
yneuron neuron183 in183 0 segParams
R183184 in183 in184 {rInterSeg}
yneuron neuron184 in184 0 segParams
R184185 in184 in185 {rInterSeg}
yneuron neuron185 in185 0 segParams
R185186 in185 in186 {rInterSeg}
yneuron neuron186 in186 0 segParams
R186187 in186 in187 {rInterSeg}
yneuron neuron187 in187 0 segParams
R187188 in187 in188 {rInterSeg}
yneuron neuron188 in188 0 segParams
R188189 in188 in189 {rInterSeg}
yneuron neuron189 in189 0 segParams
R189190 in189 in190 {rInterSeg}
yneuron neuron190 in190 0 segParams
R190191 in190 in191 {rInterSeg}
yneuron neuron191 in191 0 segParams
R191192 in191 in192 {rInterSeg}
yneuron neuron192 in192 0 segParams
R192193 in192 in193 {rInterSeg}
yneuron neuron193 in193 0 segParams
R193194 in193 in194 {rInterSeg}
yneuron neuron194 in194 0 segParams
R194195 in194 in195 {rInterSeg}
yneuron neuron195 in195 0 segParams
R195196 in195 in196 {rInterSeg}
yneuron neuron196 in196 0 segParams
R196197 in196 in197 {rInterSeg}
yneuron neuron197 in197 0 segParams
R197198 in197 in198 {rInterSeg}
yneuron neuron198 in198 0 segParams
R198199 in198 in199 {rInterSeg}
yneuron neuron199 in199 0 segParams
R199200 in199 in200 {rInterSeg}
yneuron neuron200 in200 0 segParams
R200201 in200 in201 {rInterSeg}
yneuron neuron201 in201 0 segParams
R201202 in201 in202 {rInterSeg}
yneuron neuron202 in202 0 segParams
R202203 in202 in203 {rInterSeg}
yneuron neuron203 in203 0 segParams
R203204 in203 in204 {rInterSeg}
yneuron neuron204 in204 0 segParams
R204205 in204 in205 {rInterSeg}
yneuron neuron205 in205 0 segParams
R205206 in205 in206 {rInterSeg}
yneuron neuron206 in206 0 segParams
R206207 in206 in207 {rInterSeg}
yneuron neuron207 in207 0 segParams
R207208 in207 in208 {rInterSeg}
yneuron neuron208 in208 0 segParams
R208209 in208 in209 {rInterSeg}
yneuron neuron209 in209 0 segParams
R209210 in209 in210 {rInterSeg}
yneuron neuron210 in210 0 segParams
R210211 in210 in211 {rInterSeg}
yneuron neuron211 in211 0 segParams
R211212 in211 in212 {rInterSeg}
yneuron neuron212 in212 0 segParams
R212213 in212 in213 {rInterSeg}
yneuron neuron213 in213 0 segParams
R213214 in213 in214 {rInterSeg}
yneuron neuron214 in214 0 segParams
R214215 in214 in215 {rInterSeg}
yneuron neuron215 in215 0 segParams
R215216 in215 in216 {rInterSeg}
yneuron neuron216 in216 0 segParams
R216217 in216 in217 {rInterSeg}
yneuron neuron217 in217 0 segParams
R217218 in217 in218 {rInterSeg}
yneuron neuron218 in218 0 segParams
R218219 in218 in219 {rInterSeg}
yneuron neuron219 in219 0 segParams
R219220 in219 in220 {rInterSeg}
yneuron neuron220 in220 0 segParams
R220221 in220 in221 {rInterSeg}
yneuron neuron221 in221 0 segParams
R221222 in221 in222 {rInterSeg}
yneuron neuron222 in222 0 segParams
R222223 in222 in223 {rInterSeg}
yneuron neuron223 in223 0 segParams
R223224 in223 in224 {rInterSeg}
yneuron neuron224 in224 0 segParams
R224225 in224 in225 {rInterSeg}
yneuron neuron225 in225 0 segParams
R225226 in225 in226 {rInterSeg}
yneuron neuron226 in226 0 segParams
R226227 in226 in227 {rInterSeg}
yneuron neuron227 in227 0 segParams
R227228 in227 in228 {rInterSeg}
yneuron neuron228 in228 0 segParams
R228229 in228 in229 {rInterSeg}
yneuron neuron229 in229 0 segParams
R229230 in229 in230 {rInterSeg}
yneuron neuron230 in230 0 segParams
R230231 in230 in231 {rInterSeg}
yneuron neuron231 in231 0 segParams
R231232 in231 in232 {rInterSeg}
yneuron neuron232 in232 0 segParams
R232233 in232 in233 {rInterSeg}
yneuron neuron233 in233 0 segParams
R233234 in233 in234 {rInterSeg}
yneuron neuron234 in234 0 segParams
R234235 in234 in235 {rInterSeg}
yneuron neuron235 in235 0 segParams
R235236 in235 in236 {rInterSeg}
yneuron neuron236 in236 0 segParams
R236237 in236 in237 {rInterSeg}
yneuron neuron237 in237 0 segParams
R237238 in237 in238 {rInterSeg}
yneuron neuron238 in238 0 segParams
R238239 in238 in239 {rInterSeg}
yneuron neuron239 in239 0 segParams
R239240 in239 in240 {rInterSeg}
yneuron neuron240 in240 0 segParams
R240241 in240 in241 {rInterSeg}
yneuron neuron241 in241 0 segParams
R241242 in241 in242 {rInterSeg}
yneuron neuron242 in242 0 segParams
R242243 in242 in243 {rInterSeg}
yneuron neuron243 in243 0 segParams
R243244 in243 in244 {rInterSeg}
yneuron neuron244 in244 0 segParams
R244245 in244 in245 {rInterSeg}
yneuron neuron245 in245 0 segParams
R245246 in245 in246 {rInterSeg}
yneuron neuron246 in246 0 segParams
R246247 in246 in247 {rInterSeg}
yneuron neuron247 in247 0 segParams
R247248 in247 in248 {rInterSeg}
yneuron neuron248 in248 0 segParams
R248249 in248 in249 {rInterSeg}
yneuron neuron249 in249 0 segParams
R249250 in249 in250 {rInterSeg}
yneuron neuron250 in250 0 segParams
R250251 in250 in251 {rInterSeg}
yneuron neuron251 in251 0 segParams
R251252 in251 in252 {rInterSeg}
yneuron neuron252 in252 0 segParams
R252253 in252 in253 {rInterSeg}
yneuron neuron253 in253 0 segParams
R253254 in253 in254 {rInterSeg}
yneuron neuron254 in254 0 segParams
R254255 in254 in255 {rInterSeg}
yneuron neuron255 in255 0 segParams
R255256 in255 in256 {rInterSeg}
yneuron neuron256 in256 0 segParams
R256257 in256 in257 {rInterSeg}
yneuron neuron257 in257 0 segParams
R257258 in257 in258 {rInterSeg}
yneuron neuron258 in258 0 segParams
R258259 in258 in259 {rInterSeg}
yneuron neuron259 in259 0 segParams
R259260 in259 in260 {rInterSeg}
yneuron neuron260 in260 0 segParams
R260261 in260 in261 {rInterSeg}
yneuron neuron261 in261 0 segParams
R261262 in261 in262 {rInterSeg}
yneuron neuron262 in262 0 segParams
R262263 in262 in263 {rInterSeg}
yneuron neuron263 in263 0 segParams
R263264 in263 in264 {rInterSeg}
yneuron neuron264 in264 0 segParams
R264265 in264 in265 {rInterSeg}
yneuron neuron265 in265 0 segParams
R265266 in265 in266 {rInterSeg}
yneuron neuron266 in266 0 segParams
R266267 in266 in267 {rInterSeg}
yneuron neuron267 in267 0 segParams
R267268 in267 in268 {rInterSeg}
yneuron neuron268 in268 0 segParams
R268269 in268 in269 {rInterSeg}
yneuron neuron269 in269 0 segParams
R269270 in269 in270 {rInterSeg}
yneuron neuron270 in270 0 segParams
R270271 in270 in271 {rInterSeg}
yneuron neuron271 in271 0 segParams
R271272 in271 in272 {rInterSeg}
yneuron neuron272 in272 0 segParams
R272273 in272 in273 {rInterSeg}
yneuron neuron273 in273 0 segParams
R273274 in273 in274 {rInterSeg}
yneuron neuron274 in274 0 segParams
R274275 in274 in275 {rInterSeg}
yneuron neuron275 in275 0 segParams
R275276 in275 in276 {rInterSeg}
yneuron neuron276 in276 0 segParams
R276277 in276 in277 {rInterSeg}
yneuron neuron277 in277 0 segParams
R277278 in277 in278 {rInterSeg}
yneuron neuron278 in278 0 segParams
R278279 in278 in279 {rInterSeg}
yneuron neuron279 in279 0 segParams
R279280 in279 in280 {rInterSeg}
yneuron neuron280 in280 0 segParams
R280281 in280 in281 {rInterSeg}
yneuron neuron281 in281 0 segParams
R281282 in281 in282 {rInterSeg}
yneuron neuron282 in282 0 segParams
R282283 in282 in283 {rInterSeg}
yneuron neuron283 in283 0 segParams
R283284 in283 in284 {rInterSeg}
yneuron neuron284 in284 0 segParams
R284285 in284 in285 {rInterSeg}
yneuron neuron285 in285 0 segParams
R285286 in285 in286 {rInterSeg}
yneuron neuron286 in286 0 segParams
R286287 in286 in287 {rInterSeg}
yneuron neuron287 in287 0 segParams
R287288 in287 in288 {rInterSeg}
yneuron neuron288 in288 0 segParams
R288289 in288 in289 {rInterSeg}
yneuron neuron289 in289 0 segParams
R289290 in289 in290 {rInterSeg}
yneuron neuron290 in290 0 segParams
R290291 in290 in291 {rInterSeg}
yneuron neuron291 in291 0 segParams
R291292 in291 in292 {rInterSeg}
yneuron neuron292 in292 0 segParams
R292293 in292 in293 {rInterSeg}
yneuron neuron293 in293 0 segParams
R293294 in293 in294 {rInterSeg}
yneuron neuron294 in294 0 segParams
R294295 in294 in295 {rInterSeg}
yneuron neuron295 in295 0 segParams
R295296 in295 in296 {rInterSeg}
yneuron neuron296 in296 0 segParams
R296297 in296 in297 {rInterSeg}
yneuron neuron297 in297 0 segParams
R297298 in297 in298 {rInterSeg}
yneuron neuron298 in298 0 segParams
R298299 in298 in299 {rInterSeg}
yneuron neuron299 in299 0 segParams
R299300 in299 in300 {rInterSeg}
yneuron neuron300 in300 0 segParams
R300301 in300 in301 {rInterSeg}
yneuron neuron301 in301 0 segParams
R301302 in301 in302 {rInterSeg}
yneuron neuron302 in302 0 segParams
R302303 in302 in303 {rInterSeg}
yneuron neuron303 in303 0 segParams
R303304 in303 in304 {rInterSeg}
yneuron neuron304 in304 0 segParams
R304305 in304 in305 {rInterSeg}
yneuron neuron305 in305 0 segParams
R305306 in305 in306 {rInterSeg}
yneuron neuron306 in306 0 segParams
R306307 in306 in307 {rInterSeg}
yneuron neuron307 in307 0 segParams
R307308 in307 in308 {rInterSeg}
yneuron neuron308 in308 0 segParams
R308309 in308 in309 {rInterSeg}
yneuron neuron309 in309 0 segParams
R309310 in309 in310 {rInterSeg}
yneuron neuron310 in310 0 segParams
R310311 in310 in311 {rInterSeg}
yneuron neuron311 in311 0 segParams
R311312 in311 in312 {rInterSeg}
yneuron neuron312 in312 0 segParams
R312313 in312 in313 {rInterSeg}
yneuron neuron313 in313 0 segParams
R313314 in313 in314 {rInterSeg}
yneuron neuron314 in314 0 segParams
R314315 in314 in315 {rInterSeg}
yneuron neuron315 in315 0 segParams
R315316 in315 in316 {rInterSeg}
yneuron neuron316 in316 0 segParams
R316317 in316 in317 {rInterSeg}
yneuron neuron317 in317 0 segParams
R317318 in317 in318 {rInterSeg}
yneuron neuron318 in318 0 segParams
R318319 in318 in319 {rInterSeg}
yneuron neuron319 in319 0 segParams
R319320 in319 in320 {rInterSeg}
yneuron neuron320 in320 0 segParams
R320321 in320 in321 {rInterSeg}
yneuron neuron321 in321 0 segParams
R321322 in321 in322 {rInterSeg}
yneuron neuron322 in322 0 segParams
R322323 in322 in323 {rInterSeg}
yneuron neuron323 in323 0 segParams
R323324 in323 in324 {rInterSeg}
yneuron neuron324 in324 0 segParams
R324325 in324 in325 {rInterSeg}
yneuron neuron325 in325 0 segParams
R325326 in325 in326 {rInterSeg}
yneuron neuron326 in326 0 segParams
R326327 in326 in327 {rInterSeg}
yneuron neuron327 in327 0 segParams
R327328 in327 in328 {rInterSeg}
yneuron neuron328 in328 0 segParams
R328329 in328 in329 {rInterSeg}
yneuron neuron329 in329 0 segParams
R329330 in329 in330 {rInterSeg}
yneuron neuron330 in330 0 segParams
R330331 in330 in331 {rInterSeg}
yneuron neuron331 in331 0 segParams
R331332 in331 in332 {rInterSeg}
yneuron neuron332 in332 0 segParams
R332333 in332 in333 {rInterSeg}
yneuron neuron333 in333 0 segParams
R333334 in333 in334 {rInterSeg}
yneuron neuron334 in334 0 segParams
R334335 in334 in335 {rInterSeg}
yneuron neuron335 in335 0 segParams
R335336 in335 in336 {rInterSeg}
yneuron neuron336 in336 0 segParams
R336337 in336 in337 {rInterSeg}
yneuron neuron337 in337 0 segParams
R337338 in337 in338 {rInterSeg}
yneuron neuron338 in338 0 segParams
R338339 in338 in339 {rInterSeg}
yneuron neuron339 in339 0 segParams
R339340 in339 in340 {rInterSeg}
yneuron neuron340 in340 0 segParams
R340341 in340 in341 {rInterSeg}
yneuron neuron341 in341 0 segParams
R341342 in341 in342 {rInterSeg}
yneuron neuron342 in342 0 segParams
R342343 in342 in343 {rInterSeg}
yneuron neuron343 in343 0 segParams
R343344 in343 in344 {rInterSeg}
yneuron neuron344 in344 0 segParams
R344345 in344 in345 {rInterSeg}
yneuron neuron345 in345 0 segParams
R345346 in345 in346 {rInterSeg}
yneuron neuron346 in346 0 segParams
R346347 in346 in347 {rInterSeg}
yneuron neuron347 in347 0 segParams
R347348 in347 in348 {rInterSeg}
yneuron neuron348 in348 0 segParams
R348349 in348 in349 {rInterSeg}
yneuron neuron349 in349 0 segParams
R349350 in349 in350 {rInterSeg}
yneuron neuron350 in350 0 segParams
R350351 in350 in351 {rInterSeg}
yneuron neuron351 in351 0 segParams
R351352 in351 in352 {rInterSeg}
yneuron neuron352 in352 0 segParams
R352353 in352 in353 {rInterSeg}
yneuron neuron353 in353 0 segParams
R353354 in353 in354 {rInterSeg}
yneuron neuron354 in354 0 segParams
R354355 in354 in355 {rInterSeg}
yneuron neuron355 in355 0 segParams
R355356 in355 in356 {rInterSeg}
yneuron neuron356 in356 0 segParams
R356357 in356 in357 {rInterSeg}
yneuron neuron357 in357 0 segParams
R357358 in357 in358 {rInterSeg}
yneuron neuron358 in358 0 segParams
R358359 in358 in359 {rInterSeg}
yneuron neuron359 in359 0 segParams
R359360 in359 in360 {rInterSeg}
yneuron neuron360 in360 0 segParams
R360361 in360 in361 {rInterSeg}
yneuron neuron361 in361 0 segParams
R361362 in361 in362 {rInterSeg}
yneuron neuron362 in362 0 segParams
R362363 in362 in363 {rInterSeg}
yneuron neuron363 in363 0 segParams
R363364 in363 in364 {rInterSeg}
yneuron neuron364 in364 0 segParams
R364365 in364 in365 {rInterSeg}
yneuron neuron365 in365 0 segParams
R365366 in365 in366 {rInterSeg}
yneuron neuron366 in366 0 segParams
R366367 in366 in367 {rInterSeg}
yneuron neuron367 in367 0 segParams
R367368 in367 in368 {rInterSeg}
yneuron neuron368 in368 0 segParams
R368369 in368 in369 {rInterSeg}
yneuron neuron369 in369 0 segParams
R369370 in369 in370 {rInterSeg}
yneuron neuron370 in370 0 segParams
R370371 in370 in371 {rInterSeg}
yneuron neuron371 in371 0 segParams
R371372 in371 in372 {rInterSeg}
yneuron neuron372 in372 0 segParams
R372373 in372 in373 {rInterSeg}
yneuron neuron373 in373 0 segParams
R373374 in373 in374 {rInterSeg}
yneuron neuron374 in374 0 segParams
R374375 in374 in375 {rInterSeg}
yneuron neuron375 in375 0 segParams
R375376 in375 in376 {rInterSeg}
yneuron neuron376 in376 0 segParams
R376377 in376 in377 {rInterSeg}
yneuron neuron377 in377 0 segParams
R377378 in377 in378 {rInterSeg}
yneuron neuron378 in378 0 segParams
R378379 in378 in379 {rInterSeg}
yneuron neuron379 in379 0 segParams
R379380 in379 in380 {rInterSeg}
yneuron neuron380 in380 0 segParams
R380381 in380 in381 {rInterSeg}
yneuron neuron381 in381 0 segParams
R381382 in381 in382 {rInterSeg}
yneuron neuron382 in382 0 segParams
R382383 in382 in383 {rInterSeg}
yneuron neuron383 in383 0 segParams
R383384 in383 in384 {rInterSeg}
yneuron neuron384 in384 0 segParams
R384385 in384 in385 {rInterSeg}
yneuron neuron385 in385 0 segParams
R385386 in385 in386 {rInterSeg}
yneuron neuron386 in386 0 segParams
R386387 in386 in387 {rInterSeg}
yneuron neuron387 in387 0 segParams
R387388 in387 in388 {rInterSeg}
yneuron neuron388 in388 0 segParams
R388389 in388 in389 {rInterSeg}
yneuron neuron389 in389 0 segParams
R389390 in389 in390 {rInterSeg}
yneuron neuron390 in390 0 segParams
R390391 in390 in391 {rInterSeg}
yneuron neuron391 in391 0 segParams
R391392 in391 in392 {rInterSeg}
yneuron neuron392 in392 0 segParams
R392393 in392 in393 {rInterSeg}
yneuron neuron393 in393 0 segParams
R393394 in393 in394 {rInterSeg}
yneuron neuron394 in394 0 segParams
R394395 in394 in395 {rInterSeg}
yneuron neuron395 in395 0 segParams
R395396 in395 in396 {rInterSeg}
yneuron neuron396 in396 0 segParams
R396397 in396 in397 {rInterSeg}
yneuron neuron397 in397 0 segParams
R397398 in397 in398 {rInterSeg}
yneuron neuron398 in398 0 segParams
R398399 in398 in399 {rInterSeg}
yneuron neuron399 in399 0 segParams
R399400 in399 in400 {rInterSeg}
yneuron neuron400 in400 0 segParams
R400401 in400 in401 {rInterSeg}
yneuron neuron401 in401 0 segParams
R401402 in401 in402 {rInterSeg}
yneuron neuron402 in402 0 segParams
R402403 in402 in403 {rInterSeg}
yneuron neuron403 in403 0 segParams
R403404 in403 in404 {rInterSeg}
yneuron neuron404 in404 0 segParams
R404405 in404 in405 {rInterSeg}
yneuron neuron405 in405 0 segParams
R405406 in405 in406 {rInterSeg}
yneuron neuron406 in406 0 segParams
R406407 in406 in407 {rInterSeg}
yneuron neuron407 in407 0 segParams
R407408 in407 in408 {rInterSeg}
yneuron neuron408 in408 0 segParams
R408409 in408 in409 {rInterSeg}
yneuron neuron409 in409 0 segParams
R409410 in409 in410 {rInterSeg}
yneuron neuron410 in410 0 segParams
R410411 in410 in411 {rInterSeg}
yneuron neuron411 in411 0 segParams
R411412 in411 in412 {rInterSeg}
yneuron neuron412 in412 0 segParams
R412413 in412 in413 {rInterSeg}
yneuron neuron413 in413 0 segParams
R413414 in413 in414 {rInterSeg}
yneuron neuron414 in414 0 segParams
R414415 in414 in415 {rInterSeg}
yneuron neuron415 in415 0 segParams
R415416 in415 in416 {rInterSeg}
yneuron neuron416 in416 0 segParams
R416417 in416 in417 {rInterSeg}
yneuron neuron417 in417 0 segParams
R417418 in417 in418 {rInterSeg}
yneuron neuron418 in418 0 segParams
R418419 in418 in419 {rInterSeg}
yneuron neuron419 in419 0 segParams
R419420 in419 in420 {rInterSeg}
yneuron neuron420 in420 0 segParams
R420421 in420 in421 {rInterSeg}
yneuron neuron421 in421 0 segParams
R421422 in421 in422 {rInterSeg}
yneuron neuron422 in422 0 segParams
R422423 in422 in423 {rInterSeg}
yneuron neuron423 in423 0 segParams
R423424 in423 in424 {rInterSeg}
yneuron neuron424 in424 0 segParams
R424425 in424 in425 {rInterSeg}
yneuron neuron425 in425 0 segParams
R425426 in425 in426 {rInterSeg}
yneuron neuron426 in426 0 segParams
R426427 in426 in427 {rInterSeg}
yneuron neuron427 in427 0 segParams
R427428 in427 in428 {rInterSeg}
yneuron neuron428 in428 0 segParams
R428429 in428 in429 {rInterSeg}
yneuron neuron429 in429 0 segParams
R429430 in429 in430 {rInterSeg}
yneuron neuron430 in430 0 segParams
R430431 in430 in431 {rInterSeg}
yneuron neuron431 in431 0 segParams
R431432 in431 in432 {rInterSeg}
yneuron neuron432 in432 0 segParams
R432433 in432 in433 {rInterSeg}
yneuron neuron433 in433 0 segParams
R433434 in433 in434 {rInterSeg}
yneuron neuron434 in434 0 segParams
R434435 in434 in435 {rInterSeg}
yneuron neuron435 in435 0 segParams
R435436 in435 in436 {rInterSeg}
yneuron neuron436 in436 0 segParams
R436437 in436 in437 {rInterSeg}
yneuron neuron437 in437 0 segParams
R437438 in437 in438 {rInterSeg}
yneuron neuron438 in438 0 segParams
R438439 in438 in439 {rInterSeg}
yneuron neuron439 in439 0 segParams
R439440 in439 in440 {rInterSeg}
yneuron neuron440 in440 0 segParams
R440441 in440 in441 {rInterSeg}
yneuron neuron441 in441 0 segParams
R441442 in441 in442 {rInterSeg}
yneuron neuron442 in442 0 segParams
R442443 in442 in443 {rInterSeg}
yneuron neuron443 in443 0 segParams
R443444 in443 in444 {rInterSeg}
yneuron neuron444 in444 0 segParams
R444445 in444 in445 {rInterSeg}
yneuron neuron445 in445 0 segParams
R445446 in445 in446 {rInterSeg}
yneuron neuron446 in446 0 segParams
R446447 in446 in447 {rInterSeg}
yneuron neuron447 in447 0 segParams
R447448 in447 in448 {rInterSeg}
yneuron neuron448 in448 0 segParams
R448449 in448 in449 {rInterSeg}
yneuron neuron449 in449 0 segParams
R449450 in449 in450 {rInterSeg}
yneuron neuron450 in450 0 segParams
R450451 in450 in451 {rInterSeg}
yneuron neuron451 in451 0 segParams
R451452 in451 in452 {rInterSeg}
yneuron neuron452 in452 0 segParams
R452453 in452 in453 {rInterSeg}
yneuron neuron453 in453 0 segParams
R453454 in453 in454 {rInterSeg}
yneuron neuron454 in454 0 segParams
R454455 in454 in455 {rInterSeg}
yneuron neuron455 in455 0 segParams
R455456 in455 in456 {rInterSeg}
yneuron neuron456 in456 0 segParams
R456457 in456 in457 {rInterSeg}
yneuron neuron457 in457 0 segParams
R457458 in457 in458 {rInterSeg}
yneuron neuron458 in458 0 segParams
R458459 in458 in459 {rInterSeg}
yneuron neuron459 in459 0 segParams
R459460 in459 in460 {rInterSeg}
yneuron neuron460 in460 0 segParams
R460461 in460 in461 {rInterSeg}
yneuron neuron461 in461 0 segParams
R461462 in461 in462 {rInterSeg}
yneuron neuron462 in462 0 segParams
R462463 in462 in463 {rInterSeg}
yneuron neuron463 in463 0 segParams
R463464 in463 in464 {rInterSeg}
yneuron neuron464 in464 0 segParams
R464465 in464 in465 {rInterSeg}
yneuron neuron465 in465 0 segParams
R465466 in465 in466 {rInterSeg}
yneuron neuron466 in466 0 segParams
R466467 in466 in467 {rInterSeg}
yneuron neuron467 in467 0 segParams
R467468 in467 in468 {rInterSeg}
yneuron neuron468 in468 0 segParams
R468469 in468 in469 {rInterSeg}
yneuron neuron469 in469 0 segParams
R469470 in469 in470 {rInterSeg}
yneuron neuron470 in470 0 segParams
R470471 in470 in471 {rInterSeg}
yneuron neuron471 in471 0 segParams
R471472 in471 in472 {rInterSeg}
yneuron neuron472 in472 0 segParams
R472473 in472 in473 {rInterSeg}
yneuron neuron473 in473 0 segParams
R473474 in473 in474 {rInterSeg}
yneuron neuron474 in474 0 segParams
R474475 in474 in475 {rInterSeg}
yneuron neuron475 in475 0 segParams
R475476 in475 in476 {rInterSeg}
yneuron neuron476 in476 0 segParams
R476477 in476 in477 {rInterSeg}
yneuron neuron477 in477 0 segParams
R477478 in477 in478 {rInterSeg}
yneuron neuron478 in478 0 segParams
R478479 in478 in479 {rInterSeg}
yneuron neuron479 in479 0 segParams
R479480 in479 in480 {rInterSeg}
yneuron neuron480 in480 0 segParams
R480481 in480 in481 {rInterSeg}
yneuron neuron481 in481 0 segParams
R481482 in481 in482 {rInterSeg}
yneuron neuron482 in482 0 segParams
R482483 in482 in483 {rInterSeg}
yneuron neuron483 in483 0 segParams
R483484 in483 in484 {rInterSeg}
yneuron neuron484 in484 0 segParams
R484485 in484 in485 {rInterSeg}
yneuron neuron485 in485 0 segParams
R485486 in485 in486 {rInterSeg}
yneuron neuron486 in486 0 segParams
R486487 in486 in487 {rInterSeg}
yneuron neuron487 in487 0 segParams
R487488 in487 in488 {rInterSeg}
yneuron neuron488 in488 0 segParams
R488489 in488 in489 {rInterSeg}
yneuron neuron489 in489 0 segParams
R489490 in489 in490 {rInterSeg}
yneuron neuron490 in490 0 segParams
R490491 in490 in491 {rInterSeg}
yneuron neuron491 in491 0 segParams
R491492 in491 in492 {rInterSeg}
yneuron neuron492 in492 0 segParams
R492493 in492 in493 {rInterSeg}
yneuron neuron493 in493 0 segParams
R493494 in493 in494 {rInterSeg}
yneuron neuron494 in494 0 segParams
R494495 in494 in495 {rInterSeg}
yneuron neuron495 in495 0 segParams
R495496 in495 in496 {rInterSeg}
yneuron neuron496 in496 0 segParams
R496497 in496 in497 {rInterSeg}
yneuron neuron497 in497 0 segParams
R497498 in497 in498 {rInterSeg}
yneuron neuron498 in498 0 segParams
R498499 in498 in499 {rInterSeg}
yneuron neuron499 in499 0 segParams
R499500 in499 in500 {rInterSeg}
yneuron neuron500 in500 0 segParams
R500501 in500 in501 {rInterSeg}
yneuron neuron501 in501 0 segParams
R501502 in501 in502 {rInterSeg}
yneuron neuron502 in502 0 segParams
R502503 in502 in503 {rInterSeg}
yneuron neuron503 in503 0 segParams
R503504 in503 in504 {rInterSeg}
yneuron neuron504 in504 0 segParams
R504505 in504 in505 {rInterSeg}
yneuron neuron505 in505 0 segParams
R505506 in505 in506 {rInterSeg}
yneuron neuron506 in506 0 segParams
R506507 in506 in507 {rInterSeg}
yneuron neuron507 in507 0 segParams
R507508 in507 in508 {rInterSeg}
yneuron neuron508 in508 0 segParams
R508509 in508 in509 {rInterSeg}
yneuron neuron509 in509 0 segParams
R509510 in509 in510 {rInterSeg}
yneuron neuron510 in510 0 segParams
R510511 in510 in511 {rInterSeg}
yneuron neuron511 in511 0 segParams
R511512 in511 in512 {rInterSeg}
yneuron neuron512 in512 0 segParams
R512513 in512 in513 {rInterSeg}
yneuron neuron513 in513 0 segParams
R513514 in513 in514 {rInterSeg}
yneuron neuron514 in514 0 segParams
R514515 in514 in515 {rInterSeg}
yneuron neuron515 in515 0 segParams
R515516 in515 in516 {rInterSeg}
yneuron neuron516 in516 0 segParams
R516517 in516 in517 {rInterSeg}
yneuron neuron517 in517 0 segParams
R517518 in517 in518 {rInterSeg}
yneuron neuron518 in518 0 segParams
R518519 in518 in519 {rInterSeg}
yneuron neuron519 in519 0 segParams
R519520 in519 in520 {rInterSeg}
yneuron neuron520 in520 0 segParams
R520521 in520 in521 {rInterSeg}
yneuron neuron521 in521 0 segParams
R521522 in521 in522 {rInterSeg}
yneuron neuron522 in522 0 segParams
R522523 in522 in523 {rInterSeg}
yneuron neuron523 in523 0 segParams
R523524 in523 in524 {rInterSeg}
yneuron neuron524 in524 0 segParams
R524525 in524 in525 {rInterSeg}
yneuron neuron525 in525 0 segParams
R525526 in525 in526 {rInterSeg}
yneuron neuron526 in526 0 segParams
R526527 in526 in527 {rInterSeg}
yneuron neuron527 in527 0 segParams
R527528 in527 in528 {rInterSeg}
yneuron neuron528 in528 0 segParams
R528529 in528 in529 {rInterSeg}
yneuron neuron529 in529 0 segParams
R529530 in529 in530 {rInterSeg}
yneuron neuron530 in530 0 segParams
R530531 in530 in531 {rInterSeg}
yneuron neuron531 in531 0 segParams
R531532 in531 in532 {rInterSeg}
yneuron neuron532 in532 0 segParams
R532533 in532 in533 {rInterSeg}
yneuron neuron533 in533 0 segParams
R533534 in533 in534 {rInterSeg}
yneuron neuron534 in534 0 segParams
R534535 in534 in535 {rInterSeg}
yneuron neuron535 in535 0 segParams
R535536 in535 in536 {rInterSeg}
yneuron neuron536 in536 0 segParams
R536537 in536 in537 {rInterSeg}
yneuron neuron537 in537 0 segParams
R537538 in537 in538 {rInterSeg}
yneuron neuron538 in538 0 segParams
R538539 in538 in539 {rInterSeg}
yneuron neuron539 in539 0 segParams
R539540 in539 in540 {rInterSeg}
yneuron neuron540 in540 0 segParams
R540541 in540 in541 {rInterSeg}
yneuron neuron541 in541 0 segParams
R541542 in541 in542 {rInterSeg}
yneuron neuron542 in542 0 segParams
R542543 in542 in543 {rInterSeg}
yneuron neuron543 in543 0 segParams
R543544 in543 in544 {rInterSeg}
yneuron neuron544 in544 0 segParams
R544545 in544 in545 {rInterSeg}
yneuron neuron545 in545 0 segParams
R545546 in545 in546 {rInterSeg}
yneuron neuron546 in546 0 segParams
R546547 in546 in547 {rInterSeg}
yneuron neuron547 in547 0 segParams
R547548 in547 in548 {rInterSeg}
yneuron neuron548 in548 0 segParams
R548549 in548 in549 {rInterSeg}
yneuron neuron549 in549 0 segParams
R549550 in549 in550 {rInterSeg}
yneuron neuron550 in550 0 segParams
R550551 in550 in551 {rInterSeg}
yneuron neuron551 in551 0 segParams
R551552 in551 in552 {rInterSeg}
yneuron neuron552 in552 0 segParams
R552553 in552 in553 {rInterSeg}
yneuron neuron553 in553 0 segParams
R553554 in553 in554 {rInterSeg}
yneuron neuron554 in554 0 segParams
R554555 in554 in555 {rInterSeg}
yneuron neuron555 in555 0 segParams
R555556 in555 in556 {rInterSeg}
yneuron neuron556 in556 0 segParams
R556557 in556 in557 {rInterSeg}
yneuron neuron557 in557 0 segParams
R557558 in557 in558 {rInterSeg}
yneuron neuron558 in558 0 segParams
R558559 in558 in559 {rInterSeg}
yneuron neuron559 in559 0 segParams
R559560 in559 in560 {rInterSeg}
yneuron neuron560 in560 0 segParams
R560561 in560 in561 {rInterSeg}
yneuron neuron561 in561 0 segParams
R561562 in561 in562 {rInterSeg}
yneuron neuron562 in562 0 segParams
R562563 in562 in563 {rInterSeg}
yneuron neuron563 in563 0 segParams
R563564 in563 in564 {rInterSeg}
yneuron neuron564 in564 0 segParams
R564565 in564 in565 {rInterSeg}
yneuron neuron565 in565 0 segParams
R565566 in565 in566 {rInterSeg}
yneuron neuron566 in566 0 segParams
R566567 in566 in567 {rInterSeg}
yneuron neuron567 in567 0 segParams
R567568 in567 in568 {rInterSeg}
yneuron neuron568 in568 0 segParams
R568569 in568 in569 {rInterSeg}
yneuron neuron569 in569 0 segParams
R569570 in569 in570 {rInterSeg}
yneuron neuron570 in570 0 segParams
R570571 in570 in571 {rInterSeg}
yneuron neuron571 in571 0 segParams
R571572 in571 in572 {rInterSeg}
yneuron neuron572 in572 0 segParams
R572573 in572 in573 {rInterSeg}
yneuron neuron573 in573 0 segParams
R573574 in573 in574 {rInterSeg}
yneuron neuron574 in574 0 segParams
R574575 in574 in575 {rInterSeg}
yneuron neuron575 in575 0 segParams
R575576 in575 in576 {rInterSeg}
yneuron neuron576 in576 0 segParams
R576577 in576 in577 {rInterSeg}
yneuron neuron577 in577 0 segParams
R577578 in577 in578 {rInterSeg}
yneuron neuron578 in578 0 segParams
R578579 in578 in579 {rInterSeg}
yneuron neuron579 in579 0 segParams
R579580 in579 in580 {rInterSeg}
yneuron neuron580 in580 0 segParams
R580581 in580 in581 {rInterSeg}
yneuron neuron581 in581 0 segParams
R581582 in581 in582 {rInterSeg}
yneuron neuron582 in582 0 segParams
R582583 in582 in583 {rInterSeg}
yneuron neuron583 in583 0 segParams
R583584 in583 in584 {rInterSeg}
yneuron neuron584 in584 0 segParams
R584585 in584 in585 {rInterSeg}
yneuron neuron585 in585 0 segParams
R585586 in585 in586 {rInterSeg}
yneuron neuron586 in586 0 segParams
R586587 in586 in587 {rInterSeg}
yneuron neuron587 in587 0 segParams
R587588 in587 in588 {rInterSeg}
yneuron neuron588 in588 0 segParams
R588589 in588 in589 {rInterSeg}
yneuron neuron589 in589 0 segParams
R589590 in589 in590 {rInterSeg}
yneuron neuron590 in590 0 segParams
R590591 in590 in591 {rInterSeg}
yneuron neuron591 in591 0 segParams
R591592 in591 in592 {rInterSeg}
yneuron neuron592 in592 0 segParams
R592593 in592 in593 {rInterSeg}
yneuron neuron593 in593 0 segParams
R593594 in593 in594 {rInterSeg}
yneuron neuron594 in594 0 segParams
R594595 in594 in595 {rInterSeg}
yneuron neuron595 in595 0 segParams
R595596 in595 in596 {rInterSeg}
yneuron neuron596 in596 0 segParams
R596597 in596 in597 {rInterSeg}
yneuron neuron597 in597 0 segParams
R597598 in597 in598 {rInterSeg}
yneuron neuron598 in598 0 segParams
R598599 in598 in599 {rInterSeg}
yneuron neuron599 in599 0 segParams
R599600 in599 in600 {rInterSeg}
yneuron neuron600 in600 0 segParams
R600601 in600 in601 {rInterSeg}
yneuron neuron601 in601 0 segParams
R601602 in601 in602 {rInterSeg}
yneuron neuron602 in602 0 segParams
R602603 in602 in603 {rInterSeg}
yneuron neuron603 in603 0 segParams
R603604 in603 in604 {rInterSeg}
yneuron neuron604 in604 0 segParams
R604605 in604 in605 {rInterSeg}
yneuron neuron605 in605 0 segParams
R605606 in605 in606 {rInterSeg}
yneuron neuron606 in606 0 segParams
R606607 in606 in607 {rInterSeg}
yneuron neuron607 in607 0 segParams
R607608 in607 in608 {rInterSeg}
yneuron neuron608 in608 0 segParams
R608609 in608 in609 {rInterSeg}
yneuron neuron609 in609 0 segParams
R609610 in609 in610 {rInterSeg}
yneuron neuron610 in610 0 segParams
R610611 in610 in611 {rInterSeg}
yneuron neuron611 in611 0 segParams
R611612 in611 in612 {rInterSeg}
yneuron neuron612 in612 0 segParams
R612613 in612 in613 {rInterSeg}
yneuron neuron613 in613 0 segParams
R613614 in613 in614 {rInterSeg}
yneuron neuron614 in614 0 segParams
R614615 in614 in615 {rInterSeg}
yneuron neuron615 in615 0 segParams
R615616 in615 in616 {rInterSeg}
yneuron neuron616 in616 0 segParams
R616617 in616 in617 {rInterSeg}
yneuron neuron617 in617 0 segParams
R617618 in617 in618 {rInterSeg}
yneuron neuron618 in618 0 segParams
R618619 in618 in619 {rInterSeg}
yneuron neuron619 in619 0 segParams
R619620 in619 in620 {rInterSeg}
yneuron neuron620 in620 0 segParams
R620621 in620 in621 {rInterSeg}
yneuron neuron621 in621 0 segParams
R621622 in621 in622 {rInterSeg}
yneuron neuron622 in622 0 segParams
R622623 in622 in623 {rInterSeg}
yneuron neuron623 in623 0 segParams
R623624 in623 in624 {rInterSeg}
yneuron neuron624 in624 0 segParams
R624625 in624 in625 {rInterSeg}
yneuron neuron625 in625 0 segParams
R625626 in625 in626 {rInterSeg}
yneuron neuron626 in626 0 segParams
R626627 in626 in627 {rInterSeg}
yneuron neuron627 in627 0 segParams
R627628 in627 in628 {rInterSeg}
yneuron neuron628 in628 0 segParams
R628629 in628 in629 {rInterSeg}
yneuron neuron629 in629 0 segParams
R629630 in629 in630 {rInterSeg}
yneuron neuron630 in630 0 segParams
R630631 in630 in631 {rInterSeg}
yneuron neuron631 in631 0 segParams
R631632 in631 in632 {rInterSeg}
yneuron neuron632 in632 0 segParams
R632633 in632 in633 {rInterSeg}
yneuron neuron633 in633 0 segParams
R633634 in633 in634 {rInterSeg}
yneuron neuron634 in634 0 segParams
R634635 in634 in635 {rInterSeg}
yneuron neuron635 in635 0 segParams
R635636 in635 in636 {rInterSeg}
yneuron neuron636 in636 0 segParams
R636637 in636 in637 {rInterSeg}
yneuron neuron637 in637 0 segParams
R637638 in637 in638 {rInterSeg}
yneuron neuron638 in638 0 segParams
R638639 in638 in639 {rInterSeg}
yneuron neuron639 in639 0 segParams
R639640 in639 in640 {rInterSeg}
yneuron neuron640 in640 0 segParams
R640641 in640 in641 {rInterSeg}
yneuron neuron641 in641 0 segParams
R641642 in641 in642 {rInterSeg}
yneuron neuron642 in642 0 segParams
R642643 in642 in643 {rInterSeg}
yneuron neuron643 in643 0 segParams
R643644 in643 in644 {rInterSeg}
yneuron neuron644 in644 0 segParams
R644645 in644 in645 {rInterSeg}
yneuron neuron645 in645 0 segParams
R645646 in645 in646 {rInterSeg}
yneuron neuron646 in646 0 segParams
R646647 in646 in647 {rInterSeg}
yneuron neuron647 in647 0 segParams
R647648 in647 in648 {rInterSeg}
yneuron neuron648 in648 0 segParams
R648649 in648 in649 {rInterSeg}
yneuron neuron649 in649 0 segParams
R649650 in649 in650 {rInterSeg}
yneuron neuron650 in650 0 segParams
R650651 in650 in651 {rInterSeg}
yneuron neuron651 in651 0 segParams
R651652 in651 in652 {rInterSeg}
yneuron neuron652 in652 0 segParams
R652653 in652 in653 {rInterSeg}
yneuron neuron653 in653 0 segParams
R653654 in653 in654 {rInterSeg}
yneuron neuron654 in654 0 segParams
R654655 in654 in655 {rInterSeg}
yneuron neuron655 in655 0 segParams
R655656 in655 in656 {rInterSeg}
yneuron neuron656 in656 0 segParams
R656657 in656 in657 {rInterSeg}
yneuron neuron657 in657 0 segParams
R657658 in657 in658 {rInterSeg}
yneuron neuron658 in658 0 segParams
R658659 in658 in659 {rInterSeg}
yneuron neuron659 in659 0 segParams
R659660 in659 in660 {rInterSeg}
yneuron neuron660 in660 0 segParams
R660661 in660 in661 {rInterSeg}
yneuron neuron661 in661 0 segParams
R661662 in661 in662 {rInterSeg}
yneuron neuron662 in662 0 segParams
R662663 in662 in663 {rInterSeg}
yneuron neuron663 in663 0 segParams
R663664 in663 in664 {rInterSeg}
yneuron neuron664 in664 0 segParams
R664665 in664 in665 {rInterSeg}
yneuron neuron665 in665 0 segParams
R665666 in665 in666 {rInterSeg}
yneuron neuron666 in666 0 segParams
R666667 in666 in667 {rInterSeg}
yneuron neuron667 in667 0 segParams
R667668 in667 in668 {rInterSeg}
yneuron neuron668 in668 0 segParams
R668669 in668 in669 {rInterSeg}
yneuron neuron669 in669 0 segParams
R669670 in669 in670 {rInterSeg}
yneuron neuron670 in670 0 segParams
R670671 in670 in671 {rInterSeg}
yneuron neuron671 in671 0 segParams
R671672 in671 in672 {rInterSeg}
yneuron neuron672 in672 0 segParams
R672673 in672 in673 {rInterSeg}
yneuron neuron673 in673 0 segParams
R673674 in673 in674 {rInterSeg}
yneuron neuron674 in674 0 segParams
R674675 in674 in675 {rInterSeg}
yneuron neuron675 in675 0 segParams
R675676 in675 in676 {rInterSeg}
yneuron neuron676 in676 0 segParams
R676677 in676 in677 {rInterSeg}
yneuron neuron677 in677 0 segParams
R677678 in677 in678 {rInterSeg}
yneuron neuron678 in678 0 segParams
R678679 in678 in679 {rInterSeg}
yneuron neuron679 in679 0 segParams
R679680 in679 in680 {rInterSeg}
yneuron neuron680 in680 0 segParams
R680681 in680 in681 {rInterSeg}
yneuron neuron681 in681 0 segParams
R681682 in681 in682 {rInterSeg}
yneuron neuron682 in682 0 segParams
R682683 in682 in683 {rInterSeg}
yneuron neuron683 in683 0 segParams
R683684 in683 in684 {rInterSeg}
yneuron neuron684 in684 0 segParams
R684685 in684 in685 {rInterSeg}
yneuron neuron685 in685 0 segParams
R685686 in685 in686 {rInterSeg}
yneuron neuron686 in686 0 segParams
R686687 in686 in687 {rInterSeg}
yneuron neuron687 in687 0 segParams
R687688 in687 in688 {rInterSeg}
yneuron neuron688 in688 0 segParams
R688689 in688 in689 {rInterSeg}
yneuron neuron689 in689 0 segParams
R689690 in689 in690 {rInterSeg}
yneuron neuron690 in690 0 segParams
R690691 in690 in691 {rInterSeg}
yneuron neuron691 in691 0 segParams
R691692 in691 in692 {rInterSeg}
yneuron neuron692 in692 0 segParams
R692693 in692 in693 {rInterSeg}
yneuron neuron693 in693 0 segParams
R693694 in693 in694 {rInterSeg}
yneuron neuron694 in694 0 segParams
R694695 in694 in695 {rInterSeg}
yneuron neuron695 in695 0 segParams
R695696 in695 in696 {rInterSeg}
yneuron neuron696 in696 0 segParams
R696697 in696 in697 {rInterSeg}
yneuron neuron697 in697 0 segParams
R697698 in697 in698 {rInterSeg}
yneuron neuron698 in698 0 segParams
R698699 in698 in699 {rInterSeg}
yneuron neuron699 in699 0 segParams
R699700 in699 in700 {rInterSeg}
yneuron neuron700 in700 0 segParams
R700701 in700 in701 {rInterSeg}
yneuron neuron701 in701 0 segParams
R701702 in701 in702 {rInterSeg}
yneuron neuron702 in702 0 segParams
R702703 in702 in703 {rInterSeg}
yneuron neuron703 in703 0 segParams
R703704 in703 in704 {rInterSeg}
yneuron neuron704 in704 0 segParams
R704705 in704 in705 {rInterSeg}
yneuron neuron705 in705 0 segParams
R705706 in705 in706 {rInterSeg}
yneuron neuron706 in706 0 segParams
R706707 in706 in707 {rInterSeg}
yneuron neuron707 in707 0 segParams
R707708 in707 in708 {rInterSeg}
yneuron neuron708 in708 0 segParams
R708709 in708 in709 {rInterSeg}
yneuron neuron709 in709 0 segParams
R709710 in709 in710 {rInterSeg}
yneuron neuron710 in710 0 segParams
R710711 in710 in711 {rInterSeg}
yneuron neuron711 in711 0 segParams
R711712 in711 in712 {rInterSeg}
yneuron neuron712 in712 0 segParams
R712713 in712 in713 {rInterSeg}
yneuron neuron713 in713 0 segParams
R713714 in713 in714 {rInterSeg}
yneuron neuron714 in714 0 segParams
R714715 in714 in715 {rInterSeg}
yneuron neuron715 in715 0 segParams
R715716 in715 in716 {rInterSeg}
yneuron neuron716 in716 0 segParams
R716717 in716 in717 {rInterSeg}
yneuron neuron717 in717 0 segParams
R717718 in717 in718 {rInterSeg}
yneuron neuron718 in718 0 segParams
R718719 in718 in719 {rInterSeg}
yneuron neuron719 in719 0 segParams
R719720 in719 in720 {rInterSeg}
yneuron neuron720 in720 0 segParams
R720721 in720 in721 {rInterSeg}
yneuron neuron721 in721 0 segParams
R721722 in721 in722 {rInterSeg}
yneuron neuron722 in722 0 segParams
R722723 in722 in723 {rInterSeg}
yneuron neuron723 in723 0 segParams
R723724 in723 in724 {rInterSeg}
yneuron neuron724 in724 0 segParams
R724725 in724 in725 {rInterSeg}
yneuron neuron725 in725 0 segParams
R725726 in725 in726 {rInterSeg}
yneuron neuron726 in726 0 segParams
R726727 in726 in727 {rInterSeg}
yneuron neuron727 in727 0 segParams
R727728 in727 in728 {rInterSeg}
yneuron neuron728 in728 0 segParams
R728729 in728 in729 {rInterSeg}
yneuron neuron729 in729 0 segParams
R729730 in729 in730 {rInterSeg}
yneuron neuron730 in730 0 segParams
R730731 in730 in731 {rInterSeg}
yneuron neuron731 in731 0 segParams
R731732 in731 in732 {rInterSeg}
yneuron neuron732 in732 0 segParams
R732733 in732 in733 {rInterSeg}
yneuron neuron733 in733 0 segParams
R733734 in733 in734 {rInterSeg}
yneuron neuron734 in734 0 segParams
R734735 in734 in735 {rInterSeg}
yneuron neuron735 in735 0 segParams
R735736 in735 in736 {rInterSeg}
yneuron neuron736 in736 0 segParams
R736737 in736 in737 {rInterSeg}
yneuron neuron737 in737 0 segParams
R737738 in737 in738 {rInterSeg}
yneuron neuron738 in738 0 segParams
R738739 in738 in739 {rInterSeg}
yneuron neuron739 in739 0 segParams
R739740 in739 in740 {rInterSeg}
yneuron neuron740 in740 0 segParams
R740741 in740 in741 {rInterSeg}
yneuron neuron741 in741 0 segParams
R741742 in741 in742 {rInterSeg}
yneuron neuron742 in742 0 segParams
R742743 in742 in743 {rInterSeg}
yneuron neuron743 in743 0 segParams
R743744 in743 in744 {rInterSeg}
yneuron neuron744 in744 0 segParams
R744745 in744 in745 {rInterSeg}
yneuron neuron745 in745 0 segParams
R745746 in745 in746 {rInterSeg}
yneuron neuron746 in746 0 segParams
R746747 in746 in747 {rInterSeg}
yneuron neuron747 in747 0 segParams
R747748 in747 in748 {rInterSeg}
yneuron neuron748 in748 0 segParams
R748749 in748 in749 {rInterSeg}
yneuron neuron749 in749 0 segParams
R749750 in749 in750 {rInterSeg}
yneuron neuron750 in750 0 segParams
R750751 in750 in751 {rInterSeg}
yneuron neuron751 in751 0 segParams
R751752 in751 in752 {rInterSeg}
yneuron neuron752 in752 0 segParams
R752753 in752 in753 {rInterSeg}
yneuron neuron753 in753 0 segParams
R753754 in753 in754 {rInterSeg}
yneuron neuron754 in754 0 segParams
R754755 in754 in755 {rInterSeg}
yneuron neuron755 in755 0 segParams
R755756 in755 in756 {rInterSeg}
yneuron neuron756 in756 0 segParams
R756757 in756 in757 {rInterSeg}
yneuron neuron757 in757 0 segParams
R757758 in757 in758 {rInterSeg}
yneuron neuron758 in758 0 segParams
R758759 in758 in759 {rInterSeg}
yneuron neuron759 in759 0 segParams
R759760 in759 in760 {rInterSeg}
yneuron neuron760 in760 0 segParams
R760761 in760 in761 {rInterSeg}
yneuron neuron761 in761 0 segParams
R761762 in761 in762 {rInterSeg}
yneuron neuron762 in762 0 segParams
R762763 in762 in763 {rInterSeg}
yneuron neuron763 in763 0 segParams
R763764 in763 in764 {rInterSeg}
yneuron neuron764 in764 0 segParams
R764765 in764 in765 {rInterSeg}
yneuron neuron765 in765 0 segParams
R765766 in765 in766 {rInterSeg}
yneuron neuron766 in766 0 segParams
R766767 in766 in767 {rInterSeg}
yneuron neuron767 in767 0 segParams
R767768 in767 in768 {rInterSeg}
yneuron neuron768 in768 0 segParams
R768769 in768 in769 {rInterSeg}
yneuron neuron769 in769 0 segParams
R769770 in769 in770 {rInterSeg}
yneuron neuron770 in770 0 segParams
R770771 in770 in771 {rInterSeg}
yneuron neuron771 in771 0 segParams
R771772 in771 in772 {rInterSeg}
yneuron neuron772 in772 0 segParams
R772773 in772 in773 {rInterSeg}
yneuron neuron773 in773 0 segParams
R773774 in773 in774 {rInterSeg}
yneuron neuron774 in774 0 segParams
R774775 in774 in775 {rInterSeg}
yneuron neuron775 in775 0 segParams
R775776 in775 in776 {rInterSeg}
yneuron neuron776 in776 0 segParams
R776777 in776 in777 {rInterSeg}
yneuron neuron777 in777 0 segParams
R777778 in777 in778 {rInterSeg}
yneuron neuron778 in778 0 segParams
R778779 in778 in779 {rInterSeg}
yneuron neuron779 in779 0 segParams
R779780 in779 in780 {rInterSeg}
yneuron neuron780 in780 0 segParams
R780781 in780 in781 {rInterSeg}
yneuron neuron781 in781 0 segParams
R781782 in781 in782 {rInterSeg}
yneuron neuron782 in782 0 segParams
R782783 in782 in783 {rInterSeg}
yneuron neuron783 in783 0 segParams
R783784 in783 in784 {rInterSeg}
yneuron neuron784 in784 0 segParams
R784785 in784 in785 {rInterSeg}
yneuron neuron785 in785 0 segParams
R785786 in785 in786 {rInterSeg}
yneuron neuron786 in786 0 segParams
R786787 in786 in787 {rInterSeg}
yneuron neuron787 in787 0 segParams
R787788 in787 in788 {rInterSeg}
yneuron neuron788 in788 0 segParams
R788789 in788 in789 {rInterSeg}
yneuron neuron789 in789 0 segParams
R789790 in789 in790 {rInterSeg}
yneuron neuron790 in790 0 segParams
R790791 in790 in791 {rInterSeg}
yneuron neuron791 in791 0 segParams
R791792 in791 in792 {rInterSeg}
yneuron neuron792 in792 0 segParams
R792793 in792 in793 {rInterSeg}
yneuron neuron793 in793 0 segParams
R793794 in793 in794 {rInterSeg}
yneuron neuron794 in794 0 segParams
R794795 in794 in795 {rInterSeg}
yneuron neuron795 in795 0 segParams
R795796 in795 in796 {rInterSeg}
yneuron neuron796 in796 0 segParams
R796797 in796 in797 {rInterSeg}
yneuron neuron797 in797 0 segParams
R797798 in797 in798 {rInterSeg}
yneuron neuron798 in798 0 segParams
R798799 in798 in799 {rInterSeg}
yneuron neuron799 in799 0 segParams
R799800 in799 in800 {rInterSeg}
yneuron neuron800 in800 0 segParams
R800801 in800 in801 {rInterSeg}
yneuron neuron801 in801 0 segParams
R801802 in801 in802 {rInterSeg}
yneuron neuron802 in802 0 segParams
R802803 in802 in803 {rInterSeg}
yneuron neuron803 in803 0 segParams
R803804 in803 in804 {rInterSeg}
yneuron neuron804 in804 0 segParams
R804805 in804 in805 {rInterSeg}
yneuron neuron805 in805 0 segParams
R805806 in805 in806 {rInterSeg}
yneuron neuron806 in806 0 segParams
R806807 in806 in807 {rInterSeg}
yneuron neuron807 in807 0 segParams
R807808 in807 in808 {rInterSeg}
yneuron neuron808 in808 0 segParams
R808809 in808 in809 {rInterSeg}
yneuron neuron809 in809 0 segParams
R809810 in809 in810 {rInterSeg}
yneuron neuron810 in810 0 segParams
R810811 in810 in811 {rInterSeg}
yneuron neuron811 in811 0 segParams
R811812 in811 in812 {rInterSeg}
yneuron neuron812 in812 0 segParams
R812813 in812 in813 {rInterSeg}
yneuron neuron813 in813 0 segParams
R813814 in813 in814 {rInterSeg}
yneuron neuron814 in814 0 segParams
R814815 in814 in815 {rInterSeg}
yneuron neuron815 in815 0 segParams
R815816 in815 in816 {rInterSeg}
yneuron neuron816 in816 0 segParams
R816817 in816 in817 {rInterSeg}
yneuron neuron817 in817 0 segParams
R817818 in817 in818 {rInterSeg}
yneuron neuron818 in818 0 segParams
R818819 in818 in819 {rInterSeg}
yneuron neuron819 in819 0 segParams
R819820 in819 in820 {rInterSeg}
yneuron neuron820 in820 0 segParams
R820821 in820 in821 {rInterSeg}
yneuron neuron821 in821 0 segParams
R821822 in821 in822 {rInterSeg}
yneuron neuron822 in822 0 segParams
R822823 in822 in823 {rInterSeg}
yneuron neuron823 in823 0 segParams
R823824 in823 in824 {rInterSeg}
yneuron neuron824 in824 0 segParams
R824825 in824 in825 {rInterSeg}
yneuron neuron825 in825 0 segParams
R825826 in825 in826 {rInterSeg}
yneuron neuron826 in826 0 segParams
R826827 in826 in827 {rInterSeg}
yneuron neuron827 in827 0 segParams
R827828 in827 in828 {rInterSeg}
yneuron neuron828 in828 0 segParams
R828829 in828 in829 {rInterSeg}
yneuron neuron829 in829 0 segParams
R829830 in829 in830 {rInterSeg}
yneuron neuron830 in830 0 segParams
R830831 in830 in831 {rInterSeg}
yneuron neuron831 in831 0 segParams
R831832 in831 in832 {rInterSeg}
yneuron neuron832 in832 0 segParams
R832833 in832 in833 {rInterSeg}
yneuron neuron833 in833 0 segParams
R833834 in833 in834 {rInterSeg}
yneuron neuron834 in834 0 segParams
R834835 in834 in835 {rInterSeg}
yneuron neuron835 in835 0 segParams
R835836 in835 in836 {rInterSeg}
yneuron neuron836 in836 0 segParams
R836837 in836 in837 {rInterSeg}
yneuron neuron837 in837 0 segParams
R837838 in837 in838 {rInterSeg}
yneuron neuron838 in838 0 segParams
R838839 in838 in839 {rInterSeg}
yneuron neuron839 in839 0 segParams
R839840 in839 in840 {rInterSeg}
yneuron neuron840 in840 0 segParams
R840841 in840 in841 {rInterSeg}
yneuron neuron841 in841 0 segParams
R841842 in841 in842 {rInterSeg}
yneuron neuron842 in842 0 segParams
R842843 in842 in843 {rInterSeg}
yneuron neuron843 in843 0 segParams
R843844 in843 in844 {rInterSeg}
yneuron neuron844 in844 0 segParams
R844845 in844 in845 {rInterSeg}
yneuron neuron845 in845 0 segParams
R845846 in845 in846 {rInterSeg}
yneuron neuron846 in846 0 segParams
R846847 in846 in847 {rInterSeg}
yneuron neuron847 in847 0 segParams
R847848 in847 in848 {rInterSeg}
yneuron neuron848 in848 0 segParams
R848849 in848 in849 {rInterSeg}
yneuron neuron849 in849 0 segParams
R849850 in849 in850 {rInterSeg}
yneuron neuron850 in850 0 segParams
R850851 in850 in851 {rInterSeg}
yneuron neuron851 in851 0 segParams
R851852 in851 in852 {rInterSeg}
yneuron neuron852 in852 0 segParams
R852853 in852 in853 {rInterSeg}
yneuron neuron853 in853 0 segParams
R853854 in853 in854 {rInterSeg}
yneuron neuron854 in854 0 segParams
R854855 in854 in855 {rInterSeg}
yneuron neuron855 in855 0 segParams
R855856 in855 in856 {rInterSeg}
yneuron neuron856 in856 0 segParams
R856857 in856 in857 {rInterSeg}
yneuron neuron857 in857 0 segParams
R857858 in857 in858 {rInterSeg}
yneuron neuron858 in858 0 segParams
R858859 in858 in859 {rInterSeg}
yneuron neuron859 in859 0 segParams
R859860 in859 in860 {rInterSeg}
yneuron neuron860 in860 0 segParams
R860861 in860 in861 {rInterSeg}
yneuron neuron861 in861 0 segParams
R861862 in861 in862 {rInterSeg}
yneuron neuron862 in862 0 segParams
R862863 in862 in863 {rInterSeg}
yneuron neuron863 in863 0 segParams
R863864 in863 in864 {rInterSeg}
yneuron neuron864 in864 0 segParams
R864865 in864 in865 {rInterSeg}
yneuron neuron865 in865 0 segParams
R865866 in865 in866 {rInterSeg}
yneuron neuron866 in866 0 segParams
R866867 in866 in867 {rInterSeg}
yneuron neuron867 in867 0 segParams
R867868 in867 in868 {rInterSeg}
yneuron neuron868 in868 0 segParams
R868869 in868 in869 {rInterSeg}
yneuron neuron869 in869 0 segParams
R869870 in869 in870 {rInterSeg}
yneuron neuron870 in870 0 segParams
R870871 in870 in871 {rInterSeg}
yneuron neuron871 in871 0 segParams
R871872 in871 in872 {rInterSeg}
yneuron neuron872 in872 0 segParams
R872873 in872 in873 {rInterSeg}
yneuron neuron873 in873 0 segParams
R873874 in873 in874 {rInterSeg}
yneuron neuron874 in874 0 segParams
R874875 in874 in875 {rInterSeg}
yneuron neuron875 in875 0 segParams
R875876 in875 in876 {rInterSeg}
yneuron neuron876 in876 0 segParams
R876877 in876 in877 {rInterSeg}
yneuron neuron877 in877 0 segParams
R877878 in877 in878 {rInterSeg}
yneuron neuron878 in878 0 segParams
R878879 in878 in879 {rInterSeg}
yneuron neuron879 in879 0 segParams
R879880 in879 in880 {rInterSeg}
yneuron neuron880 in880 0 segParams
R880881 in880 in881 {rInterSeg}
yneuron neuron881 in881 0 segParams
R881882 in881 in882 {rInterSeg}
yneuron neuron882 in882 0 segParams
R882883 in882 in883 {rInterSeg}
yneuron neuron883 in883 0 segParams
R883884 in883 in884 {rInterSeg}
yneuron neuron884 in884 0 segParams
R884885 in884 in885 {rInterSeg}
yneuron neuron885 in885 0 segParams
R885886 in885 in886 {rInterSeg}
yneuron neuron886 in886 0 segParams
R886887 in886 in887 {rInterSeg}
yneuron neuron887 in887 0 segParams
R887888 in887 in888 {rInterSeg}
yneuron neuron888 in888 0 segParams
R888889 in888 in889 {rInterSeg}
yneuron neuron889 in889 0 segParams
R889890 in889 in890 {rInterSeg}
yneuron neuron890 in890 0 segParams
R890891 in890 in891 {rInterSeg}
yneuron neuron891 in891 0 segParams
R891892 in891 in892 {rInterSeg}
yneuron neuron892 in892 0 segParams
R892893 in892 in893 {rInterSeg}
yneuron neuron893 in893 0 segParams
R893894 in893 in894 {rInterSeg}
yneuron neuron894 in894 0 segParams
R894895 in894 in895 {rInterSeg}
yneuron neuron895 in895 0 segParams
R895896 in895 in896 {rInterSeg}
yneuron neuron896 in896 0 segParams
R896897 in896 in897 {rInterSeg}
yneuron neuron897 in897 0 segParams
R897898 in897 in898 {rInterSeg}
yneuron neuron898 in898 0 segParams
R898899 in898 in899 {rInterSeg}
yneuron neuron899 in899 0 segParams
R899900 in899 in900 {rInterSeg}
yneuron neuron900 in900 0 segParams
R900901 in900 in901 {rInterSeg}
yneuron neuron901 in901 0 segParams
R901902 in901 in902 {rInterSeg}
yneuron neuron902 in902 0 segParams
R902903 in902 in903 {rInterSeg}
yneuron neuron903 in903 0 segParams
R903904 in903 in904 {rInterSeg}
yneuron neuron904 in904 0 segParams
R904905 in904 in905 {rInterSeg}
yneuron neuron905 in905 0 segParams
R905906 in905 in906 {rInterSeg}
yneuron neuron906 in906 0 segParams
R906907 in906 in907 {rInterSeg}
yneuron neuron907 in907 0 segParams
R907908 in907 in908 {rInterSeg}
yneuron neuron908 in908 0 segParams
R908909 in908 in909 {rInterSeg}
yneuron neuron909 in909 0 segParams
R909910 in909 in910 {rInterSeg}
yneuron neuron910 in910 0 segParams
R910911 in910 in911 {rInterSeg}
yneuron neuron911 in911 0 segParams
R911912 in911 in912 {rInterSeg}
yneuron neuron912 in912 0 segParams
R912913 in912 in913 {rInterSeg}
yneuron neuron913 in913 0 segParams
R913914 in913 in914 {rInterSeg}
yneuron neuron914 in914 0 segParams
R914915 in914 in915 {rInterSeg}
yneuron neuron915 in915 0 segParams
R915916 in915 in916 {rInterSeg}
yneuron neuron916 in916 0 segParams
R916917 in916 in917 {rInterSeg}
yneuron neuron917 in917 0 segParams
R917918 in917 in918 {rInterSeg}
yneuron neuron918 in918 0 segParams
R918919 in918 in919 {rInterSeg}
yneuron neuron919 in919 0 segParams
R919920 in919 in920 {rInterSeg}
yneuron neuron920 in920 0 segParams
R920921 in920 in921 {rInterSeg}
yneuron neuron921 in921 0 segParams
R921922 in921 in922 {rInterSeg}
yneuron neuron922 in922 0 segParams
R922923 in922 in923 {rInterSeg}
yneuron neuron923 in923 0 segParams
R923924 in923 in924 {rInterSeg}
yneuron neuron924 in924 0 segParams
R924925 in924 in925 {rInterSeg}
yneuron neuron925 in925 0 segParams
R925926 in925 in926 {rInterSeg}
yneuron neuron926 in926 0 segParams
R926927 in926 in927 {rInterSeg}
yneuron neuron927 in927 0 segParams
R927928 in927 in928 {rInterSeg}
yneuron neuron928 in928 0 segParams
R928929 in928 in929 {rInterSeg}
yneuron neuron929 in929 0 segParams
R929930 in929 in930 {rInterSeg}
yneuron neuron930 in930 0 segParams
R930931 in930 in931 {rInterSeg}
yneuron neuron931 in931 0 segParams
R931932 in931 in932 {rInterSeg}
yneuron neuron932 in932 0 segParams
R932933 in932 in933 {rInterSeg}
yneuron neuron933 in933 0 segParams
R933934 in933 in934 {rInterSeg}
yneuron neuron934 in934 0 segParams
R934935 in934 in935 {rInterSeg}
yneuron neuron935 in935 0 segParams
R935936 in935 in936 {rInterSeg}
yneuron neuron936 in936 0 segParams
R936937 in936 in937 {rInterSeg}
yneuron neuron937 in937 0 segParams
R937938 in937 in938 {rInterSeg}
yneuron neuron938 in938 0 segParams
R938939 in938 in939 {rInterSeg}
yneuron neuron939 in939 0 segParams
R939940 in939 in940 {rInterSeg}
yneuron neuron940 in940 0 segParams
R940941 in940 in941 {rInterSeg}
yneuron neuron941 in941 0 segParams
R941942 in941 in942 {rInterSeg}
yneuron neuron942 in942 0 segParams
R942943 in942 in943 {rInterSeg}
yneuron neuron943 in943 0 segParams
R943944 in943 in944 {rInterSeg}
yneuron neuron944 in944 0 segParams
R944945 in944 in945 {rInterSeg}
yneuron neuron945 in945 0 segParams
R945946 in945 in946 {rInterSeg}
yneuron neuron946 in946 0 segParams
R946947 in946 in947 {rInterSeg}
yneuron neuron947 in947 0 segParams
R947948 in947 in948 {rInterSeg}
yneuron neuron948 in948 0 segParams
R948949 in948 in949 {rInterSeg}
yneuron neuron949 in949 0 segParams
R949950 in949 in950 {rInterSeg}
yneuron neuron950 in950 0 segParams
R950951 in950 in951 {rInterSeg}
yneuron neuron951 in951 0 segParams
R951952 in951 in952 {rInterSeg}
yneuron neuron952 in952 0 segParams
R952953 in952 in953 {rInterSeg}
yneuron neuron953 in953 0 segParams
R953954 in953 in954 {rInterSeg}
yneuron neuron954 in954 0 segParams
R954955 in954 in955 {rInterSeg}
yneuron neuron955 in955 0 segParams
R955956 in955 in956 {rInterSeg}
yneuron neuron956 in956 0 segParams
R956957 in956 in957 {rInterSeg}
yneuron neuron957 in957 0 segParams
R957958 in957 in958 {rInterSeg}
yneuron neuron958 in958 0 segParams
R958959 in958 in959 {rInterSeg}
yneuron neuron959 in959 0 segParams
R959960 in959 in960 {rInterSeg}
yneuron neuron960 in960 0 segParams
R960961 in960 in961 {rInterSeg}
yneuron neuron961 in961 0 segParams
R961962 in961 in962 {rInterSeg}
yneuron neuron962 in962 0 segParams
R962963 in962 in963 {rInterSeg}
yneuron neuron963 in963 0 segParams
R963964 in963 in964 {rInterSeg}
yneuron neuron964 in964 0 segParams
R964965 in964 in965 {rInterSeg}
yneuron neuron965 in965 0 segParams
R965966 in965 in966 {rInterSeg}
yneuron neuron966 in966 0 segParams
R966967 in966 in967 {rInterSeg}
yneuron neuron967 in967 0 segParams
R967968 in967 in968 {rInterSeg}
yneuron neuron968 in968 0 segParams
R968969 in968 in969 {rInterSeg}
yneuron neuron969 in969 0 segParams
R969970 in969 in970 {rInterSeg}
yneuron neuron970 in970 0 segParams
R970971 in970 in971 {rInterSeg}
yneuron neuron971 in971 0 segParams
R971972 in971 in972 {rInterSeg}
yneuron neuron972 in972 0 segParams
R972973 in972 in973 {rInterSeg}
yneuron neuron973 in973 0 segParams
R973974 in973 in974 {rInterSeg}
yneuron neuron974 in974 0 segParams
R974975 in974 in975 {rInterSeg}
yneuron neuron975 in975 0 segParams
R975976 in975 in976 {rInterSeg}
yneuron neuron976 in976 0 segParams
R976977 in976 in977 {rInterSeg}
yneuron neuron977 in977 0 segParams
R977978 in977 in978 {rInterSeg}
yneuron neuron978 in978 0 segParams
R978979 in978 in979 {rInterSeg}
yneuron neuron979 in979 0 segParams
R979980 in979 in980 {rInterSeg}
yneuron neuron980 in980 0 segParams
R980981 in980 in981 {rInterSeg}
yneuron neuron981 in981 0 segParams
R981982 in981 in982 {rInterSeg}
yneuron neuron982 in982 0 segParams
R982983 in982 in983 {rInterSeg}
yneuron neuron983 in983 0 segParams
R983984 in983 in984 {rInterSeg}
yneuron neuron984 in984 0 segParams
R984985 in984 in985 {rInterSeg}
yneuron neuron985 in985 0 segParams
R985986 in985 in986 {rInterSeg}
yneuron neuron986 in986 0 segParams
R986987 in986 in987 {rInterSeg}
yneuron neuron987 in987 0 segParams
R987988 in987 in988 {rInterSeg}
yneuron neuron988 in988 0 segParams
R988989 in988 in989 {rInterSeg}
yneuron neuron989 in989 0 segParams
R989990 in989 in990 {rInterSeg}
yneuron neuron990 in990 0 segParams
R990991 in990 in991 {rInterSeg}
yneuron neuron991 in991 0 segParams
R991992 in991 in992 {rInterSeg}
yneuron neuron992 in992 0 segParams
R992993 in992 in993 {rInterSeg}
yneuron neuron993 in993 0 segParams
R993994 in993 in994 {rInterSeg}
yneuron neuron994 in994 0 segParams
R994995 in994 in995 {rInterSeg}
yneuron neuron995 in995 0 segParams
R995996 in995 in996 {rInterSeg}
yneuron neuron996 in996 0 segParams
R996997 in996 in997 {rInterSeg}
yneuron neuron997 in997 0 segParams
R997998 in997 in998 {rInterSeg}
yneuron neuron998 in998 0 segParams
R998999 in998 in999 {rInterSeg}
yneuron neuron999 in999 0 segParams
R9991000 in999 in1000 {rInterSeg}
yneuron neuron1000 in1000 0 segParams
* final resistor
Rend in1000 out {rInterSeg/2.0}

.print tran 
*+ i(Iin) 
+ v(in0) 
*+ v(in1) 
*+ v(in2) 
*+ v(in500) 
*+ v(in999) 
*+ v(in1000) 
+ v(out) 

.end
