*Sample netlist for BSIM6 with sensitivity
*Drain current symmetry
.options nonlin abstol=1e-6 reltol=1e-6 
.options device temp=25

* --- Voltage Sources ---
vdrain drain 0 dc 0
esource source 0 drain 0 -1
vgate gate  0 dc -0.5
vbulk bulk 0 dc 0


* --- Transistor ---
M1 drain gate source bulk pmos W=10e-6 L=10e-6 

* --- DC Analysis ---
.dc vdrain -0.1 0.1 0.001 vgate -1 -0.4 0.3
*.probe dc ids=par'-i(vdrain)'
*.probe dc gx=deriv(ids)
*.probe dc gx2=deriv(gx)
*.probe dc gx3=deriv(gx2)
*.probe dc gx4=deriv(gx3)
*.print dc par'ids' par'gx' par'gx2' par'gx3' par 'gx4'
.print dc v(drain) v(gate) {-i(vdrain)}
*comp  d{i(vdrain)}/d(pmos:vfb)_dir reltol=0.02 abstol=1e-6
.print sens v(drain) v(gate)

.sens param=pmos:vfb,m1:l,m1:w objfunc={I(vdrain)}
.options sensitivity direct=1 adjoint=0


*modelcard for BSIM6_BD
.model pmos pmos level=77 ; bsim6
+TYPE	 = -1.0	; this is actually redundant with the model type in Xyce
+toxe    = 2.34e-009       
+toxp    = 1.925e-009       
+dtox    = 0               
+epsrox  = 3.9           
+tnom    = 25              
+xl      = 0               
+xw      = 0               
+lint    = 0             
+llong   = 1000000         
+ll      = 0               
+lw      = 0               
+lwl     = 0             
+lln     = 1               
+lwn     = 1               
+wint    = -9.0134104e-009  
+wl      = 0             
+ww      = 0               
+wwl     = 0               
+wln     = 1               
+wwn     = 1             
+wwide   = 1000000         
+dlc     = 0               
+llc     = 0               
+lwc     = 0             
+lwlc    = 0               
+dwc     = 0               
+wlc     = 0               
+wwc     = 0             
+wwlc    = 0               
+geomod  = 0               
+rgeomod = 0             
+rgatemod= 0               
+rbodymod= 0               
+igcmod  = 0               
+igbmod  = 0             
+covmod  = 1               
+rdsmod  = 0               
+gidlmod = 0               
+tnoimod = 0             
+gmin    = 1e-012          
+jss     = 0.0001          
+jsd     = 0.0001          
+jsws    = 0               
+jswd    = 0             
+jswgs   = 0               
+jswgd   = 0               
+njs     = 1               
+njd     = 1             
+ijthsfwd= 0.1             
+ijthdfwd= 0.1             
+ijthsrev= 0.1             
+ijthdrev= 0.1           
+bvs     = 10              
+bvd     = 10              
+xjbvs   = 1               
+xjbvd   = 1             
+jtss    = 0               
+jtsd    = 0               
+jtssws  = 0               
+jtsswd  = 0             
+jtsswgs = 0               
+jtsswgd = 0               
+jtweff  = 0               
+njts    = 20            
+njtsd   = 20              
+njtssw  = 20              
+njtsswd = 20              
+njtsswg = 20            
+njtsswgd= 20              
+vtss    = 10              
+vtsd    = 10              
+vtssws  = 10            
+vtsswd  = 10              
+vtsswgs = 10              
+vtsswgd = 10              
+cjs     = 0.0005        
+cjd     = 0.0005          
+cjsws   = 5e-010          
+cjswd   = 5e-010          
+cjswgs  = 0             
+cjswgd  = 0               
+pbs     = 1               
+pbd     = 1               
+pbsws   = 1             
+pbswd   = 1               
+pbswgs  = 1               
+pbswgd  = 1               
+mjs     = 0.5           
+mjd     = 0.5             
+mjsws   = 0.33            
+mjswd   = 0.33            
+mjswgs  = 0.33          
+mjswgd  = 0.33            
+tpb     = 0               
+tcj     = 0               
+tpbsw   = 0             
+tcjsw   = 0               
+tpbswg  = 0               
+tcjswg  = 0               
+xtis    = 3             
+xtid    = 3               
+xtss    = 0.02            
+xtsd    = 0.02            
+xtssws  = 0.02          
+xtsswd  = 0.02            
+xtsswgs = 0.02            
+xtsswgd = 0.02            
+tnjts   = 0             
+tnjtsd  = 0               
+tnjtssw = 0               
+tnjtsswd= 0               
+tnjtsswg= 0             
+tnjtsswgd= 0             
+noia    = 6.25e+040       
+noib    = 3.125e+025      
+noic    = 8.75e+008       
+em      = 41000000      
+ef      = 1               
+lintnoi = 0               
+ntnoi   = 1               
+tnoia   = 0             
+tnoib   = 0               
+tnoic   = 0               
+rnoia   = 0.577           
+rnoib   = 0.5164        
+rnoic   = 0.395         
+dwj     = 0               
+dmcg    = 0               
+dmci    = 0               
+dmdg    = 0             
+dmcgt   = 0               
+xgw     = 0               
+xgl     = 0             
+gbmin   = 1e-012          
+rshg    = 0.1             
+rbpb    = 50              
+rbpd    = 50            
+rbps    = 50              
+rbdb    = 50              
+rbsb    = 50              
+rbps0   = 50            
+rbpsl   = 0               
+rbpsw   = 0               
+rbpsnf  = 0               
+rbpd0   = 50            
+rbpdl   = 0               
+rbpdw   = 0               
+rbpdnf  = 0               
+rbpbx0  = 100           
+rbpbxl  = 0               
+rbpbxw  = 0               
+rbpbxnf = 0               
+rbpby0  = 100           
+rbpbyl  = 0               
+rbpbyw  = 0               
+rbpbynf = 0               
+rbsbx0  = 100           
+rbsby0  = 100             
+rbdbx0  = 100             
+rbdby0  = 100             
+rbsdbxl = 0             
+rbsdbxw = 0               
+rbsdbxnf= 0               
+rbsdbyl = 0               
+rbsdbyw = 0             
+rbsdbynf= 0               
+xrcrg1  = 12              
+xrcrg2  = 1               
+ngcon   = 1             
+ndep    = 8.062e+023      
+ndepl1  = 1.2139          
+ndeplexp1= 1.9088         
+ndepl2  = -1.1825       
+ndeplexp2= 1.9173         
+ndepw   = 0.065035        
+ndepwexp= 0.48882         
+ndepwl  = 0.00040893    
+ndepwlexp= 1.3273          
+easub   = 4.05            
+ni0sub  = 1.1e+016      
+bg0sub  = 1.17            
+epsrsub = 11.9            
+xj      = 1.5e-007        
+vfb     = -1.2108       
+vfbsdoff= 0               
+nsd     = 1e+026          
+dvtp0   = 1.8335e-007     
+dvtp1   = 220.59        
+dvtp2   = 9.6351e-010     
+dvtp3   = 0.89017         
+dvtp4   = 98.728          
+dvtp5   = 5.1435e-017   
+phin    = 0.045           
+eta0    = 0.0051075       
+etab    = -0.010908157    
+etabexp = 0.09999       
+dsub    = 1.0667          
+k2      = -0.093146       
+k2l     = 0.065574        
+k2lexp  = 0.79778       
+k2w     = 0.030809        
+k2wexp  = 0.87253         
+cit     = 1.0136148e-005  
+cdscd   = 0.0011509049  
+cdscdl  = -0.00048388809  
+cdscdlexp= 0.13963388      
+cdscb   = 9.9995516e-006  
+cdscbl  = 1.4756534e-009
+cdscblexp= 1               
+nfactor = 0.0017201       
+nfactorl= 1.7832e-006     
+nfactorlexp= 0.99988       
+nfactorw= 0.11149         
+nfactorwexp= 0.8993          
+nfactorwl= -0.01386        
+u0      = 0.04004       
+u0l     = 0.58676         
+u0lexp  = 0.11151         
+etamob  = 4.0947          
+ua      = 0.4298        
+ual     = -0.0087246      
+ualexp  = 1.3647          
+uaw     = 0.11575         
+uawexp  = 0.4385        
+uawl    = -7.027e-005     
+eu      = 1.3371          
+eul     = 0.0021948       
+eulexp  = 1.4769        
+euw     = -0.0031666      
+euwexp  = 1.9366          
+euwl    = -0.00013929     
+ud      = 0.0093995     
+udl     = 0.067484        
+udlexp  = 0.099452        
+ucs     = 0.9999          
+uc      = 4.91e-006     
+ucl     = 0.001096        
+uclexp  = 0.0015937       
+vsat    = 9609100         
+vsatl   = 6.8282        
+vsatlexp= 0.086396        
+vsatw   = 0.016834        
+vsatwexp= 3.0172          
+vsatcvl = 0             
+vsatcvlexp= 1               
+vsatcvw = 0               
+vsatcvwexp= 1               
+delta   = 0.1779        
+deltal  = 0.1269          
+deltalexp= 0.18156         
+pclm    = 0               
+pclml   = 0             
+pclmlexp= 1e-013          
+pclmg   = 0               
+pclmcvl = 0               
+pclmcvlexp= 1             
+pscbe1  = 4.24e+008       
+pscbe2  = 1e-008          
+pdits   = 0.85536         
+pditsl  = 8473.9        
+pditsd  = 0               
+pdiblc  = 0.005           
+pdiblcl = 0               
+pdiblclexp= 1             
+pdiblcb = -0.49995        
+pvag    = 1               
+fprout  = 0               
+fproutl = 0             
+fproutlexp= 1               
+ptwg    = 0.09999        
+ptwgl   = 0.069993        
+ptwglexp= 0.0009999     
+psat    = 1e-013          
+psatl   = 0               
+psatlexp= 1               
+psatb   = 0.9999        
+psatx   = 1e-013          
+rsh     = 0               
+prwg    = 1               
+prwb    = 0.010098993   
+prwbl   = 0.00070000265   
+prwblexp= 1               
+wr      = 1               
+rswmin  = 0             
+rsw     = 10              
+rswl    = 0               
+rswlexp = 1               
+rdwmin  = 0             
+rdw     = 10              
+rdwl    = 0               
+rdwlexp = 1               
+rdswmin = 0             
+rdsw    = 0               
+rdswl   = 0.0007          
+rdswlexp= 1e-007          
+alpha0  = 0             
+alpha0l = 0               
+alpha0lexp= 1               
+beta0   = 0               
+agidl   = 0             
+agidll  = 0               
+agidlw  = 0               
+bgidl   = 2.3e+009        
+cgidl   = 0.5           
+egidl   = 0.8             
+agisl   = 0               
+agisll  = 0               
+agislw  = 0             
+bgisl   = 2.3e+009        
+cgisl   = 0.5             
+egisl   = 0.00171         
+aigbacc = 0.00171       
+bigbacc = 0.00171         
+cigbacc = 0.075           
+nigbacc = 1               
+aigbinv = 0.0111        
+bigbinv = 0.000949        
+cigbinv = 0.006           
+eigbinv = 1.1             
+nigbinv = 3             
+aigc    = 0.0136          
+aigcl   = 3               
+aigcw   = 0.0136          
+bigc    = 0.00171       
+cigc    = 0.075           
+aigs    = 0.0136          
+aigsl   = 0.075           
+aigsw   = 0.0136        
+aigd    = 0.0136          
+aigdl   = 0               
+aigdw   = 0.0136          
+bigs    = 0.00171       
+bigd    = 0.00171         
+cigs    = 0.075           
+cigd    = 0.075           
+toxref  = 0.075         
+ntox    = 1               
+poxedge = 1               
+pigcd   = 1               
+pigcdl  = 1             
+ndepcv = 4.598e+23	   
+ndepcvl1= 0               
+ndepcvlexp1= 1               
+ndepcvl2= 0             
+ndepcvlexp2= 2            
+ndepcvw = 0               
+ndepcvwexp= 1               
+ndepcvwl= 0             
+ndepcvwlexp= 1            
+ngate   = 7.764e+25       
+cf      = 0               
+cfrcoeff= 1               
+cgso    = 187.0e-12       
+cgdo    = 187.0e-12             
+cgbo    = 0               
+cgsl    = 130.0e-12       
+cgdl    = 130.0e-12       
+ckappas = 1.6           
+ckappad = 1.6             
+ados    = 221.4           
+bdos    = 1.350           
+qm0     = 405.7e-6         
+etaqm   = 848.5e-3        
+vfbcv   = -996.0e-3       
+vfbcvl  = 0               
+vfbcvlexp= 1             
+vfbcvw  = 0               
+vfbcvwexp= 1               
+vfbcvwl = 0               
+vfbcvwlexp= 1             
+tbgasub = 0.000473        
+tbgbsub = 636            
+tdelta  = 0               
+ptwgt   = 0             
+iit     = 0               
+tgidl   = 0               
+igt     = 0               
+kt1     = -0.11         
+kt1l    = 0               
+kt2     = 0.022           
+kt1exp  = 1               
+ute     = -1.5          
+ua1     = 0.001           
+ud1     = 0               
+uc1     = -5.6e-011       
+ucste   = -0.004775     
+prt     = 0               
+at      = -0.00156      
+sca     = 0               
+scb     = 0               
+scc     = 0               
+sc      = 0             
+ku0we   = 0               
+kvth0we = 0               
+k2we    = 0               
+web     = 0             
+wec     = 0               
+scref   = 1e-006          
+sa      = 0               
+sb      = 0             
+sd      = 0               
+saref   = 1e-006          
+sbref   = 1e-006          
+wlod    = 0             
+kvsat   = 0               
+ku0     = 0               
+tku0    = 0               
+lku0    = 0             
+wku0    = 0               
+pku0    = 0               
+llodku0 = 0               
+wlodku0 = 0             
+kvth0   = 0               
+lkvth0  = 0               
+wkvth0  = 0               
+pkvth0  = 0             
+llodvth = 0               
+wlodvth = 0               
+stk2    = 0               
+lodk2   = 1             
+steta0  = 0               
+lodeta0 = 1             

.end
