RES_NOISE.CIR - NOISE ANALYSIS: RESISTOR DIVIDER, AMP, AND LP FILTER
*
* RESISTOR DIVIDER
*V1  1 0 AC  1 DC  5
V1  1 0 DC 5.0 AC  1.0   
R1  1 2 100K
R2  2 0 100K
*
* AMP AND LP FILTER
EAMP  3 0 2 0 1
RLP1  3 4 100
CLP1  4 0 1.59NF
* 

.NOISE  V(4)  V1  DEC   5 100 100MEG 1
.PRINT NOISE {log(ONOISE)} {log(INOISE)}
+ {log(DNO(RLP1))} {log(dno(r2))} {log(DNO(R1))}
+ {log(DNI(RLP1))} {log(DNI(R2))} {log(dni(r1))}

.options device debuglevel=-100
.options timeint debuglevel=-100

.END
