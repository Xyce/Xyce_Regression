A simple netlist to test user defined functions on the print line
*******************************************************************************
*
* a few sources of different types
VS  1  0  SIN(0 1.0 1KHZ 0 0)
VP  2  0  PULSE( 0 100 0.2ms 0.2ms 0.2ms 1ms 2ms )

R1  1  0  100
R2  2  0  100

.func f(x) {abs(x)}
.func g(x) {3*x + 1}

.TRAN 0  10ms
.PRINT TRAN  V(1) {f(v(1))} V(2) {g(v(2))}

.END

