*Trivial sweep of diode to produce I/V curve, DTEMP version

.param diodeDtemp = -82
.options device temp = 27.0

.tran 0 1 0 100m
.step diodeDtemp list -82 -2 45

.print tran V(2) 
*{TEMP+diodeDtemp}

*COMP V(2) reltol=0.005

VIN 1 0 pulse ( 7.5 10 1m 1 1 3 6)
R1  1 2 1k
DZR 0 2 DZR   DTEMP=diodeDtemp
.MODEL DZR D( level=2
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 1P
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 7.255;7.25 yields vout=5V @25C;6.9504;Vref determines Vout
+        IBV = .001
+ tbv1 = 0.00013
+ tbv2 = -5e-8
+        
+ )
