$special variables
* Xyce netlist for corresponding HSPICE netlist.
* Netlist tests XDM recognizes special variables 
* in source & target languages, and makes the
* appropriate translation if possible or comments
* out the line if not. Only the HSPICE special
* variable "temper" can be translated, into "temp"
* in Xyce. Expressions using "hertz" will
* have warnings and be commented out.
* A parameter name of "vt" or an expression
* that uses a parameter "vt" in HSPICE will 
* have warnings and be commented out (see issue
* #69 on XDM gitlab).

.GLOBAL_PARAM XYCE_TEMP = 'TEMP'
.PARAM KTQ='1.38e-23*XYCE_TEMP/1.602e-19'
.PARAM USESVT1='2'

VA 1 0 DC 0.8 AC 1
R1 1 2 R='XYCE_TEMP'
C1 2 0 C=1n
.AC dec 2 1000 100000

.PRINT AC FORMAT=PROBE 'XYCE_TEMP' 'ktq' 

