A simple test case of a resistor with zero resistance

* test case for when resistance is near zero
V1 a 0 5V
R1 a b {1.0e-101}
R2 b 0 1K

.DC V1 0 5V 1V
.PRINT dc V(a) I(R1) 

.END
