AC test of FORMAT=CSV output format with .OP
*

* Trivial high-pass filter
R1 b 0 2
C1 a b 1u
V1 a 0 DC 0V AC 1

.print AC FORMAT=CSV R1:R vm(b)
.ac dec 5 100Hz 1e6
.op

.end
