* Xyce netlist for testing various syntaxes for H-Sources

* source that provides the controlling current
R1 1 0  1 
V1 1 0  SIN(0V 1V 1e3 0 0 0)

* linear form
H2 2 0 V1 2
R2 2 0 1

* poly form
H3 3 0 poly(1) V1 0 3
R3 3 0 1

.TRAN 10us 1ms
.PRINT TRAN format=probe V(1) V(2) V(3)
.END
