Basic dual diode circuit for baseline calculation
* All this does is provide a standard against which alternate versions
* of the circuit can be compared

V1 1 0 DC 5V
R1 1 2 2K
Vmon1 2 3 0V
D1 3 0 DMOD1
Vmon2 2 4 0V
D2 4 0 DMOD2

.model DMOD1 D (IS=100FA)
.model DMOD2 D (IS=200FA)
.dc V1 0 5 1
.print DC v(1) I(v1) I(vmon1) I(vmon2)
.end
