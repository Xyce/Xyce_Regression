Test Circuit for the Inductor 
********************************************************************************
* Tier No.:  1
* Description: Circuit netlist to verify calculation 
*              accuracy of the inductor model. 
* Analysis:
*       A small resistor and a zero volt source, VMON, is placed in series with
*       the inductor.  The input current, defined by a nonlinear dependent 
*       source, B1, is:
*
*         B1 = I = 10*t*exp(-5t)   for t>0
*
*       The voltage generated by the inductor is given by:
*
*         V(3) = L*dI/dt 
*              = L * d(10*t*exp(-5t))/dt 
*              = 10 * L * exp(-5t) * (1 - 5t)
*
*       where L is calculated from the temperature model:
*
*         L = baseL*factor;
*         baseL = 10mH = 0.01;
*
*         tdel = (temp - tnom) = 363.15 - 300.15 = 63;
*         TC1 = 0.01;
*         TC2 = 0.926e-4;
*
*         factor = 1.0 + (TC1)*tdel + (TC2)*tdel*tdel = 1.99753;
*
*         L = 0.0199753 H;
*
* The values for I(VMON) and V(3) can be calculated analytically, using
* the perl script tempind.cir.prn.gs.pl.  This script must be run after
* Xyce has been run on this netlist to produce a *prn file.
*
********************************************************************************
B1 0 1  I = {10 * TIME * EXP( - 5*TIME)}
VMON 1 2 0
R1 2 3  0.000001
L1 3 0 IND1 10mH TEMP=90
.MODEL IND1 L  ( TC1=0.010 TC2=0.926e-4 )
*
.TRAN 0.1MS 20MS
.PRINT TRAN I(VMON) V(3)
.END

