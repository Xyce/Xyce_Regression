Netlist to Test Xyce with RLC
*********************************************************************
* Tier No.:     1
* Description: Solution verfication circuit containing the linear
*              resistor, capacitor, and inductor models implemented
*              in Xyce.
* Creator:  Ben Long
*
* Input: VIN=10V DC
* Output: Current through V1
* Circuit Elements: R1, L1, C1
* Analysis:
*       The solution is the zero state response of the circuit below:
*       A DC voltage source in series with a 3 Ohm resistor,
*       a 1H inductor, and a .5F capacitor.  The measured output
*       is the current through the loop.
*
*        1___/\/\/\___2___ccccc__3
*        |       R1             L1   |
*        |      --> I                   ---
*       (V1)                       C1 ---
*        |                               |
*        |                               |
*        |_______________________|
*                       0
*
***********************************************************************
r1 1 2 3
l1 2 3 1
c1 3 0 .5
v1 1 0 1

* Note: the current has 1 subtracted from it to help with xyce_verify.
.print tran v(1)
.options timeint reltol=1.0e-3

* Analysis
.TRAN 0 2e-07
.OPTIONS OUTPUT outputtimepoints=0.000000e+00,7.014409e-08,7.750647e-08,8.185960e-08,8.496698e-08,8.738731e-08,8.937110e-08,9.105258e-08,9.251216e-08,9.380187e-08,9.495731e-08,9.600394e-08,9.696058e-08,9.784155e-08,9.865800e-08,9.941878e-08,1.001310e-07,1.008006e-07,1.014323e-07,1.020303e-07,1.025979e-07,1.031381e-07,1.036535e-07,1.041462e-07,1.046182e-07,1.050712e-07,1.055065e-07,1.059256e-07,1.063297e-07,1.067197e-07,1.070966e-07,1.074613e-07,1.078145e-07,1.081570e-07,1.084893e-07,1.088121e-07,1.091260e-07,1.094313e-07,1.097285e-07,1.100181e-07,1.103005e-07,1.105759e-07,1.108448e-07,1.111074e-07,1.113641e-07,1.116150e-07,1.118604e-07,1.121007e-07,1.123359e-07,1.125663e-07,1.127922e-07,1.130135e-07,1.132307e-07,1.134437e-07,1.136528e-07,1.138581e-07,1.140597e-07,1.142578e-07,1.144525e-07,1.146439e-07,1.148321e-07,1.150172e-07,1.151993e-07,1.153786e-07,1.155550e-07,1.157288e-07,1.158999e-07,1.160684e-07,1.162345e-07,1.163982e-07,1.165596e-07,1.167186e-07,1.168755e-07,1.170303e-07,1.171829e-07,1.173335e-07,1.174822e-07,1.176289e-07,1.177737e-07,1.179167e-07,1.180580e-07,1.181975e-07,1.183353e-07,1.184714e-07,1.186059e-07,1.187389e-07,1.188703e-07,1.190002e-07,1.191286e-07,1.192556e-07,1.193812e-07,1.195054e-07,1.196282e-07,1.197498e-07,1.198700e-07,1.199890e-07,1.201068e-07,1.202233e-07,1.203387e-07,1.204529e-07,1.205660e-07,1.206779e-07,1.207888e-07,1.208986e-07,1.210073e-07,1.211150e-07,1.212217e-07,1.213274e-07,1.214321e-07,1.215359e-07,1.216387e-07,1.217406e-07,1.218416e-07,1.219417e-07,1.220410e-07,1.221393e-07,1.222369e-07,1.223336e-07,1.224294e-07,1.225245e-07,1.226188e-07,1.227123e-07,1.228051e-07,1.228971e-07,1.229883e-07,1.230789e-07,1.231687e-07,1.232578e-07,1.233462e-07,1.234340e-07,1.235210e-07,1.236075e-07,1.236932e-07,1.237783e-07,1.238628e-07,1.239467e-07,1.240299e-07,1.241125e-07,1.241946e-07,1.242760e-07,1.243569e-07,1.244372e-07,1.245170e-07,1.245962e-07,1.246748e-07,1.247529e-07,1.248305e-07,1.249075e-07,1.249840e-07,1.250601e-07,1.251356e-07,1.252106e-07,1.252851e-07,1.253591e-07,1.254327e-07,1.255058e-07,1.255784e-07,1.256506e-07,1.257223e-07,1.257935e-07,1.258643e-07,1.259347e-07,1.260047e-07,1.260742e-07,1.261433e-07,1.262119e-07,1.262802e-07,1.263481e-07,1.264155e-07,1.264826e-07,1.265492e-07,1.266155e-07,1.266814e-07,1.267469e-07,1.268121e-07,1.268769e-07,1.269413e-07,1.270053e-07,1.270690e-07,1.271323e-07,1.271953e-07,1.272579e-07,1.273202e-07,1.273822e-07,1.274438e-07,1.275051e-07,1.275661e-07,1.276267e-07,1.276870e-07,1.277470e-07,1.278067e-07,1.278661e-07,1.279251e-07,1.279839e-07,1.280424e-07,1.281005e-07,1.281584e-07,1.282160e-07,1.282732e-07,1.283302e-07,1.283870e-07,1.284434e-07,1.284995e-07,1.285554e-07,1.286110e-07,1.286664e-07,1.287214e-07,1.287763e-07,1.288308e-07,1.288851e-07,1.289391e-07,1.289929e-07,1.290464e-07,1.290997e-07,1.291527e-07,1.292055e-07,1.292580e-07,1.293103e-07,1.293624e-07,1.294142e-07,1.294658e-07,1.295171e-07,1.295682e-07,1.296191e-07,1.296698e-07,1.297203e-07,1.297705e-07,1.298205e-07,1.298703e-07,1.299198e-07,1.299692e-07,1.300183e-07,1.300673e-07,1.301160e-07,1.301645e-07,1.302128e-07,1.302609e-07,1.303088e-07,1.303565e-07,1.304040e-07,1.304513e-07,1.304985e-07,1.305454e-07,1.305921e-07,1.306386e-07,1.306850e-07,1.307312e-07,1.307771e-07,1.308229e-07,1.308685e-07,1.309140e-07,1.309592e-07,1.310043e-07,1.310492e-07,1.310939e-07,1.311384e-07,1.311828e-07,1.312270e-07,1.312710e-07,1.313149e-07,1.313586e-07,1.314021e-07,1.314454e-07,1.314886e-07,1.315317e-07,1.315745e-07,1.316172e-07,1.316598e-07,1.317022e-07,1.317444e-07,1.317865e-07,1.318284e-07,1.318702e-07,1.319118e-07,1.319533e-07,1.319946e-07,1.320358e-07,1.320768e-07,1.321177e-07,1.321584e-07,1.321990e-07,1.322394e-07,1.322797e-07,1.323199e-07,1.323599e-07,1.323998e-07,1.324395e-07,1.324791e-07,1.325186e-07,1.325579e-07,1.325971e-07,1.326362e-07,1.326751e-07,1.327139e-07,1.327525e-07,1.327911e-07,1.328295e-07,1.328677e-07,1.329059e-07,1.329439e-07,1.329818e-07,1.330196e-07,1.330572e-07,1.330947e-07,1.331321e-07,1.331694e-07,1.332066e-07,1.332436e-07,1.332805e-07,1.333173e-07,1.333540e-07,1.333906e-07,1.334270e-07,1.334633e-07,1.334995e-07,1.335356e-07,1.335716e-07,1.336075e-07,1.336433e-07,1.336789e-07,1.337145e-07,1.337499e-07,1.337852e-07,1.338204e-07,1.338555e-07,1.338905e-07,1.339254e-07,1.339602e-07,1.339949e-07,1.340294e-07,1.340639e-07,1.340983e-07,1.341325e-07,1.341667e-07,1.342007e-07,1.342347e-07,1.342686e-07,1.343023e-07,1.343360e-07,1.343695e-07,1.344030e-07,1.344363e-07,1.344696e-07,1.345028e-07,1.345359e-07,1.345688e-07,1.346017e-07,1.346345e-07,1.346672e-07,1.346998e-07,1.347323e-07,1.347647e-07,1.347970e-07,1.348293e-07,1.348614e-07,1.348935e-07,1.349254e-07,1.349573e-07,1.349891e-07,1.350208e-07,1.350524e-07,1.350839e-07,1.351154e-07,1.351467e-07,1.351780e-07,1.352092e-07,1.352403e-07,1.352713e-07,1.353022e-07,1.353331e-07,1.353638e-07,1.353945e-07,1.354251e-07,1.354556e-07,1.354860e-07,1.355164e-07,1.355467e-07,1.355769e-07,1.356070e-07,1.356370e-07,1.356670e-07,1.356968e-07,1.357266e-07,1.357564e-07,1.357860e-07,1.358156e-07,1.358451e-07,1.358745e-07,1.359038e-07,1.359331e-07,1.359623e-07,1.359914e-07,1.360205e-07,1.360494e-07,1.360783e-07,1.361072e-07,1.361359e-07,1.361646e-07,1.361932e-07,1.362217e-07,1.362502e-07,1.362786e-07,1.363069e-07,1.363352e-07,1.363634e-07,1.363915e-07,1.364195e-07,1.364475e-07,1.364754e-07,1.365033e-07,1.365311e-07,1.365588e-07,1.365864e-07,1.366140e-07,1.366415e-07,1.366689e-07,1.366963e-07,1.367236e-07,1.367509e-07,1.367781e-07,1.368052e-07,1.368322e-07,1.368592e-07,1.368861e-07,1.369130e-07,1.369398e-07,1.369666e-07,1.369932e-07,1.370198e-07,1.370464e-07,1.370729e-07,1.370993e-07,1.371257e-07,1.371520e-07,1.371783e-07,1.372044e-07,1.372306e-07,1.372566e-07,1.372827e-07,1.373086e-07,1.373345e-07,1.373603e-07,1.373861e-07,1.374118e-07,1.374375e-07,1.374631e-07,1.374886e-07,1.375141e-07,1.375396e-07,1.375649e-07,1.375903e-07,1.376155e-07,1.376407e-07,1.376659e-07,1.376910e-07,1.377160e-07,1.377410e-07,1.377660e-07,1.377908e-07,1.378157e-07,1.378404e-07,1.378652e-07,1.378898e-07,1.379144e-07,1.379390e-07,1.379635e-07,1.379880e-07,1.380124e-07,1.380367e-07,1.380610e-07,1.380853e-07,1.381095e-07,1.381336e-07,1.381577e-07,1.381818e-07,1.382058e-07,1.382297e-07,1.382536e-07,1.382775e-07,1.383012e-07,1.383250e-07,1.383487e-07,1.383723e-07,1.383959e-07,1.384195e-07,1.384430e-07,1.384665e-07,1.384899e-07,1.385132e-07,1.385365e-07,1.385598e-07,1.385830e-07,1.386062e-07,1.386293e-07,1.386524e-07,1.386754e-07,1.386984e-07,1.387214e-07,1.387442e-07,1.387671e-07,1.387899e-07,1.388127e-07,1.388354e-07,1.388580e-07,1.388807e-07,1.389032e-07,1.389258e-07,1.389483e-07,1.389707e-07,1.389931e-07,1.390155e-07,1.390378e-07,1.390601e-07,1.390823e-07,1.391045e-07,1.391266e-07,1.391487e-07,1.391708e-07,1.391928e-07,1.392148e-07,1.392367e-07,1.392586e-07,1.392804e-07,1.393022e-07,1.393240e-07,1.393457e-07,1.393674e-07,1.393890e-07,1.394106e-07,1.394322e-07,1.394537e-07,1.394752e-07,1.394966e-07,1.395180e-07,1.395394e-07,1.395607e-07,1.395820e-07,1.396032e-07,1.396244e-07,1.396456e-07,1.396667e-07,1.396878e-07,1.397088e-07,1.397299e-07,1.397508e-07,1.397718e-07,1.397926e-07,1.398135e-07,1.398343e-07,1.398551e-07,1.398758e-07,1.398965e-07,1.399172e-07,1.399378e-07,1.399584e-07,1.399790e-07,1.399995e-07,1.400200e-07,1.400404e-07,1.400608e-07,1.400812e-07,1.401016e-07,1.401219e-07,1.401421e-07,1.401623e-07,1.401825e-07,1.402027e-07,1.402228e-07,1.402429e-07,1.402630e-07,1.402830e-07,1.403030e-07,1.403229e-07,1.403428e-07,1.403627e-07,1.403825e-07,1.404024e-07,1.404221e-07,1.404419e-07,1.404616e-07,1.404813e-07,1.405009e-07,1.405205e-07,1.405401e-07,1.405596e-07,1.405791e-07,1.405986e-07,1.406180e-07,1.406374e-07,1.406568e-07,1.406762e-07,1.406955e-07,1.407148e-07,1.407340e-07,1.407532e-07,1.407724e-07,1.407915e-07,1.408107e-07,1.408297e-07,1.408488e-07,1.408678e-07,1.408868e-07,1.409058e-07,1.409247e-07,1.409436e-07,1.409625e-07,1.409813e-07,1.410001e-07,1.410189e-07,1.410376e-07,1.410563e-07,1.410750e-07,1.410937e-07,1.411123e-07,1.411309e-07,1.411494e-07,1.411680e-07,1.411865e-07,1.412049e-07,1.412234e-07,1.412418e-07,1.412602e-07,1.412785e-07,1.412969e-07,1.413151e-07,1.413334e-07,1.413517e-07,1.413699e-07,1.413880e-07,1.414062e-07,1.414243e-07,1.414424e-07,1.414605e-07,1.414785e-07,1.414965e-07,1.415145e-07,1.415324e-07,1.415504e-07,1.415683e-07,1.415861e-07,1.416040e-07,1.416218e-07,1.416396e-07,1.416573e-07,1.416751e-07,1.416928e-07,1.417104e-07,1.417281e-07,1.417457e-07,1.417633e-07,1.417809e-07,1.417984e-07,1.418159e-07,1.418334e-07,1.418509e-07,1.418683e-07,1.418857e-07,1.419031e-07,1.419204e-07,1.419378e-07,1.419551e-07,1.419723e-07,1.419896e-07,1.420068e-07,1.420240e-07,1.420412e-07,1.420583e-07,1.420755e-07,1.420926e-07,1.421096e-07,1.421267e-07,1.421437e-07,1.421607e-07,1.421777e-07,1.421946e-07,1.422115e-07,1.422284e-07,1.422453e-07,1.422621e-07,1.422790e-07,1.422958e-07,1.423125e-07,1.423293e-07,1.423460e-07,1.423627e-07,1.423794e-07,1.423960e-07,1.424126e-07,1.424292e-07,1.424458e-07,1.424624e-07,1.424789e-07,1.424954e-07,1.425119e-07,1.425284e-07,1.425448e-07,1.425612e-07,1.425776e-07,1.425940e-07,1.426103e-07,1.426266e-07,1.426429e-07,1.426592e-07,1.426754e-07,1.426917e-07,1.427079e-07,1.427241e-07,1.427402e-07,1.427563e-07,1.427725e-07,1.427886e-07,1.428046e-07,1.428207e-07,1.428367e-07,1.428527e-07,1.428687e-07,1.428846e-07,1.429006e-07,1.429165e-07,1.429324e-07,1.429482e-07,1.429641e-07,1.429799e-07,1.429957e-07,1.430115e-07,1.430272e-07,1.430430e-07,1.430587e-07,1.430744e-07,1.430901e-07,1.431057e-07,1.431214e-07,1.431370e-07,1.431525e-07,1.431681e-07,1.431837e-07,1.431992e-07,1.432147e-07,1.432302e-07,1.432456e-07,1.432611e-07,1.432765e-07,1.432919e-07,1.433073e-07,1.433226e-07,1.433380e-07,1.433533e-07,1.433686e-07,1.433839e-07,1.433991e-07,1.434144e-07,1.434296e-07,1.434448e-07,1.434600e-07,1.434751e-07,1.434903e-07,1.435054e-07,1.435205e-07,1.435355e-07,1.435506e-07,1.435656e-07,1.435807e-07,1.435957e-07,1.436106e-07,1.436256e-07,1.436405e-07,1.436555e-07,1.436704e-07,1.436852e-07,1.437001e-07,1.437149e-07,1.437298e-07,1.437446e-07,1.437594e-07,1.437741e-07,1.437889e-07,1.438036e-07,1.438183e-07,1.438330e-07,1.438477e-07,1.438623e-07,1.438770e-07,1.438916e-07,1.439062e-07,1.439208e-07,1.439353e-07,1.439499e-07,1.439644e-07,1.439789e-07,1.439934e-07,1.440079e-07,1.440223e-07,1.440367e-07,1.440512e-07,1.440656e-07,1.440799e-07,1.440943e-07,1.441086e-07,1.441230e-07,1.441373e-07,1.441516e-07,1.441658e-07,1.441801e-07,1.441943e-07,1.442086e-07,1.442228e-07,1.442369e-07,1.442511e-07,1.442653e-07,1.442794e-07,1.442935e-07,1.443076e-07,1.443217e-07,1.443357e-07,1.443498e-07,1.443638e-07,1.443778e-07,1.443918e-07,1.444058e-07,1.444198e-07,1.444337e-07,1.444476e-07,1.444615e-07,1.444754e-07,1.444893e-07,1.445032e-07,1.445170e-07,1.445308e-07,1.445446e-07,1.445584e-07,1.445722e-07,1.445860e-07,1.445997e-07,1.446134e-07,1.446272e-07,1.446409e-07,1.446545e-07,1.446682e-07,1.446818e-07,1.446955e-07,1.447091e-07,1.447227e-07,1.447363e-07,1.447498e-07,1.447634e-07,1.447769e-07,1.447904e-07,1.448039e-07,1.448174e-07,1.448309e-07,1.448443e-07,1.448578e-07,1.448712e-07,1.448846e-07,1.448980e-07,1.449114e-07,1.449247e-07,1.449381e-07,1.449514e-07,1.449647e-07,1.449780e-07,1.449913e-07,1.450046e-07,1.450178e-07,1.450311e-07,1.450443e-07,1.450575e-07,1.450707e-07,1.450839e-07,1.450970e-07,1.451102e-07,1.451233e-07,1.451364e-07,1.451495e-07,1.451626e-07,1.451757e-07,1.451887e-07,1.452018e-07,1.452148e-07,1.452278e-07,1.452408e-07,1.452538e-07,1.452668e-07,1.452797e-07,1.452927e-07,1.453056e-07,1.453185e-07,1.453314e-07,1.453443e-07,1.453571e-07,1.453700e-07,1.453828e-07,1.453957e-07,1.454085e-07,1.454213e-07,1.454340e-07,1.454468e-07,1.454596e-07,1.454723e-07,1.454850e-07,1.454977e-07,1.455104e-07,1.455231e-07,1.455358e-07,1.455484e-07,1.455611e-07,1.455737e-07,1.455863e-07,1.455989e-07,1.456115e-07,1.456241e-07,1.456366e-07,1.456492e-07,1.456617e-07,1.456742e-07,1.456867e-07,1.456992e-07,1.457117e-07,1.457242e-07,1.457366e-07,1.457490e-07,1.457615e-07,1.457739e-07,1.457863e-07,1.457987e-07,1.458110e-07,1.458234e-07,1.458357e-07,1.458480e-07,1.458604e-07,1.458727e-07,1.458850e-07,1.458972e-07,1.459095e-07,1.459217e-07,1.459340e-07,1.459462e-07,1.459584e-07,1.459706e-07,1.459828e-07,1.459950e-07,1.460071e-07,1.460193e-07,1.460314e-07,1.460435e-07,1.460557e-07,1.460677e-07,1.460798e-07,1.460919e-07,1.461040e-07,1.461160e-07,1.461280e-07,1.461401e-07,1.461521e-07,1.461641e-07,1.461760e-07,1.461880e-07,1.462000e-07,1.462119e-07,1.462238e-07,1.462358e-07,1.462477e-07,1.462596e-07,1.462715e-07,1.462833e-07,1.462952e-07,1.463070e-07,1.463189e-07,1.463307e-07,1.463425e-07,1.463543e-07,1.463661e-07,1.463779e-07,1.463896e-07,1.464014e-07,1.464131e-07,1.464248e-07,1.464366e-07,1.464483e-07,1.464599e-07,1.464716e-07,1.464833e-07,1.464949e-07,1.465066e-07,1.465182e-07,1.465298e-07,1.465415e-07,1.465530e-07,1.465646e-07,1.465762e-07,1.465878e-07,1.465993e-07,1.466109e-07,1.466224e-07,1.466339e-07,1.466454e-07,1.466569e-07,1.466684e-07,1.466798e-07,1.466913e-07,1.467027e-07,1.467142e-07,1.467256e-07,1.467370e-07,1.467484e-07,1.467598e-07,1.467712e-07,1.467826e-07,1.467939e-07,1.468053e-07,1.468166e-07,1.468279e-07,1.468392e-07,1.468505e-07,1.468618e-07,1.468731e-07,1.468844e-07,1.468956e-07,1.469069e-07,1.469181e-07,1.469293e-07,1.469405e-07,1.469517e-07,1.469629e-07,1.469741e-07,1.469853e-07,1.469964e-07,1.470076e-07,1.470187e-07,1.470298e-07,1.470410e-07,1.470521e-07,1.470631e-07,1.470742e-07,1.470853e-07,1.470964e-07,1.471074e-07,1.471185e-07,1.471295e-07,1.471405e-07,1.471515e-07,1.471625e-07,1.471735e-07,1.471845e-07,1.471954e-07,1.472064e-07,1.472173e-07,1.472283e-07,1.472392e-07,1.472501e-07,1.472610e-07,1.472719e-07,1.472828e-07,1.472937e-07,1.473045e-07,1.473154e-07,1.473262e-07,1.473371e-07,1.473479e-07,1.473587e-07,1.473695e-07,1.473803e-07,1.473911e-07,1.474018e-07,1.474126e-07,1.474234e-07,1.474341e-07,1.474448e-07,1.474556e-07,1.474663e-07,1.474770e-07,1.474877e-07,1.474983e-07,1.475090e-07,1.475197e-07,1.475303e-07,1.475410e-07,1.475516e-07,1.475622e-07,1.475728e-07,1.475834e-07,1.475940e-07,1.476046e-07,1.476152e-07,1.476258e-07,1.476363e-07,1.476469e-07,1.476574e-07,1.476679e-07,1.476784e-07,1.476889e-07,1.476994e-07,1.477099e-07,1.477204e-07,1.477309e-07,1.477413e-07,1.477518e-07,1.477622e-07,1.477726e-07,1.477831e-07,1.477935e-07,1.478039e-07,1.478143e-07,1.478247e-07,1.478350e-07,1.478454e-07,1.478557e-07,1.478661e-07,1.478764e-07,1.478868e-07,1.478971e-07,1.479074e-07,1.479177e-07,1.479280e-07,1.479383e-07,1.479485e-07,1.479588e-07,1.479690e-07,1.479793e-07,1.479895e-07,1.479998e-07,1.480100e-07,1.480202e-07,1.480304e-07,1.480406e-07,1.480507e-07,1.480609e-07,1.480711e-07,1.480812e-07,1.480914e-07,1.481015e-07,1.481116e-07,1.481218e-07,1.481319e-07,1.481420e-07,1.481521e-07,1.481622e-07,1.481722e-07,1.481823e-07,1.481924e-07,1.482024e-07,1.482124e-07,1.482225e-07,1.482325e-07,1.482425e-07,1.482525e-07,1.482625e-07,1.482725e-07,1.482825e-07,1.482924e-07,1.483024e-07,1.483124e-07,1.483223e-07,1.483322e-07,1.483422e-07,1.483521e-07,1.483620e-07,1.483719e-07,1.483818e-07,1.483917e-07,1.484015e-07,1.484114e-07,1.484213e-07,1.484311e-07,1.484410e-07,1.484508e-07,1.484606e-07,1.484704e-07,1.484802e-07,1.484900e-07,1.484998e-07,1.485096e-07,1.485194e-07,1.485292e-07,1.485389e-07,1.485487e-07,1.485584e-07,1.485681e-07,1.485779e-07,1.485876e-07,1.485973e-07,1.486070e-07,1.486167e-07,1.486264e-07,1.486361e-07,1.486457e-07,1.486554e-07,1.486650e-07,1.486747e-07,1.486843e-07,1.486939e-07,1.487036e-07,1.487132e-07,1.487228e-07,1.487324e-07,1.487420e-07,1.487515e-07,1.487611e-07,1.487707e-07,1.487802e-07,1.487898e-07,1.487993e-07,1.488089e-07,1.488184e-07,1.488279e-07,1.488374e-07,1.488469e-07,1.488564e-07,1.488659e-07,1.488754e-07,1.488848e-07,1.488943e-07,1.489038e-07,1.489132e-07,1.489226e-07,1.489321e-07,1.489415e-07,1.489509e-07,1.489603e-07,1.489697e-07,1.489791e-07,1.489885e-07,1.489979e-07,1.490072e-07,1.490166e-07,1.490260e-07,1.490353e-07,1.490446e-07,1.490540e-07,1.490633e-07,1.490726e-07,1.490819e-07,1.490912e-07,1.491005e-07,1.491098e-07,1.491191e-07,1.491284e-07,1.491376e-07,1.491469e-07,1.491561e-07,1.491654e-07,1.491746e-07,1.491838e-07,1.491931e-07,1.492023e-07,1.492115e-07,1.492207e-07,1.492299e-07,1.492390e-07,1.492482e-07,1.492574e-07,1.492665e-07,1.492757e-07,1.492848e-07,1.492940e-07,1.493031e-07,1.493122e-07,1.493214e-07,1.493305e-07,1.493396e-07,1.493487e-07,1.493578e-07,1.493668e-07,1.493759e-07,1.493850e-07,1.493940e-07,1.494031e-07,1.494121e-07,1.494212e-07,1.494302e-07,1.494392e-07,1.494483e-07,1.494573e-07,1.494663e-07,1.494753e-07,1.494843e-07,1.494932e-07,1.495022e-07,1.495112e-07,1.495201e-07,1.495291e-07,1.495381e-07,1.495470e-07,1.495559e-07,1.495649e-07,1.495738e-07,1.495827e-07,1.495916e-07,1.496005e-07,1.496094e-07,1.496183e-07,1.496271e-07,1.496360e-07,1.496449e-07,1.496537e-07,1.496626e-07,1.496714e-07,1.496803e-07,1.496891e-07,1.496979e-07,1.497068e-07,1.497156e-07,1.497244e-07,1.497332e-07,1.497420e-07,1.497507e-07,1.497595e-07,1.497683e-07,1.497771e-07,1.497858e-07,1.497946e-07,1.498033e-07,1.498120e-07,1.498208e-07,1.498295e-07,1.498382e-07,1.498469e-07,1.498556e-07,1.498643e-07,1.498730e-07,1.498817e-07,1.498904e-07,1.498991e-07,1.499077e-07,1.499164e-07,1.499250e-07,1.499337e-07,1.499423e-07,1.499509e-07,1.499596e-07,1.499682e-07,1.499768e-07,1.499854e-07,1.499940e-07,1.500026e-07,1.500112e-07,1.500198e-07,1.500284e-07,1.500369e-07,1.500455e-07,1.500540e-07,1.500626e-07,1.500711e-07,1.500797e-07,1.500882e-07,1.500967e-07,1.501052e-07,1.501138e-07,1.501223e-07,1.501308e-07,1.501393e-07,1.501477e-07,1.501562e-07,1.501647e-07,1.501732e-07,1.501816e-07,1.501901e-07,1.501985e-07,1.502070e-07,1.502154e-07,1.502238e-07,1.502323e-07,1.502407e-07,1.502491e-07,1.502575e-07,1.502659e-07,1.502743e-07,1.502827e-07,1.502911e-07,1.502994e-07,1.503078e-07,1.503162e-07,1.503245e-07,1.503329e-07,1.503412e-07,1.503496e-07,1.503579e-07,1.503662e-07,1.503745e-07,1.503829e-07,1.503912e-07,1.503995e-07,1.504078e-07,1.504161e-07,1.504244e-07,1.504326e-07,1.504409e-07,1.504492e-07,1.504574e-07,1.504657e-07,1.504739e-07,1.504822e-07,1.504904e-07,1.504987e-07,1.505069e-07,1.505151e-07,1.505233e-07,1.505315e-07,1.505397e-07,1.505479e-07,1.505561e-07,1.505643e-07,1.505725e-07,1.505807e-07,1.505888e-07,1.505970e-07,1.506051e-07,1.506133e-07,1.506214e-07,1.506296e-07,1.506377e-07,1.506458e-07,1.506540e-07,1.506621e-07,1.506702e-07,1.506783e-07,1.506864e-07,1.506945e-07,1.507026e-07,1.507107e-07,1.507187e-07,1.507268e-07,1.507349e-07,1.507429e-07,1.507510e-07,1.507590e-07,1.507671e-07,1.507751e-07,1.507831e-07,1.507912e-07,1.507992e-07,1.508072e-07,1.508152e-07,1.508232e-07,1.508312e-07,1.508392e-07,1.508472e-07,1.508552e-07,1.508631e-07,1.508711e-07,1.508791e-07,1.508870e-07,1.508950e-07,1.509029e-07,1.509109e-07,1.509188e-07,1.509268e-07,1.509347e-07,1.509426e-07,1.509505e-07,1.509584e-07,1.509663e-07,1.509742e-07,1.509821e-07,1.509900e-07,1.509979e-07,1.510058e-07,1.510136e-07,1.510215e-07,1.510294e-07,1.510372e-07,1.510451e-07,1.510529e-07,1.510608e-07,1.510686e-07,1.510764e-07,1.510843e-07,1.510921e-07,1.510999e-07,1.511077e-07,1.511155e-07,1.511233e-07,1.511311e-07,1.511389e-07,1.511467e-07,1.511544e-07,1.511622e-07,1.511700e-07,1.511777e-07,1.511855e-07,1.511932e-07,1.512010e-07,1.512087e-07,1.512165e-07,1.512242e-07,1.512319e-07,1.512396e-07,1.512474e-07,1.512551e-07,1.512628e-07,1.512705e-07,1.512782e-07,1.512859e-07,1.512935e-07,1.513012e-07,1.513089e-07,1.513166e-07,1.513242e-07,1.513319e-07,1.513395e-07,1.513472e-07,1.513548e-07,1.513625e-07,1.513701e-07,1.513777e-07,1.513853e-07,1.513930e-07,1.514006e-07,1.514082e-07,1.514158e-07,1.514234e-07,1.514310e-07,1.514386e-07,1.514461e-07,1.514537e-07,1.514613e-07,1.514689e-07,1.514764e-07,1.514840e-07,1.514915e-07,1.514991e-07,1.515066e-07,1.515142e-07,1.515217e-07,1.515292e-07,1.515367e-07,1.515443e-07,1.515518e-07,1.515593e-07,1.515668e-07,1.515743e-07,1.515818e-07,1.515893e-07,1.515968e-07,1.516042e-07,1.516117e-07,1.516192e-07,1.516266e-07,1.516341e-07,1.516416e-07,1.516490e-07,1.516565e-07,1.516639e-07,1.516713e-07,1.516788e-07,1.516862e-07,1.516936e-07,1.517010e-07,1.517084e-07,1.517159e-07,1.517233e-07,1.517307e-07,1.517380e-07,1.517454e-07,1.517528e-07,1.517602e-07,1.517676e-07,1.517749e-07,1.517823e-07,1.517897e-07,1.517970e-07,1.518044e-07,1.518117e-07,1.518191e-07,1.518264e-07,1.518337e-07,1.518411e-07,1.518484e-07,1.518557e-07,1.518630e-07,1.518703e-07,1.518776e-07,1.518849e-07,1.518922e-07,1.518995e-07,1.519068e-07,1.519141e-07,1.519213e-07,1.519286e-07,1.519359e-07,1.519432e-07,1.519504e-07,1.519577e-07,1.519649e-07,1.519722e-07,1.519794e-07,1.519866e-07,1.519939e-07,1.520011e-07,1.520083e-07,1.520155e-07,1.520227e-07,1.520299e-07,1.520372e-07,1.520444e-07,1.520515e-07,1.520587e-07,1.520659e-07,1.520731e-07,1.520803e-07,1.520875e-07,1.520946e-07,1.521018e-07,1.521089e-07,1.521161e-07,1.521233e-07,1.521304e-07,1.521375e-07,1.521447e-07,1.521518e-07,1.521589e-07,1.521661e-07,1.521732e-07,1.521803e-07,1.521874e-07,1.521945e-07,1.522016e-07,1.522087e-07,1.522158e-07,1.522229e-07,1.522300e-07,1.522371e-07,1.522441e-07,1.522512e-07,1.522583e-07,1.522653e-07,1.522724e-07,1.522794e-07,1.522865e-07,1.522935e-07,1.523006e-07,1.523076e-07,1.523147e-07,1.523217e-07,1.523287e-07,1.523357e-07,1.523427e-07,1.523498e-07,1.523568e-07,1.523638e-07,1.523708e-07,1.523778e-07,1.523847e-07,1.523917e-07,1.523987e-07,1.524057e-07,1.524127e-07,1.524196e-07,1.524266e-07,1.524336e-07,1.524405e-07,1.524475e-07,1.524544e-07,1.524614e-07,1.524683e-07,1.524752e-07,1.524822e-07,1.524891e-07,1.524960e-07,1.525029e-07,1.525098e-07,1.525168e-07,1.525237e-07,1.525306e-07,1.525375e-07,1.525444e-07,1.525512e-07,1.525581e-07,1.525650e-07,1.525719e-07,1.525788e-07,1.525856e-07,1.525925e-07,1.525994e-07,1.526062e-07,1.526131e-07,1.526199e-07,1.526268e-07,1.526336e-07,1.526404e-07,1.526473e-07,1.526541e-07,1.526609e-07,1.526677e-07,1.526746e-07,1.526814e-07,1.526882e-07,1.526950e-07,1.527018e-07,1.527086e-07,1.527154e-07,1.527222e-07,1.527290e-07,1.527357e-07,1.527425e-07,1.527493e-07,1.527561e-07,1.527628e-07,1.527696e-07,1.527763e-07,1.527831e-07,1.527898e-07,1.527966e-07,1.528033e-07,1.528101e-07,1.528168e-07,1.528235e-07,1.528302e-07,1.528370e-07,1.528437e-07,1.528504e-07,1.528571e-07,1.528638e-07,1.528705e-07,1.528772e-07,1.528839e-07,1.528906e-07,1.528973e-07,1.529040e-07,1.529106e-07,1.529173e-07,1.529240e-07,1.529307e-07,1.529373e-07,1.529440e-07,1.529506e-07,1.529573e-07,1.529639e-07,1.529706e-07,1.529772e-07,1.529839e-07,1.529905e-07,1.529971e-07,1.530037e-07,1.530104e-07,1.530170e-07,1.530236e-07,1.530302e-07,1.530368e-07,1.530434e-07,1.530500e-07,1.530566e-07,1.530632e-07,1.530698e-07,1.530764e-07,1.530829e-07,1.530895e-07,1.530961e-07,1.531027e-07,1.531092e-07,1.531158e-07,1.531223e-07,1.531289e-07,1.531354e-07,1.531420e-07,1.531485e-07,1.531551e-07,1.531616e-07,1.531681e-07,1.531747e-07,1.531812e-07,1.531877e-07,1.531942e-07,1.532007e-07,1.532072e-07,1.532138e-07,1.532203e-07,1.532268e-07,1.532332e-07,1.532397e-07,1.532462e-07,1.532527e-07,1.532592e-07,1.532657e-07,1.532721e-07,1.532786e-07,1.532851e-07,1.532915e-07,1.532980e-07,1.533044e-07,1.533109e-07,1.533173e-07,1.533238e-07,1.533302e-07,1.533367e-07,1.533431e-07,1.533495e-07,1.533560e-07,1.533624e-07,1.533688e-07,1.533752e-07,1.533816e-07,1.533880e-07,1.533944e-07,1.534008e-07,1.534072e-07,1.534136e-07,1.534200e-07,1.534264e-07,1.534328e-07,1.534392e-07,1.534455e-07,1.534519e-07,1.534583e-07,1.534646e-07,1.534710e-07,1.534774e-07,1.534837e-07,1.534901e-07,1.534964e-07,1.535028e-07,1.535091e-07,1.535154e-07,1.535218e-07,1.535281e-07,1.535344e-07,1.535408e-07,1.535471e-07,1.535534e-07,1.535597e-07,1.535660e-07,1.535723e-07,1.535786e-07,1.535849e-07,1.535912e-07,1.535975e-07,1.536038e-07,1.536101e-07,1.536164e-07,1.536227e-07,1.536289e-07,1.536352e-07,1.536415e-07,1.536477e-07,1.536540e-07,1.536603e-07,1.536665e-07,1.536728e-07,1.536790e-07,1.536853e-07,1.536915e-07,1.536977e-07,1.537040e-07,1.537102e-07,1.537164e-07,1.537227e-07,1.537289e-07,1.537351e-07,1.537413e-07,1.537475e-07,1.537537e-07,1.537599e-07,1.537661e-07,1.537723e-07,1.537785e-07,1.537847e-07,1.537909e-07,1.537971e-07,1.538033e-07,1.538094e-07,1.538156e-07,1.538218e-07,1.538280e-07,1.538341e-07,1.538403e-07,1.538464e-07,1.538526e-07,1.538588e-07,1.538649e-07,1.538710e-07,1.538772e-07,1.538833e-07,1.538895e-07,1.538956e-07,1.539017e-07,1.539079e-07,1.539140e-07,1.539201e-07,1.539262e-07,1.539323e-07,1.539384e-07,1.539445e-07,1.539506e-07,1.539567e-07,1.539628e-07,1.539689e-07,1.539750e-07,1.539811e-07,1.539872e-07,1.539933e-07,1.539994e-07,1.540054e-07,1.540115e-07,1.540176e-07,1.540236e-07,1.540297e-07,1.540357e-07,1.540418e-07,1.540479e-07,1.540539e-07,1.540599e-07,1.540660e-07,1.540720e-07,1.540781e-07,1.540841e-07,1.540901e-07,1.540962e-07,1.541022e-07,1.541082e-07,1.541142e-07,1.541202e-07,1.541262e-07,1.541322e-07,1.541383e-07,1.541443e-07,1.541503e-07,1.541562e-07,1.541622e-07,1.541682e-07,1.541742e-07,1.541802e-07,1.541862e-07,1.541922e-07,1.541981e-07,1.542041e-07,1.542101e-07,1.542160e-07,1.542220e-07,1.542280e-07,1.542339e-07,1.542399e-07,1.542458e-07,1.542518e-07,1.542577e-07,1.542636e-07,1.542696e-07,1.542755e-07,1.542814e-07,1.542874e-07,1.542933e-07,1.542992e-07,1.543051e-07,1.543110e-07,1.543170e-07,1.543229e-07,1.543288e-07,1.543347e-07,1.543406e-07,1.543465e-07,1.543524e-07,1.543583e-07,1.543641e-07,1.543700e-07,1.543759e-07,1.543818e-07,1.543877e-07,1.543935e-07,1.543994e-07,1.544053e-07,1.544111e-07,1.544170e-07,1.544229e-07,1.544287e-07,1.544346e-07,1.544404e-07,1.544463e-07,1.544521e-07,1.544580e-07,1.544638e-07,1.544696e-07,1.544755e-07,1.544813e-07,1.544871e-07,1.544929e-07,1.544988e-07,1.545046e-07,1.545104e-07,1.545162e-07,1.545220e-07,1.545278e-07,1.545336e-07,1.545394e-07,1.545452e-07,1.545510e-07,1.545568e-07,1.545626e-07,1.545684e-07,1.545742e-07,1.545799e-07,1.545857e-07,1.545915e-07,1.545973e-07,1.546030e-07,1.546088e-07,1.546145e-07,1.546203e-07,1.546261e-07,1.546318e-07,1.546376e-07,1.546433e-07,1.546491e-07,1.546548e-07,1.546605e-07,1.546663e-07,1.546720e-07,1.546777e-07,1.546835e-07,1.546892e-07,1.546949e-07,1.547006e-07,1.547064e-07,1.547121e-07,1.547178e-07,1.547235e-07,1.547292e-07,1.547349e-07,1.547406e-07,1.547463e-07,1.547520e-07,1.547577e-07,1.547634e-07,1.547690e-07,1.547747e-07,1.547804e-07,1.547861e-07,1.547918e-07,1.547974e-07,1.548031e-07,1.548088e-07,1.548144e-07,1.548201e-07,1.548257e-07,1.548314e-07,1.548371e-07,1.548427e-07,1.548483e-07,1.548540e-07,1.548596e-07,1.548653e-07,1.548709e-07,1.548765e-07,1.548822e-07,1.548878e-07,1.548934e-07,1.548990e-07,1.549047e-07,1.549103e-07,1.549159e-07,1.549215e-07,1.549271e-07,1.549327e-07,1.549383e-07,1.549439e-07,1.549495e-07,1.549551e-07,1.549607e-07,1.549663e-07,1.549719e-07,1.549775e-07,1.549830e-07,1.549886e-07,1.549942e-07,1.549998e-07,1.550053e-07,1.550109e-07,1.550165e-07,1.550220e-07,1.550276e-07,1.550332e-07,1.550387e-07,1.550443e-07,1.550498e-07,1.550554e-07,1.550609e-07,1.550664e-07,1.550720e-07,1.550775e-07,1.550830e-07,1.550886e-07,1.550941e-07,1.550996e-07,1.551051e-07,1.551107e-07,1.551162e-07,1.551217e-07,1.551272e-07,1.551327e-07,1.551382e-07,1.551437e-07,1.551492e-07,1.551547e-07,1.551602e-07,1.551657e-07,1.551712e-07,1.551767e-07,1.551822e-07,1.551877e-07,1.551931e-07,1.551986e-07,1.552041e-07,1.552096e-07,1.552150e-07,1.552205e-07,1.552260e-07,1.552314e-07,1.552369e-07,1.552424e-07,1.552478e-07,1.552533e-07,1.552587e-07,1.552642e-07,1.552696e-07,1.552750e-07,1.552805e-07,1.552859e-07,1.552914e-07,1.552968e-07,1.553022e-07,1.553076e-07,1.553131e-07,1.553185e-07,1.553239e-07,1.553293e-07,1.553347e-07,1.553401e-07,1.553456e-07,1.553510e-07,1.553564e-07,1.553618e-07,1.553672e-07,1.553726e-07,1.553780e-07,1.553833e-07,1.553887e-07,1.553941e-07,1.553995e-07,1.554049e-07,1.554103e-07,1.554156e-07,1.554210e-07,1.554264e-07,1.554318e-07,1.554371e-07,1.554425e-07,1.554478e-07,1.554532e-07,1.554586e-07,1.554639e-07,1.554693e-07,1.554746e-07,1.554800e-07,1.554853e-07,1.554906e-07,1.554960e-07,1.555013e-07,1.555066e-07,1.555120e-07,1.555173e-07,1.555226e-07,1.555280e-07,1.555333e-07,1.555386e-07,1.555439e-07,1.555492e-07,1.555545e-07,1.555598e-07,1.555652e-07,1.555705e-07,1.555758e-07,1.555811e-07,1.555864e-07,1.555917e-07,1.555969e-07,1.556022e-07,1.556075e-07,1.556128e-07,1.556181e-07,1.556234e-07,1.556286e-07,1.556339e-07,1.556392e-07,1.556445e-07,1.556497e-07,1.556550e-07,1.556603e-07,1.556655e-07,1.556708e-07,1.556760e-07,1.556813e-07,1.556865e-07,1.556918e-07,1.556970e-07,1.557023e-07,1.557075e-07,1.557128e-07,1.557180e-07,1.557232e-07,1.557285e-07,1.557337e-07,1.557389e-07,1.557442e-07,1.557494e-07,1.557546e-07,1.557598e-07,1.557650e-07,1.557702e-07,1.557755e-07,1.557807e-07,1.557859e-07,1.557911e-07,1.557963e-07,1.558015e-07,1.558067e-07,1.558119e-07,1.558171e-07,1.558222e-07,1.558274e-07,1.558326e-07,1.558378e-07,1.558430e-07,1.558482e-07,1.558533e-07,1.558585e-07,1.558637e-07,1.558689e-07,1.558740e-07,1.558792e-07,1.558843e-07,1.558895e-07,1.558947e-07,1.558998e-07,1.559050e-07,1.559101e-07,1.559153e-07,1.559204e-07,1.559256e-07,1.559307e-07,1.559358e-07,1.559410e-07,1.559461e-07,1.559512e-07,1.559564e-07,1.559615e-07,1.559666e-07,1.559717e-07,1.559769e-07,1.559820e-07,1.559871e-07,1.559922e-07,1.559973e-07,1.560024e-07,1.560075e-07,1.560127e-07,1.560178e-07,1.560229e-07,1.560280e-07,1.560331e-07,1.560381e-07,1.560432e-07,1.560483e-07,1.560534e-07,1.560585e-07,1.560636e-07,1.560687e-07,1.560737e-07,1.560788e-07,1.560839e-07,1.560890e-07,1.560940e-07,1.560991e-07,1.561042e-07,1.561092e-07,1.561143e-07,1.561193e-07,1.561244e-07,1.561295e-07,1.561345e-07,1.561396e-07,1.561446e-07,1.561496e-07,1.561547e-07,1.561597e-07,1.561648e-07,1.561698e-07,1.561748e-07,1.561799e-07,1.561849e-07,1.561899e-07,1.561950e-07,1.562000e-07,1.562050e-07,1.562100e-07,1.562150e-07,1.562200e-07,1.562251e-07,1.562301e-07,1.562351e-07,1.562401e-07,1.562451e-07,1.562501e-07,1.562551e-07,1.562601e-07,1.562651e-07,1.562701e-07,1.562751e-07,1.562800e-07,1.562850e-07,1.562900e-07,1.562950e-07,1.563000e-07,1.563050e-07,1.563099e-07,1.563149e-07,1.563199e-07,1.563248e-07,1.563298e-07,1.563348e-07,1.563397e-07,1.563447e-07,1.563497e-07,1.563546e-07,1.563596e-07,1.563645e-07,1.563695e-07,1.563744e-07,1.563794e-07,1.563843e-07,1.563893e-07,1.563942e-07,1.563991e-07,1.564041e-07,1.564090e-07,1.564139e-07,1.564189e-07,1.564238e-07,1.564287e-07,1.564336e-07,1.564386e-07,1.564435e-07,1.564484e-07,1.564533e-07,1.564582e-07,1.564631e-07,1.564680e-07,1.564729e-07,1.564778e-07,1.564827e-07,1.564876e-07,1.564925e-07,1.564974e-07,1.565023e-07,1.565072e-07,1.565121e-07,1.565170e-07,1.565219e-07,1.565268e-07,1.565316e-07,1.565365e-07,1.565414e-07,1.565463e-07,1.565511e-07,1.565560e-07,1.565609e-07,1.565658e-07,1.565706e-07,1.565755e-07,1.565803e-07,1.565852e-07,1.565901e-07,1.565949e-07,1.565998e-07,1.566046e-07,1.566095e-07,1.566143e-07,1.566191e-07,1.566240e-07,1.566288e-07,1.566337e-07,1.566385e-07,1.566433e-07,1.566482e-07,1.566530e-07,1.566578e-07,1.566627e-07,1.566675e-07,1.566723e-07,1.566771e-07,1.566819e-07,1.566868e-07,1.566916e-07,1.566964e-07,1.567012e-07,1.567060e-07,1.567108e-07,1.567156e-07,1.567204e-07,1.567252e-07,1.567300e-07,1.567348e-07,1.567396e-07,1.567444e-07,1.567492e-07,1.567540e-07,1.567588e-07,1.567635e-07,1.567683e-07,1.567731e-07,1.567779e-07,1.567827e-07,1.567874e-07,1.567922e-07,1.567970e-07,1.568017e-07,1.568065e-07,1.568113e-07,1.568160e-07,1.568208e-07,1.568255e-07,1.568303e-07,1.568351e-07,1.568398e-07,1.568446e-07,1.568493e-07,1.568541e-07,1.568588e-07,1.568635e-07,1.568683e-07,1.568730e-07,1.568778e-07,1.568825e-07,1.568872e-07,1.568920e-07,1.568967e-07,1.569014e-07,1.569061e-07,1.569109e-07,1.569156e-07,1.569203e-07,1.569250e-07,1.569297e-07,1.569345e-07,1.569392e-07,1.569439e-07,1.569486e-07,1.569533e-07,1.569580e-07,1.569627e-07,1.569674e-07,1.569721e-07,1.569768e-07,1.569815e-07,1.569862e-07,1.569909e-07,1.569956e-07,1.570002e-07,1.570049e-07,1.570096e-07,1.570143e-07,1.570190e-07,1.570237e-07,1.570283e-07,1.570330e-07,1.570377e-07,1.570423e-07,1.570470e-07,1.570517e-07,1.570563e-07,1.570610e-07,1.570657e-07,1.570703e-07,1.570750e-07,1.570796e-07,1.570843e-07,1.570889e-07,1.570936e-07,1.570982e-07,1.571029e-07,1.571075e-07,1.571122e-07,1.571168e-07,1.571214e-07,1.571261e-07,1.571307e-07,1.571353e-07,1.571400e-07,1.571446e-07,1.571492e-07,1.571539e-07,1.571585e-07,1.571631e-07,1.571677e-07,1.571723e-07,1.571770e-07,1.571816e-07,1.571862e-07,1.571908e-07,1.571954e-07,1.572000e-07,1.572046e-07,1.572092e-07,1.572138e-07,1.572184e-07,1.572230e-07,1.572276e-07,1.572322e-07,1.572368e-07,1.572414e-07,1.572460e-07,1.572506e-07,1.572551e-07,1.572597e-07,1.572643e-07,1.572689e-07,1.572735e-07,1.572780e-07,1.572826e-07,1.572872e-07,1.572918e-07,1.572963e-07,1.573009e-07,1.573055e-07,1.573100e-07,1.573146e-07,1.573191e-07,1.573237e-07,1.573283e-07,1.573328e-07,1.573374e-07,1.573419e-07,1.573465e-07,1.573510e-07,1.573556e-07,1.573601e-07,1.573646e-07,1.573692e-07,1.573737e-07,1.573783e-07,1.573828e-07,1.573873e-07,1.573919e-07,1.573964e-07,1.574009e-07,1.574054e-07,1.574100e-07,1.574145e-07,1.574190e-07,1.574235e-07,1.574280e-07,1.574325e-07,1.574371e-07,1.574416e-07,1.574461e-07,1.574506e-07,1.574551e-07,1.574596e-07,1.574641e-07,1.574686e-07,1.574731e-07,1.574776e-07,1.574821e-07,1.574866e-07,1.574911e-07,1.574956e-07,1.575001e-07,1.575046e-07,1.575090e-07,1.575135e-07,1.575180e-07,1.575225e-07,1.575270e-07,1.575314e-07,1.575359e-07,1.575404e-07,1.575449e-07,1.575493e-07,1.575538e-07,1.575583e-07,1.575627e-07,1.575672e-07,1.575716e-07,1.575761e-07,1.575806e-07,1.575850e-07,1.575895e-07,1.575939e-07,1.575984e-07,1.576028e-07,1.576073e-07,1.576117e-07,1.576162e-07,1.576206e-07,1.576250e-07,1.576295e-07,1.576339e-07,1.576384e-07,1.576428e-07,1.576472e-07,1.576517e-07,1.576561e-07,1.576605e-07,1.576649e-07,1.576694e-07,1.576738e-07,1.576782e-07,1.576826e-07,1.576870e-07,1.576914e-07,1.576959e-07,1.577003e-07,1.577047e-07,1.577091e-07,1.577135e-07,1.577179e-07,1.577223e-07,1.577267e-07,1.577311e-07,1.577355e-07,1.577399e-07,1.577443e-07,1.577487e-07,1.577531e-07,1.577575e-07,1.577619e-07,1.577662e-07,1.577706e-07,1.577750e-07,1.577794e-07,1.577838e-07,1.577882e-07,1.577925e-07,1.577969e-07,1.578013e-07,1.578056e-07,1.578100e-07,1.578144e-07,1.578188e-07,1.578231e-07,1.578275e-07,1.578318e-07,1.578362e-07,1.578406e-07,1.578449e-07,1.578493e-07,1.578536e-07,1.578580e-07,1.578623e-07,1.578667e-07,1.578710e-07,1.578754e-07,1.578797e-07,1.578841e-07,1.578884e-07,1.578927e-07,1.578971e-07,1.579014e-07,1.579057e-07,1.579101e-07,1.579144e-07,1.579187e-07,1.579231e-07,1.579274e-07,1.579317e-07,1.579360e-07,1.579404e-07,1.579447e-07,1.579490e-07,1.579533e-07,1.579576e-07,1.579619e-07,1.579662e-07,1.579706e-07,1.579749e-07,1.579792e-07,1.579835e-07,1.579878e-07,1.579921e-07,1.579964e-07,1.580007e-07,1.580050e-07,1.580093e-07,1.580136e-07,1.580179e-07,1.580221e-07,1.580264e-07,1.580307e-07,1.580350e-07,1.580393e-07,1.580436e-07,1.580479e-07,1.580521e-07,1.580564e-07,1.580607e-07,1.580650e-07,1.580692e-07,1.580735e-07,1.580778e-07,1.580820e-07,1.580863e-07,1.580906e-07,1.580948e-07,1.580991e-07,1.581034e-07,1.581076e-07,1.581119e-07,1.581161e-07,1.581204e-07,1.581246e-07,1.581289e-07,1.581331e-07,1.581374e-07,1.581416e-07,1.581459e-07,1.581501e-07,1.581544e-07,1.581586e-07,1.581628e-07,1.581671e-07,1.581713e-07,1.581756e-07,1.581798e-07,1.581840e-07,1.581882e-07,1.581925e-07,1.581967e-07,1.582009e-07,1.582051e-07,1.582094e-07,1.582136e-07,1.582178e-07,1.582220e-07,1.582262e-07,1.582305e-07,1.582347e-07,1.582389e-07,1.582431e-07,1.582473e-07,1.582515e-07,1.582557e-07,1.582599e-07,1.582641e-07,1.582683e-07,1.582725e-07,1.582767e-07,1.582809e-07,1.582851e-07,1.582893e-07,1.582935e-07,1.582977e-07,1.583019e-07,1.583060e-07,1.583102e-07,1.583144e-07,1.583186e-07,1.583228e-07,1.583270e-07,1.583311e-07,1.583353e-07,1.583395e-07,1.583437e-07,1.583478e-07,1.583520e-07,1.583562e-07,1.583603e-07,1.583645e-07,1.583687e-07,1.583728e-07,1.583770e-07,1.583811e-07,1.583853e-07,1.583895e-07,1.583936e-07,1.583978e-07,1.584019e-07,1.584061e-07,1.584102e-07,1.584144e-07,1.584185e-07,1.584227e-07,1.584268e-07,1.584309e-07,1.584351e-07,1.584392e-07,1.584434e-07,1.584475e-07,1.584516e-07,1.584558e-07,1.584599e-07,1.584640e-07,1.584681e-07,1.584723e-07,1.584764e-07,1.584805e-07,1.584846e-07,1.584888e-07,1.584929e-07,1.584970e-07,1.585011e-07,1.585052e-07,1.585093e-07,1.585135e-07,1.585176e-07,1.585217e-07,1.585258e-07,1.585299e-07,1.585340e-07,1.585381e-07,1.585422e-07,1.585463e-07,1.585504e-07,1.585545e-07,1.585586e-07,1.585627e-07,1.585668e-07,1.585709e-07,1.585750e-07,1.585791e-07,1.585831e-07,1.585872e-07,1.585913e-07,1.585954e-07,1.585995e-07,1.586036e-07,1.586076e-07,1.586117e-07,1.586158e-07,1.586199e-07,1.586239e-07,1.586280e-07,1.586321e-07,1.586361e-07,1.586402e-07,1.586443e-07,1.586483e-07,1.586524e-07,1.586565e-07,1.586605e-07,1.586646e-07,1.586686e-07,1.586727e-07,1.586768e-07,1.586808e-07,1.586849e-07,1.586889e-07,1.586930e-07,1.586970e-07,1.587011e-07,1.587051e-07,1.587091e-07,1.587132e-07,1.587172e-07,1.587213e-07,1.587253e-07,1.587293e-07,1.587334e-07,1.587374e-07,1.587414e-07,1.587455e-07,1.587495e-07,1.587535e-07,1.587575e-07,1.587616e-07,1.587656e-07,1.587696e-07,1.587736e-07,1.587777e-07,1.587817e-07,1.587857e-07,1.587897e-07,1.587937e-07,1.587977e-07,1.588017e-07,1.588058e-07,1.588098e-07,1.588138e-07,1.588178e-07,1.588218e-07,1.588258e-07,1.588298e-07,1.588338e-07,1.588378e-07,1.588418e-07,1.588458e-07,1.588498e-07,1.588538e-07,1.588577e-07,1.588617e-07,1.588657e-07,1.588697e-07,1.588737e-07,1.588777e-07,1.588817e-07,1.588857e-07,1.588896e-07,1.588936e-07,1.588976e-07,1.589016e-07,1.589055e-07,1.589095e-07,1.589135e-07,1.589175e-07,1.589214e-07,1.589254e-07,1.589294e-07,1.589333e-07,1.589373e-07,1.589413e-07,1.589452e-07,1.589492e-07,1.589531e-07,1.589571e-07,1.589610e-07,1.589650e-07,1.589690e-07,1.589729e-07,1.589769e-07,1.589808e-07,1.589848e-07,1.589887e-07,1.589926e-07,1.589966e-07,1.590005e-07,1.590045e-07,1.590084e-07,1.590124e-07,1.590163e-07,1.590202e-07,1.590242e-07,1.590281e-07,1.590320e-07,1.590360e-07,1.590399e-07,1.590438e-07,1.590477e-07,1.590517e-07,1.590556e-07,1.590595e-07,1.590634e-07,1.590673e-07,1.590713e-07,1.590752e-07,1.590791e-07,1.590830e-07,1.590869e-07,1.590908e-07,1.590948e-07,1.590987e-07,1.591026e-07,1.591065e-07,1.591104e-07,1.591143e-07,1.591182e-07,1.591221e-07,1.591260e-07,1.591299e-07,1.591338e-07,1.591377e-07,1.591416e-07,1.591455e-07,1.591494e-07,1.591533e-07,1.591571e-07,1.591610e-07,1.591649e-07,1.591688e-07,1.591727e-07,1.591766e-07,1.591805e-07,1.591843e-07,1.591882e-07,1.591921e-07,1.591960e-07,1.591998e-07,1.592037e-07,1.592076e-07,1.592115e-07,1.592153e-07,1.592192e-07,1.592231e-07,1.592269e-07,1.592308e-07,1.592347e-07,1.592385e-07,1.592424e-07,1.592462e-07,1.592501e-07,1.592540e-07,1.592578e-07,1.592617e-07,1.592655e-07,1.592694e-07,1.592732e-07,1.592771e-07,1.592809e-07,1.592848e-07,1.592886e-07,1.592925e-07,1.592963e-07,1.593001e-07,1.593040e-07,1.593078e-07,1.593117e-07,1.593155e-07,1.593193e-07,1.593232e-07,1.593270e-07,1.593308e-07,1.593347e-07,1.593385e-07,1.593423e-07,1.593461e-07,1.593500e-07,1.593538e-07,1.593576e-07,1.593614e-07,1.593653e-07,1.593691e-07,1.593729e-07,1.593767e-07,1.593805e-07,1.593843e-07,1.593882e-07,1.593920e-07,1.593958e-07,1.593996e-07,1.594034e-07,1.594072e-07,1.594110e-07,1.594148e-07,1.594186e-07,1.594224e-07,1.594262e-07,1.594300e-07,1.594338e-07,1.594376e-07,1.594414e-07,1.594452e-07,1.594490e-07,1.594528e-07,1.594566e-07,1.594604e-07,1.594641e-07,1.594679e-07,1.594717e-07,1.594755e-07,1.594793e-07,1.594831e-07,1.594868e-07,1.594906e-07,1.594944e-07,1.594982e-07,1.595019e-07,1.595057e-07,1.595095e-07,1.595133e-07,1.595170e-07,1.595208e-07,1.595246e-07,1.595283e-07,1.595321e-07,1.595359e-07,1.595396e-07,1.595434e-07,1.595472e-07,1.595509e-07,1.595547e-07,1.595584e-07,1.595622e-07,1.595659e-07,1.595697e-07,1.595734e-07,1.595772e-07,1.595809e-07,1.595847e-07,1.595884e-07,1.595922e-07,1.595959e-07,1.595997e-07,1.596034e-07,1.596072e-07,1.596109e-07,1.596146e-07,1.596184e-07,1.596221e-07,1.596258e-07,1.596296e-07,1.596333e-07,1.596370e-07,1.596408e-07,1.596445e-07,1.596482e-07,1.596520e-07,1.596557e-07,1.596594e-07,1.596631e-07,1.596669e-07,1.596706e-07,1.596743e-07,1.596780e-07,1.596817e-07,1.596854e-07,1.596892e-07,1.596929e-07,1.596966e-07,1.597003e-07,1.597040e-07,1.597077e-07,1.597114e-07,1.597151e-07,1.597188e-07,1.597225e-07,1.597262e-07,1.597299e-07,1.597336e-07,1.597373e-07,1.597410e-07,1.597447e-07,1.597484e-07,1.597521e-07,1.597558e-07,1.597595e-07,1.597632e-07,1.597669e-07,1.597706e-07,1.597743e-07,1.597780e-07,1.597816e-07,1.597853e-07,1.597890e-07,1.597927e-07,1.597964e-07,1.598001e-07,1.598037e-07,1.598074e-07,1.598111e-07,1.598148e-07,1.598184e-07,1.598221e-07,1.598258e-07,1.598294e-07,1.598331e-07,1.598368e-07,1.598404e-07,1.598441e-07,1.598478e-07,1.598514e-07,1.598551e-07,1.598588e-07,1.598624e-07,1.598661e-07,1.598697e-07,1.598734e-07,1.598770e-07,1.598807e-07,1.598844e-07,1.598880e-07,1.598917e-07,1.598953e-07,1.598990e-07,1.599026e-07,1.599062e-07,1.599099e-07,1.599135e-07,1.599172e-07,1.599208e-07,1.599245e-07,1.599281e-07,1.599317e-07,1.599354e-07,1.599390e-07,1.599426e-07,1.599463e-07,1.599499e-07,1.599535e-07,1.599572e-07,1.599608e-07,1.599644e-07,1.599680e-07,1.599717e-07,1.599753e-07,1.599789e-07,1.599825e-07,1.599862e-07,1.599898e-07,1.599934e-07,1.599970e-07,1.600006e-07,1.600042e-07,1.600079e-07,1.600115e-07,1.600151e-07,1.600187e-07,1.600223e-07,1.600259e-07,1.600295e-07,1.600331e-07,1.600367e-07,1.600403e-07,1.600439e-07,1.600475e-07,1.600511e-07,1.600547e-07,1.600583e-07,1.600619e-07,1.600655e-07,1.600691e-07,1.600727e-07,1.600763e-07,1.600799e-07,1.600835e-07,1.600871e-07,1.600907e-07,1.600943e-07,1.600978e-07,1.601014e-07,1.601050e-07,1.601086e-07,1.601122e-07,1.601158e-07,1.601193e-07,1.601229e-07,1.601265e-07,1.601301e-07,1.601336e-07,1.601372e-07,1.601408e-07,1.601444e-07,1.601479e-07,1.601515e-07,1.601551e-07,1.601586e-07,1.601622e-07,1.601658e-07,1.601693e-07,1.601729e-07,1.601764e-07,1.601800e-07,1.601836e-07,1.601871e-07,1.601907e-07,1.601942e-07,1.601978e-07,1.602013e-07,1.602049e-07,1.602085e-07,1.602120e-07,1.602156e-07,1.602191e-07,1.602226e-07,1.602262e-07,1.602297e-07,1.602333e-07,1.602368e-07,1.602404e-07,1.602439e-07,1.602475e-07,1.602510e-07,1.602545e-07,1.602581e-07,1.602616e-07,1.602651e-07,1.602687e-07,1.602722e-07,1.602757e-07,1.602793e-07,1.602828e-07,1.602863e-07,1.602898e-07,1.602934e-07,1.602969e-07,1.603004e-07,1.603039e-07,1.603075e-07,1.603110e-07,1.603145e-07,1.603180e-07,1.603215e-07,1.603251e-07,1.603286e-07,1.603321e-07,1.603356e-07,1.603391e-07,1.603426e-07,1.603461e-07,1.603496e-07,1.603531e-07,1.603566e-07,1.603602e-07,1.603637e-07,1.603672e-07,1.603707e-07,1.603742e-07,1.603777e-07,1.603812e-07,1.603847e-07,1.603882e-07,1.603917e-07,1.603952e-07,1.603986e-07,1.604021e-07,1.604056e-07,1.604091e-07,1.604126e-07,1.604161e-07,1.604196e-07,1.604231e-07,1.604266e-07,1.604300e-07,1.604335e-07,1.604370e-07,1.604405e-07,1.604440e-07,1.604474e-07,1.604509e-07,1.604544e-07,1.604579e-07,1.604614e-07,1.604648e-07,1.604683e-07,1.604718e-07,1.604752e-07,1.604787e-07,1.604822e-07,1.604857e-07,1.604891e-07,1.604926e-07,1.604960e-07,1.604995e-07,1.605030e-07,1.605064e-07,1.605099e-07,1.605134e-07,1.605168e-07,1.605203e-07,1.605237e-07,1.605272e-07,1.605306e-07,1.605341e-07,1.605375e-07,1.605410e-07,1.605444e-07,1.605479e-07,1.605513e-07,1.605548e-07,1.605582e-07,1.605617e-07,1.605651e-07,1.605686e-07,1.605720e-07,1.605754e-07,1.605789e-07,1.605823e-07,1.605858e-07,1.605892e-07,1.605926e-07,1.605961e-07,1.605995e-07,1.606029e-07,1.606064e-07,1.606098e-07,1.606132e-07,1.606167e-07,1.606201e-07,1.606235e-07,1.606269e-07,1.606304e-07,1.606338e-07,1.606372e-07,1.606406e-07,1.606441e-07,1.606475e-07,1.606509e-07,1.606543e-07,1.606577e-07,1.606611e-07,1.606646e-07,1.606680e-07,1.606714e-07,1.606748e-07,1.606782e-07,1.606816e-07,1.606850e-07,1.606884e-07,1.606918e-07,1.606952e-07,1.606986e-07,1.607020e-07,1.607054e-07,1.607088e-07,1.607123e-07,1.607156e-07,1.607190e-07,1.607224e-07,1.607258e-07,1.607292e-07,1.607326e-07,1.607360e-07,1.607394e-07,1.607428e-07,1.607462e-07,1.607496e-07,1.607530e-07,1.607564e-07,1.607598e-07,1.607631e-07,1.607665e-07,1.607699e-07,1.607733e-07,1.607767e-07,1.607801e-07,1.607834e-07,1.607868e-07,1.607902e-07,1.607936e-07,1.607969e-07,1.608003e-07,1.608037e-07,1.608071e-07,1.608104e-07,1.608138e-07,1.608172e-07,1.608205e-07,1.608239e-07,1.608273e-07,1.608306e-07,1.608340e-07,1.608374e-07,1.608407e-07,1.608441e-07,1.608475e-07,1.608508e-07,1.608542e-07,1.608575e-07,1.608609e-07,1.608642e-07,1.608676e-07,1.608710e-07,1.608743e-07,1.608777e-07,1.608810e-07,1.608844e-07,1.608877e-07,1.608911e-07,1.608944e-07,1.608978e-07,1.609011e-07,1.609044e-07,1.609078e-07,1.609111e-07,1.609145e-07,1.609178e-07,1.609212e-07,1.609245e-07,1.609278e-07,1.609312e-07,1.609345e-07,1.609378e-07,1.609412e-07,1.609445e-07,1.609478e-07,1.609512e-07,1.609545e-07,1.609578e-07,1.609612e-07,1.609645e-07,1.609678e-07,1.609711e-07,1.609745e-07,1.609778e-07,1.609811e-07,1.609844e-07,1.609877e-07,1.609911e-07,1.609944e-07,1.609977e-07,1.610010e-07,1.610043e-07,1.610076e-07,1.610110e-07,1.610143e-07,1.610176e-07,1.610209e-07,1.610242e-07,1.610275e-07,1.610308e-07,1.610341e-07,1.610374e-07,1.610407e-07,1.610440e-07,1.610473e-07,1.610507e-07,1.610540e-07,1.610573e-07,1.610606e-07,1.610639e-07,1.610672e-07,1.610704e-07,1.610737e-07,1.610770e-07,1.610803e-07,1.610836e-07,1.610869e-07,1.610902e-07,1.610935e-07,1.610968e-07,1.611001e-07,1.611034e-07,1.611067e-07,1.611099e-07,1.611132e-07,1.611165e-07,1.611198e-07,1.611231e-07,1.611264e-07,1.611296e-07,1.611329e-07,1.611362e-07,1.611395e-07,1.611427e-07,1.611460e-07,1.611493e-07,1.611526e-07,1.611558e-07,1.611591e-07,1.611624e-07,1.611657e-07,1.611689e-07,1.611722e-07,1.611755e-07,1.611787e-07,1.611820e-07,1.611852e-07,1.611885e-07,1.611918e-07,1.611950e-07,1.611983e-07,1.612016e-07,1.612048e-07,1.612081e-07,1.612113e-07,1.612146e-07,1.612178e-07,1.612211e-07,1.612244e-07,1.612276e-07,1.612309e-07,1.612341e-07,1.612374e-07,1.612406e-07,1.612439e-07,1.612471e-07,1.612503e-07,1.612536e-07,1.612568e-07,1.612601e-07,1.612633e-07,1.612666e-07,1.612698e-07,1.612730e-07,1.612763e-07,1.612795e-07,1.612828e-07,1.612860e-07,1.612892e-07,1.612925e-07,1.612957e-07,1.612989e-07,1.613022e-07,1.613054e-07,1.613086e-07,1.613118e-07,1.613151e-07,1.613183e-07,1.613215e-07,1.613248e-07,1.613280e-07,1.613312e-07,1.613344e-07,1.613376e-07,1.613409e-07,1.613441e-07,1.613473e-07,1.613505e-07,1.613537e-07,1.613570e-07,1.613602e-07,1.613634e-07,1.613666e-07,1.613698e-07,1.613730e-07,1.613762e-07,1.613794e-07,1.613827e-07,1.613859e-07,1.613891e-07,1.613923e-07,1.613955e-07,1.613987e-07,1.614019e-07,1.614051e-07,1.614083e-07,1.614115e-07,1.614147e-07,1.614179e-07,1.614211e-07,1.614243e-07,1.614275e-07,1.614307e-07,1.614339e-07,1.614371e-07,1.614403e-07,1.614435e-07,1.614467e-07,1.614498e-07,1.614530e-07,1.614562e-07,1.614594e-07,1.614626e-07,1.614658e-07,1.614690e-07,1.614722e-07,1.614753e-07,1.614785e-07,1.614817e-07,1.614849e-07,1.614881e-07,1.614912e-07,1.614944e-07,1.614976e-07,1.615008e-07,1.615039e-07,1.615071e-07,1.615103e-07,1.615135e-07,1.615166e-07,1.615198e-07,1.615230e-07,1.615262e-07,1.615293e-07,1.615325e-07,1.615357e-07,1.615388e-07,1.615420e-07,1.615452e-07,1.615483e-07,1.615515e-07,1.615546e-07,1.615578e-07,1.615610e-07,1.615641e-07,1.615673e-07,1.615704e-07,1.615736e-07,1.615767e-07,1.615799e-07,1.615831e-07,1.615862e-07,1.615894e-07,1.615925e-07,1.615957e-07,1.615988e-07,1.616020e-07,1.616051e-07,1.616083e-07,1.616114e-07,1.616146e-07,1.616177e-07,1.616208e-07,1.616240e-07,1.616271e-07,1.616303e-07,1.616334e-07,1.616365e-07,1.616397e-07,1.616428e-07,1.616460e-07,1.616491e-07,1.616522e-07,1.616554e-07,1.616585e-07,1.616616e-07,1.616648e-07,1.616679e-07,1.616710e-07,1.616742e-07,1.616773e-07,1.616804e-07,1.616835e-07,1.616867e-07,1.616898e-07,1.616929e-07,1.616960e-07,1.616992e-07,1.617023e-07,1.617054e-07,1.617085e-07,1.617116e-07,1.617148e-07,1.617179e-07,1.617210e-07,1.617241e-07,1.617272e-07,1.617303e-07,1.617335e-07,1.617366e-07,1.617397e-07,1.617428e-07,1.617459e-07,1.617490e-07,1.617521e-07,1.617552e-07,1.617583e-07,1.617614e-07,1.617645e-07,1.617676e-07,1.617707e-07,1.617739e-07,1.617770e-07,1.617801e-07,1.617832e-07,1.617863e-07,1.617894e-07,1.617925e-07,1.617955e-07,1.617986e-07,1.618017e-07,1.618048e-07,1.618079e-07,1.618110e-07,1.618141e-07,1.618172e-07,1.618203e-07,1.618234e-07,1.618265e-07,1.618296e-07,1.618326e-07,1.618357e-07,1.618388e-07,1.618419e-07,1.618450e-07,1.618481e-07,1.618511e-07,1.618542e-07,1.618573e-07,1.618604e-07,1.618635e-07,1.618665e-07,1.618696e-07,1.618727e-07,1.618758e-07,1.618788e-07,1.618819e-07,1.618850e-07,1.618881e-07,1.618911e-07,1.618942e-07,1.618973e-07,1.619003e-07,1.619034e-07,1.619065e-07,1.619095e-07,1.619126e-07,1.619157e-07,1.619187e-07,1.619218e-07,1.619249e-07,1.619279e-07,1.619310e-07,1.619341e-07,1.619371e-07,1.619402e-07,1.619432e-07,1.619463e-07,1.619493e-07,1.619524e-07,1.619554e-07,1.619585e-07,1.619616e-07,1.619646e-07,1.619677e-07,1.619707e-07,1.619738e-07,1.619768e-07,1.619799e-07,1.619829e-07,1.619859e-07,1.619890e-07,1.619920e-07,1.619951e-07,1.619981e-07,1.620012e-07,1.620042e-07,1.620072e-07,1.620103e-07,1.620133e-07,1.620164e-07,1.620194e-07,1.620224e-07,1.620255e-07,1.620285e-07,1.620315e-07,1.620346e-07,1.620376e-07,1.620406e-07,1.620437e-07,1.620467e-07,1.620497e-07,1.620528e-07,1.620558e-07,1.620588e-07,1.620618e-07,1.620649e-07,1.620679e-07,1.620709e-07,1.620739e-07,1.620770e-07,1.620800e-07,1.620830e-07,1.620860e-07,1.620890e-07,1.620921e-07,1.620951e-07,1.620981e-07,1.621011e-07,1.621041e-07,1.621071e-07,1.621102e-07,1.621132e-07,1.621162e-07,1.621192e-07,1.621222e-07,1.621252e-07,1.621282e-07,1.621312e-07,1.621342e-07,1.621372e-07,1.621403e-07,1.621433e-07,1.621463e-07,1.621493e-07,1.621523e-07,1.621553e-07,1.621583e-07,1.621613e-07,1.621643e-07,1.621673e-07,1.621703e-07,1.621733e-07,1.621763e-07,1.621793e-07,1.621823e-07,1.621852e-07,1.621882e-07,1.621912e-07,1.621942e-07,1.621972e-07,1.622002e-07,1.622032e-07,1.622062e-07,1.622092e-07,1.622122e-07,1.622151e-07,1.622181e-07,1.622211e-07,1.622241e-07,1.622271e-07,1.622301e-07,1.622331e-07,1.622360e-07,1.622390e-07,1.622420e-07,1.622450e-07,1.622480e-07,1.622509e-07,1.622539e-07,1.622569e-07,1.622599e-07,1.622628e-07,1.622658e-07,1.622688e-07,1.622717e-07,1.622747e-07,1.622777e-07,1.622807e-07,1.622836e-07,1.622866e-07,1.622896e-07,1.622925e-07,1.622955e-07,1.622985e-07,1.623014e-07,1.623044e-07,1.623074e-07,1.623103e-07,1.623133e-07,1.623162e-07,1.623192e-07,1.623222e-07,1.623251e-07,1.623281e-07,1.623310e-07,1.623340e-07,1.623369e-07,1.623399e-07,1.623428e-07,1.623458e-07,1.623488e-07,1.623517e-07,1.623547e-07,1.623576e-07,1.623606e-07,1.623635e-07,1.623665e-07,1.623694e-07,1.623723e-07,1.623753e-07,1.623782e-07,1.623812e-07,1.623841e-07,1.623871e-07,1.623900e-07,1.623929e-07,1.623959e-07,1.623988e-07,1.624018e-07,1.624047e-07,1.624076e-07,1.624106e-07,1.624135e-07,1.624165e-07,1.624194e-07,1.624223e-07,1.624253e-07,1.624282e-07,1.624311e-07,1.624340e-07,1.624370e-07,1.624399e-07,1.624428e-07,1.624458e-07,1.624487e-07,1.624516e-07,1.624545e-07,1.624575e-07,1.624604e-07,1.624633e-07,1.624662e-07,1.624692e-07,1.624721e-07,1.624750e-07,1.624779e-07,1.624808e-07,1.624838e-07,1.624867e-07,1.624896e-07,1.624925e-07,1.624954e-07,1.624983e-07,1.625012e-07,1.625042e-07,1.625071e-07,1.625100e-07,1.625129e-07,1.625158e-07,1.625187e-07,1.625216e-07,1.625245e-07,1.625274e-07,1.625303e-07,1.625333e-07,1.625362e-07,1.625391e-07,1.625420e-07,1.625449e-07,1.625478e-07,1.625507e-07,1.625536e-07,1.625565e-07,1.625594e-07,1.625623e-07,1.625652e-07,1.625681e-07,1.625710e-07,1.625739e-07,1.625767e-07,1.625796e-07,1.625825e-07,1.625854e-07,1.625883e-07,1.625912e-07,1.625941e-07,1.625970e-07,1.625999e-07,1.626028e-07,1.626057e-07,1.626085e-07,1.626114e-07,1.626143e-07,1.626172e-07,1.626201e-07,1.626230e-07,1.626259e-07,1.626287e-07,1.626316e-07,1.626345e-07,1.626374e-07,1.626403e-07,1.626431e-07,1.626460e-07,1.626489e-07,1.626518e-07,1.626546e-07,1.626575e-07,1.626604e-07,1.626633e-07,1.626661e-07,1.626690e-07,1.626719e-07,1.626747e-07,1.626776e-07,1.626805e-07,1.626834e-07,1.626862e-07,1.626891e-07,1.626920e-07,1.626948e-07,1.626977e-07,1.627005e-07,1.627034e-07,1.627063e-07,1.627091e-07,1.627120e-07,1.627149e-07,1.627177e-07,1.627206e-07,1.627234e-07,1.627263e-07,1.627291e-07,1.627320e-07,1.627349e-07,1.627377e-07,1.627406e-07,1.627434e-07,1.627463e-07,1.627491e-07,1.627520e-07,1.627548e-07,1.627577e-07,1.627605e-07,1.627634e-07,1.627662e-07,1.627691e-07,1.627719e-07,1.627748e-07,1.627776e-07,1.627805e-07,1.627833e-07,1.627861e-07,1.627890e-07,1.627918e-07,1.627947e-07,1.627975e-07,1.628003e-07,1.628032e-07,1.628060e-07,1.628089e-07,1.628117e-07,1.628145e-07,1.628174e-07,1.628202e-07,1.628230e-07,1.628259e-07,1.628287e-07,1.628315e-07,1.628344e-07,1.628372e-07,1.628400e-07,1.628429e-07,1.628457e-07,1.628485e-07,1.628513e-07,1.628542e-07,1.628570e-07,1.628598e-07,1.628626e-07,1.628655e-07,1.628683e-07,1.628711e-07,1.628739e-07,1.628767e-07,1.628796e-07,1.628824e-07,1.628852e-07,1.628880e-07,1.628908e-07,1.628937e-07,1.628965e-07,1.628993e-07,1.629021e-07,1.629049e-07,1.629077e-07,1.629105e-07,1.629134e-07,1.629162e-07,1.629190e-07,1.629218e-07,1.629246e-07,1.629274e-07,1.629302e-07,1.629330e-07,1.629358e-07,1.629386e-07,1.629414e-07,1.629442e-07,1.629470e-07,1.629498e-07,1.629527e-07,1.629555e-07,1.629583e-07,1.629611e-07,1.629639e-07,1.629667e-07,1.629695e-07,1.629722e-07,1.629750e-07,1.629778e-07,1.629806e-07,1.629834e-07,1.629862e-07,1.629890e-07,1.629918e-07,1.629946e-07,1.629974e-07,1.630002e-07,1.630030e-07,1.630058e-07,1.630086e-07,1.630113e-07,1.630141e-07,1.630169e-07,1.630197e-07,1.630225e-07,1.630253e-07,1.630281e-07,1.630308e-07,1.630336e-07,1.630364e-07,1.630392e-07,1.630420e-07,1.630448e-07,1.630475e-07,1.630503e-07,1.630531e-07,1.630559e-07,1.630586e-07,1.630614e-07,1.630642e-07,1.630670e-07,1.630697e-07,1.630725e-07,1.630753e-07,1.630781e-07,1.630808e-07,1.630836e-07,1.630864e-07,1.630891e-07,1.630919e-07,1.630947e-07,1.630974e-07,1.631002e-07,1.631030e-07,1.631057e-07,1.631085e-07,1.631113e-07,1.631140e-07,1.631168e-07,1.631196e-07,1.631223e-07,1.631251e-07,1.631278e-07,1.631306e-07,1.631334e-07,1.631361e-07,1.631389e-07,1.631416e-07,1.631444e-07,1.631472e-07,1.631499e-07,1.631527e-07,1.631554e-07,1.631582e-07,1.631609e-07,1.631637e-07,1.631664e-07,1.631692e-07,1.631719e-07,1.631747e-07,1.631774e-07,1.631802e-07,1.631829e-07,1.631857e-07,1.631884e-07,1.631912e-07,1.631939e-07,1.631966e-07,1.631994e-07,1.632021e-07,1.632049e-07,1.632076e-07,1.632104e-07,1.632131e-07,1.632158e-07,1.632186e-07,1.632213e-07,1.632240e-07,1.632268e-07,1.632295e-07,1.632323e-07,1.632350e-07,1.632377e-07,1.632405e-07,1.632432e-07,1.632459e-07,1.632487e-07,1.632514e-07,1.632541e-07,1.632568e-07,1.632596e-07,1.632623e-07,1.632650e-07,1.632678e-07,1.632705e-07,1.632732e-07,1.632759e-07,1.632787e-07,1.632814e-07,1.632841e-07,1.632868e-07,1.632896e-07,1.632923e-07,1.632950e-07,1.632977e-07,1.633004e-07,1.633032e-07,1.633059e-07,1.633086e-07,1.633113e-07,1.633140e-07,1.633167e-07,1.633195e-07,1.633222e-07,1.633249e-07,1.633276e-07,1.633303e-07,1.633330e-07,1.633357e-07,1.633384e-07,1.633412e-07,1.633439e-07,1.633466e-07,1.633493e-07,1.633520e-07,1.633547e-07,1.633574e-07,1.633601e-07,1.633628e-07,1.633655e-07,1.633682e-07,1.633709e-07,1.633736e-07,1.633763e-07,1.633790e-07,1.633817e-07,1.633844e-07,1.633871e-07,1.633898e-07,1.633925e-07,1.633952e-07,1.633979e-07,1.634006e-07,1.634033e-07,1.634060e-07,1.634087e-07,1.634114e-07,1.634141e-07,1.634168e-07,1.634195e-07,1.634222e-07,1.634248e-07,1.634275e-07,1.634302e-07,1.634329e-07,1.634356e-07,1.634383e-07,1.634410e-07,1.634437e-07,1.634464e-07,1.634490e-07,1.634517e-07,1.634544e-07,1.634571e-07,1.634598e-07,1.634625e-07,1.634651e-07,1.634678e-07,1.634705e-07,1.634732e-07,1.634759e-07,1.634785e-07,1.634812e-07,1.634839e-07,1.634866e-07,1.634892e-07,1.634919e-07,1.634946e-07,1.634973e-07,1.634999e-07,1.635026e-07,1.635053e-07,1.635079e-07,1.635106e-07,1.635133e-07,1.635160e-07,1.635186e-07,1.635213e-07,1.635240e-07,1.635266e-07,1.635293e-07,1.635320e-07,1.635346e-07,1.635373e-07,1.635400e-07,1.635426e-07,1.635453e-07,1.635479e-07,1.635506e-07,1.635533e-07,1.635559e-07,1.635586e-07,1.635612e-07,1.635639e-07,1.635666e-07,1.635692e-07,1.635719e-07,1.635745e-07,1.635772e-07,1.635798e-07,1.635825e-07,1.635851e-07,1.635878e-07,1.635905e-07,1.635931e-07,1.635958e-07,1.635984e-07,1.636011e-07,1.636037e-07,1.636064e-07,1.636090e-07,1.636116e-07,1.636143e-07,1.636169e-07,1.636196e-07,1.636222e-07,1.636249e-07,1.636275e-07,1.636302e-07,1.636328e-07,1.636354e-07,1.636381e-07,1.636407e-07,1.636434e-07,1.636460e-07,1.636486e-07,1.636513e-07,1.636539e-07,1.636566e-07,1.636592e-07,1.636618e-07,1.636645e-07,1.636671e-07,1.636697e-07,1.636724e-07,1.636750e-07,1.636776e-07,1.636803e-07,1.636829e-07,1.636855e-07,1.636882e-07,1.636908e-07,1.636934e-07,1.636960e-07,1.636987e-07,1.637013e-07,1.637039e-07,1.637066e-07,1.637092e-07,1.637118e-07,1.637144e-07,1.637171e-07,1.637197e-07,1.637223e-07,1.637249e-07,1.637275e-07,1.637302e-07,1.637328e-07,1.637354e-07,1.637380e-07,1.637406e-07,1.637433e-07,1.637459e-07,1.637485e-07,1.637511e-07,1.637537e-07,1.637563e-07,1.637589e-07,1.637616e-07,1.637642e-07,1.637668e-07,1.637694e-07,1.637720e-07,1.637746e-07,1.637772e-07,1.637798e-07,1.637824e-07,1.637851e-07,1.637877e-07,1.637903e-07,1.637929e-07,1.637955e-07,1.637981e-07,1.638007e-07,1.638033e-07,1.638059e-07,1.638085e-07,1.638111e-07,1.638137e-07,1.638163e-07,1.638189e-07,1.638215e-07,1.638241e-07,1.638267e-07,1.638293e-07,1.638319e-07,1.638345e-07,1.638371e-07,1.638397e-07,1.638423e-07,1.638449e-07,1.638475e-07,1.638501e-07,1.638527e-07,1.638553e-07,1.638578e-07,1.638604e-07,1.638630e-07,1.638656e-07,1.638682e-07,1.638708e-07,1.638734e-07,1.638760e-07,1.638786e-07,1.638811e-07,1.638837e-07,1.638863e-07,1.638889e-07,1.638915e-07,1.638941e-07,1.638967e-07,1.638992e-07,1.639018e-07,1.639044e-07,1.639070e-07,1.639096e-07,1.639121e-07,1.639147e-07,1.639173e-07,1.639199e-07,1.639225e-07,1.639250e-07,1.639276e-07,1.639302e-07,1.639328e-07,1.639353e-07,1.639379e-07,1.639405e-07,1.639431e-07,1.639456e-07,1.639482e-07,1.639508e-07,1.639533e-07,1.639559e-07,1.639585e-07,1.639610e-07,1.639636e-07,1.639662e-07,1.639688e-07,1.639713e-07,1.639739e-07,1.639764e-07,1.639790e-07,1.639816e-07,1.639841e-07,1.639867e-07,1.639893e-07,1.639918e-07,1.639944e-07,1.639970e-07,1.639995e-07,1.640021e-07,1.640046e-07,1.640072e-07,1.640097e-07,1.640123e-07,1.640149e-07,1.640174e-07,1.640200e-07,1.640225e-07,1.640251e-07,1.640276e-07,1.640302e-07,1.640327e-07,1.640353e-07,1.640379e-07,1.640404e-07,1.640430e-07,1.640455e-07,1.640481e-07,1.640506e-07,1.640532e-07,1.640557e-07,1.640582e-07,1.640608e-07,1.640633e-07,1.640659e-07,1.640684e-07,1.640710e-07,1.640735e-07,1.640761e-07,1.640786e-07,1.640811e-07,1.640837e-07,1.640862e-07,1.640888e-07,1.640913e-07,1.640939e-07,1.640964e-07,1.640989e-07,1.641015e-07,1.641040e-07,1.641065e-07,1.641091e-07,1.641116e-07,1.641141e-07,1.641167e-07,1.641192e-07,1.641217e-07,1.641243e-07,1.641268e-07,1.641293e-07,1.641319e-07,1.641344e-07,1.641369e-07,1.641395e-07,1.641420e-07,1.641445e-07,1.641471e-07,1.641496e-07,1.641521e-07,1.641546e-07,1.641572e-07,1.641597e-07,1.641622e-07,1.641647e-07,1.641673e-07,1.641698e-07,1.641723e-07,1.641748e-07,1.641773e-07,1.641799e-07,1.641824e-07,1.641849e-07,1.641874e-07,1.641899e-07,1.641925e-07,1.641950e-07,1.641975e-07,1.642000e-07,1.642025e-07,1.642050e-07,1.642076e-07,1.642101e-07,1.642126e-07,1.642151e-07,1.642176e-07,1.642201e-07,1.642226e-07,1.642251e-07,1.642277e-07,1.642302e-07,1.642327e-07,1.642352e-07,1.642377e-07,1.642402e-07,1.642427e-07,1.642452e-07,1.642477e-07,1.642502e-07,1.642527e-07,1.642552e-07,1.642577e-07,1.642602e-07,1.642627e-07,1.642653e-07,1.642678e-07,1.642703e-07,1.642728e-07,1.642753e-07,1.642778e-07,1.642803e-07,1.642828e-07,1.642852e-07,1.642877e-07,1.642902e-07,1.642927e-07,1.642952e-07,1.642977e-07,1.643002e-07,1.643027e-07,1.643052e-07,1.643077e-07,1.643102e-07,1.643127e-07,1.643152e-07,1.643177e-07,1.643202e-07,1.643227e-07,1.643251e-07,1.643276e-07,1.643301e-07,1.643326e-07,1.643351e-07,1.643376e-07,1.643401e-07,1.643426e-07,1.643450e-07,1.643475e-07,1.643500e-07,1.643525e-07,1.643550e-07,1.643575e-07,1.643599e-07,1.643624e-07,1.643649e-07,1.643674e-07,1.643699e-07,1.643723e-07,1.643748e-07,1.643773e-07,1.643798e-07,1.643823e-07,1.643847e-07,1.643872e-07,1.643897e-07,1.643922e-07,1.643946e-07,1.643971e-07,1.643996e-07,1.644021e-07,1.644045e-07,1.644070e-07,1.644095e-07,1.644119e-07,1.644144e-07,1.644169e-07,1.644193e-07,1.644218e-07,1.644243e-07,1.644268e-07,1.644292e-07,1.644317e-07,1.644342e-07,1.644366e-07,1.644391e-07,1.644415e-07,1.644440e-07,1.644465e-07,1.644489e-07,1.644514e-07,1.644539e-07,1.644563e-07,1.644588e-07,1.644612e-07,1.644637e-07,1.644662e-07,1.644686e-07,1.644711e-07,1.644735e-07,1.644760e-07,1.644785e-07,1.644809e-07,1.644834e-07,1.644858e-07,1.644883e-07,1.644907e-07,1.644932e-07,1.644956e-07,1.644981e-07,1.645005e-07,1.645030e-07,1.645054e-07,1.645079e-07,1.645103e-07,1.645128e-07,1.645152e-07,1.645177e-07,1.645201e-07,1.645226e-07,1.645250e-07,1.645275e-07,1.645299e-07,1.645324e-07,1.645348e-07,1.645373e-07,1.645397e-07,1.645421e-07,1.645446e-07,1.645470e-07,1.645495e-07,1.645519e-07,1.645544e-07,1.645568e-07,1.645592e-07,1.645617e-07,1.645641e-07,1.645666e-07,1.645690e-07,1.645714e-07,1.645739e-07,1.645763e-07,1.645787e-07,1.645812e-07,1.645836e-07,1.645860e-07,1.645885e-07,1.645909e-07,1.645933e-07,1.645958e-07,1.645982e-07,1.646006e-07,1.646031e-07,1.646055e-07,1.646079e-07,1.646103e-07,1.646128e-07,1.646152e-07,1.646176e-07,1.646201e-07,1.646225e-07,1.646249e-07,1.646273e-07,1.646298e-07,1.646322e-07,1.646346e-07,1.646370e-07,1.646395e-07,1.646419e-07,1.646443e-07,1.646467e-07,1.646491e-07,1.646516e-07,1.646540e-07,1.646564e-07,1.646588e-07,1.646612e-07,1.646637e-07,1.646661e-07,1.646685e-07,1.646709e-07,1.646733e-07,1.646757e-07,1.646782e-07,1.646806e-07,1.646830e-07,1.646854e-07,1.646878e-07,1.646902e-07,1.646926e-07,1.646950e-07,1.646975e-07,1.646999e-07,1.647023e-07,1.647047e-07,1.647071e-07,1.647095e-07,1.647119e-07,1.647143e-07,1.647167e-07,1.647191e-07,1.647215e-07,1.647239e-07,1.647263e-07,1.647287e-07,1.647312e-07,1.647336e-07,1.647360e-07,1.647384e-07,1.647408e-07,1.647432e-07,1.647456e-07,1.647480e-07,1.647504e-07,1.647528e-07,1.647552e-07,1.647576e-07,1.647600e-07,1.647624e-07,1.647648e-07,1.647671e-07,1.647695e-07,1.647719e-07,1.647743e-07,1.647767e-07,1.647791e-07,1.647815e-07,1.647839e-07,1.647863e-07,1.647887e-07,1.647911e-07,1.647935e-07,1.647959e-07,1.647983e-07,1.648006e-07,1.648030e-07,1.648054e-07,1.648078e-07,1.648102e-07,1.648126e-07,1.648150e-07,1.648174e-07,1.648197e-07,1.648221e-07,1.648245e-07,1.648269e-07,1.648293e-07,1.648317e-07,1.648340e-07,1.648364e-07,1.648388e-07,1.648412e-07,1.648436e-07,1.648459e-07,1.648483e-07,1.648507e-07,1.648531e-07,1.648555e-07,1.648578e-07,1.648602e-07,1.648626e-07,1.648650e-07,1.648673e-07,1.648697e-07,1.648721e-07,1.648745e-07,1.648768e-07,1.648792e-07,1.648816e-07,1.648840e-07,1.648863e-07,1.648887e-07,1.648911e-07,1.648934e-07,1.648958e-07,1.648982e-07,1.649006e-07,1.649029e-07,1.649053e-07,1.649077e-07,1.649100e-07,1.649124e-07,1.649148e-07,1.649171e-07,1.649195e-07,1.649219e-07,1.649242e-07,1.649266e-07,1.649289e-07,1.649313e-07,1.649337e-07,1.649360e-07,1.649384e-07,1.649408e-07,1.649431e-07,1.649455e-07,1.649478e-07,1.649502e-07,1.649526e-07,1.649549e-07,1.649573e-07,1.649596e-07,1.649620e-07,1.649643e-07,1.649667e-07,1.649690e-07,1.649714e-07,1.649738e-07,1.649761e-07,1.649785e-07,1.649808e-07,1.649832e-07,1.649855e-07,1.649879e-07,1.649902e-07,1.649926e-07,1.649949e-07,1.649973e-07,1.649996e-07,1.650020e-07,1.650043e-07,1.650067e-07,1.650090e-07,1.650114e-07,1.650137e-07,1.650160e-07,1.650184e-07,1.650207e-07,1.650231e-07,1.650254e-07,1.650278e-07,1.650301e-07,1.650324e-07,1.650348e-07,1.650371e-07,1.650395e-07,1.650418e-07,1.650442e-07,1.650465e-07,1.650488e-07,1.650512e-07,1.650535e-07,1.650558e-07,1.650582e-07,1.650605e-07,1.650629e-07,1.650652e-07,1.650675e-07,1.650699e-07,1.650722e-07,1.650745e-07,1.650769e-07,1.650792e-07,1.650815e-07,1.650839e-07,1.650862e-07,1.650885e-07,1.650908e-07,1.650932e-07,1.650955e-07,1.650978e-07,1.651002e-07,1.651025e-07,1.651048e-07,1.651071e-07,1.651095e-07,1.651118e-07,1.651141e-07,1.651165e-07,1.651188e-07,1.651211e-07,1.651234e-07,1.651257e-07,1.651281e-07,1.651304e-07,1.651327e-07,1.651350e-07,1.651374e-07,1.651397e-07,1.651420e-07,1.651443e-07,1.651466e-07,1.651490e-07,1.651513e-07,1.651536e-07,1.651559e-07,1.651582e-07,1.651605e-07,1.651629e-07,1.651652e-07,1.651675e-07,1.651698e-07,1.651721e-07,1.651744e-07,1.651767e-07,1.651791e-07,1.651814e-07,1.651837e-07,1.651860e-07,1.651883e-07,1.651906e-07,1.651929e-07,1.651952e-07,1.651975e-07,1.651998e-07,1.652022e-07,1.652045e-07,1.652068e-07,1.652091e-07,1.652114e-07,1.652137e-07,1.652160e-07,1.652183e-07,1.652206e-07,1.652229e-07,1.652252e-07,1.652275e-07,1.652298e-07,1.652321e-07,1.652344e-07,1.652367e-07,1.652390e-07,1.652413e-07,1.652436e-07,1.652459e-07,1.652482e-07,1.652505e-07,1.652528e-07,1.652551e-07,1.652574e-07,1.652597e-07,1.652620e-07,1.652643e-07,1.652666e-07,1.652689e-07,1.652712e-07,1.652735e-07,1.652758e-07,1.652781e-07,1.652804e-07,1.652827e-07,1.652849e-07,1.652872e-07,1.652895e-07,1.652918e-07,1.652941e-07,1.652964e-07,1.652987e-07,1.653010e-07,1.653033e-07,1.653055e-07,1.653078e-07,1.653101e-07,1.653124e-07,1.653147e-07,1.653170e-07,1.653193e-07,1.653215e-07,1.653238e-07,1.653261e-07,1.653284e-07,1.653307e-07,1.653330e-07,1.653352e-07,1.653375e-07,1.653398e-07,1.653421e-07,1.653444e-07,1.653466e-07,1.653489e-07,1.653512e-07,1.653535e-07,1.653558e-07,1.653580e-07,1.653603e-07,1.653626e-07,1.653649e-07,1.653671e-07,1.653694e-07,1.653717e-07,1.653740e-07,1.653762e-07,1.653785e-07,1.653808e-07,1.653831e-07,1.653853e-07,1.653876e-07,1.653899e-07,1.653921e-07,1.653944e-07,1.653967e-07,1.653990e-07,1.654012e-07,1.654035e-07,1.654058e-07,1.654080e-07,1.654103e-07,1.654126e-07,1.654148e-07,1.654171e-07,1.654194e-07,1.654216e-07,1.654239e-07,1.654261e-07,1.654284e-07,1.654307e-07,1.654329e-07,1.654352e-07,1.654375e-07,1.654397e-07,1.654420e-07,1.654442e-07,1.654465e-07,1.654488e-07,1.654510e-07,1.654533e-07,1.654555e-07,1.654578e-07,1.654601e-07,1.654623e-07,1.654646e-07,1.654668e-07,1.654691e-07,1.654713e-07,1.654736e-07,1.654758e-07,1.654781e-07,1.654804e-07,1.654826e-07,1.654849e-07,1.654871e-07,1.654894e-07,1.654916e-07,1.654939e-07,1.654961e-07,1.654984e-07,1.655006e-07,1.655029e-07,1.655051e-07,1.655074e-07,1.655096e-07,1.655119e-07,1.655141e-07,1.655163e-07,1.655186e-07,1.655208e-07,1.655231e-07,1.655253e-07,1.655276e-07,1.655298e-07,1.655321e-07,1.655343e-07,1.655365e-07,1.655388e-07,1.655410e-07,1.655433e-07,1.655455e-07,1.655477e-07,1.655500e-07,1.655522e-07,1.655545e-07,1.655567e-07,1.655589e-07,1.655612e-07,1.655634e-07,1.655657e-07,1.655679e-07,1.655701e-07,1.655724e-07,1.655746e-07,1.655768e-07,1.655791e-07,1.655813e-07,1.655835e-07,1.655858e-07,1.655880e-07,1.655902e-07,1.655925e-07,1.655947e-07,1.655969e-07,1.655992e-07,1.656014e-07,1.656036e-07,1.656058e-07,1.656081e-07,1.656103e-07,1.656125e-07,1.656148e-07,1.656170e-07,1.656192e-07,1.656214e-07,1.656237e-07,1.656259e-07,1.656281e-07,1.656303e-07,1.656326e-07,1.656348e-07,1.656370e-07,1.656392e-07,1.656415e-07,1.656437e-07,1.656459e-07,1.656481e-07,1.656503e-07,1.656526e-07,1.656548e-07,1.656570e-07,1.656592e-07,1.656614e-07,1.656637e-07,1.656659e-07,1.656681e-07,1.656703e-07,1.656725e-07,1.656747e-07,1.656770e-07,1.656792e-07,1.656814e-07,1.656836e-07,1.656858e-07,1.656880e-07,1.656902e-07,1.656924e-07,1.656947e-07,1.656969e-07,1.656991e-07,1.657013e-07,1.657035e-07,1.657057e-07,1.657079e-07,1.657101e-07,1.657123e-07,1.657146e-07,1.657168e-07,1.657190e-07,1.657212e-07,1.657234e-07,1.657256e-07,1.657278e-07,1.657300e-07,1.657322e-07,1.657344e-07,1.657366e-07,1.657388e-07,1.657410e-07,1.657432e-07,1.657454e-07,1.657476e-07,1.657498e-07,1.657520e-07,1.657542e-07,1.657564e-07,1.657586e-07,1.657608e-07,1.657630e-07,1.657652e-07,1.657674e-07,1.657696e-07,1.657718e-07,1.657740e-07,1.657762e-07,1.657784e-07,1.657806e-07,1.657828e-07,1.657850e-07,1.657872e-07,1.657894e-07,1.657916e-07,1.657938e-07,1.657960e-07,1.657982e-07,1.658003e-07,1.658025e-07,1.658047e-07,1.658069e-07,1.658091e-07,1.658113e-07,1.658135e-07,1.658157e-07,1.658179e-07,1.658201e-07,1.658222e-07,1.658244e-07,1.658266e-07,1.658288e-07,1.658310e-07,1.658332e-07,1.658354e-07,1.658376e-07,1.658397e-07,1.658419e-07,1.658441e-07,1.658463e-07,1.658485e-07,1.658507e-07,1.658528e-07,1.658550e-07,1.658572e-07,1.658594e-07,1.658616e-07,1.658637e-07,1.658659e-07,1.658681e-07,1.658703e-07,1.658725e-07,1.658746e-07,1.658768e-07,1.658790e-07,1.658812e-07,1.658833e-07,1.658855e-07,1.658877e-07,1.658899e-07,1.658920e-07,1.658942e-07,1.658964e-07,1.658986e-07,1.659007e-07,1.659029e-07,1.659051e-07,1.659073e-07,1.659094e-07,1.659116e-07,1.659138e-07,1.659159e-07,1.659181e-07,1.659203e-07,1.659224e-07,1.659246e-07,1.659268e-07,1.659290e-07,1.659311e-07,1.659333e-07,1.659355e-07,1.659376e-07,1.659398e-07,1.659420e-07,1.659441e-07,1.659463e-07,1.659484e-07,1.659506e-07,1.659528e-07,1.659549e-07,1.659571e-07,1.659593e-07,1.659614e-07,1.659636e-07,1.659657e-07,1.659679e-07,1.659701e-07,1.659722e-07,1.659744e-07,1.659765e-07,1.659787e-07,1.659809e-07,1.659830e-07,1.659852e-07,1.659873e-07,1.659895e-07,1.659916e-07,1.659938e-07,1.659960e-07,1.659981e-07,1.660003e-07,1.660024e-07,1.660046e-07,1.660067e-07,1.660089e-07,1.660110e-07,1.660132e-07,1.660153e-07,1.660175e-07,1.660196e-07,1.660218e-07,1.660239e-07,1.660261e-07,1.660282e-07,1.660304e-07,1.660325e-07,1.660347e-07,1.660368e-07,1.660390e-07,1.660411e-07,1.660433e-07,1.660454e-07,1.660476e-07,1.660497e-07,1.660519e-07,1.660540e-07,1.660561e-07,1.660583e-07,1.660604e-07,1.660626e-07,1.660647e-07,1.660669e-07,1.660690e-07,1.660711e-07,1.660733e-07,1.660754e-07,1.660776e-07,1.660797e-07,1.660818e-07,1.660840e-07,1.660861e-07,1.660883e-07,1.660904e-07,1.660925e-07,1.660947e-07,1.660968e-07,1.660989e-07,1.661011e-07,1.661032e-07,1.661054e-07,1.661075e-07,1.661096e-07,1.661118e-07,1.661139e-07,1.661160e-07,1.661182e-07,1.661203e-07,1.661224e-07,1.661246e-07,1.661267e-07,1.661288e-07,1.661309e-07,1.661331e-07,1.661352e-07,1.661373e-07,1.661395e-07,1.661416e-07,1.661437e-07,1.661458e-07,1.661480e-07,1.661501e-07,1.661522e-07,1.661544e-07,1.661565e-07,1.661586e-07,1.661607e-07,1.661629e-07,1.661650e-07,1.661671e-07,1.661692e-07,1.661713e-07,1.661735e-07,1.661756e-07,1.661777e-07,1.661798e-07,1.661820e-07,1.661841e-07,1.661862e-07,1.661883e-07,1.661904e-07,1.661926e-07,1.661947e-07,1.661968e-07,1.661989e-07,1.662010e-07,1.662031e-07,1.662053e-07,1.662074e-07,1.662095e-07,1.662116e-07,1.662137e-07,1.662158e-07,1.662180e-07,1.662201e-07,1.662222e-07,1.662243e-07,1.662264e-07,1.662285e-07,1.662306e-07,1.662328e-07,1.662349e-07,1.662370e-07,1.662391e-07,1.662412e-07,1.662433e-07,1.662454e-07,1.662475e-07,1.662496e-07,1.662517e-07,1.662538e-07,1.662560e-07,1.662581e-07,1.662602e-07,1.662623e-07,1.662644e-07,1.662665e-07,1.662686e-07,1.662707e-07,1.662728e-07,1.662749e-07,1.662770e-07,1.662791e-07,1.662812e-07,1.662833e-07,1.662854e-07,1.662875e-07,1.662896e-07,1.662917e-07,1.662938e-07,1.662959e-07,1.662980e-07,1.663001e-07,1.663022e-07,1.663043e-07,1.663064e-07,1.663085e-07,1.663106e-07,1.663127e-07,1.663148e-07,1.663169e-07,1.663190e-07,1.663211e-07,1.663232e-07,1.663253e-07,1.663274e-07,1.663295e-07,1.663316e-07,1.663337e-07,1.663358e-07,1.663379e-07,1.663399e-07,1.663420e-07,1.663441e-07,1.663462e-07,1.663483e-07,1.663504e-07,1.663525e-07,1.663546e-07,1.663567e-07,1.663588e-07,1.663609e-07,1.663629e-07,1.663650e-07,1.663671e-07,1.663692e-07,1.663713e-07,1.663734e-07,1.663755e-07,1.663775e-07,1.663796e-07,1.663817e-07,1.663838e-07,1.663859e-07,1.663880e-07,1.663901e-07,1.663921e-07,1.663942e-07,1.663963e-07,1.663984e-07,1.664005e-07,1.664025e-07,1.664046e-07,1.664067e-07,1.664088e-07,1.664109e-07,1.664129e-07,1.664150e-07,1.664171e-07,1.664192e-07,1.664213e-07,1.664233e-07,1.664254e-07,1.664275e-07,1.664296e-07,1.664316e-07,1.664337e-07,1.664358e-07,1.664379e-07,1.664399e-07,1.664420e-07,1.664441e-07,1.664462e-07,1.664482e-07,1.664503e-07,1.664524e-07,1.664545e-07,1.664565e-07,1.664586e-07,1.664607e-07,1.664627e-07,1.664648e-07,1.664669e-07,1.664689e-07,1.664710e-07,1.664731e-07,1.664752e-07,1.664772e-07,1.664793e-07,1.664814e-07,1.664834e-07,1.664855e-07,1.664876e-07,1.664896e-07,1.664917e-07,1.664937e-07,1.664958e-07,1.664979e-07,1.664999e-07,1.665020e-07,1.665041e-07,1.665061e-07,1.665082e-07,1.665103e-07,1.665123e-07,1.665144e-07,1.665164e-07,1.665185e-07,1.665206e-07,1.665226e-07,1.665247e-07,1.665267e-07,1.665288e-07,1.665309e-07,1.665329e-07,1.665350e-07,1.665370e-07,1.665391e-07,1.665411e-07,1.665432e-07,1.665453e-07,1.665473e-07,1.665494e-07,1.665514e-07,1.665535e-07,1.665555e-07,1.665576e-07,1.665596e-07,1.665617e-07,1.665637e-07,1.665658e-07,1.665678e-07,1.665699e-07,1.665719e-07,1.665740e-07,1.665760e-07,1.665781e-07,1.665801e-07,1.665822e-07,1.665842e-07,1.665863e-07,1.665883e-07,1.665904e-07,1.665924e-07,1.665945e-07,1.665965e-07,1.665986e-07,1.666006e-07,1.666027e-07,1.666047e-07,1.666068e-07,1.666088e-07,1.666108e-07,1.666129e-07,1.666149e-07,1.666170e-07,1.666190e-07,1.666211e-07,1.666231e-07,1.666251e-07,1.666272e-07,1.666292e-07,1.666313e-07,1.666333e-07,1.666353e-07,1.666374e-07,1.666394e-07,1.666415e-07,1.666435e-07,1.666455e-07,1.666476e-07,1.666496e-07,1.666517e-07,1.666537e-07,1.666557e-07,1.666578e-07,1.666598e-07,1.666618e-07,1.666639e-07,1.666659e-07,1.666679e-07,1.666700e-07,1.666720e-07,1.666740e-07,1.666761e-07,1.666781e-07,1.666801e-07,1.666822e-07,1.666842e-07,1.666862e-07,1.666883e-07,1.666903e-07,1.666923e-07,1.666943e-07,1.666964e-07,1.666984e-07,1.667004e-07,1.667025e-07,1.667045e-07,1.667065e-07,1.667085e-07,1.667106e-07,1.667126e-07,1.667146e-07,1.667166e-07,1.667187e-07,1.667207e-07,1.667227e-07,1.667247e-07,1.667268e-07,1.667288e-07,1.667308e-07,1.667328e-07,1.667349e-07,1.667369e-07,1.667389e-07,1.667409e-07,1.667429e-07,1.667450e-07,1.667470e-07,1.667490e-07,1.667510e-07,1.667530e-07,1.667551e-07,1.667571e-07,1.667591e-07,1.667611e-07,1.667631e-07,1.667652e-07,1.667672e-07,1.667692e-07,1.667712e-07,1.667732e-07,1.667752e-07,1.667772e-07,1.667793e-07,1.667813e-07,1.667833e-07,1.667853e-07,1.667873e-07,1.667893e-07,1.667913e-07,1.667934e-07,1.667954e-07,1.667974e-07,1.667994e-07,1.668014e-07,1.668034e-07,1.668054e-07,1.668074e-07,1.668094e-07,1.668115e-07,1.668135e-07,1.668155e-07,1.668175e-07,1.668195e-07,1.668215e-07,1.668235e-07,1.668255e-07,1.668275e-07,1.668295e-07,1.668315e-07,1.668335e-07,1.668355e-07,1.668375e-07,1.668395e-07,1.668415e-07,1.668435e-07,1.668456e-07,1.668476e-07,1.668496e-07,1.668516e-07,1.668536e-07,1.668556e-07,1.668576e-07,1.668596e-07,1.668616e-07,1.668636e-07,1.668656e-07,1.668676e-07,1.668696e-07,1.668716e-07,1.668736e-07,1.668756e-07,1.668776e-07,1.668796e-07,1.668816e-07,1.668835e-07,1.668855e-07,1.668875e-07,1.668895e-07,1.668915e-07,1.668935e-07,1.668955e-07,1.668975e-07,1.668995e-07,1.669015e-07,1.669035e-07,1.669055e-07,1.669075e-07,1.669095e-07,1.669115e-07,1.669135e-07,1.669154e-07,1.669174e-07,1.669194e-07,1.669214e-07,1.669234e-07,1.669254e-07,1.669274e-07,1.669294e-07,1.669314e-07,1.669334e-07,1.669353e-07,1.669373e-07,1.669393e-07,1.669413e-07,1.669433e-07,1.669453e-07,1.669473e-07,1.669492e-07,1.669512e-07,1.669532e-07,1.669552e-07,1.669572e-07,1.669592e-07,1.669612e-07,1.669631e-07,1.669651e-07,1.669671e-07,1.669691e-07,1.669711e-07,1.669730e-07,1.669750e-07,1.669770e-07,1.669790e-07,1.669810e-07,1.669829e-07,1.669849e-07,1.669869e-07,1.669889e-07,1.669909e-07,1.669928e-07,1.669948e-07,1.669968e-07,1.669988e-07,1.670007e-07,1.670027e-07,1.670047e-07,1.670067e-07,1.670086e-07,1.670106e-07,1.670126e-07,1.670146e-07,1.670165e-07,1.670185e-07,1.670205e-07,1.670225e-07,1.670244e-07,1.670264e-07,1.670284e-07,1.670304e-07,1.670323e-07,1.670343e-07,1.670363e-07,1.670382e-07,1.670402e-07,1.670422e-07,1.670441e-07,1.670461e-07,1.670481e-07,1.670501e-07,1.670520e-07,1.670540e-07,1.670560e-07,1.670579e-07,1.670599e-07,1.670619e-07,1.670638e-07,1.670658e-07,1.670678e-07,1.670697e-07,1.670717e-07,1.670736e-07,1.670756e-07,1.670776e-07,1.670795e-07,1.670815e-07,1.670835e-07,1.670854e-07,1.670874e-07,1.670893e-07,1.670913e-07,1.670933e-07,1.670952e-07,1.670972e-07,1.670991e-07,1.671011e-07,1.671031e-07,1.671050e-07,1.671070e-07,1.671089e-07,1.671109e-07,1.671129e-07,1.671148e-07,1.671168e-07,1.671187e-07,1.671207e-07,1.671226e-07,1.671246e-07,1.671266e-07,1.671285e-07,1.671305e-07,1.671324e-07,1.671344e-07,1.671363e-07,1.671383e-07,1.671402e-07,1.671422e-07,1.671441e-07,1.671461e-07,1.671480e-07,1.671500e-07,1.671519e-07,1.671539e-07,1.671558e-07,1.671578e-07,1.671597e-07,1.671617e-07,1.671636e-07,1.671656e-07,1.671675e-07,1.671695e-07,1.671714e-07,1.671734e-07,1.671753e-07,1.671773e-07,1.671792e-07,1.671812e-07,1.671831e-07,1.671851e-07,1.671870e-07,1.671889e-07,1.671909e-07,1.671928e-07,1.671948e-07,1.671967e-07,1.671987e-07,1.672006e-07,1.672026e-07,1.672045e-07,1.672064e-07,1.672084e-07,1.672103e-07,1.672123e-07,1.672142e-07,1.672161e-07,1.672181e-07,1.672200e-07,1.672220e-07,1.672239e-07,1.672258e-07,1.672278e-07,1.672297e-07,1.672317e-07,1.672336e-07,1.672355e-07,1.672375e-07,1.672394e-07,1.672413e-07,1.672433e-07,1.672452e-07,1.672471e-07,1.672491e-07,1.672510e-07,1.672529e-07,1.672549e-07,1.672568e-07,1.672587e-07,1.672607e-07,1.672626e-07,1.672645e-07,1.672665e-07,1.672684e-07,1.672703e-07,1.672723e-07,1.672742e-07,1.672761e-07,1.672781e-07,1.672800e-07,1.672819e-07,1.672838e-07,1.672858e-07,1.672877e-07,1.672896e-07,1.672916e-07,1.672935e-07,1.672954e-07,1.672973e-07,1.672993e-07,1.673012e-07,1.673031e-07,1.673050e-07,1.673070e-07,1.673089e-07,1.673108e-07,1.673127e-07,1.673147e-07,1.673166e-07,1.673185e-07,1.673204e-07,1.673224e-07,1.673243e-07,1.673262e-07,1.673281e-07,1.673300e-07,1.673320e-07,1.673339e-07,1.673358e-07,1.673377e-07,1.673396e-07,1.673416e-07,1.673435e-07,1.673454e-07,1.673473e-07,1.673492e-07,1.673512e-07,1.673531e-07,1.673550e-07,1.673569e-07,1.673588e-07,1.673607e-07,1.673627e-07,1.673646e-07,1.673665e-07,1.673684e-07,1.673703e-07,1.673722e-07,1.673741e-07,1.673761e-07,1.673780e-07,1.673799e-07,1.673818e-07,1.673837e-07,1.673856e-07,1.673875e-07,1.673894e-07,1.673914e-07,1.673933e-07,1.673952e-07,1.673971e-07,1.673990e-07,1.674009e-07,1.674028e-07,1.674047e-07,1.674066e-07,1.674085e-07,1.674105e-07,1.674124e-07,1.674143e-07,1.674162e-07,1.674181e-07,1.674200e-07,1.674219e-07,1.674238e-07,1.674257e-07,1.674276e-07,1.674295e-07,1.674314e-07,1.674333e-07,1.674352e-07,1.674371e-07,1.674390e-07,1.674409e-07,1.674428e-07,1.674447e-07,1.674466e-07,1.674485e-07,1.674505e-07,1.674524e-07,1.674543e-07,1.674562e-07,1.674581e-07,1.674600e-07,1.674619e-07,1.674638e-07,1.674657e-07,1.674676e-07,1.674694e-07,1.674713e-07,1.674732e-07,1.674751e-07,1.674770e-07,1.674789e-07,1.674808e-07,1.674827e-07,1.674846e-07,1.674865e-07,1.674884e-07,1.674903e-07,1.674922e-07,1.674941e-07,1.674960e-07,1.674979e-07,1.674998e-07,1.675017e-07,1.675036e-07,1.675055e-07,1.675074e-07,1.675092e-07,1.675111e-07,1.675130e-07,1.675149e-07,1.675168e-07,1.675187e-07,1.675206e-07,1.675225e-07,1.675244e-07,1.675263e-07,1.675281e-07,1.675300e-07,1.675319e-07,1.675338e-07,1.675357e-07,1.675376e-07,1.675395e-07,1.675414e-07,1.675432e-07,1.675451e-07,1.675470e-07,1.675489e-07,1.675508e-07,1.675527e-07,1.675546e-07,1.675564e-07,1.675583e-07,1.675602e-07,1.675621e-07,1.675640e-07,1.675659e-07,1.675677e-07,1.675696e-07,1.675715e-07,1.675734e-07,1.675753e-07,1.675771e-07,1.675790e-07,1.675809e-07,1.675828e-07,1.675847e-07,1.675865e-07,1.675884e-07,1.675903e-07,1.675922e-07,1.675941e-07,1.675959e-07,1.675978e-07,1.675997e-07,1.676016e-07,1.676034e-07,1.676053e-07,1.676072e-07,1.676091e-07,1.676109e-07,1.676128e-07,1.676147e-07,1.676166e-07,1.676184e-07,1.676203e-07,1.676222e-07,1.676241e-07,1.676259e-07,1.676278e-07,1.676297e-07,1.676316e-07,1.676334e-07,1.676353e-07,1.676372e-07,1.676390e-07,1.676409e-07,1.676428e-07,1.676447e-07,1.676465e-07,1.676484e-07,1.676503e-07,1.676521e-07,1.676540e-07,1.676559e-07,1.676577e-07,1.676596e-07,1.676615e-07,1.676633e-07,1.676652e-07,1.676671e-07,1.676689e-07,1.676708e-07,1.676727e-07,1.676745e-07,1.676764e-07,1.676783e-07,1.676801e-07,1.676820e-07,1.676839e-07,1.676857e-07,1.676876e-07,1.676894e-07,1.676913e-07,1.676932e-07,1.676950e-07,1.676969e-07,1.676987e-07,1.677006e-07,1.677025e-07,1.677043e-07,1.677062e-07,1.677081e-07,1.677099e-07,1.677118e-07,1.677136e-07,1.677155e-07,1.677173e-07,1.677192e-07,1.677211e-07,1.677229e-07,1.677248e-07,1.677266e-07,1.677285e-07,1.677303e-07,1.677322e-07,1.677341e-07,1.677359e-07,1.677378e-07,1.677396e-07,1.677415e-07,1.677433e-07,1.677452e-07,1.677470e-07,1.677489e-07,1.677507e-07,1.677526e-07,1.677544e-07,1.677563e-07,1.677582e-07,1.677600e-07,1.677619e-07,1.677637e-07,1.677656e-07,1.677674e-07,1.677693e-07,1.677711e-07,1.677730e-07,1.677748e-07,1.677767e-07,1.677785e-07,1.677803e-07,1.677822e-07,1.677840e-07,1.677859e-07,1.677877e-07,1.677896e-07,1.677914e-07,1.677933e-07,1.677951e-07,1.677970e-07,1.677988e-07,1.678007e-07,1.678025e-07,1.678043e-07,1.678062e-07,1.678080e-07,1.678099e-07,1.678117e-07,1.678136e-07,1.678154e-07,1.678173e-07,1.678191e-07,1.678209e-07,1.678228e-07,1.678246e-07,1.678265e-07,1.678283e-07,1.678301e-07,1.678320e-07,1.678338e-07,1.678357e-07,1.678375e-07,1.678393e-07,1.678412e-07,1.678430e-07,1.678449e-07,1.678467e-07,1.678485e-07,1.678504e-07,1.678522e-07,1.678540e-07,1.678559e-07,1.678577e-07,1.678595e-07,1.678614e-07,1.678632e-07,1.678650e-07,1.678669e-07,1.678687e-07,1.678706e-07,1.678724e-07,1.678742e-07,1.678761e-07,1.678779e-07,1.678797e-07,1.678815e-07,1.678834e-07,1.678852e-07,1.678870e-07,1.678889e-07,1.678907e-07,1.678925e-07,1.678944e-07,1.678962e-07,1.678980e-07,1.678999e-07,1.679017e-07,1.679035e-07,1.679053e-07,1.679072e-07,1.679090e-07,1.679108e-07,1.679127e-07,1.679145e-07,1.679163e-07,1.679181e-07,1.679200e-07,1.679218e-07,1.679236e-07,1.679254e-07,1.679273e-07,1.679291e-07,1.679309e-07,1.679327e-07,1.679346e-07,1.679364e-07,1.679382e-07,1.679400e-07,1.679418e-07,1.679437e-07,1.679455e-07,1.679473e-07,1.679491e-07,1.679510e-07,1.679528e-07,1.679546e-07,1.679564e-07,1.679582e-07,1.679601e-07,1.679619e-07,1.679637e-07,1.679655e-07,1.679673e-07,1.679692e-07,1.679710e-07,1.679728e-07,1.679746e-07,1.679764e-07,1.679782e-07,1.679801e-07,1.679819e-07,1.679837e-07,1.679855e-07,1.679873e-07,1.679891e-07,1.679910e-07,1.679928e-07,1.679946e-07,1.679964e-07,1.679982e-07,1.680000e-07,1.680018e-07,1.680036e-07,1.680055e-07,1.680073e-07,1.680091e-07,1.680109e-07,1.680127e-07,1.680145e-07,1.680163e-07,1.680181e-07,1.680200e-07,1.680218e-07,1.680236e-07,1.680254e-07,1.680272e-07,1.680290e-07,1.680308e-07,1.680326e-07,1.680344e-07,1.680362e-07,1.680380e-07,1.680398e-07,1.680417e-07,1.680435e-07,1.680453e-07,1.680471e-07,1.680489e-07,1.680507e-07,1.680525e-07,1.680543e-07,1.680561e-07,1.680579e-07,1.680597e-07,1.680615e-07,1.680633e-07,1.680651e-07,1.680669e-07,1.680687e-07,1.680705e-07,1.680723e-07,1.680741e-07,1.680759e-07,1.680777e-07,1.680795e-07,1.680813e-07,1.680831e-07,1.680849e-07,1.680867e-07,1.680885e-07,1.680903e-07,1.680921e-07,1.680939e-07,1.680957e-07,1.680975e-07,1.680993e-07,1.681011e-07,1.681029e-07,1.681047e-07,1.681065e-07,1.681083e-07,1.681101e-07,1.681119e-07,1.681137e-07,1.681155e-07,1.681173e-07,1.681191e-07,1.681209e-07,1.681227e-07,1.681245e-07,1.681263e-07,1.681281e-07,1.681299e-07,1.681317e-07,1.681334e-07,1.681352e-07,1.681370e-07,1.681388e-07,1.681406e-07,1.681424e-07,1.681442e-07,1.681460e-07,1.681478e-07,1.681496e-07,1.681514e-07,1.681531e-07,1.681549e-07,1.681567e-07,1.681585e-07,1.681603e-07,1.681621e-07,1.681639e-07,1.681657e-07,1.681675e-07,1.681692e-07,1.681710e-07,1.681728e-07,1.681746e-07,1.681764e-07,1.681782e-07,1.681800e-07,1.681817e-07,1.681835e-07,1.681853e-07,1.681871e-07,1.681889e-07,1.681907e-07,1.681925e-07,1.681942e-07,1.681960e-07,1.681978e-07,1.681996e-07,1.682014e-07,1.682031e-07,1.682049e-07,1.682067e-07,1.682085e-07,1.682103e-07,1.682121e-07,1.682138e-07,1.682156e-07,1.682174e-07,1.682192e-07,1.682210e-07,1.682227e-07,1.682245e-07,1.682263e-07,1.682281e-07,1.682298e-07,1.682316e-07,1.682334e-07,1.682352e-07,1.682370e-07,1.682387e-07,1.682405e-07,1.682423e-07,1.682441e-07,1.682458e-07,1.682476e-07,1.682494e-07,1.682512e-07,1.682529e-07,1.682547e-07,1.682565e-07,1.682583e-07,1.682600e-07,1.682618e-07,1.682636e-07,1.682653e-07,1.682671e-07,1.682689e-07,1.682707e-07,1.682724e-07,1.682742e-07,1.682760e-07,1.682778e-07,1.682795e-07,1.682813e-07,1.682831e-07,1.682848e-07,1.682866e-07,1.682884e-07,1.682901e-07,1.682919e-07,1.682937e-07,1.682954e-07,1.682972e-07,1.682990e-07,1.683007e-07,1.683025e-07,1.683043e-07,1.683060e-07,1.683078e-07,1.683096e-07,1.683113e-07,1.683131e-07,1.683149e-07,1.683166e-07,1.683184e-07,1.683202e-07,1.683219e-07,1.683237e-07,1.683255e-07,1.683272e-07,1.683290e-07,1.683307e-07,1.683325e-07,1.683343e-07,1.683360e-07,1.683378e-07,1.683396e-07,1.683413e-07,1.683431e-07,1.683448e-07,1.683466e-07,1.683484e-07,1.683501e-07,1.683519e-07,1.683536e-07,1.683554e-07,1.683572e-07,1.683589e-07,1.683607e-07,1.683624e-07,1.683642e-07,1.683659e-07,1.683677e-07,1.683695e-07,1.683712e-07,1.683730e-07,1.683747e-07,1.683765e-07,1.683782e-07,1.683800e-07,1.683817e-07,1.683835e-07,1.683853e-07,1.683870e-07,1.683888e-07,1.683905e-07,1.683923e-07,1.683940e-07,1.683958e-07,1.683975e-07,1.683993e-07,1.684010e-07,1.684028e-07,1.684045e-07,1.684063e-07,1.684080e-07,1.684098e-07,1.684115e-07,1.684133e-07,1.684150e-07,1.684168e-07,1.684185e-07,1.684203e-07,1.684220e-07,1.684238e-07,1.684255e-07,1.684273e-07,1.684290e-07,1.684308e-07,1.684325e-07,1.684343e-07,1.684360e-07,1.684378e-07,1.684395e-07,1.684413e-07,1.684430e-07,1.684447e-07,1.684465e-07,1.684482e-07,1.684500e-07,1.684517e-07,1.684535e-07,1.684552e-07,1.684570e-07,1.684587e-07,1.684604e-07,1.684622e-07,1.684639e-07,1.684657e-07,1.684674e-07,1.684692e-07,1.684709e-07,1.684726e-07,1.684744e-07,1.684761e-07,1.684779e-07,1.684796e-07,1.684813e-07,1.684831e-07,1.684848e-07,1.684866e-07,1.684883e-07,1.684900e-07,1.684918e-07,1.684935e-07,1.684952e-07,1.684970e-07,1.684987e-07,1.685005e-07,1.685022e-07,1.685039e-07,1.685057e-07,1.685074e-07,1.685091e-07,1.685109e-07,1.685126e-07,1.685143e-07,1.685161e-07,1.685178e-07,1.685195e-07,1.685213e-07,1.685230e-07,1.685247e-07,1.685265e-07,1.685282e-07,1.685299e-07,1.685317e-07,1.685334e-07,1.685351e-07,1.685369e-07,1.685386e-07,1.685403e-07,1.685421e-07,1.685438e-07,1.685455e-07,1.685473e-07,1.685490e-07,1.685507e-07,1.685524e-07,1.685542e-07,1.685559e-07,1.685576e-07,1.685594e-07,1.685611e-07,1.685628e-07,1.685645e-07,1.685663e-07,1.685680e-07,1.685697e-07,1.685715e-07,1.685732e-07,1.685749e-07,1.685766e-07,1.685784e-07,1.685801e-07,1.685818e-07,1.685835e-07,1.685853e-07,1.685870e-07,1.685887e-07,1.685904e-07,1.685922e-07,1.685939e-07,1.685956e-07,1.685973e-07,1.685990e-07,1.686008e-07,1.686025e-07,1.686042e-07,1.686059e-07,1.686077e-07,1.686094e-07,1.686111e-07,1.686128e-07,1.686145e-07,1.686163e-07,1.686180e-07,1.686197e-07,1.686214e-07,1.686231e-07,1.686248e-07,1.686266e-07,1.686283e-07,1.686300e-07,1.686317e-07,1.686334e-07,1.686352e-07,1.686369e-07,1.686386e-07,1.686403e-07,1.686420e-07,1.686437e-07,1.686454e-07,1.686472e-07,1.686489e-07,1.686506e-07,1.686523e-07,1.686540e-07,1.686557e-07,1.686575e-07,1.686592e-07,1.686609e-07,1.686626e-07,1.686643e-07,1.686660e-07,1.686677e-07,1.686694e-07,1.686712e-07,1.686729e-07,1.686746e-07,1.686763e-07,1.686780e-07,1.686797e-07,1.686814e-07,1.686831e-07,1.686848e-07,1.686865e-07,1.686883e-07,1.686900e-07,1.686917e-07,1.686934e-07,1.686951e-07,1.686968e-07,1.686985e-07,1.687002e-07,1.687019e-07,1.687036e-07,1.687053e-07,1.687070e-07,1.687087e-07,1.687105e-07,1.687122e-07,1.687139e-07,1.687156e-07,1.687173e-07,1.687190e-07,1.687207e-07,1.687224e-07,1.687241e-07,1.687258e-07,1.687275e-07,1.687292e-07,1.687309e-07,1.687326e-07,1.687343e-07,1.687360e-07,1.687377e-07,1.687394e-07,1.687411e-07,1.687428e-07,1.687445e-07,1.687462e-07,1.687479e-07,1.687496e-07,1.687513e-07,1.687530e-07,1.687547e-07,1.687564e-07,1.687581e-07,1.687598e-07,1.687615e-07,1.687632e-07,1.687649e-07,1.687666e-07,1.687683e-07,1.687700e-07,1.687717e-07,1.687734e-07,1.687751e-07,1.687768e-07,1.687785e-07,1.687802e-07,1.687819e-07,1.687836e-07,1.687853e-07,1.687870e-07,1.687887e-07,1.687903e-07,1.687920e-07,1.687937e-07,1.687954e-07,1.687971e-07,1.687988e-07,1.688005e-07,1.688022e-07,1.688039e-07,1.688056e-07,1.688073e-07,1.688090e-07,1.688107e-07,1.688123e-07,1.688140e-07,1.688157e-07,1.688174e-07,1.688191e-07,1.688208e-07,1.688225e-07,1.688242e-07,1.688259e-07,1.688276e-07,1.688292e-07,1.688309e-07,1.688326e-07,1.688343e-07,1.688360e-07,1.688377e-07,1.688394e-07,1.688411e-07,1.688427e-07,1.688444e-07,1.688461e-07,1.688478e-07,1.688495e-07,1.688512e-07,1.688529e-07,1.688545e-07,1.688562e-07,1.688579e-07,1.688596e-07,1.688613e-07,1.688630e-07,1.688646e-07,1.688663e-07,1.688680e-07,1.688697e-07,1.688714e-07,1.688731e-07,1.688747e-07,1.688764e-07,1.688781e-07,1.688798e-07,1.688815e-07,1.688831e-07,1.688848e-07,1.688865e-07,1.688882e-07,1.688899e-07,1.688915e-07,1.688932e-07,1.688949e-07,1.688966e-07,1.688983e-07,1.688999e-07,1.689016e-07,1.689033e-07,1.689050e-07,1.689067e-07,1.689083e-07,1.689100e-07,1.689117e-07,1.689134e-07,1.689150e-07,1.689167e-07,1.689184e-07,1.689201e-07,1.689217e-07,1.689234e-07,1.689251e-07,1.689268e-07,1.689284e-07,1.689301e-07,1.689318e-07,1.689335e-07,1.689351e-07,1.689368e-07,1.689385e-07,1.689401e-07,1.689418e-07,1.689435e-07,1.689452e-07,1.689468e-07,1.689485e-07,1.689502e-07,1.689518e-07,1.689535e-07,1.689552e-07,1.689569e-07,1.689585e-07,1.689602e-07,1.689619e-07,1.689635e-07,1.689652e-07,1.689669e-07,1.689685e-07,1.689702e-07,1.689719e-07,1.689735e-07,1.689752e-07,1.689769e-07,1.689785e-07,1.689802e-07,1.689819e-07,1.689835e-07,1.689852e-07,1.689869e-07,1.689885e-07,1.689902e-07,1.689919e-07,1.689935e-07,1.689952e-07,1.689969e-07,1.689985e-07,1.690002e-07,1.690019e-07,1.690035e-07,1.690052e-07,1.690069e-07,1.690085e-07,1.690102e-07,1.690118e-07,1.690135e-07,1.690152e-07,1.690168e-07,1.690185e-07,1.690201e-07,1.690218e-07,1.690235e-07,1.690251e-07,1.690268e-07,1.690284e-07,1.690301e-07,1.690318e-07,1.690334e-07,1.690351e-07,1.690367e-07,1.690384e-07,1.690401e-07,1.690417e-07,1.690434e-07,1.690450e-07,1.690467e-07,1.690483e-07,1.690500e-07,1.690517e-07,1.690533e-07,1.690550e-07,1.690566e-07,1.690583e-07,1.690599e-07,1.690616e-07,1.690632e-07,1.690649e-07,1.690666e-07,1.690682e-07,1.690699e-07,1.690715e-07,1.690732e-07,1.690748e-07,1.690765e-07,1.690781e-07,1.690798e-07,1.690814e-07,1.690831e-07,1.690847e-07,1.690864e-07,1.690880e-07,1.690897e-07,1.690913e-07,1.690930e-07,1.690946e-07,1.690963e-07,1.690979e-07,1.690996e-07,1.691012e-07,1.691029e-07,1.691045e-07,1.691062e-07,1.691078e-07,1.691095e-07,1.691111e-07,1.691128e-07,1.691144e-07,1.691161e-07,1.691177e-07,1.691194e-07,1.691210e-07,1.691227e-07,1.691243e-07,1.691260e-07,1.691276e-07,1.691293e-07,1.691309e-07,1.691325e-07,1.691342e-07,1.691358e-07,1.691375e-07,1.691391e-07,1.691408e-07,1.691424e-07,1.691440e-07,1.691457e-07,1.691473e-07,1.691490e-07,1.691506e-07,1.691523e-07,1.691539e-07,1.691555e-07,1.691572e-07,1.691588e-07,1.691605e-07,1.691621e-07,1.691638e-07,1.691654e-07,1.691670e-07,1.691687e-07,1.691703e-07,1.691720e-07,1.691736e-07,1.691752e-07,1.691769e-07,1.691785e-07,1.691801e-07,1.691818e-07,1.691834e-07,1.691851e-07,1.691867e-07,1.691883e-07,1.691900e-07,1.691916e-07,1.691932e-07,1.691949e-07,1.691965e-07,1.691982e-07,1.691998e-07,1.692014e-07,1.692031e-07,1.692047e-07,1.692063e-07,1.692080e-07,1.692096e-07,1.692112e-07,1.692129e-07,1.692145e-07,1.692161e-07,1.692178e-07,1.692194e-07,1.692210e-07,1.692227e-07,1.692243e-07,1.692259e-07,1.692276e-07,1.692292e-07,1.692308e-07,1.692324e-07,1.692341e-07,1.692357e-07,1.692373e-07,1.692390e-07,1.692406e-07,1.692422e-07,1.692439e-07,1.692455e-07,1.692471e-07,1.692487e-07,1.692504e-07,1.692520e-07,1.692536e-07,1.692553e-07,1.692569e-07,1.692585e-07,1.692601e-07,1.692618e-07,1.692634e-07,1.692650e-07,1.692666e-07,1.692683e-07,1.692699e-07,1.692715e-07,1.692731e-07,1.692748e-07,1.692764e-07,1.692780e-07,1.692796e-07,1.692813e-07,1.692829e-07,1.692845e-07,1.692861e-07,1.692878e-07,1.692894e-07,1.692910e-07,1.692926e-07,1.692943e-07,1.692959e-07,1.692975e-07,1.692991e-07,1.693007e-07,1.693024e-07,1.693040e-07,1.693056e-07,1.693072e-07,1.693088e-07,1.693105e-07,1.693121e-07,1.693137e-07,1.693153e-07,1.693169e-07,1.693186e-07,1.693202e-07,1.693218e-07,1.693234e-07,1.693250e-07,1.693267e-07,1.693283e-07,1.693299e-07,1.693315e-07,1.693331e-07,1.693347e-07,1.693364e-07,1.693380e-07,1.693396e-07,1.693412e-07,1.693428e-07,1.693444e-07,1.693460e-07,1.693477e-07,1.693493e-07,1.693509e-07,1.693525e-07,1.693541e-07,1.693557e-07,1.693573e-07,1.693590e-07,1.693606e-07,1.693622e-07,1.693638e-07,1.693654e-07,1.693670e-07,1.693686e-07,1.693702e-07,1.693719e-07,1.693735e-07,1.693751e-07,1.693767e-07,1.693783e-07,1.693799e-07,1.693815e-07,1.693831e-07,1.693847e-07,1.693864e-07,1.693880e-07,1.693896e-07,1.693912e-07,1.693928e-07,1.693944e-07,1.693960e-07,1.693976e-07,1.693992e-07,1.694008e-07,1.694024e-07,1.694040e-07,1.694056e-07,1.694073e-07,1.694089e-07,1.694105e-07,1.694121e-07,1.694137e-07,1.694153e-07,1.694169e-07,1.694185e-07,1.694201e-07,1.694217e-07,1.694233e-07,1.694249e-07,1.694265e-07,1.694281e-07,1.694297e-07,1.694313e-07,1.694329e-07,1.694345e-07,1.694361e-07,1.694377e-07,1.694393e-07,1.694409e-07,1.694425e-07,1.694441e-07,1.694457e-07,1.694473e-07,1.694489e-07,1.694505e-07,1.694521e-07,1.694537e-07,1.694553e-07,1.694569e-07,1.694585e-07,1.694601e-07,1.694617e-07,1.694633e-07,1.694649e-07,1.694665e-07,1.694681e-07,1.694697e-07,1.694713e-07,1.694729e-07,1.694745e-07,1.694761e-07,1.694777e-07,1.694793e-07,1.694809e-07,1.694825e-07,1.694841e-07,1.694857e-07,1.694873e-07,1.694889e-07,1.694905e-07,1.694921e-07,1.694937e-07,1.694953e-07,1.694969e-07,1.694985e-07,1.695001e-07,1.695016e-07,1.695032e-07,1.695048e-07,1.695064e-07,1.695080e-07,1.695096e-07,1.695112e-07,1.695128e-07,1.695144e-07,1.695160e-07,1.695176e-07,1.695192e-07,1.695208e-07,1.695223e-07,1.695239e-07,1.695255e-07,1.695271e-07,1.695287e-07,1.695303e-07,1.695319e-07,1.695335e-07,1.695351e-07,1.695367e-07,1.695382e-07,1.695398e-07,1.695414e-07,1.695430e-07,1.695446e-07,1.695462e-07,1.695478e-07,1.695494e-07,1.695509e-07,1.695525e-07,1.695541e-07,1.695557e-07,1.695573e-07,1.695589e-07,1.695605e-07,1.695620e-07,1.695636e-07,1.695652e-07,1.695668e-07,1.695684e-07,1.695700e-07,1.695715e-07,1.695731e-07,1.695747e-07,1.695763e-07,1.695779e-07,1.695795e-07,1.695810e-07,1.695826e-07,1.695842e-07,1.695858e-07,1.695874e-07,1.695890e-07,1.695905e-07,1.695921e-07,1.695937e-07,1.695953e-07,1.695969e-07,1.695984e-07,1.696000e-07,1.696016e-07,1.696032e-07,1.696048e-07,1.696063e-07,1.696079e-07,1.696095e-07,1.696111e-07,1.696127e-07,1.696142e-07,1.696158e-07,1.696174e-07,1.696190e-07,1.696205e-07,1.696221e-07,1.696237e-07,1.696253e-07,1.696269e-07,1.696284e-07,1.696300e-07,1.696316e-07,1.696332e-07,1.696347e-07,1.696363e-07,1.696379e-07,1.696395e-07,1.696410e-07,1.696426e-07,1.696442e-07,1.696458e-07,1.696473e-07,1.696489e-07,1.696505e-07,1.696520e-07,1.696536e-07,1.696552e-07,1.696568e-07,1.696583e-07,1.696599e-07,1.696615e-07,1.696631e-07,1.696646e-07,1.696662e-07,1.696678e-07,1.696693e-07,1.696709e-07,1.696725e-07,1.696740e-07,1.696756e-07,1.696772e-07,1.696788e-07,1.696803e-07,1.696819e-07,1.696835e-07,1.696850e-07,1.696866e-07,1.696882e-07,1.696897e-07,1.696913e-07,1.696929e-07,1.696944e-07,1.696960e-07,1.696976e-07,1.696991e-07,1.697007e-07,1.697023e-07,1.697038e-07,1.697054e-07,1.697070e-07,1.697085e-07,1.697101e-07,1.697117e-07,1.697132e-07,1.697148e-07,1.697164e-07,1.697179e-07,1.697195e-07,1.697211e-07,1.697226e-07,1.697242e-07,1.697257e-07,1.697273e-07,1.697289e-07,1.697304e-07,1.697320e-07,1.697336e-07,1.697351e-07,1.697367e-07,1.697382e-07,1.697398e-07,1.697414e-07,1.697429e-07,1.697445e-07,1.697460e-07,1.697476e-07,1.697492e-07,1.697507e-07,1.697523e-07,1.697538e-07,1.697554e-07,1.697570e-07,1.697585e-07,1.697601e-07,1.697616e-07,1.697632e-07,1.697648e-07,1.697663e-07,1.697679e-07,1.697694e-07,1.697710e-07,1.697725e-07,1.697741e-07,1.697757e-07,1.697772e-07,1.697788e-07,1.697803e-07,1.697819e-07,1.697834e-07,1.697850e-07,1.697865e-07,1.697881e-07,1.697896e-07,1.697912e-07,1.697928e-07,1.697943e-07,1.697959e-07,1.697974e-07,1.697990e-07,1.698005e-07,1.698021e-07,1.698036e-07,1.698052e-07,1.698067e-07,1.698083e-07,1.698098e-07,1.698114e-07,1.698129e-07,1.698145e-07,1.698160e-07,1.698176e-07,1.698191e-07,1.698207e-07,1.698222e-07,1.698238e-07,1.698253e-07,1.698269e-07,1.698284e-07,1.698300e-07,1.698315e-07,1.698331e-07,1.698346e-07,1.698362e-07,1.698377e-07,1.698393e-07,1.698408e-07,1.698424e-07,1.698439e-07,1.698455e-07,1.698470e-07,1.698486e-07,1.698501e-07,1.698517e-07,1.698532e-07,1.698548e-07,1.698563e-07,1.698578e-07,1.698594e-07,1.698609e-07,1.698625e-07,1.698640e-07,1.698656e-07,1.698671e-07,1.698687e-07,1.698702e-07,1.698717e-07,1.698733e-07,1.698748e-07,1.698764e-07,1.698779e-07,1.698795e-07,1.698810e-07,1.698825e-07,1.698841e-07,1.698856e-07,1.698872e-07,1.698887e-07,1.698902e-07,1.698918e-07,1.698933e-07,1.698949e-07,1.698964e-07,1.698980e-07,1.698995e-07,1.699010e-07,1.699026e-07,1.699041e-07,1.699056e-07,1.699072e-07,1.699087e-07,1.699103e-07,1.699118e-07,1.699133e-07,1.699149e-07,1.699164e-07,1.699180e-07,1.699195e-07,1.699210e-07,1.699226e-07,1.699241e-07,1.699256e-07,1.699272e-07,1.699287e-07,1.699302e-07,1.699318e-07,1.699333e-07,1.699349e-07,1.699364e-07,1.699379e-07,1.699395e-07,1.699410e-07,1.699425e-07,1.699441e-07,1.699456e-07,1.699471e-07,1.699487e-07,1.699502e-07,1.699517e-07,1.699533e-07,1.699548e-07,1.699563e-07,1.699579e-07,1.699594e-07,1.699609e-07,1.699625e-07,1.699640e-07,1.699655e-07,1.699670e-07,1.699686e-07,1.699701e-07,1.699716e-07,1.699732e-07,1.699747e-07,1.699762e-07,1.699778e-07,1.699793e-07,1.699808e-07,1.699823e-07,1.699839e-07,1.699854e-07,1.699869e-07,1.699885e-07,1.699900e-07,1.699915e-07,1.699930e-07,1.699946e-07,1.699961e-07,1.699976e-07,1.699991e-07,1.700007e-07,1.700022e-07,1.700037e-07,1.700053e-07,1.700068e-07,1.700083e-07,1.700098e-07,1.700114e-07,1.700129e-07,1.700144e-07,1.700159e-07,1.700175e-07,1.700190e-07,1.700205e-07,1.700220e-07,1.700236e-07,1.700251e-07,1.700266e-07,1.700281e-07,1.700296e-07,1.700312e-07,1.700327e-07,1.700342e-07,1.700357e-07,1.700373e-07,1.700388e-07,1.700403e-07,1.700418e-07,1.700433e-07,1.700449e-07,1.700464e-07,1.700479e-07,1.700494e-07,1.700509e-07,1.700525e-07,1.700540e-07,1.700555e-07,1.700570e-07,1.700585e-07,1.700601e-07,1.700616e-07,1.700631e-07,1.700646e-07,1.700661e-07,1.700676e-07,1.700692e-07,1.700707e-07,1.700722e-07,1.700737e-07,1.700752e-07,1.700767e-07,1.700783e-07,1.700798e-07,1.700813e-07,1.700828e-07,1.700843e-07,1.700858e-07,1.700874e-07,1.700889e-07,1.700904e-07,1.700919e-07,1.700934e-07,1.700949e-07,1.700964e-07,1.700980e-07,1.700995e-07,1.701010e-07,1.701025e-07,1.701040e-07,1.701055e-07,1.701070e-07,1.701086e-07,1.701101e-07,1.701116e-07,1.701131e-07,1.701146e-07,1.701161e-07,1.701176e-07,1.701191e-07,1.701206e-07,1.701222e-07,1.701237e-07,1.701252e-07,1.701267e-07,1.701282e-07,1.701297e-07,1.701312e-07,1.701327e-07,1.701342e-07,1.701357e-07,1.701372e-07,1.701388e-07,1.701403e-07,1.701418e-07,1.701433e-07,1.701448e-07,1.701463e-07,1.701478e-07,1.701493e-07,1.701508e-07,1.701523e-07,1.701538e-07,1.701553e-07,1.701568e-07,1.701584e-07,1.701599e-07,1.701614e-07,1.701629e-07,1.701644e-07,1.701659e-07,1.701674e-07,1.701689e-07,1.701704e-07,1.701719e-07,1.701734e-07,1.701749e-07,1.701764e-07,1.701779e-07,1.701794e-07,1.701809e-07,1.701824e-07,1.701839e-07,1.701854e-07,1.701869e-07,1.701884e-07,1.701899e-07,1.701914e-07,1.701929e-07,1.701944e-07,1.701959e-07,1.701974e-07,1.701989e-07,1.702004e-07,1.702019e-07,1.702034e-07,1.702049e-07,1.702064e-07,1.702079e-07,1.702094e-07,1.702109e-07,1.702124e-07,1.702139e-07,1.702154e-07,1.702169e-07,1.702184e-07,1.702199e-07,1.702214e-07,1.702229e-07,1.702244e-07,1.702259e-07,1.702274e-07,1.702289e-07,1.702304e-07,1.702319e-07,1.702334e-07,1.702349e-07,1.702364e-07,1.702379e-07,1.702394e-07,1.702409e-07,1.702424e-07,1.702439e-07,1.702454e-07,1.702469e-07,1.702484e-07,1.702498e-07,1.702513e-07,1.702528e-07,1.702543e-07,1.702558e-07,1.702573e-07,1.702588e-07,1.702603e-07,1.702618e-07,1.702633e-07,1.702648e-07,1.702663e-07,1.702678e-07,1.702693e-07,1.702707e-07,1.702722e-07,1.702737e-07,1.702752e-07,1.702767e-07,1.702782e-07,1.702797e-07,1.702812e-07,1.702827e-07,1.702842e-07,1.702856e-07,1.702871e-07,1.702886e-07,1.702901e-07,1.702916e-07,1.702931e-07,1.702946e-07,1.702961e-07,1.702976e-07,1.702990e-07,1.703005e-07,1.703020e-07,1.703035e-07,1.703050e-07,1.703065e-07,1.703080e-07,1.703095e-07,1.703109e-07,1.703124e-07,1.703139e-07,1.703154e-07,1.703169e-07,1.703184e-07,1.703199e-07,1.703213e-07,1.703228e-07,1.703243e-07,1.703258e-07,1.703273e-07,1.703288e-07,1.703302e-07,1.703317e-07,1.703332e-07,1.703347e-07,1.703362e-07,1.703377e-07,1.703391e-07,1.703406e-07,1.703421e-07,1.703436e-07,1.703451e-07,1.703466e-07,1.703480e-07,1.703495e-07,1.703510e-07,1.703525e-07,1.703540e-07,1.703554e-07,1.703569e-07,1.703584e-07,1.703599e-07,1.703614e-07,1.703628e-07,1.703643e-07,1.703658e-07,1.703673e-07,1.703688e-07,1.703702e-07,1.703717e-07,1.703732e-07,1.703747e-07,1.703762e-07,1.703776e-07,1.703791e-07,1.703806e-07,1.703821e-07,1.703835e-07,1.703850e-07,1.703865e-07,1.703880e-07,1.703894e-07,1.703909e-07,1.703924e-07,1.703939e-07,1.703954e-07,1.703968e-07,1.703983e-07,1.703998e-07,1.704013e-07,1.704027e-07,1.704042e-07,1.704057e-07,1.704071e-07,1.704086e-07,1.704101e-07,1.704116e-07,1.704130e-07,1.704145e-07,1.704160e-07,1.704175e-07,1.704189e-07,1.704204e-07,1.704219e-07,1.704234e-07,1.704248e-07,1.704263e-07,1.704278e-07,1.704292e-07,1.704307e-07,1.704322e-07,1.704336e-07,1.704351e-07,1.704366e-07,1.704381e-07,1.704395e-07,1.704410e-07,1.704425e-07,1.704439e-07,1.704454e-07,1.704469e-07,1.704483e-07,1.704498e-07,1.704513e-07,1.704528e-07,1.704542e-07,1.704557e-07,1.704572e-07,1.704586e-07,1.704601e-07,1.704616e-07,1.704630e-07,1.704645e-07,1.704660e-07,1.704674e-07,1.704689e-07,1.704704e-07,1.704718e-07,1.704733e-07,1.704748e-07,1.704762e-07,1.704777e-07,1.704791e-07,1.704806e-07,1.704821e-07,1.704835e-07,1.704850e-07,1.704865e-07,1.704879e-07,1.704894e-07,1.704909e-07,1.704923e-07,1.704938e-07,1.704953e-07,1.704967e-07,1.704982e-07,1.704996e-07,1.705011e-07,1.705026e-07,1.705040e-07,1.705055e-07,1.705069e-07,1.705084e-07,1.705099e-07,1.705113e-07,1.705128e-07,1.705143e-07,1.705157e-07,1.705172e-07,1.705186e-07,1.705201e-07,1.705216e-07,1.705230e-07,1.705245e-07,1.705259e-07,1.705274e-07,1.705288e-07,1.705303e-07,1.705318e-07,1.705332e-07,1.705347e-07,1.705361e-07,1.705376e-07,1.705391e-07,1.705405e-07,1.705420e-07,1.705434e-07,1.705449e-07,1.705463e-07,1.705478e-07,1.705493e-07,1.705507e-07,1.705522e-07,1.705536e-07,1.705551e-07,1.705565e-07,1.705580e-07,1.705594e-07,1.705609e-07,1.705623e-07,1.705638e-07,1.705653e-07,1.705667e-07,1.705682e-07,1.705696e-07,1.705711e-07,1.705725e-07,1.705740e-07,1.705754e-07,1.705769e-07,1.705783e-07,1.705798e-07,1.705812e-07,1.705827e-07,1.705841e-07,1.705856e-07,1.705870e-07,1.705885e-07,1.705899e-07,1.705914e-07,1.705928e-07,1.705943e-07,1.705958e-07,1.705972e-07,1.705987e-07,1.706001e-07,1.706016e-07,1.706030e-07,1.706044e-07,1.706059e-07,1.706073e-07,1.706088e-07,1.706102e-07,1.706117e-07,1.706131e-07,1.706146e-07,1.706160e-07,1.706175e-07,1.706189e-07,1.706204e-07,1.706218e-07,1.706233e-07,1.706247e-07,1.706262e-07,1.706276e-07,1.706291e-07,1.706305e-07,1.706320e-07,1.706334e-07,1.706348e-07,1.706363e-07,1.706377e-07,1.706392e-07,1.706406e-07,1.706421e-07,1.706435e-07,1.706450e-07,1.706464e-07,1.706478e-07,1.706493e-07,1.706507e-07,1.706522e-07,1.706536e-07,1.706551e-07,1.706565e-07,1.706579e-07,1.706594e-07,1.706608e-07,1.706623e-07,1.706637e-07,1.706652e-07,1.706666e-07,1.706680e-07,1.706695e-07,1.706709e-07,1.706724e-07,1.706738e-07,1.706752e-07,1.706767e-07,1.706781e-07,1.706796e-07,1.706810e-07,1.706824e-07,1.706839e-07,1.706853e-07,1.706868e-07,1.706882e-07,1.706896e-07,1.706911e-07,1.706925e-07,1.706940e-07,1.706954e-07,1.706968e-07,1.706983e-07,1.706997e-07,1.707011e-07,1.707026e-07,1.707040e-07,1.707054e-07,1.707069e-07,1.707083e-07,1.707098e-07,1.707112e-07,1.707126e-07,1.707141e-07,1.707155e-07,1.707169e-07,1.707184e-07,1.707198e-07,1.707212e-07,1.707227e-07,1.707241e-07,1.707255e-07,1.707270e-07,1.707284e-07,1.707298e-07,1.707313e-07,1.707327e-07,1.707341e-07,1.707356e-07,1.707370e-07,1.707384e-07,1.707399e-07,1.707413e-07,1.707427e-07,1.707442e-07,1.707456e-07,1.707470e-07,1.707485e-07,1.707499e-07,1.707513e-07,1.707528e-07,1.707542e-07,1.707556e-07,1.707571e-07,1.707585e-07,1.707599e-07,1.707613e-07,1.707628e-07,1.707642e-07,1.707656e-07,1.707671e-07,1.707685e-07,1.707699e-07,1.707713e-07,1.707728e-07,1.707742e-07,1.707756e-07,1.707771e-07,1.707785e-07,1.707799e-07,1.707813e-07,1.707828e-07,1.707842e-07,1.707856e-07,1.707870e-07,1.707885e-07,1.707899e-07,1.707913e-07,1.707928e-07,1.707942e-07,1.707956e-07,1.707970e-07,1.707985e-07,1.707999e-07,1.708013e-07,1.708027e-07,1.708042e-07,1.708056e-07,1.708070e-07,1.708084e-07,1.708099e-07,1.708113e-07,1.708127e-07,1.708141e-07,1.708155e-07,1.708170e-07,1.708184e-07,1.708198e-07,1.708212e-07,1.708227e-07,1.708241e-07,1.708255e-07,1.708269e-07,1.708283e-07,1.708298e-07,1.708312e-07,1.708326e-07,1.708340e-07,1.708355e-07,1.708369e-07,1.708383e-07,1.708397e-07,1.708411e-07,1.708426e-07,1.708440e-07,1.708454e-07,1.708468e-07,1.708482e-07,1.708496e-07,1.708511e-07,1.708525e-07,1.708539e-07,1.708553e-07,1.708567e-07,1.708582e-07,1.708596e-07,1.708610e-07,1.708624e-07,1.708638e-07,1.708652e-07,1.708667e-07,1.708681e-07,1.708695e-07,1.708709e-07,1.708723e-07,1.708737e-07,1.708752e-07,1.708766e-07,1.708780e-07,1.708794e-07,1.708808e-07,1.708822e-07,1.708837e-07,1.708851e-07,1.708865e-07,1.708879e-07,1.708893e-07,1.708907e-07,1.708921e-07,1.708936e-07,1.708950e-07,1.708964e-07,1.708978e-07,1.708992e-07,1.709006e-07,1.709020e-07,1.709034e-07,1.709049e-07,1.709063e-07,1.709077e-07,1.709091e-07,1.709105e-07,1.709119e-07,1.709133e-07,1.709147e-07,1.709161e-07,1.709176e-07,1.709190e-07,1.709204e-07,1.709218e-07,1.709232e-07,1.709246e-07,1.709260e-07,1.709274e-07,1.709288e-07,1.709302e-07,1.709317e-07,1.709331e-07,1.709345e-07,1.709359e-07,1.709373e-07,1.709387e-07,1.709401e-07,1.709415e-07,1.709429e-07,1.709443e-07,1.709457e-07,1.709471e-07,1.709485e-07,1.709500e-07,1.709514e-07,1.709528e-07,1.709542e-07,1.709556e-07,1.709570e-07,1.709584e-07,1.709598e-07,1.709612e-07,1.709626e-07,1.709640e-07,1.709654e-07,1.709668e-07,1.709682e-07,1.709696e-07,1.709710e-07,1.709724e-07,1.709738e-07,1.709752e-07,1.709767e-07,1.709781e-07,1.709795e-07,1.709809e-07,1.709823e-07,1.709837e-07,1.709851e-07,1.709865e-07,1.709879e-07,1.709893e-07,1.709907e-07,1.709921e-07,1.709935e-07,1.709949e-07,1.709963e-07,1.709977e-07,1.709991e-07,1.710005e-07,1.710019e-07,1.710033e-07,1.710047e-07,1.710061e-07,1.710075e-07,1.710089e-07,1.710103e-07,1.710117e-07,1.710131e-07,1.710145e-07,1.710159e-07,1.710173e-07,1.710187e-07,1.710201e-07,1.710215e-07,1.710229e-07,1.710243e-07,1.710257e-07,1.710271e-07,1.710285e-07,1.710299e-07,1.710313e-07,1.710327e-07,1.710341e-07,1.710354e-07,1.710368e-07,1.710382e-07,1.710396e-07,1.710410e-07,1.710424e-07,1.710438e-07,1.710452e-07,1.710466e-07,1.710480e-07,1.710494e-07,1.710508e-07,1.710522e-07,1.710536e-07,1.710550e-07,1.710564e-07,1.710578e-07,1.710592e-07,1.710606e-07,1.710620e-07,1.710633e-07,1.710647e-07,1.710661e-07,1.710675e-07,1.710689e-07,1.710703e-07,1.710717e-07,1.710731e-07,1.710745e-07,1.710759e-07,1.710773e-07,1.710787e-07,1.710800e-07,1.710814e-07,1.710828e-07,1.710842e-07,1.710856e-07,1.710870e-07,1.710884e-07,1.710898e-07,1.710912e-07,1.710926e-07,1.710940e-07,1.710953e-07,1.710967e-07,1.710981e-07,1.710995e-07,1.711009e-07,1.711023e-07,1.711037e-07,1.711051e-07,1.711064e-07,1.711078e-07,1.711092e-07,1.711106e-07,1.711120e-07,1.711134e-07,1.711148e-07,1.711162e-07,1.711175e-07,1.711189e-07,1.711203e-07,1.711217e-07,1.711231e-07,1.711245e-07,1.711259e-07,1.711272e-07,1.711286e-07,1.711300e-07,1.711314e-07,1.711328e-07,1.711342e-07,1.711356e-07,1.711369e-07,1.711383e-07,1.711397e-07,1.711411e-07,1.711425e-07,1.711439e-07,1.711452e-07,1.711466e-07,1.711480e-07,1.711494e-07,1.711508e-07,1.711522e-07,1.711535e-07,1.711549e-07,1.711563e-07,1.711577e-07,1.711591e-07,1.711604e-07,1.711618e-07,1.711632e-07,1.711646e-07,1.711660e-07,1.711674e-07,1.711687e-07,1.711701e-07,1.711715e-07,1.711729e-07,1.711743e-07,1.711756e-07,1.711770e-07,1.711784e-07,1.711798e-07,1.711812e-07,1.711825e-07,1.711839e-07,1.711853e-07,1.711867e-07,1.711880e-07,1.711894e-07,1.711908e-07,1.711922e-07,1.711936e-07,1.711949e-07,1.711963e-07,1.711977e-07,1.711991e-07,1.712004e-07,1.712018e-07,1.712032e-07,1.712046e-07,1.712059e-07,1.712073e-07,1.712087e-07,1.712101e-07,1.712115e-07,1.712128e-07,1.712142e-07,1.712156e-07,1.712170e-07,1.712183e-07,1.712197e-07,1.712211e-07,1.712224e-07,1.712238e-07,1.712252e-07,1.712266e-07,1.712279e-07,1.712293e-07,1.712307e-07,1.712321e-07,1.712334e-07,1.712348e-07,1.712362e-07,1.712376e-07,1.712389e-07,1.712403e-07,1.712417e-07,1.712430e-07,1.712444e-07,1.712458e-07,1.712472e-07,1.712485e-07,1.712499e-07,1.712513e-07,1.712526e-07,1.712540e-07,1.712554e-07,1.712568e-07,1.712581e-07,1.712595e-07,1.712609e-07,1.712622e-07,1.712636e-07,1.712650e-07,1.712663e-07,1.712677e-07,1.712691e-07,1.712704e-07,1.712718e-07,1.712732e-07,1.712745e-07,1.712759e-07,1.712773e-07,1.712787e-07,1.712800e-07,1.712814e-07,1.712828e-07,1.712841e-07,1.712855e-07,1.712869e-07,1.712882e-07,1.712896e-07,1.712910e-07,1.712923e-07,1.712937e-07,1.712950e-07,1.712964e-07,1.712978e-07,1.712991e-07,1.713005e-07,1.713019e-07,1.713032e-07,1.713046e-07,1.713060e-07,1.713073e-07,1.713087e-07,1.713101e-07,1.713114e-07,1.713128e-07,1.713142e-07,1.713155e-07,1.713169e-07,1.713182e-07,1.713196e-07,1.713210e-07,1.713223e-07,1.713237e-07,1.713251e-07,1.713264e-07,1.713278e-07,1.713291e-07,1.713305e-07,1.713319e-07,1.713332e-07,1.713346e-07,1.713359e-07,1.713373e-07,1.713387e-07,1.713400e-07,1.713414e-07,1.713427e-07,1.713441e-07,1.713455e-07,1.713468e-07,1.713482e-07,1.713495e-07,1.713509e-07,1.713523e-07,1.713536e-07,1.713550e-07,1.713563e-07,1.713577e-07,1.713591e-07,1.713604e-07,1.713618e-07,1.713631e-07,1.713645e-07,1.713658e-07,1.713672e-07,1.713686e-07,1.713699e-07,1.713713e-07,1.713726e-07,1.713740e-07,1.713753e-07,1.713767e-07,1.713781e-07,1.713794e-07,1.713808e-07,1.713821e-07,1.713835e-07,1.713848e-07,1.713862e-07,1.713875e-07,1.713889e-07,1.713902e-07,1.713916e-07,1.713930e-07,1.713943e-07,1.713957e-07,1.713970e-07,1.713984e-07,1.713997e-07,1.714011e-07,1.714024e-07,1.714038e-07,1.714051e-07,1.714065e-07,1.714078e-07,1.714092e-07,1.714105e-07,1.714119e-07,1.714132e-07,1.714146e-07,1.714160e-07,1.714173e-07,1.714187e-07,1.714200e-07,1.714214e-07,1.714227e-07,1.714241e-07,1.714254e-07,1.714268e-07,1.714281e-07,1.714295e-07,1.714308e-07,1.714322e-07,1.714335e-07,1.714349e-07,1.714362e-07,1.714376e-07,1.714389e-07,1.714403e-07,1.714416e-07,1.714429e-07,1.714443e-07,1.714456e-07,1.714470e-07,1.714483e-07,1.714497e-07,1.714510e-07,1.714524e-07,1.714537e-07,1.714551e-07,1.714564e-07,1.714578e-07,1.714591e-07,1.714605e-07,1.714618e-07,1.714632e-07,1.714645e-07,1.714658e-07,1.714672e-07,1.714685e-07,1.714699e-07,1.714712e-07,1.714726e-07,1.714739e-07,1.714753e-07,1.714766e-07,1.714780e-07,1.714793e-07,1.714806e-07,1.714820e-07,1.714833e-07,1.714847e-07,1.714860e-07,1.714874e-07,1.714887e-07,1.714900e-07,1.714914e-07,1.714927e-07,1.714941e-07,1.714954e-07,1.714968e-07,1.714981e-07,1.714994e-07,1.715008e-07,1.715021e-07,1.715035e-07,1.715048e-07,1.715061e-07,1.715075e-07,1.715088e-07,1.715102e-07,1.715115e-07,1.715128e-07,1.715142e-07,1.715155e-07,1.715169e-07,1.715182e-07,1.715195e-07,1.715209e-07,1.715222e-07,1.715236e-07,1.715249e-07,1.715262e-07,1.715276e-07,1.715289e-07,1.715303e-07,1.715316e-07,1.715329e-07,1.715343e-07,1.715356e-07,1.715369e-07,1.715383e-07,1.715396e-07,1.715410e-07,1.715423e-07,1.715436e-07,1.715450e-07,1.715463e-07,1.715476e-07,1.715490e-07,1.715503e-07,1.715517e-07,1.715530e-07,1.715543e-07,1.715557e-07,1.715570e-07,1.715583e-07,1.715597e-07,1.715610e-07,1.715623e-07,1.715637e-07,1.715650e-07,1.715663e-07,1.715677e-07,1.715690e-07,1.715703e-07,1.715717e-07,1.715730e-07,1.715743e-07,1.715757e-07,1.715770e-07,1.715783e-07,1.715797e-07,1.715810e-07,1.715823e-07,1.715837e-07,1.715850e-07,1.715863e-07,1.715877e-07,1.715890e-07,1.715903e-07,1.715917e-07,1.715930e-07,1.715943e-07,1.715956e-07,1.715970e-07,1.715983e-07,1.715996e-07,1.716010e-07,1.716023e-07,1.716036e-07,1.716050e-07,1.716063e-07,1.716076e-07,1.716089e-07,1.716103e-07,1.716116e-07,1.716129e-07,1.716143e-07,1.716156e-07,1.716169e-07,1.716182e-07,1.716196e-07,1.716209e-07,1.716222e-07,1.716236e-07,1.716249e-07,1.716262e-07,1.716275e-07,1.716289e-07,1.716302e-07,1.716315e-07,1.716328e-07,1.716342e-07,1.716355e-07,1.716368e-07,1.716382e-07,1.716395e-07,1.716408e-07,1.716421e-07,1.716435e-07,1.716448e-07,1.716461e-07,1.716474e-07,1.716488e-07,1.716501e-07,1.716514e-07,1.716527e-07,1.716540e-07,1.716554e-07,1.716567e-07,1.716580e-07,1.716593e-07,1.716607e-07,1.716620e-07,1.716633e-07,1.716646e-07,1.716660e-07,1.716673e-07,1.716686e-07,1.716699e-07,1.716712e-07,1.716726e-07,1.716739e-07,1.716752e-07,1.716765e-07,1.716779e-07,1.716792e-07,1.716805e-07,1.716818e-07,1.716831e-07,1.716845e-07,1.716858e-07,1.716871e-07,1.716884e-07,1.716897e-07,1.716911e-07,1.716924e-07,1.716937e-07,1.716950e-07,1.716963e-07,1.716977e-07,1.716990e-07,1.717003e-07,1.717016e-07,1.717029e-07,1.717043e-07,1.717056e-07,1.717069e-07,1.717082e-07,1.717095e-07,1.717108e-07,1.717122e-07,1.717135e-07,1.717148e-07,1.717161e-07,1.717174e-07,1.717187e-07,1.717201e-07,1.717214e-07,1.717227e-07,1.717240e-07,1.717253e-07,1.717266e-07,1.717280e-07,1.717293e-07,1.717306e-07,1.717319e-07,1.717332e-07,1.717345e-07,1.717358e-07,1.717372e-07,1.717385e-07,1.717398e-07,1.717411e-07,1.717424e-07,1.717437e-07,1.717450e-07,1.717464e-07,1.717477e-07,1.717490e-07,1.717503e-07,1.717516e-07,1.717529e-07,1.717542e-07,1.717556e-07,1.717569e-07,1.717582e-07,1.717595e-07,1.717608e-07,1.717621e-07,1.717634e-07,1.717647e-07,1.717660e-07,1.717674e-07,1.717687e-07,1.717700e-07,1.717713e-07,1.717726e-07,1.717739e-07,1.717752e-07,1.717765e-07,1.717778e-07,1.717792e-07,1.717805e-07,1.717818e-07,1.717831e-07,1.717844e-07,1.717857e-07,1.717870e-07,1.717883e-07,1.717896e-07,1.717909e-07,1.717922e-07,1.717936e-07,1.717949e-07,1.717962e-07,1.717975e-07,1.717988e-07,1.718001e-07,1.718014e-07,1.718027e-07,1.718040e-07,1.718053e-07,1.718066e-07,1.718079e-07,1.718092e-07,1.718105e-07,1.718119e-07,1.718132e-07,1.718145e-07,1.718158e-07,1.718171e-07,1.718184e-07,1.718197e-07,1.718210e-07,1.718223e-07,1.718236e-07,1.718249e-07,1.718262e-07,1.718275e-07,1.718288e-07,1.718301e-07,1.718314e-07,1.718327e-07,1.718340e-07,1.718353e-07,1.718366e-07,1.718379e-07,1.718393e-07,1.718406e-07,1.718419e-07,1.718432e-07,1.718445e-07,1.718458e-07,1.718471e-07,1.718484e-07,1.718497e-07,1.718510e-07,1.718523e-07,1.718536e-07,1.718549e-07,1.718562e-07,1.718575e-07,1.718588e-07,1.718601e-07,1.718614e-07,1.718627e-07,1.718640e-07,1.718653e-07,1.718666e-07,1.718679e-07,1.718692e-07,1.718705e-07,1.718718e-07,1.718731e-07,1.718744e-07,1.718757e-07,1.718770e-07,1.718783e-07,1.718796e-07,1.718809e-07,1.718822e-07,1.718835e-07,1.718848e-07,1.718861e-07,1.718874e-07,1.718887e-07,1.718900e-07,1.718913e-07,1.718926e-07,1.718939e-07,1.718952e-07,1.718964e-07,1.718977e-07,1.718990e-07,1.719003e-07,1.719016e-07,1.719029e-07,1.719042e-07,1.719055e-07,1.719068e-07,1.719081e-07,1.719094e-07,1.719107e-07,1.719120e-07,1.719133e-07,1.719146e-07,1.719159e-07,1.719172e-07,1.719185e-07,1.719198e-07,1.719211e-07,1.719224e-07,1.719236e-07,1.719249e-07,1.719262e-07,1.719275e-07,1.719288e-07,1.719301e-07,1.719314e-07,1.719327e-07,1.719340e-07,1.719353e-07,1.719366e-07,1.719379e-07,1.719392e-07,1.719405e-07,1.719417e-07,1.719430e-07,1.719443e-07,1.719456e-07,1.719469e-07,1.719482e-07,1.719495e-07,1.719508e-07,1.719521e-07,1.719534e-07,1.719547e-07,1.719559e-07,1.719572e-07,1.719585e-07,1.719598e-07,1.719611e-07,1.719624e-07,1.719637e-07,1.719650e-07,1.719663e-07,1.719675e-07,1.719688e-07,1.719701e-07,1.719714e-07,1.719727e-07,1.719740e-07,1.719753e-07,1.719766e-07,1.719779e-07,1.719791e-07,1.719804e-07,1.719817e-07,1.719830e-07,1.719843e-07,1.719856e-07,1.719869e-07,1.719882e-07,1.719894e-07,1.719907e-07,1.719920e-07,1.719933e-07,1.719946e-07,1.719959e-07,1.719972e-07,1.719984e-07,1.719997e-07,1.720010e-07,1.720023e-07,1.720036e-07,1.720049e-07,1.720061e-07,1.720074e-07,1.720087e-07,1.720100e-07,1.720113e-07,1.720126e-07,1.720139e-07,1.720151e-07,1.720164e-07,1.720177e-07,1.720190e-07,1.720203e-07,1.720216e-07,1.720228e-07,1.720241e-07,1.720254e-07,1.720267e-07,1.720280e-07,1.720292e-07,1.720305e-07,1.720318e-07,1.720331e-07,1.720344e-07,1.720357e-07,1.720369e-07,1.720382e-07,1.720395e-07,1.720408e-07,1.720421e-07,1.720433e-07,1.720446e-07,1.720459e-07,1.720472e-07,1.720485e-07,1.720497e-07,1.720510e-07,1.720523e-07,1.720536e-07,1.720549e-07,1.720561e-07,1.720574e-07,1.720587e-07,1.720600e-07,1.720613e-07,1.720625e-07,1.720638e-07,1.720651e-07,1.720664e-07,1.720676e-07,1.720689e-07,1.720702e-07,1.720715e-07,1.720728e-07,1.720740e-07,1.720753e-07,1.720766e-07,1.720779e-07,1.720791e-07,1.720804e-07,1.720817e-07,1.720830e-07,1.720842e-07,1.720855e-07,1.720868e-07,1.720881e-07,1.720893e-07,1.720906e-07,1.720919e-07,1.720932e-07,1.720944e-07,1.720957e-07,1.720970e-07,1.720983e-07,1.720995e-07,1.721008e-07,1.721021e-07,1.721034e-07,1.721046e-07,1.721059e-07,1.721072e-07,1.721085e-07,1.721097e-07,1.721110e-07,1.721123e-07,1.721135e-07,1.721148e-07,1.721161e-07,1.721174e-07,1.721186e-07,1.721199e-07,1.721212e-07,1.721225e-07,1.721237e-07,1.721250e-07,1.721263e-07,1.721275e-07,1.721288e-07,1.721301e-07,1.721314e-07,1.721326e-07,1.721339e-07,1.721352e-07,1.721364e-07,1.721377e-07,1.721390e-07,1.721402e-07,1.721415e-07,1.721428e-07,1.721441e-07,1.721453e-07,1.721466e-07,1.721479e-07,1.721491e-07,1.721504e-07,1.721517e-07,1.721529e-07,1.721542e-07,1.721555e-07,1.721567e-07,1.721580e-07,1.721593e-07,1.721605e-07,1.721618e-07,1.721631e-07,1.721643e-07,1.721656e-07,1.721669e-07,1.721681e-07,1.721694e-07,1.721707e-07,1.721719e-07,1.721732e-07,1.721745e-07,1.721757e-07,1.721770e-07,1.721783e-07,1.721795e-07,1.721808e-07,1.721821e-07,1.721833e-07,1.721846e-07,1.721859e-07,1.721871e-07,1.721884e-07,1.721897e-07,1.721909e-07,1.721922e-07,1.721935e-07,1.721947e-07,1.721960e-07,1.721972e-07,1.721985e-07,1.721998e-07,1.722010e-07,1.722023e-07,1.722036e-07,1.722048e-07,1.722061e-07,1.722074e-07,1.722086e-07,1.722099e-07,1.722111e-07,1.722124e-07,1.722137e-07,1.722149e-07,1.722162e-07,1.722174e-07,1.722187e-07,1.722200e-07,1.722212e-07,1.722225e-07,1.722238e-07,1.722250e-07,1.722263e-07,1.722275e-07,1.722288e-07,1.722301e-07,1.722313e-07,1.722326e-07,1.722338e-07,1.722351e-07,1.722364e-07,1.722376e-07,1.722389e-07,1.722401e-07,1.722414e-07,1.722426e-07,1.722439e-07,1.722452e-07,1.722464e-07,1.722477e-07,1.722489e-07,1.722502e-07,1.722515e-07,1.722527e-07,1.722540e-07,1.722552e-07,1.722565e-07,1.722577e-07,1.722590e-07,1.722603e-07,1.722615e-07,1.722628e-07,1.722640e-07,1.722653e-07,1.722665e-07,1.722678e-07,1.722690e-07,1.722703e-07,1.722716e-07,1.722728e-07,1.722741e-07,1.722753e-07,1.722766e-07,1.722778e-07,1.722791e-07,1.722803e-07,1.722816e-07,1.722829e-07,1.722841e-07,1.722854e-07,1.722866e-07,1.722879e-07,1.722891e-07,1.722904e-07,1.722916e-07,1.722929e-07,1.722941e-07,1.722954e-07,1.722966e-07,1.722979e-07,1.722991e-07,1.723004e-07,1.723017e-07,1.723029e-07,1.723042e-07,1.723054e-07,1.723067e-07,1.723079e-07,1.723092e-07,1.723104e-07,1.723117e-07,1.723129e-07,1.723142e-07,1.723154e-07,1.723167e-07,1.723179e-07,1.723192e-07,1.723204e-07,1.723217e-07,1.723229e-07,1.723242e-07,1.723254e-07,1.723267e-07,1.723279e-07,1.723292e-07,1.723304e-07,1.723317e-07,1.723329e-07,1.723342e-07,1.723354e-07,1.723367e-07,1.723379e-07,1.723392e-07,1.723404e-07,1.723417e-07,1.723429e-07,1.723442e-07,1.723454e-07,1.723466e-07,1.723479e-07,1.723491e-07,1.723504e-07,1.723516e-07,1.723529e-07,1.723541e-07,1.723554e-07,1.723566e-07,1.723579e-07,1.723591e-07,1.723604e-07,1.723616e-07,1.723629e-07,1.723641e-07,1.723653e-07,1.723666e-07,1.723678e-07,1.723691e-07,1.723703e-07,1.723716e-07,1.723728e-07,1.723741e-07,1.723753e-07,1.723765e-07,1.723778e-07,1.723790e-07,1.723803e-07,1.723815e-07,1.723828e-07,1.723840e-07,1.723853e-07,1.723865e-07,1.723877e-07,1.723890e-07,1.723902e-07,1.723915e-07,1.723927e-07,1.723940e-07,1.723952e-07,1.723964e-07,1.723977e-07,1.723989e-07,1.724002e-07,1.724014e-07,1.724026e-07,1.724039e-07,1.724051e-07,1.724064e-07,1.724076e-07,1.724089e-07,1.724101e-07,1.724113e-07,1.724126e-07,1.724138e-07,1.724151e-07,1.724163e-07,1.724175e-07,1.724188e-07,1.724200e-07,1.724213e-07,1.724225e-07,1.724237e-07,1.724250e-07,1.724262e-07,1.724275e-07,1.724287e-07,1.724299e-07,1.724312e-07,1.724324e-07,1.724336e-07,1.724349e-07,1.724361e-07,1.724374e-07,1.724386e-07,1.724398e-07,1.724411e-07,1.724423e-07,1.724435e-07,1.724448e-07,1.724460e-07,1.724473e-07,1.724485e-07,1.724497e-07,1.724510e-07,1.724522e-07,1.724534e-07,1.724547e-07,1.724559e-07,1.724571e-07,1.724584e-07,1.724596e-07,1.724609e-07,1.724621e-07,1.724633e-07,1.724646e-07,1.724658e-07,1.724670e-07,1.724683e-07,1.724695e-07,1.724707e-07,1.724720e-07,1.724732e-07,1.724744e-07,1.724757e-07,1.724769e-07,1.724781e-07,1.724794e-07,1.724806e-07,1.724818e-07,1.724831e-07,1.724843e-07,1.724855e-07,1.724868e-07,1.724880e-07,1.724892e-07,1.724905e-07,1.724917e-07,1.724929e-07,1.724942e-07,1.724954e-07,1.724966e-07,1.724978e-07,1.724991e-07,1.725003e-07,1.725015e-07,1.725028e-07,1.725040e-07,1.725052e-07,1.725065e-07,1.725077e-07,1.725089e-07,1.725102e-07,1.725114e-07,1.725126e-07,1.725138e-07,1.725151e-07,1.725163e-07,1.725175e-07,1.725188e-07,1.725200e-07,1.725212e-07,1.725224e-07,1.725237e-07,1.725249e-07,1.725261e-07,1.725274e-07,1.725286e-07,1.725298e-07,1.725310e-07,1.725323e-07,1.725335e-07,1.725347e-07,1.725360e-07,1.725372e-07,1.725384e-07,1.725396e-07,1.725409e-07,1.725421e-07,1.725433e-07,1.725445e-07,1.725458e-07,1.725470e-07,1.725482e-07,1.725494e-07,1.725507e-07,1.725519e-07,1.725531e-07,1.725544e-07,1.725556e-07,1.725568e-07,1.725580e-07,1.725593e-07,1.725605e-07,1.725617e-07,1.725629e-07,1.725642e-07,1.725654e-07,1.725666e-07,1.725678e-07,1.725690e-07,1.725703e-07,1.725715e-07,1.725727e-07,1.725739e-07,1.725752e-07,1.725764e-07,1.725776e-07,1.725788e-07,1.725801e-07,1.725813e-07,1.725825e-07,1.725837e-07,1.725849e-07,1.725862e-07,1.725874e-07,1.725886e-07,1.725898e-07,1.725911e-07,1.725923e-07,1.725935e-07,1.725947e-07,1.725959e-07,1.725972e-07,1.725984e-07,1.725996e-07,1.726008e-07,1.726020e-07,1.726033e-07,1.726045e-07,1.726057e-07,1.726069e-07,1.726081e-07,1.726094e-07,1.726106e-07,1.726118e-07,1.726130e-07,1.726142e-07,1.726155e-07,1.726167e-07,1.726179e-07,1.726191e-07,1.726203e-07,1.726216e-07,1.726228e-07,1.726240e-07,1.726252e-07,1.726264e-07,1.726276e-07,1.726289e-07,1.726301e-07,1.726313e-07,1.726325e-07,1.726337e-07,1.726349e-07,1.726362e-07,1.726374e-07,1.726386e-07,1.726398e-07,1.726410e-07,1.726422e-07,1.726435e-07,1.726447e-07,1.726459e-07,1.726471e-07,1.726483e-07,1.726495e-07,1.726508e-07,1.726520e-07,1.726532e-07,1.726544e-07,1.726556e-07,1.726568e-07,1.726580e-07,1.726593e-07,1.726605e-07,1.726617e-07,1.726629e-07,1.726641e-07,1.726653e-07,1.726665e-07,1.726678e-07,1.726690e-07,1.726702e-07,1.726714e-07,1.726726e-07,1.726738e-07,1.726750e-07,1.726762e-07,1.726775e-07,1.726787e-07,1.726799e-07,1.726811e-07,1.726823e-07,1.726835e-07,1.726847e-07,1.726859e-07,1.726872e-07,1.726884e-07,1.726896e-07,1.726908e-07,1.726920e-07,1.726932e-07,1.726944e-07,1.726956e-07,1.726968e-07,1.726981e-07,1.726993e-07,1.727005e-07,1.727017e-07,1.727029e-07,1.727041e-07,1.727053e-07,1.727065e-07,1.727077e-07,1.727089e-07,1.727102e-07,1.727114e-07,1.727126e-07,1.727138e-07,1.727150e-07,1.727162e-07,1.727174e-07,1.727186e-07,1.727198e-07,1.727210e-07,1.727222e-07,1.727234e-07,1.727246e-07,1.727259e-07,1.727271e-07,1.727283e-07,1.727295e-07,1.727307e-07,1.727319e-07,1.727331e-07,1.727343e-07,1.727355e-07,1.727367e-07,1.727379e-07,1.727391e-07,1.727403e-07,1.727415e-07,1.727427e-07,1.727440e-07,1.727452e-07,1.727464e-07,1.727476e-07,1.727488e-07,1.727500e-07,1.727512e-07,1.727524e-07,1.727536e-07,1.727548e-07,1.727560e-07,1.727572e-07,1.727584e-07,1.727596e-07,1.727608e-07,1.727620e-07,1.727632e-07,1.727644e-07,1.727656e-07,1.727668e-07,1.727680e-07,1.727692e-07,1.727704e-07,1.727716e-07,1.727729e-07,1.727741e-07,1.727753e-07,1.727765e-07,1.727777e-07,1.727789e-07,1.727801e-07,1.727813e-07,1.727825e-07,1.727837e-07,1.727849e-07,1.727861e-07,1.727873e-07,1.727885e-07,1.727897e-07,1.727909e-07,1.727921e-07,1.727933e-07,1.727945e-07,1.727957e-07,1.727969e-07,1.727981e-07,1.727993e-07,1.728005e-07,1.728017e-07,1.728029e-07,1.728041e-07,1.728053e-07,1.728065e-07,1.728077e-07,1.728089e-07,1.728101e-07,1.728113e-07,1.728125e-07,1.728137e-07,1.728149e-07,1.728161e-07,1.728173e-07,1.728185e-07,1.728197e-07,1.728209e-07,1.728221e-07,1.728232e-07,1.728244e-07,1.728256e-07,1.728268e-07,1.728280e-07,1.728292e-07,1.728304e-07,1.728316e-07,1.728328e-07,1.728340e-07,1.728352e-07,1.728364e-07,1.728376e-07,1.728388e-07,1.728400e-07,1.728412e-07,1.728424e-07,1.728436e-07,1.728448e-07,1.728460e-07,1.728472e-07,1.728484e-07,1.728496e-07,1.728508e-07,1.728520e-07,1.728531e-07,1.728543e-07,1.728555e-07,1.728567e-07,1.728579e-07,1.728591e-07,1.728603e-07,1.728615e-07,1.728627e-07,1.728639e-07,1.728651e-07,1.728663e-07,1.728675e-07,1.728687e-07,1.728699e-07,1.728710e-07,1.728722e-07,1.728734e-07,1.728746e-07,1.728758e-07,1.728770e-07,1.728782e-07,1.728794e-07,1.728806e-07,1.728818e-07,1.728830e-07,1.728842e-07,1.728853e-07,1.728865e-07,1.728877e-07,1.728889e-07,1.728901e-07,1.728913e-07,1.728925e-07,1.728937e-07,1.728949e-07,1.728961e-07,1.728972e-07,1.728984e-07,1.728996e-07,1.729008e-07,1.729020e-07,1.729032e-07,1.729044e-07,1.729056e-07,1.729068e-07,1.729080e-07,1.729091e-07,1.729103e-07,1.729115e-07,1.729127e-07,1.729139e-07,1.729151e-07,1.729163e-07,1.729175e-07,1.729186e-07,1.729198e-07,1.729210e-07,1.729222e-07,1.729234e-07,1.729246e-07,1.729258e-07,1.729270e-07,1.729281e-07,1.729293e-07,1.729305e-07,1.729317e-07,1.729329e-07,1.729341e-07,1.729353e-07,1.729364e-07,1.729376e-07,1.729388e-07,1.729400e-07,1.729412e-07,1.729424e-07,1.729436e-07,1.729447e-07,1.729459e-07,1.729471e-07,1.729483e-07,1.729495e-07,1.729507e-07,1.729518e-07,1.729530e-07,1.729542e-07,1.729554e-07,1.729566e-07,1.729578e-07,1.729590e-07,1.729601e-07,1.729613e-07,1.729625e-07,1.729637e-07,1.729649e-07,1.729661e-07,1.729672e-07,1.729684e-07,1.729696e-07,1.729708e-07,1.729720e-07,1.729731e-07,1.729743e-07,1.729755e-07,1.729767e-07,1.729779e-07,1.729791e-07,1.729802e-07,1.729814e-07,1.729826e-07,1.729838e-07,1.729850e-07,1.729861e-07,1.729873e-07,1.729885e-07,1.729897e-07,1.729909e-07,1.729920e-07,1.729932e-07,1.729944e-07,1.729956e-07,1.729968e-07,1.729979e-07,1.729991e-07,1.730003e-07,1.730015e-07,1.730027e-07,1.730038e-07,1.730050e-07,1.730062e-07,1.730074e-07,1.730086e-07,1.730097e-07,1.730109e-07,1.730121e-07,1.730133e-07,1.730144e-07,1.730156e-07,1.730168e-07,1.730180e-07,1.730192e-07,1.730203e-07,1.730215e-07,1.730227e-07,1.730239e-07,1.730250e-07,1.730262e-07,1.730274e-07,1.730286e-07,1.730297e-07,1.730309e-07,1.730321e-07,1.730333e-07,1.730344e-07,1.730356e-07,1.730368e-07,1.730380e-07,1.730392e-07,1.730403e-07,1.730415e-07,1.730427e-07,1.730439e-07,1.730450e-07,1.730462e-07,1.730474e-07,1.730485e-07,1.730497e-07,1.730509e-07,1.730521e-07,1.730532e-07,1.730544e-07,1.730556e-07,1.730568e-07,1.730579e-07,1.730591e-07,1.730603e-07,1.730615e-07,1.730626e-07,1.730638e-07,1.730650e-07,1.730662e-07,1.730673e-07,1.730685e-07,1.730697e-07,1.730708e-07,1.730720e-07,1.730732e-07,1.730744e-07,1.730755e-07,1.730767e-07,1.730779e-07,1.730790e-07,1.730802e-07,1.730814e-07,1.730826e-07,1.730837e-07,1.730849e-07,1.730861e-07,1.730872e-07,1.730884e-07,1.730896e-07,1.730908e-07,1.730919e-07,1.730931e-07,1.730943e-07,1.730954e-07,1.730966e-07,1.730978e-07,1.730989e-07,1.731001e-07,1.731013e-07,1.731024e-07,1.731036e-07,1.731048e-07,1.731060e-07,1.731071e-07,1.731083e-07,1.731095e-07,1.731106e-07,1.731118e-07,1.731130e-07,1.731141e-07,1.731153e-07,1.731165e-07,1.731176e-07,1.731188e-07,1.731200e-07,1.731211e-07,1.731223e-07,1.731235e-07,1.731246e-07,1.731258e-07,1.731270e-07,1.731281e-07,1.731293e-07,1.731305e-07,1.731316e-07,1.731328e-07,1.731340e-07,1.731351e-07,1.731363e-07,1.731375e-07,1.731386e-07,1.731398e-07,1.731410e-07,1.731421e-07,1.731433e-07,1.731445e-07,1.731456e-07,1.731468e-07,1.731479e-07,1.731491e-07,1.731503e-07,1.731514e-07,1.731526e-07,1.731538e-07,1.731549e-07,1.731561e-07,1.731573e-07,1.731584e-07,1.731596e-07,1.731607e-07,1.731619e-07,1.731631e-07,1.731642e-07,1.731654e-07,1.731666e-07,1.731677e-07,1.731689e-07,1.731700e-07,1.731712e-07,1.731724e-07,1.731735e-07,1.731747e-07,1.731759e-07,1.731770e-07,1.731782e-07,1.731793e-07,1.731805e-07,1.731817e-07,1.731828e-07,1.731840e-07,1.731851e-07,1.731863e-07,1.731875e-07,1.731886e-07,1.731898e-07,1.731909e-07,1.731921e-07,1.731933e-07,1.731944e-07,1.731956e-07,1.731967e-07,1.731979e-07,1.731991e-07,1.732002e-07,1.732014e-07,1.732025e-07,1.732037e-07,1.732049e-07,1.732060e-07,1.732072e-07,1.732083e-07,1.732095e-07,1.732107e-07,1.732118e-07,1.732130e-07,1.732141e-07,1.732153e-07,1.732164e-07,1.732176e-07,1.732188e-07,1.732199e-07,1.732211e-07,1.732222e-07,1.732234e-07,1.732245e-07,1.732257e-07,1.732269e-07,1.732280e-07,1.732292e-07,1.732303e-07,1.732315e-07,1.732326e-07,1.732338e-07,1.732349e-07,1.732361e-07,1.732373e-07,1.732384e-07,1.732396e-07,1.732407e-07,1.732419e-07,1.732430e-07,1.732442e-07,1.732453e-07,1.732465e-07,1.732477e-07,1.732488e-07,1.732500e-07,1.732511e-07,1.732523e-07,1.732534e-07,1.732546e-07,1.732557e-07,1.732569e-07,1.732580e-07,1.732592e-07,1.732603e-07,1.732615e-07,1.732627e-07,1.732638e-07,1.732650e-07,1.732661e-07,1.732673e-07,1.732684e-07,1.732696e-07,1.732707e-07,1.732719e-07,1.732730e-07,1.732742e-07,1.732753e-07,1.732765e-07,1.732776e-07,1.732788e-07,1.732799e-07,1.732811e-07,1.732822e-07,1.732834e-07,1.732845e-07,1.732857e-07,1.732868e-07,1.732880e-07,1.732891e-07,1.732903e-07,1.732914e-07,1.732926e-07,1.732937e-07,1.732949e-07,1.732960e-07,1.732972e-07,1.732983e-07,1.732995e-07,1.733006e-07,1.733018e-07,1.733029e-07,1.733041e-07,1.733052e-07,1.733064e-07,1.733075e-07,1.733087e-07,1.733098e-07,1.733110e-07,1.733121e-07,1.733133e-07,1.733144e-07,1.733156e-07,1.733167e-07,1.733179e-07,1.733190e-07,1.733202e-07,1.733213e-07,1.733225e-07,1.733236e-07,1.733247e-07,1.733259e-07,1.733270e-07,1.733282e-07,1.733293e-07,1.733305e-07,1.733316e-07,1.733328e-07,1.733339e-07,1.733351e-07,1.733362e-07,1.733374e-07,1.733385e-07,1.733396e-07,1.733408e-07,1.733419e-07,1.733431e-07,1.733442e-07,1.733454e-07,1.733465e-07,1.733477e-07,1.733488e-07,1.733499e-07,1.733511e-07,1.733522e-07,1.733534e-07,1.733545e-07,1.733557e-07,1.733568e-07,1.733580e-07,1.733591e-07,1.733602e-07,1.733614e-07,1.733625e-07,1.733637e-07,1.733648e-07,1.733660e-07,1.733671e-07,1.733682e-07,1.733694e-07,1.733705e-07,1.733717e-07,1.733728e-07,1.733740e-07,1.733751e-07,1.733762e-07,1.733774e-07,1.733785e-07,1.733797e-07,1.733808e-07,1.733819e-07,1.733831e-07,1.733842e-07,1.733854e-07,1.733865e-07,1.733877e-07,1.733888e-07,1.733899e-07,1.733911e-07,1.733922e-07,1.733934e-07,1.733945e-07,1.733956e-07,1.733968e-07,1.733979e-07,1.733991e-07,1.734002e-07,1.734013e-07,1.734025e-07,1.734036e-07,1.734047e-07,1.734059e-07,1.734070e-07,1.734082e-07,1.734093e-07,1.734104e-07,1.734116e-07,1.734127e-07,1.734139e-07,1.734150e-07,1.734161e-07,1.734173e-07,1.734184e-07,1.734195e-07,1.734207e-07,1.734218e-07,1.734230e-07,1.734241e-07,1.734252e-07,1.734264e-07,1.734275e-07,1.734286e-07,1.734298e-07,1.734309e-07,1.734321e-07,1.734332e-07,1.734343e-07,1.734355e-07,1.734366e-07,1.734377e-07,1.734389e-07,1.734400e-07,1.734411e-07,1.734423e-07,1.734434e-07,1.734445e-07,1.734457e-07,1.734468e-07,1.734479e-07,1.734491e-07,1.734502e-07,1.734514e-07,1.734525e-07,1.734536e-07,1.734548e-07,1.734559e-07,1.734570e-07,1.734582e-07,1.734593e-07,1.734604e-07,1.734616e-07,1.734627e-07,1.734638e-07,1.734650e-07,1.734661e-07,1.734672e-07,1.734684e-07,1.734695e-07,1.734706e-07,1.734718e-07,1.734729e-07,1.734740e-07,1.734751e-07,1.734763e-07,1.734774e-07,1.734785e-07,1.734797e-07,1.734808e-07,1.734819e-07,1.734831e-07,1.734842e-07,1.734853e-07,1.734865e-07,1.734876e-07,1.734887e-07,1.734899e-07,1.734910e-07,1.734921e-07,1.734932e-07,1.734944e-07,1.734955e-07,1.734966e-07,1.734978e-07,1.734989e-07,1.735000e-07,1.735012e-07,1.735023e-07,1.735034e-07,1.735045e-07,1.735057e-07,1.735068e-07,1.735079e-07,1.735091e-07,1.735102e-07,1.735113e-07,1.735124e-07,1.735136e-07,1.735147e-07,1.735158e-07,1.735170e-07,1.735181e-07,1.735192e-07,1.735203e-07,1.735215e-07,1.735226e-07,1.735237e-07,1.735249e-07,1.735260e-07,1.735271e-07,1.735282e-07,1.735294e-07,1.735305e-07,1.735316e-07,1.735327e-07,1.735339e-07,1.735350e-07,1.735361e-07,1.735372e-07,1.735384e-07,1.735395e-07,1.735406e-07,1.735418e-07,1.735429e-07,1.735440e-07,1.735451e-07,1.735463e-07,1.735474e-07,1.735485e-07,1.735496e-07,1.735508e-07,1.735519e-07,1.735530e-07,1.735541e-07,1.735553e-07,1.735564e-07,1.735575e-07,1.735586e-07,1.735597e-07,1.735609e-07,1.735620e-07,1.735631e-07,1.735642e-07,1.735654e-07,1.735665e-07,1.735676e-07,1.735687e-07,1.735699e-07,1.735710e-07,1.735721e-07,1.735732e-07,1.735743e-07,1.735755e-07,1.735766e-07,1.735777e-07,1.735788e-07,1.735800e-07,1.735811e-07,1.735822e-07,1.735833e-07,1.735844e-07,1.735856e-07,1.735867e-07,1.735878e-07,1.735889e-07,1.735901e-07,1.735912e-07,1.735923e-07,1.735934e-07,1.735945e-07,1.735957e-07,1.735968e-07,1.735979e-07,1.735990e-07,1.736001e-07,1.736013e-07,1.736024e-07,1.736035e-07,1.736046e-07,1.736057e-07,1.736069e-07,1.736080e-07,1.736091e-07,1.736102e-07,1.736113e-07,1.736125e-07,1.736136e-07,1.736147e-07,1.736158e-07,1.736169e-07,1.736180e-07,1.736192e-07,1.736203e-07,1.736214e-07,1.736225e-07,1.736236e-07,1.736248e-07,1.736259e-07,1.736270e-07,1.736281e-07,1.736292e-07,1.736303e-07,1.736315e-07,1.736326e-07,1.736337e-07,1.736348e-07,1.736359e-07,1.736370e-07,1.736382e-07,1.736393e-07,1.736404e-07,1.736415e-07,1.736426e-07,1.736437e-07,1.736449e-07,1.736460e-07,1.736471e-07,1.736482e-07,1.736493e-07,1.736504e-07,1.736515e-07,1.736527e-07,1.736538e-07,1.736549e-07,1.736560e-07,1.736571e-07,1.736582e-07,1.736593e-07,1.736605e-07,1.736616e-07,1.736627e-07,1.736638e-07,1.736649e-07,1.736660e-07,1.736671e-07,1.736683e-07,1.736694e-07,1.736705e-07,1.736716e-07,1.736727e-07,1.736738e-07,1.736749e-07,1.736760e-07,1.736772e-07,1.736783e-07,1.736794e-07,1.736805e-07,1.736816e-07,1.736827e-07,1.736838e-07,1.736849e-07,1.736861e-07,1.736872e-07,1.736883e-07,1.736894e-07,1.736905e-07,1.736916e-07,1.736927e-07,1.736938e-07,1.736949e-07,1.736961e-07,1.736972e-07,1.736983e-07,1.736994e-07,1.737005e-07,1.737016e-07,1.737027e-07,1.737038e-07,1.737049e-07,1.737061e-07,1.737072e-07,1.737083e-07,1.737094e-07,1.737105e-07,1.737116e-07,1.737127e-07,1.737138e-07,1.737149e-07,1.737160e-07,1.737171e-07,1.737183e-07,1.737194e-07,1.737205e-07,1.737216e-07,1.737227e-07,1.737238e-07,1.737249e-07,1.737260e-07,1.737271e-07,1.737282e-07,1.737293e-07,1.737304e-07,1.737316e-07,1.737327e-07,1.737338e-07,1.737349e-07,1.737360e-07,1.737371e-07,1.737382e-07,1.737393e-07,1.737404e-07,1.737415e-07,1.737426e-07,1.737437e-07,1.737448e-07,1.737459e-07,1.737470e-07,1.737482e-07,1.737493e-07,1.737504e-07,1.737515e-07,1.737526e-07,1.737537e-07,1.737548e-07,1.737559e-07,1.737570e-07,1.737581e-07,1.737592e-07,1.737603e-07,1.737614e-07,1.737625e-07,1.737636e-07,1.737647e-07,1.737658e-07,1.737669e-07,1.737680e-07,1.737691e-07,1.737702e-07,1.737713e-07,1.737725e-07,1.737736e-07,1.737747e-07,1.737758e-07,1.737769e-07,1.737780e-07,1.737791e-07,1.737802e-07,1.737813e-07,1.737824e-07,1.737835e-07,1.737846e-07,1.737857e-07,1.737868e-07,1.737879e-07,1.737890e-07,1.737901e-07,1.737912e-07,1.737923e-07,1.737934e-07,1.737945e-07,1.737956e-07,1.737967e-07,1.737978e-07,1.737989e-07,1.738000e-07,1.738011e-07,1.738022e-07,1.738033e-07,1.738044e-07,1.738055e-07,1.738066e-07,1.738077e-07,1.738088e-07,1.738099e-07,1.738110e-07,1.738121e-07,1.738132e-07,1.738143e-07,1.738154e-07,1.738165e-07,1.738176e-07,1.738187e-07,1.738198e-07,1.738209e-07,1.738220e-07,1.738231e-07,1.738242e-07,1.738253e-07,1.738264e-07,1.738275e-07,1.738286e-07,1.738297e-07,1.738308e-07,1.738319e-07,1.738330e-07,1.738341e-07,1.738352e-07,1.738363e-07,1.738374e-07,1.738385e-07,1.738396e-07,1.738407e-07,1.738418e-07,1.738429e-07,1.738440e-07,1.738451e-07,1.738462e-07,1.738473e-07,1.738483e-07,1.738494e-07,1.738505e-07,1.738516e-07,1.738527e-07,1.738538e-07,1.738549e-07,1.738560e-07,1.738571e-07,1.738582e-07,1.738593e-07,1.738604e-07,1.738615e-07,1.738626e-07,1.738637e-07,1.738648e-07,1.738659e-07,1.738670e-07,1.738681e-07,1.738692e-07,1.738703e-07,1.738713e-07,1.738724e-07,1.738735e-07,1.738746e-07,1.738757e-07,1.738768e-07,1.738779e-07,1.738790e-07,1.738801e-07,1.738812e-07,1.738823e-07,1.738834e-07,1.738845e-07,1.738856e-07,1.738867e-07,1.738877e-07,1.738888e-07,1.738899e-07,1.738910e-07,1.738921e-07,1.738932e-07,1.738943e-07,1.738954e-07,1.738965e-07,1.738976e-07,1.738987e-07,1.738998e-07,1.739009e-07,1.739019e-07,1.739030e-07,1.739041e-07,1.739052e-07,1.739063e-07,1.739074e-07,1.739085e-07,1.739096e-07,1.739107e-07,1.739118e-07,1.739129e-07,1.739139e-07,1.739150e-07,1.739161e-07,1.739172e-07,1.739183e-07,1.739194e-07,1.739205e-07,1.739216e-07,1.739227e-07,1.739238e-07,1.739248e-07,1.739259e-07,1.739270e-07,1.739281e-07,1.739292e-07,1.739303e-07,1.739314e-07,1.739325e-07,1.739335e-07,1.739346e-07,1.739357e-07,1.739368e-07,1.739379e-07,1.739390e-07,1.739401e-07,1.739412e-07,1.739423e-07,1.739433e-07,1.739444e-07,1.739455e-07,1.739466e-07,1.739477e-07,1.739488e-07,1.739499e-07,1.739509e-07,1.739520e-07,1.739531e-07,1.739542e-07,1.739553e-07,1.739564e-07,1.739575e-07,1.739586e-07,1.739596e-07,1.739607e-07,1.739618e-07,1.739629e-07,1.739640e-07,1.739651e-07,1.739662e-07,1.739672e-07,1.739683e-07,1.739694e-07,1.739705e-07,1.739716e-07,1.739727e-07,1.739737e-07,1.739748e-07,1.739759e-07,1.739770e-07,1.739781e-07,1.739792e-07,1.739803e-07,1.739813e-07,1.739824e-07,1.739835e-07,1.739846e-07,1.739857e-07,1.739868e-07,1.739878e-07,1.739889e-07,1.739900e-07,1.739911e-07,1.739922e-07,1.739933e-07,1.739943e-07,1.739954e-07,1.739965e-07,1.739976e-07,1.739987e-07,1.739997e-07,1.740008e-07,1.740019e-07,1.740030e-07,1.740041e-07,1.740052e-07,1.740062e-07,1.740073e-07,1.740084e-07,1.740095e-07,1.740106e-07,1.740116e-07,1.740127e-07,1.740138e-07,1.740149e-07,1.740160e-07,1.740171e-07,1.740181e-07,1.740192e-07,1.740203e-07,1.740214e-07,1.740225e-07,1.740235e-07,1.740246e-07,1.740257e-07,1.740268e-07,1.740279e-07,1.740289e-07,1.740300e-07,1.740311e-07,1.740322e-07,1.740332e-07,1.740343e-07,1.740354e-07,1.740365e-07,1.740376e-07,1.740386e-07,1.740397e-07,1.740408e-07,1.740419e-07,1.740430e-07,1.740440e-07,1.740451e-07,1.740462e-07,1.740473e-07,1.740483e-07,1.740494e-07,1.740505e-07,1.740516e-07,1.740527e-07,1.740537e-07,1.740548e-07,1.740559e-07,1.740570e-07,1.740580e-07,1.740591e-07,1.740602e-07,1.740613e-07,1.740623e-07,1.740634e-07,1.740645e-07,1.740656e-07,1.740667e-07,1.740677e-07,1.740688e-07,1.740699e-07,1.740710e-07,1.740720e-07,1.740731e-07,1.740742e-07,1.740753e-07,1.740763e-07,1.740774e-07,1.740785e-07,1.740796e-07,1.740806e-07,1.740817e-07,1.740828e-07,1.740839e-07,1.740849e-07,1.740860e-07,1.740871e-07,1.740882e-07,1.740892e-07,1.740903e-07,1.740914e-07,1.740924e-07,1.740935e-07,1.740946e-07,1.740957e-07,1.740967e-07,1.740978e-07,1.740989e-07,1.741000e-07,1.741010e-07,1.741021e-07,1.741032e-07,1.741042e-07,1.741053e-07,1.741064e-07,1.741075e-07,1.741085e-07,1.741096e-07,1.741107e-07,1.741118e-07,1.741128e-07,1.741139e-07,1.741150e-07,1.741160e-07,1.741171e-07,1.741182e-07,1.741193e-07,1.741203e-07,1.741214e-07,1.741225e-07,1.741235e-07,1.741246e-07,1.741257e-07,1.741267e-07,1.741278e-07,1.741289e-07,1.741300e-07,1.741310e-07,1.741321e-07,1.741332e-07,1.741342e-07,1.741353e-07,1.741364e-07,1.741374e-07,1.741385e-07,1.741396e-07,1.741407e-07,1.741417e-07,1.741428e-07,1.741439e-07,1.741449e-07,1.741460e-07,1.741471e-07,1.741481e-07,1.741492e-07,1.741503e-07,1.741513e-07,1.741524e-07,1.741535e-07,1.741545e-07,1.741556e-07,1.741567e-07,1.741578e-07,1.741588e-07,1.741599e-07,1.741610e-07,1.741620e-07,1.741631e-07,1.741642e-07,1.741652e-07,1.741663e-07,1.741674e-07,1.741684e-07,1.741695e-07,1.741706e-07,1.741716e-07,1.741727e-07,1.741738e-07,1.741748e-07,1.741759e-07,1.741770e-07,1.741780e-07,1.741791e-07,1.741801e-07,1.741812e-07,1.741823e-07,1.741833e-07,1.741844e-07,1.741855e-07,1.741865e-07,1.741876e-07,1.741887e-07,1.741897e-07,1.741908e-07,1.741919e-07,1.741929e-07,1.741940e-07,1.741951e-07,1.741961e-07,1.741972e-07,1.741982e-07,1.741993e-07,1.742004e-07,1.742014e-07,1.742025e-07,1.742036e-07,1.742046e-07,1.742057e-07,1.742068e-07,1.742078e-07,1.742089e-07,1.742099e-07,1.742110e-07,1.742121e-07,1.742131e-07,1.742142e-07,1.742153e-07,1.742163e-07,1.742174e-07,1.742184e-07,1.742195e-07,1.742206e-07,1.742216e-07,1.742227e-07,1.742238e-07,1.742248e-07,1.742259e-07,1.742269e-07,1.742280e-07,1.742291e-07,1.742301e-07,1.742312e-07,1.742322e-07,1.742333e-07,1.742344e-07,1.742354e-07,1.742365e-07,1.742375e-07,1.742386e-07,1.742397e-07,1.742407e-07,1.742418e-07,1.742428e-07,1.742439e-07,1.742450e-07,1.742460e-07,1.742471e-07,1.742481e-07,1.742492e-07,1.742503e-07,1.742513e-07,1.742524e-07,1.742534e-07,1.742545e-07,1.742556e-07,1.742566e-07,1.742577e-07,1.742587e-07,1.742598e-07,1.742608e-07,1.742619e-07,1.742630e-07,1.742640e-07,1.742651e-07,1.742661e-07,1.742672e-07,1.742683e-07,1.742693e-07,1.742704e-07,1.742714e-07,1.742725e-07,1.742735e-07,1.742746e-07,1.742757e-07,1.742767e-07,1.742778e-07,1.742788e-07,1.742799e-07,1.742809e-07,1.742820e-07,1.742830e-07,1.742841e-07,1.742852e-07,1.742862e-07,1.742873e-07,1.742883e-07,1.742894e-07,1.742904e-07,1.742915e-07,1.742925e-07,1.742936e-07,1.742947e-07,1.742957e-07,1.742968e-07,1.742978e-07,1.742989e-07,1.742999e-07,1.743010e-07,1.743020e-07,1.743031e-07,1.743042e-07,1.743052e-07,1.743063e-07,1.743073e-07,1.743084e-07,1.743094e-07,1.743105e-07,1.743115e-07,1.743126e-07,1.743136e-07,1.743147e-07,1.743157e-07,1.743168e-07,1.743178e-07,1.743189e-07,1.743200e-07,1.743210e-07,1.743221e-07,1.743231e-07,1.743242e-07,1.743252e-07,1.743263e-07,1.743273e-07,1.743284e-07,1.743294e-07,1.743305e-07,1.743315e-07,1.743326e-07,1.743336e-07,1.743347e-07,1.743357e-07,1.743368e-07,1.743378e-07,1.743389e-07,1.743399e-07,1.743410e-07,1.743420e-07,1.743431e-07,1.743441e-07,1.743452e-07,1.743462e-07,1.743473e-07,1.743483e-07,1.743494e-07,1.743504e-07,1.743515e-07,1.743525e-07,1.743536e-07,1.743546e-07,1.743557e-07,1.743567e-07,1.743578e-07,1.743588e-07,1.743599e-07,1.743609e-07,1.743620e-07,1.743630e-07,1.743641e-07,1.743651e-07,1.743662e-07,1.743672e-07,1.743683e-07,1.743693e-07,1.743704e-07,1.743714e-07,1.743725e-07,1.743735e-07,1.743746e-07,1.743756e-07,1.743767e-07,1.743777e-07,1.743788e-07,1.743798e-07,1.743809e-07,1.743819e-07,1.743829e-07,1.743840e-07,1.743850e-07,1.743861e-07,1.743871e-07,1.743882e-07,1.743892e-07,1.743903e-07,1.743913e-07,1.743924e-07,1.743934e-07,1.743945e-07,1.743955e-07,1.743966e-07,1.743976e-07,1.743986e-07,1.743997e-07,1.744007e-07,1.744018e-07,1.744028e-07,1.744039e-07,1.744049e-07,1.744060e-07,1.744070e-07,1.744081e-07,1.744091e-07,1.744101e-07,1.744112e-07,1.744122e-07,1.744133e-07,1.744143e-07,1.744154e-07,1.744164e-07,1.744175e-07,1.744185e-07,1.744195e-07,1.744206e-07,1.744216e-07,1.744227e-07,1.744237e-07,1.744248e-07,1.744258e-07,1.744268e-07,1.744279e-07,1.744289e-07,1.744300e-07,1.744310e-07,1.744321e-07,1.744331e-07,1.744341e-07,1.744352e-07,1.744362e-07,1.744373e-07,1.744383e-07,1.744394e-07,1.744404e-07,1.744414e-07,1.744425e-07,1.744435e-07,1.744446e-07,1.744456e-07,1.744466e-07,1.744477e-07,1.744487e-07,1.744498e-07,1.744508e-07,1.744519e-07,1.744529e-07,1.744539e-07,1.744550e-07,1.744560e-07,1.744571e-07,1.744581e-07,1.744591e-07,1.744602e-07,1.744612e-07,1.744623e-07,1.744633e-07,1.744643e-07,1.744654e-07,1.744664e-07,1.744675e-07,1.744685e-07,1.744695e-07,1.744706e-07,1.744716e-07,1.744727e-07,1.744737e-07,1.744747e-07,1.744758e-07,1.744768e-07,1.744778e-07,1.744789e-07,1.744799e-07,1.744810e-07,1.744820e-07,1.744830e-07,1.744841e-07,1.744851e-07,1.744862e-07,1.744872e-07,1.744882e-07,1.744893e-07,1.744903e-07,1.744913e-07,1.744924e-07,1.744934e-07,1.744945e-07,1.744955e-07,1.744965e-07,1.744976e-07,1.744986e-07,1.744996e-07,1.745007e-07,1.745017e-07,1.745027e-07,1.745038e-07,1.745048e-07,1.745059e-07,1.745069e-07,1.745079e-07,1.745090e-07,1.745100e-07,1.745110e-07,1.745121e-07,1.745131e-07,1.745141e-07,1.745152e-07,1.745162e-07,1.745172e-07,1.745183e-07,1.745193e-07,1.745204e-07,1.745214e-07,1.745224e-07,1.745235e-07,1.745245e-07,1.745255e-07,1.745266e-07,1.745276e-07,1.745286e-07,1.745297e-07,1.745307e-07,1.745317e-07,1.745328e-07,1.745338e-07,1.745348e-07,1.745359e-07,1.745369e-07,1.745379e-07,1.745390e-07,1.745400e-07,1.745410e-07,1.745421e-07,1.745431e-07,1.745441e-07,1.745452e-07,1.745462e-07,1.745472e-07,1.745483e-07,1.745493e-07,1.745503e-07,1.745514e-07,1.745524e-07,1.745534e-07,1.745545e-07,1.745555e-07,1.745565e-07,1.745575e-07,1.745586e-07,1.745596e-07,1.745606e-07,1.745617e-07,1.745627e-07,1.745637e-07,1.745648e-07,1.745658e-07,1.745668e-07,1.745679e-07,1.745689e-07,1.745699e-07,1.745709e-07,1.745720e-07,1.745730e-07,1.745740e-07,1.745751e-07,1.745761e-07,1.745771e-07,1.745782e-07,1.745792e-07,1.745802e-07,1.745812e-07,1.745823e-07,1.745833e-07,1.745843e-07,1.745854e-07,1.745864e-07,1.745874e-07,1.745885e-07,1.745895e-07,1.745905e-07,1.745915e-07,1.745926e-07,1.745936e-07,1.745946e-07,1.745957e-07,1.745967e-07,1.745977e-07,1.745987e-07,1.745998e-07,1.746008e-07,1.746018e-07,1.746028e-07,1.746039e-07,1.746049e-07,1.746059e-07,1.746070e-07,1.746080e-07,1.746090e-07,1.746100e-07,1.746111e-07,1.746121e-07,1.746131e-07,1.746141e-07,1.746152e-07,1.746162e-07,1.746172e-07,1.746182e-07,1.746193e-07,1.746203e-07,1.746213e-07,1.746224e-07,1.746234e-07,1.746244e-07,1.746254e-07,1.746265e-07,1.746275e-07,1.746285e-07,1.746295e-07,1.746306e-07,1.746316e-07,1.746326e-07,1.746336e-07,1.746347e-07,1.746357e-07,1.746367e-07,1.746377e-07,1.746388e-07,1.746398e-07,1.746408e-07,1.746418e-07,1.746428e-07,1.746439e-07,1.746449e-07,1.746459e-07,1.746469e-07,1.746480e-07,1.746490e-07,1.746500e-07,1.746510e-07,1.746521e-07,1.746531e-07,1.746541e-07,1.746551e-07,1.746562e-07,1.746572e-07,1.746582e-07,1.746592e-07,1.746602e-07,1.746613e-07,1.746623e-07,1.746633e-07,1.746643e-07,1.746654e-07,1.746664e-07,1.746674e-07,1.746684e-07,1.746694e-07,1.746705e-07,1.746715e-07,1.746725e-07,1.746735e-07,1.746745e-07,1.746756e-07,1.746766e-07,1.746776e-07,1.746786e-07,1.746797e-07,1.746807e-07,1.746817e-07,1.746827e-07,1.746837e-07,1.746848e-07,1.746858e-07,1.746868e-07,1.746878e-07,1.746888e-07,1.746899e-07,1.746909e-07,1.746919e-07,1.746929e-07,1.746939e-07,1.746950e-07,1.746960e-07,1.746970e-07,1.746980e-07,1.746990e-07,1.747001e-07,1.747011e-07,1.747021e-07,1.747031e-07,1.747041e-07,1.747051e-07,1.747062e-07,1.747072e-07,1.747082e-07,1.747092e-07,1.747102e-07,1.747113e-07,1.747123e-07,1.747133e-07,1.747143e-07,1.747153e-07,1.747163e-07,1.747174e-07,1.747184e-07,1.747194e-07,1.747204e-07,1.747214e-07,1.747224e-07,1.747235e-07,1.747245e-07,1.747255e-07,1.747265e-07,1.747275e-07,1.747285e-07,1.747296e-07,1.747306e-07,1.747316e-07,1.747326e-07,1.747336e-07,1.747346e-07,1.747357e-07,1.747367e-07,1.747377e-07,1.747387e-07,1.747397e-07,1.747407e-07,1.747418e-07,1.747428e-07,1.747438e-07,1.747448e-07,1.747458e-07,1.747468e-07,1.747478e-07,1.747489e-07,1.747499e-07,1.747509e-07,1.747519e-07,1.747529e-07,1.747539e-07,1.747549e-07,1.747560e-07,1.747570e-07,1.747580e-07,1.747590e-07,1.747600e-07,1.747610e-07,1.747620e-07,1.747631e-07,1.747641e-07,1.747651e-07,1.747661e-07,1.747671e-07,1.747681e-07,1.747691e-07,1.747701e-07,1.747712e-07,1.747722e-07,1.747732e-07,1.747742e-07,1.747752e-07,1.747762e-07,1.747772e-07,1.747782e-07,1.747793e-07,1.747803e-07,1.747813e-07,1.747823e-07,1.747833e-07,1.747843e-07,1.747853e-07,1.747863e-07,1.747874e-07,1.747884e-07,1.747894e-07,1.747904e-07,1.747914e-07,1.747924e-07,1.747934e-07,1.747944e-07,1.747954e-07,1.747965e-07,1.747975e-07,1.747985e-07,1.747995e-07,1.748005e-07,1.748015e-07,1.748025e-07,1.748035e-07,1.748045e-07,1.748055e-07,1.748066e-07,1.748076e-07,1.748086e-07,1.748096e-07,1.748106e-07,1.748116e-07,1.748126e-07,1.748136e-07,1.748146e-07,1.748156e-07,1.748166e-07,1.748177e-07,1.748187e-07,1.748197e-07,1.748207e-07,1.748217e-07,1.748227e-07,1.748237e-07,1.748247e-07,1.748257e-07,1.748267e-07,1.748277e-07,1.748287e-07,1.748298e-07,1.748308e-07,1.748318e-07,1.748328e-07,1.748338e-07,1.748348e-07,1.748358e-07,1.748368e-07,1.748378e-07,1.748388e-07,1.748398e-07,1.748408e-07,1.748418e-07,1.748428e-07,1.748439e-07,1.748449e-07,1.748459e-07,1.748469e-07,1.748479e-07,1.748489e-07,1.748499e-07,1.748509e-07,1.748519e-07,1.748529e-07,1.748539e-07,1.748549e-07,1.748559e-07,1.748569e-07,1.748579e-07,1.748589e-07,1.748599e-07,1.748609e-07,1.748620e-07,1.748630e-07,1.748640e-07,1.748650e-07,1.748660e-07,1.748670e-07,1.748680e-07,1.748690e-07,1.748700e-07,1.748710e-07,1.748720e-07,1.748730e-07,1.748740e-07,1.748750e-07,1.748760e-07,1.748770e-07,1.748780e-07,1.748790e-07,1.748800e-07,1.748810e-07,1.748820e-07,1.748830e-07,1.748840e-07,1.748850e-07,1.748860e-07,1.748870e-07,1.748880e-07,1.748891e-07,1.748901e-07,1.748911e-07,1.748921e-07,1.748931e-07,1.748941e-07,1.748951e-07,1.748961e-07,1.748971e-07,1.748981e-07,1.748991e-07,1.749001e-07,1.749011e-07,1.749021e-07,1.749031e-07,1.749041e-07,1.749051e-07,1.749061e-07,1.749071e-07,1.749081e-07,1.749091e-07,1.749101e-07,1.749111e-07,1.749121e-07,1.749131e-07,1.749141e-07,1.749151e-07,1.749161e-07,1.749171e-07,1.749181e-07,1.749191e-07,1.749201e-07,1.749211e-07,1.749221e-07,1.749231e-07,1.749241e-07,1.749251e-07,1.749261e-07,1.749271e-07,1.749281e-07,1.749291e-07,1.749301e-07,1.749311e-07,1.749321e-07,1.749331e-07,1.749341e-07,1.749351e-07,1.749361e-07,1.749371e-07,1.749381e-07,1.749391e-07,1.749401e-07,1.749411e-07,1.749421e-07,1.749431e-07,1.749441e-07,1.749451e-07,1.749461e-07,1.749471e-07,1.749481e-07,1.749490e-07,1.749500e-07,1.749510e-07,1.749520e-07,1.749530e-07,1.749540e-07,1.749550e-07,1.749560e-07,1.749570e-07,1.749580e-07,1.749590e-07,1.749600e-07,1.749610e-07,1.749620e-07,1.749630e-07,1.749640e-07,1.749650e-07,1.749660e-07,1.749670e-07,1.749680e-07,1.749690e-07,1.749700e-07,1.749710e-07,1.749720e-07,1.749730e-07,1.749740e-07,1.749750e-07,1.749759e-07,1.749769e-07,1.749779e-07,1.749789e-07,1.749799e-07,1.749809e-07,1.749819e-07,1.749829e-07,1.749839e-07,1.749849e-07,1.749859e-07,1.749869e-07,1.749879e-07,1.749889e-07,1.749899e-07,1.749909e-07,1.749919e-07,1.749929e-07,1.749938e-07,1.749948e-07,1.749958e-07,1.749968e-07,1.749978e-07,1.749988e-07,1.749998e-07,1.750008e-07,1.750018e-07,1.750028e-07,1.750038e-07,1.750048e-07,1.750058e-07,1.750068e-07,1.750077e-07,1.750087e-07,1.750097e-07,1.750107e-07,1.750117e-07,1.750127e-07,1.750137e-07,1.750147e-07,1.750157e-07,1.750167e-07,1.750177e-07,1.750187e-07,1.750196e-07,1.750206e-07,1.750216e-07,1.750226e-07,1.750236e-07,1.750246e-07,1.750256e-07,1.750266e-07,1.750276e-07,1.750286e-07,1.750296e-07,1.750305e-07,1.750315e-07,1.750325e-07,1.750335e-07,1.750345e-07,1.750355e-07,1.750365e-07,1.750375e-07,1.750385e-07,1.750395e-07,1.750404e-07,1.750414e-07,1.750424e-07,1.750434e-07,1.750444e-07,1.750454e-07,1.750464e-07,1.750474e-07,1.750484e-07,1.750494e-07,1.750503e-07,1.750513e-07,1.750523e-07,1.750533e-07,1.750543e-07,1.750553e-07,1.750563e-07,1.750573e-07,1.750582e-07,1.750592e-07,1.750602e-07,1.750612e-07,1.750622e-07,1.750632e-07,1.750642e-07,1.750652e-07,1.750662e-07,1.750671e-07,1.750681e-07,1.750691e-07,1.750701e-07,1.750711e-07,1.750721e-07,1.750731e-07,1.750740e-07,1.750750e-07,1.750760e-07,1.750770e-07,1.750780e-07,1.750790e-07,1.750800e-07,1.750810e-07,1.750819e-07,1.750829e-07,1.750839e-07,1.750849e-07,1.750859e-07,1.750869e-07,1.750879e-07,1.750888e-07,1.750898e-07,1.750908e-07,1.750918e-07,1.750928e-07,1.750938e-07,1.750947e-07,1.750957e-07,1.750967e-07,1.750977e-07,1.750987e-07,1.750997e-07,1.751007e-07,1.751016e-07,1.751026e-07,1.751036e-07,1.751046e-07,1.751056e-07,1.751066e-07,1.751075e-07,1.751085e-07,1.751095e-07,1.751105e-07,1.751115e-07,1.751125e-07,1.751134e-07,1.751144e-07,1.751154e-07,1.751164e-07,1.751174e-07,1.751184e-07,1.751193e-07,1.751203e-07,1.751213e-07,1.751223e-07,1.751233e-07,1.751243e-07,1.751252e-07,1.751262e-07,1.751272e-07,1.751282e-07,1.751292e-07,1.751302e-07,1.751311e-07,1.751321e-07,1.751331e-07,1.751341e-07,1.751351e-07,1.751360e-07,1.751370e-07,1.751380e-07,1.751390e-07,1.751400e-07,1.751410e-07,1.751419e-07,1.751429e-07,1.751439e-07,1.751449e-07,1.751459e-07,1.751468e-07,1.751478e-07,1.751488e-07,1.751498e-07,1.751508e-07,1.751517e-07,1.751527e-07,1.751537e-07,1.751547e-07,1.751557e-07,1.751566e-07,1.751576e-07,1.751586e-07,1.751596e-07,1.751606e-07,1.751615e-07,1.751625e-07,1.751635e-07,1.751645e-07,1.751655e-07,1.751664e-07,1.751674e-07,1.751684e-07,1.751694e-07,1.751703e-07,1.751713e-07,1.751723e-07,1.751733e-07,1.751743e-07,1.751752e-07,1.751762e-07,1.751772e-07,1.751782e-07,1.751792e-07,1.751801e-07,1.751811e-07,1.751821e-07,1.751831e-07,1.751840e-07,1.751850e-07,1.751860e-07,1.751870e-07,1.751879e-07,1.751889e-07,1.751899e-07,1.751909e-07,1.751919e-07,1.751928e-07,1.751938e-07,1.751948e-07,1.751958e-07,1.751967e-07,1.751977e-07,1.751987e-07,1.751997e-07,1.752006e-07,1.752016e-07,1.752026e-07,1.752036e-07,1.752045e-07,1.752055e-07,1.752065e-07,1.752075e-07,1.752084e-07,1.752094e-07,1.752104e-07,1.752114e-07,1.752124e-07,1.752133e-07,1.752143e-07,1.752153e-07,1.752163e-07,1.752172e-07,1.752182e-07,1.752192e-07,1.752201e-07,1.752211e-07,1.752221e-07,1.752231e-07,1.752240e-07,1.752250e-07,1.752260e-07,1.752270e-07,1.752279e-07,1.752289e-07,1.752299e-07,1.752309e-07,1.752318e-07,1.752328e-07,1.752338e-07,1.752348e-07,1.752357e-07,1.752367e-07,1.752377e-07,1.752386e-07,1.752396e-07,1.752406e-07,1.752416e-07,1.752425e-07,1.752435e-07,1.752445e-07,1.752455e-07,1.752464e-07,1.752474e-07,1.752484e-07,1.752493e-07,1.752503e-07,1.752513e-07,1.752523e-07,1.752532e-07,1.752542e-07,1.752552e-07,1.752561e-07,1.752571e-07,1.752581e-07,1.752591e-07,1.752600e-07,1.752610e-07,1.752620e-07,1.752629e-07,1.752639e-07,1.752649e-07,1.752659e-07,1.752668e-07,1.752678e-07,1.752688e-07,1.752697e-07,1.752707e-07,1.752717e-07,1.752726e-07,1.752736e-07,1.752746e-07,1.752756e-07,1.752765e-07,1.752775e-07,1.752785e-07,1.752794e-07,1.752804e-07,1.752814e-07,1.752823e-07,1.752833e-07,1.752843e-07,1.752853e-07,1.752862e-07,1.752872e-07,1.752882e-07,1.752891e-07,1.752901e-07,1.752911e-07,1.752920e-07,1.752930e-07,1.752940e-07,1.752949e-07,1.752959e-07,1.752969e-07,1.752978e-07,1.752988e-07,1.752998e-07,1.753007e-07,1.753017e-07,1.753027e-07,1.753036e-07,1.753046e-07,1.753056e-07,1.753066e-07,1.753075e-07,1.753085e-07,1.753095e-07,1.753104e-07,1.753114e-07,1.753124e-07,1.753133e-07,1.753143e-07,1.753153e-07,1.753162e-07,1.753172e-07,1.753182e-07,1.753191e-07,1.753201e-07,1.753210e-07,1.753220e-07,1.753230e-07,1.753239e-07,1.753249e-07,1.753259e-07,1.753268e-07,1.753278e-07,1.753288e-07,1.753297e-07,1.753307e-07,1.753317e-07,1.753326e-07,1.753336e-07,1.753346e-07,1.753355e-07,1.753365e-07,1.753375e-07,1.753384e-07,1.753394e-07,1.753404e-07,1.753413e-07,1.753423e-07,1.753432e-07,1.753442e-07,1.753452e-07,1.753461e-07,1.753471e-07,1.753481e-07,1.753490e-07,1.753500e-07,1.753510e-07,1.753519e-07,1.753529e-07,1.753538e-07,1.753548e-07,1.753558e-07,1.753567e-07,1.753577e-07,1.753587e-07,1.753596e-07,1.753606e-07,1.753616e-07,1.753625e-07,1.753635e-07,1.753644e-07,1.753654e-07,1.753664e-07,1.753673e-07,1.753683e-07,1.753693e-07,1.753702e-07,1.753712e-07,1.753721e-07,1.753731e-07,1.753741e-07,1.753750e-07,1.753760e-07,1.753769e-07,1.753779e-07,1.753789e-07,1.753798e-07,1.753808e-07,1.753817e-07,1.753827e-07,1.753837e-07,1.753846e-07,1.753856e-07,1.753866e-07,1.753875e-07,1.753885e-07,1.753894e-07,1.753904e-07,1.753914e-07,1.753923e-07,1.753933e-07,1.753942e-07,1.753952e-07,1.753962e-07,1.753971e-07,1.753981e-07,1.753990e-07,1.754000e-07,1.754010e-07,1.754019e-07,1.754029e-07,1.754038e-07,1.754048e-07,1.754057e-07,1.754067e-07,1.754077e-07,1.754086e-07,1.754096e-07,1.754105e-07,1.754115e-07,1.754125e-07,1.754134e-07,1.754144e-07,1.754153e-07,1.754163e-07,1.754173e-07,1.754182e-07,1.754192e-07,1.754201e-07,1.754211e-07,1.754220e-07,1.754230e-07,1.754240e-07,1.754249e-07,1.754259e-07,1.754268e-07,1.754278e-07,1.754287e-07,1.754297e-07,1.754307e-07,1.754316e-07,1.754326e-07,1.754335e-07,1.754345e-07,1.754354e-07,1.754364e-07,1.754374e-07,1.754383e-07,1.754393e-07,1.754402e-07,1.754412e-07,1.754421e-07,1.754431e-07,1.754440e-07,1.754450e-07,1.754460e-07,1.754469e-07,1.754479e-07,1.754488e-07,1.754498e-07,1.754507e-07,1.754517e-07,1.754526e-07,1.754536e-07,1.754546e-07,1.754555e-07,1.754565e-07,1.754574e-07,1.754584e-07,1.754593e-07,1.754603e-07,1.754612e-07,1.754622e-07,1.754631e-07,1.754641e-07,1.754651e-07,1.754660e-07,1.754670e-07,1.754679e-07,1.754689e-07,1.754698e-07,1.754708e-07,1.754717e-07,1.754727e-07,1.754736e-07,1.754746e-07,1.754755e-07,1.754765e-07,1.754775e-07,1.754784e-07,1.754794e-07,1.754803e-07,1.754813e-07,1.754822e-07,1.754832e-07,1.754841e-07,1.754851e-07,1.754860e-07,1.754870e-07,1.754879e-07,1.754889e-07,1.754898e-07,1.754908e-07,1.754917e-07,1.754927e-07,1.754936e-07,1.754946e-07,1.754955e-07,1.754965e-07,1.754975e-07,1.754984e-07,1.754994e-07,1.755003e-07,1.755013e-07,1.755022e-07,1.755032e-07,1.755041e-07,1.755051e-07,1.755060e-07,1.755070e-07,1.755079e-07,1.755089e-07,1.755098e-07,1.755108e-07,1.755117e-07,1.755127e-07,1.755136e-07,1.755146e-07,1.755155e-07,1.755165e-07,1.755174e-07,1.755184e-07,1.755193e-07,1.755203e-07,1.755212e-07,1.755222e-07,1.755231e-07,1.755241e-07,1.755250e-07,1.755260e-07,1.755269e-07,1.755279e-07,1.755288e-07,1.755298e-07,1.755307e-07,1.755317e-07,1.755326e-07,1.755336e-07,1.755345e-07,1.755354e-07,1.755364e-07,1.755373e-07,1.755383e-07,1.755392e-07,1.755402e-07,1.755411e-07,1.755421e-07,1.755430e-07,1.755440e-07,1.755449e-07,1.755459e-07,1.755468e-07,1.755478e-07,1.755487e-07,1.755497e-07,1.755506e-07,1.755516e-07,1.755525e-07,1.755535e-07,1.755544e-07,1.755553e-07,1.755563e-07,1.755572e-07,1.755582e-07,1.755591e-07,1.755601e-07,1.755610e-07,1.755620e-07,1.755629e-07,1.755639e-07,1.755648e-07,1.755658e-07,1.755667e-07,1.755676e-07,1.755686e-07,1.755695e-07,1.755705e-07,1.755714e-07,1.755724e-07,1.755733e-07,1.755743e-07,1.755752e-07,1.755762e-07,1.755771e-07,1.755780e-07,1.755790e-07,1.755799e-07,1.755809e-07,1.755818e-07,1.755828e-07,1.755837e-07,1.755847e-07,1.755856e-07,1.755865e-07,1.755875e-07,1.755884e-07,1.755894e-07,1.755903e-07,1.755913e-07,1.755922e-07,1.755932e-07,1.755941e-07,1.755950e-07,1.755960e-07,1.755969e-07,1.755979e-07,1.755988e-07,1.755998e-07,1.756007e-07,1.756016e-07,1.756026e-07,1.756035e-07,1.756045e-07,1.756054e-07,1.756064e-07,1.756073e-07,1.756082e-07,1.756092e-07,1.756101e-07,1.756111e-07,1.756120e-07,1.756130e-07,1.756139e-07,1.756148e-07,1.756158e-07,1.756167e-07,1.756177e-07,1.756186e-07,1.756196e-07,1.756205e-07,1.756214e-07,1.756224e-07,1.756233e-07,1.756243e-07,1.756252e-07,1.756261e-07,1.756271e-07,1.756280e-07,1.756290e-07,1.756299e-07,1.756308e-07,1.756318e-07,1.756327e-07,1.756337e-07,1.756346e-07,1.756355e-07,1.756365e-07,1.756374e-07,1.756384e-07,1.756393e-07,1.756402e-07,1.756412e-07,1.756421e-07,1.756431e-07,1.756440e-07,1.756449e-07,1.756459e-07,1.756468e-07,1.756478e-07,1.756487e-07,1.756496e-07,1.756506e-07,1.756515e-07,1.756525e-07,1.756534e-07,1.756543e-07,1.756553e-07,1.756562e-07,1.756572e-07,1.756581e-07,1.756590e-07,1.756600e-07,1.756609e-07,1.756618e-07,1.756628e-07,1.756637e-07,1.756647e-07,1.756656e-07,1.756665e-07,1.756675e-07,1.756684e-07,1.756693e-07,1.756703e-07,1.756712e-07,1.756722e-07,1.756731e-07,1.756740e-07,1.756750e-07,1.756759e-07,1.756768e-07,1.756778e-07,1.756787e-07,1.756797e-07,1.756806e-07,1.756815e-07,1.756825e-07,1.756834e-07,1.756843e-07,1.756853e-07,1.756862e-07,1.756871e-07,1.756881e-07,1.756890e-07,1.756900e-07,1.756909e-07,1.756918e-07,1.756928e-07,1.756937e-07,1.756946e-07,1.756956e-07,1.756965e-07,1.756974e-07,1.756984e-07,1.756993e-07,1.757002e-07,1.757012e-07,1.757021e-07,1.757030e-07,1.757040e-07,1.757049e-07,1.757059e-07,1.757068e-07,1.757077e-07,1.757087e-07,1.757096e-07,1.757105e-07,1.757115e-07,1.757124e-07,1.757133e-07,1.757143e-07,1.757152e-07,1.757161e-07,1.757171e-07,1.757180e-07,1.757189e-07,1.757199e-07,1.757208e-07,1.757217e-07,1.757227e-07,1.757236e-07,1.757245e-07,1.757255e-07,1.757264e-07,1.757273e-07,1.757283e-07,1.757292e-07,1.757301e-07,1.757311e-07,1.757320e-07,1.757329e-07,1.757339e-07,1.757348e-07,1.757357e-07,1.757367e-07,1.757376e-07,1.757385e-07,1.757394e-07,1.757404e-07,1.757413e-07,1.757422e-07,1.757432e-07,1.757441e-07,1.757450e-07,1.757460e-07,1.757469e-07,1.757478e-07,1.757488e-07,1.757497e-07,1.757506e-07,1.757516e-07,1.757525e-07,1.757534e-07,1.757543e-07,1.757553e-07,1.757562e-07,1.757571e-07,1.757581e-07,1.757590e-07,1.757599e-07,1.757609e-07,1.757618e-07,1.757627e-07,1.757637e-07,1.757646e-07,1.757655e-07,1.757664e-07,1.757674e-07,1.757683e-07,1.757692e-07,1.757702e-07,1.757711e-07,1.757720e-07,1.757729e-07,1.757739e-07,1.757748e-07,1.757757e-07,1.757767e-07,1.757776e-07,1.757785e-07,1.757795e-07,1.757804e-07,1.757813e-07,1.757822e-07,1.757832e-07,1.757841e-07,1.757850e-07,1.757860e-07,1.757869e-07,1.757878e-07,1.757887e-07,1.757897e-07,1.757906e-07,1.757915e-07,1.757924e-07,1.757934e-07,1.757943e-07,1.757952e-07,1.757962e-07,1.757971e-07,1.757980e-07,1.757989e-07,1.757999e-07,1.758008e-07,1.758017e-07,1.758026e-07,1.758036e-07,1.758045e-07,1.758054e-07,1.758064e-07,1.758073e-07,1.758082e-07,1.758091e-07,1.758101e-07,1.758110e-07,1.758119e-07,1.758128e-07,1.758138e-07,1.758147e-07,1.758156e-07,1.758165e-07,1.758175e-07,1.758184e-07,1.758193e-07,1.758202e-07,1.758212e-07,1.758221e-07,1.758230e-07,1.758239e-07,1.758249e-07,1.758258e-07,1.758267e-07,1.758276e-07,1.758286e-07,1.758295e-07,1.758304e-07,1.758313e-07,1.758323e-07,1.758332e-07,1.758341e-07,1.758350e-07,1.758360e-07,1.758369e-07,1.758378e-07,1.758387e-07,1.758397e-07,1.758406e-07,1.758415e-07,1.758424e-07,1.758434e-07,1.758443e-07,1.758452e-07,1.758461e-07,1.758471e-07,1.758480e-07,1.758489e-07,1.758498e-07,1.758507e-07,1.758517e-07,1.758526e-07,1.758535e-07,1.758544e-07,1.758554e-07,1.758563e-07,1.758572e-07,1.758581e-07,1.758590e-07,1.758600e-07,1.758609e-07,1.758618e-07,1.758627e-07,1.758637e-07,1.758646e-07,1.758655e-07,1.758664e-07,1.758673e-07,1.758683e-07,1.758692e-07,1.758701e-07,1.758710e-07,1.758720e-07,1.758729e-07,1.758738e-07,1.758747e-07,1.758756e-07,1.758766e-07,1.758775e-07,1.758784e-07,1.758793e-07,1.758802e-07,1.758812e-07,1.758821e-07,1.758830e-07,1.758839e-07,1.758848e-07,1.758858e-07,1.758867e-07,1.758876e-07,1.758885e-07,1.758894e-07,1.758904e-07,1.758913e-07,1.758922e-07,1.758931e-07,1.758940e-07,1.758950e-07,1.758959e-07,1.758968e-07,1.758977e-07,1.758986e-07,1.758996e-07,1.759005e-07,1.759014e-07,1.759023e-07,1.759032e-07,1.759042e-07,1.759051e-07,1.759060e-07,1.759069e-07,1.759078e-07,1.759088e-07,1.759097e-07,1.759106e-07,1.759115e-07,1.759124e-07,1.759133e-07,1.759143e-07,1.759152e-07,1.759161e-07,1.759170e-07,1.759179e-07,1.759188e-07,1.759198e-07,1.759207e-07,1.759216e-07,1.759225e-07,1.759234e-07,1.759244e-07,1.759253e-07,1.759262e-07,1.759271e-07,1.759280e-07,1.759289e-07,1.759299e-07,1.759308e-07,1.759317e-07,1.759326e-07,1.759335e-07,1.759344e-07,1.759354e-07,1.759363e-07,1.759372e-07,1.759381e-07,1.759390e-07,1.759399e-07,1.759409e-07,1.759418e-07,1.759427e-07,1.759436e-07,1.759445e-07,1.759454e-07,1.759463e-07,1.759473e-07,1.759482e-07,1.759491e-07,1.759500e-07,1.759509e-07,1.759518e-07,1.759528e-07,1.759537e-07,1.759546e-07,1.759555e-07,1.759564e-07,1.759573e-07,1.759582e-07,1.759592e-07,1.759601e-07,1.759610e-07,1.759619e-07,1.759628e-07,1.759637e-07,1.759646e-07,1.759656e-07,1.759665e-07,1.759674e-07,1.759683e-07,1.759692e-07,1.759701e-07,1.759710e-07,1.759720e-07,1.759729e-07,1.759738e-07,1.759747e-07,1.759756e-07,1.759765e-07,1.759774e-07,1.759783e-07,1.759793e-07,1.759802e-07,1.759811e-07,1.759820e-07,1.759829e-07,1.759838e-07,1.759847e-07,1.759856e-07,1.759866e-07,1.759875e-07,1.759884e-07,1.759893e-07,1.759902e-07,1.759911e-07,1.759920e-07,1.759929e-07,1.759939e-07,1.759948e-07,1.759957e-07,1.759966e-07,1.759975e-07,1.759984e-07,1.759993e-07,1.760002e-07,1.760011e-07,1.760021e-07,1.760030e-07,1.760039e-07,1.760048e-07,1.760057e-07,1.760066e-07,1.760075e-07,1.760084e-07,1.760093e-07,1.760103e-07,1.760112e-07,1.760121e-07,1.760130e-07,1.760139e-07,1.760148e-07,1.760157e-07,1.760166e-07,1.760175e-07,1.760184e-07,1.760194e-07,1.760203e-07,1.760212e-07,1.760221e-07,1.760230e-07,1.760239e-07,1.760248e-07,1.760257e-07,1.760266e-07,1.760275e-07,1.760284e-07,1.760294e-07,1.760303e-07,1.760312e-07,1.760321e-07,1.760330e-07,1.760339e-07,1.760348e-07,1.760357e-07,1.760366e-07,1.760375e-07,1.760384e-07,1.760394e-07,1.760403e-07,1.760412e-07,1.760421e-07,1.760430e-07,1.760439e-07,1.760448e-07,1.760457e-07,1.760466e-07,1.760475e-07,1.760484e-07,1.760493e-07,1.760502e-07,1.760512e-07,1.760521e-07,1.760530e-07,1.760539e-07,1.760548e-07,1.760557e-07,1.760566e-07,1.760575e-07,1.760584e-07,1.760593e-07,1.760602e-07,1.760611e-07,1.760620e-07,1.760629e-07,1.760638e-07,1.760648e-07,1.760657e-07,1.760666e-07,1.760675e-07,1.760684e-07,1.760693e-07,1.760702e-07,1.760711e-07,1.760720e-07,1.760729e-07,1.760738e-07,1.760747e-07,1.760756e-07,1.760765e-07,1.760774e-07,1.760783e-07,1.760792e-07,1.760802e-07,1.760811e-07,1.760820e-07,1.760829e-07,1.760838e-07,1.760847e-07,1.760856e-07,1.760865e-07,1.760874e-07,1.760883e-07,1.760892e-07,1.760901e-07,1.760910e-07,1.760919e-07,1.760928e-07,1.760937e-07,1.760946e-07,1.760955e-07,1.760964e-07,1.760973e-07,1.760982e-07,1.760991e-07,1.761000e-07,1.761009e-07,1.761019e-07,1.761028e-07,1.761037e-07,1.761046e-07,1.761055e-07,1.761064e-07,1.761073e-07,1.761082e-07,1.761091e-07,1.761100e-07,1.761109e-07,1.761118e-07,1.761127e-07,1.761136e-07,1.761145e-07,1.761154e-07,1.761163e-07,1.761172e-07,1.761181e-07,1.761190e-07,1.761199e-07,1.761208e-07,1.761217e-07,1.761226e-07,1.761235e-07,1.761244e-07,1.761253e-07,1.761262e-07,1.761271e-07,1.761280e-07,1.761289e-07,1.761298e-07,1.761307e-07,1.761316e-07,1.761325e-07,1.761334e-07,1.761343e-07,1.761352e-07,1.761361e-07,1.761370e-07,1.761379e-07,1.761388e-07,1.761397e-07,1.761406e-07,1.761415e-07,1.761424e-07,1.761433e-07,1.761442e-07,1.761451e-07,1.761460e-07,1.761469e-07,1.761478e-07,1.761487e-07,1.761496e-07,1.761505e-07,1.761514e-07,1.761523e-07,1.761532e-07,1.761541e-07,1.761550e-07,1.761559e-07,1.761568e-07,1.761577e-07,1.761586e-07,1.761595e-07,1.761604e-07,1.761613e-07,1.761622e-07,1.761631e-07,1.761640e-07,1.761649e-07,1.761658e-07,1.761667e-07,1.761676e-07,1.761685e-07,1.761694e-07,1.761703e-07,1.761712e-07,1.761721e-07,1.761730e-07,1.761739e-07,1.761748e-07,1.761757e-07,1.761766e-07,1.761775e-07,1.761784e-07,1.761793e-07,1.761802e-07,1.761811e-07,1.761820e-07,1.761829e-07,1.761838e-07,1.761847e-07,1.761856e-07,1.761865e-07,1.761874e-07,1.761882e-07,1.761891e-07,1.761900e-07,1.761909e-07,1.761918e-07,1.761927e-07,1.761936e-07,1.761945e-07,1.761954e-07,1.761963e-07,1.761972e-07,1.761981e-07,1.761990e-07,1.761999e-07,1.762008e-07,1.762017e-07,1.762026e-07,1.762035e-07,1.762044e-07,1.762053e-07,1.762062e-07,1.762071e-07,1.762080e-07,1.762089e-07,1.762097e-07,1.762106e-07,1.762115e-07,1.762124e-07,1.762133e-07,1.762142e-07,1.762151e-07,1.762160e-07,1.762169e-07,1.762178e-07,1.762187e-07,1.762196e-07,1.762205e-07,1.762214e-07,1.762223e-07,1.762232e-07,1.762241e-07,1.762250e-07,1.762258e-07,1.762267e-07,1.762276e-07,1.762285e-07,1.762294e-07,1.762303e-07,1.762312e-07,1.762321e-07,1.762330e-07,1.762339e-07,1.762348e-07,1.762357e-07,1.762366e-07,1.762375e-07,1.762384e-07,1.762392e-07,1.762401e-07,1.762410e-07,1.762419e-07,1.762428e-07,1.762437e-07,1.762446e-07,1.762455e-07,1.762464e-07,1.762473e-07,1.762482e-07,1.762491e-07,1.762500e-07,1.762508e-07,1.762517e-07,1.762526e-07,1.762535e-07,1.762544e-07,1.762553e-07,1.762562e-07,1.762571e-07,1.762580e-07,1.762589e-07,1.762598e-07,1.762607e-07,1.762615e-07,1.762624e-07,1.762633e-07,1.762642e-07,1.762651e-07,1.762660e-07,1.762669e-07,1.762678e-07,1.762687e-07,1.762696e-07,1.762705e-07,1.762713e-07,1.762722e-07,1.762731e-07,1.762740e-07,1.762749e-07,1.762758e-07,1.762767e-07,1.762776e-07,1.762785e-07,1.762794e-07,1.762802e-07,1.762811e-07,1.762820e-07,1.762829e-07,1.762838e-07,1.762847e-07,1.762856e-07,1.762865e-07,1.762874e-07,1.762882e-07,1.762891e-07,1.762900e-07,1.762909e-07,1.762918e-07,1.762927e-07,1.762936e-07,1.762945e-07,1.762954e-07,1.762962e-07,1.762971e-07,1.762980e-07,1.762989e-07,1.762998e-07,1.763007e-07,1.763016e-07,1.763025e-07,1.763033e-07,1.763042e-07,1.763051e-07,1.763060e-07,1.763069e-07,1.763078e-07,1.763087e-07,1.763096e-07,1.763104e-07,1.763113e-07,1.763122e-07,1.763131e-07,1.763140e-07,1.763149e-07,1.763158e-07,1.763167e-07,1.763175e-07,1.763184e-07,1.763193e-07,1.763202e-07,1.763211e-07,1.763220e-07,1.763229e-07,1.763238e-07,1.763246e-07,1.763255e-07,1.763264e-07,1.763273e-07,1.763282e-07,1.763291e-07,1.763300e-07,1.763308e-07,1.763317e-07,1.763326e-07,1.763335e-07,1.763344e-07,1.763353e-07,1.763362e-07,1.763370e-07,1.763379e-07,1.763388e-07,1.763397e-07,1.763406e-07,1.763415e-07,1.763423e-07,1.763432e-07,1.763441e-07,1.763450e-07,1.763459e-07,1.763468e-07,1.763477e-07,1.763485e-07,1.763494e-07,1.763503e-07,1.763512e-07,1.763521e-07,1.763530e-07,1.763538e-07,1.763547e-07,1.763556e-07,1.763565e-07,1.763574e-07,1.763583e-07,1.763591e-07,1.763600e-07,1.763609e-07,1.763618e-07,1.763627e-07,1.763636e-07,1.763644e-07,1.763653e-07,1.763662e-07,1.763671e-07,1.763680e-07,1.763689e-07,1.763697e-07,1.763706e-07,1.763715e-07,1.763724e-07,1.763733e-07,1.763742e-07,1.763750e-07,1.763759e-07,1.763768e-07,1.763777e-07,1.763786e-07,1.763795e-07,1.763803e-07,1.763812e-07,1.763821e-07,1.763830e-07,1.763839e-07,1.763847e-07,1.763856e-07,1.763865e-07,1.763874e-07,1.763883e-07,1.763892e-07,1.763900e-07,1.763909e-07,1.763918e-07,1.763927e-07,1.763936e-07,1.763944e-07,1.763953e-07,1.763962e-07,1.763971e-07,1.763980e-07,1.763988e-07,1.763997e-07,1.764006e-07,1.764015e-07,1.764024e-07,1.764032e-07,1.764041e-07,1.764050e-07,1.764059e-07,1.764068e-07,1.764076e-07,1.764085e-07,1.764094e-07,1.764103e-07,1.764112e-07,1.764120e-07,1.764129e-07,1.764138e-07,1.764147e-07,1.764156e-07,1.764164e-07,1.764173e-07,1.764182e-07,1.764191e-07,1.764200e-07,1.764208e-07,1.764217e-07,1.764226e-07,1.764235e-07,1.764244e-07,1.764252e-07,1.764261e-07,1.764270e-07,1.764279e-07,1.764287e-07,1.764296e-07,1.764305e-07,1.764314e-07,1.764323e-07,1.764331e-07,1.764340e-07,1.764349e-07,1.764358e-07,1.764366e-07,1.764375e-07,1.764384e-07,1.764393e-07,1.764402e-07,1.764410e-07,1.764419e-07,1.764428e-07,1.764437e-07,1.764445e-07,1.764454e-07,1.764463e-07,1.764472e-07,1.764481e-07,1.764489e-07,1.764498e-07,1.764507e-07,1.764516e-07,1.764524e-07,1.764533e-07,1.764542e-07,1.764551e-07,1.764559e-07,1.764568e-07,1.764577e-07,1.764586e-07,1.764594e-07,1.764603e-07,1.764612e-07,1.764621e-07,1.764629e-07,1.764638e-07,1.764647e-07,1.764656e-07,1.764665e-07,1.764673e-07,1.764682e-07,1.764691e-07,1.764700e-07,1.764708e-07,1.764717e-07,1.764726e-07,1.764735e-07,1.764743e-07,1.764752e-07,1.764761e-07,1.764770e-07,1.764778e-07,1.764787e-07,1.764796e-07,1.764805e-07,1.764813e-07,1.764822e-07,1.764831e-07,1.764839e-07,1.764848e-07,1.764857e-07,1.764866e-07,1.764874e-07,1.764883e-07,1.764892e-07,1.764901e-07,1.764909e-07,1.764918e-07,1.764927e-07,1.764936e-07,1.764944e-07,1.764953e-07,1.764962e-07,1.764971e-07,1.764979e-07,1.764988e-07,1.764997e-07,1.765005e-07,1.765014e-07,1.765023e-07,1.765032e-07,1.765040e-07,1.765049e-07,1.765058e-07,1.765067e-07,1.765075e-07,1.765084e-07,1.765093e-07,1.765101e-07,1.765110e-07,1.765119e-07,1.765128e-07,1.765136e-07,1.765145e-07,1.765154e-07,1.765162e-07,1.765171e-07,1.765180e-07,1.765189e-07,1.765197e-07,1.765206e-07,1.765215e-07,1.765223e-07,1.765232e-07,1.765241e-07,1.765250e-07,1.765258e-07,1.765267e-07,1.765276e-07,1.765284e-07,1.765293e-07,1.765302e-07,1.765311e-07,1.765319e-07,1.765328e-07,1.765337e-07,1.765345e-07,1.765354e-07,1.765363e-07,1.765372e-07,1.765380e-07,1.765389e-07,1.765398e-07,1.765406e-07,1.765415e-07,1.765424e-07,1.765432e-07,1.765441e-07,1.765450e-07,1.765458e-07,1.765467e-07,1.765476e-07,1.765485e-07,1.765493e-07,1.765502e-07,1.765511e-07,1.765519e-07,1.765528e-07,1.765537e-07,1.765545e-07,1.765554e-07,1.765563e-07,1.765571e-07,1.765580e-07,1.765589e-07,1.765598e-07,1.765606e-07,1.765615e-07,1.765624e-07,1.765632e-07,1.765641e-07,1.765650e-07,1.765658e-07,1.765667e-07,1.765676e-07,1.765684e-07,1.765693e-07,1.765702e-07,1.765710e-07,1.765719e-07,1.765728e-07,1.765736e-07,1.765745e-07,1.765754e-07,1.765762e-07,1.765771e-07,1.765780e-07,1.765788e-07,1.765797e-07,1.765806e-07,1.765814e-07,1.765823e-07,1.765832e-07,1.765840e-07,1.765849e-07,1.765858e-07,1.765866e-07,1.765875e-07,1.765884e-07,1.765892e-07,1.765901e-07,1.765910e-07,1.765918e-07,1.765927e-07,1.765936e-07,1.765944e-07,1.765953e-07,1.765962e-07,1.765970e-07,1.765979e-07,1.765988e-07,1.765996e-07,1.766005e-07,1.766014e-07,1.766022e-07,1.766031e-07,1.766040e-07,1.766048e-07,1.766057e-07,1.766066e-07,1.766074e-07,1.766083e-07,1.766092e-07,1.766100e-07,1.766109e-07,1.766117e-07,1.766126e-07,1.766135e-07,1.766143e-07,1.766152e-07,1.766161e-07,1.766169e-07,1.766178e-07,1.766187e-07,1.766195e-07,1.766204e-07,1.766213e-07,1.766221e-07,1.766230e-07,1.766238e-07,1.766247e-07,1.766256e-07,1.766264e-07,1.766273e-07,1.766282e-07,1.766290e-07,1.766299e-07,1.766308e-07,1.766316e-07,1.766325e-07,1.766333e-07,1.766342e-07,1.766351e-07,1.766359e-07,1.766368e-07,1.766377e-07,1.766385e-07,1.766394e-07,1.766402e-07,1.766411e-07,1.766420e-07,1.766428e-07,1.766437e-07,1.766446e-07,1.766454e-07,1.766463e-07,1.766471e-07,1.766480e-07,1.766489e-07,1.766497e-07,1.766506e-07,1.766515e-07,1.766523e-07,1.766532e-07,1.766540e-07,1.766549e-07,1.766558e-07,1.766566e-07,1.766575e-07,1.766583e-07,1.766592e-07,1.766601e-07,1.766609e-07,1.766618e-07,1.766626e-07,1.766635e-07,1.766644e-07,1.766652e-07,1.766661e-07,1.766670e-07,1.766678e-07,1.766687e-07,1.766695e-07,1.766704e-07,1.766713e-07,1.766721e-07,1.766730e-07,1.766738e-07,1.766747e-07,1.766756e-07,1.766764e-07,1.766773e-07,1.766781e-07,1.766790e-07,1.766799e-07,1.766807e-07,1.766816e-07,1.766824e-07,1.766833e-07,1.766842e-07,1.766850e-07,1.766859e-07,1.766867e-07,1.766876e-07,1.766884e-07,1.766893e-07,1.766902e-07,1.766910e-07,1.766919e-07,1.766927e-07,1.766936e-07,1.766945e-07,1.766953e-07,1.766962e-07,1.766970e-07,1.766979e-07,1.766987e-07,1.766996e-07,1.767005e-07,1.767013e-07,1.767022e-07,1.767030e-07,1.767039e-07,1.767048e-07,1.767056e-07,1.767065e-07,1.767073e-07,1.767082e-07,1.767090e-07,1.767099e-07,1.767108e-07,1.767116e-07,1.767125e-07,1.767133e-07,1.767142e-07,1.767150e-07,1.767159e-07,1.767168e-07,1.767176e-07,1.767185e-07,1.767193e-07,1.767202e-07,1.767210e-07,1.767219e-07,1.767228e-07,1.767236e-07,1.767245e-07,1.767253e-07,1.767262e-07,1.767270e-07,1.767279e-07,1.767287e-07,1.767296e-07,1.767305e-07,1.767313e-07,1.767322e-07,1.767330e-07,1.767339e-07,1.767347e-07,1.767356e-07,1.767364e-07,1.767373e-07,1.767382e-07,1.767390e-07,1.767399e-07,1.767407e-07,1.767416e-07,1.767424e-07,1.767433e-07,1.767441e-07,1.767450e-07,1.767459e-07,1.767467e-07,1.767476e-07,1.767484e-07,1.767493e-07,1.767501e-07,1.767510e-07,1.767518e-07,1.767527e-07,1.767535e-07,1.767544e-07,1.767553e-07,1.767561e-07,1.767570e-07,1.767578e-07,1.767587e-07,1.767595e-07,1.767604e-07,1.767612e-07,1.767621e-07,1.767629e-07,1.767638e-07,1.767646e-07,1.767655e-07,1.767663e-07,1.767672e-07,1.767681e-07,1.767689e-07,1.767698e-07,1.767706e-07,1.767715e-07,1.767723e-07,1.767732e-07,1.767740e-07,1.767749e-07,1.767757e-07,1.767766e-07,1.767774e-07,1.767783e-07,1.767791e-07,1.767800e-07,1.767808e-07,1.767817e-07,1.767825e-07,1.767834e-07,1.767843e-07,1.767851e-07,1.767860e-07,1.767868e-07,1.767877e-07,1.767885e-07,1.767894e-07,1.767902e-07,1.767911e-07,1.767919e-07,1.767928e-07,1.767936e-07,1.767945e-07,1.767953e-07,1.767962e-07,1.767970e-07,1.767979e-07,1.767987e-07,1.767996e-07,1.768004e-07,1.768013e-07,1.768021e-07,1.768030e-07,1.768038e-07,1.768047e-07,1.768055e-07,1.768064e-07,1.768072e-07,1.768081e-07,1.768089e-07,1.768098e-07,1.768106e-07,1.768115e-07,1.768123e-07,1.768132e-07,1.768140e-07,1.768149e-07,1.768157e-07,1.768166e-07,1.768174e-07,1.768183e-07,1.768191e-07,1.768200e-07,1.768208e-07,1.768217e-07,1.768225e-07,1.768234e-07,1.768242e-07,1.768251e-07,1.768259e-07,1.768268e-07,1.768276e-07,1.768285e-07,1.768293e-07,1.768302e-07,1.768310e-07,1.768319e-07,1.768327e-07,1.768336e-07,1.768344e-07,1.768353e-07,1.768361e-07,1.768370e-07,1.768378e-07,1.768386e-07,1.768395e-07,1.768403e-07,1.768412e-07,1.768420e-07,1.768429e-07,1.768437e-07,1.768446e-07,1.768454e-07,1.768463e-07,1.768471e-07,1.768480e-07,1.768488e-07,1.768497e-07,1.768505e-07,1.768514e-07,1.768522e-07,1.768531e-07,1.768539e-07,1.768547e-07,1.768556e-07,1.768564e-07,1.768573e-07,1.768581e-07,1.768590e-07,1.768598e-07,1.768607e-07,1.768615e-07,1.768624e-07,1.768632e-07,1.768641e-07,1.768649e-07,1.768658e-07,1.768666e-07,1.768674e-07,1.768683e-07,1.768691e-07,1.768700e-07,1.768708e-07,1.768717e-07,1.768725e-07,1.768734e-07,1.768742e-07,1.768751e-07,1.768759e-07,1.768767e-07,1.768776e-07,1.768784e-07,1.768793e-07,1.768801e-07,1.768810e-07,1.768818e-07,1.768827e-07,1.768835e-07,1.768843e-07,1.768852e-07,1.768860e-07,1.768869e-07,1.768877e-07,1.768886e-07,1.768894e-07,1.768903e-07,1.768911e-07,1.768919e-07,1.768928e-07,1.768936e-07,1.768945e-07,1.768953e-07,1.768962e-07,1.768970e-07,1.768979e-07,1.768987e-07,1.768995e-07,1.769004e-07,1.769012e-07,1.769021e-07,1.769029e-07,1.769038e-07,1.769046e-07,1.769054e-07,1.769063e-07,1.769071e-07,1.769080e-07,1.769088e-07,1.769097e-07,1.769105e-07,1.769113e-07,1.769122e-07,1.769130e-07,1.769139e-07,1.769147e-07,1.769156e-07,1.769164e-07,1.769172e-07,1.769181e-07,1.769189e-07,1.769198e-07,1.769206e-07,1.769215e-07,1.769223e-07,1.769231e-07,1.769240e-07,1.769248e-07,1.769257e-07,1.769265e-07,1.769273e-07,1.769282e-07,1.769290e-07,1.769299e-07,1.769307e-07,1.769316e-07,1.769324e-07,1.769332e-07,1.769341e-07,1.769349e-07,1.769358e-07,1.769366e-07,1.769374e-07,1.769383e-07,1.769391e-07,1.769400e-07,1.769408e-07,1.769416e-07,1.769425e-07,1.769433e-07,1.769442e-07,1.769450e-07,1.769458e-07,1.769467e-07,1.769475e-07,1.769484e-07,1.769492e-07,1.769500e-07,1.769509e-07,1.769517e-07,1.769526e-07,1.769534e-07,1.769542e-07,1.769551e-07,1.769559e-07,1.769568e-07,1.769576e-07,1.769584e-07,1.769593e-07,1.769601e-07,1.769610e-07,1.769618e-07,1.769626e-07,1.769635e-07,1.769643e-07,1.769652e-07,1.769660e-07,1.769668e-07,1.769677e-07,1.769685e-07,1.769693e-07,1.769702e-07,1.769710e-07,1.769719e-07,1.769727e-07,1.769735e-07,1.769744e-07,1.769752e-07,1.769761e-07,1.769769e-07,1.769777e-07,1.769786e-07,1.769794e-07,1.769802e-07,1.769811e-07,1.769819e-07,1.769828e-07,1.769836e-07,1.769844e-07,1.769853e-07,1.769861e-07,1.769869e-07,1.769878e-07,1.769886e-07,1.769895e-07,1.769903e-07,1.769911e-07,1.769920e-07,1.769928e-07,1.769936e-07,1.769945e-07,1.769953e-07,1.769961e-07,1.769970e-07,1.769978e-07,1.769987e-07,1.769995e-07,1.770003e-07,1.770012e-07,1.770020e-07,1.770028e-07,1.770037e-07,1.770045e-07,1.770053e-07,1.770062e-07,1.770070e-07,1.770079e-07,1.770087e-07,1.770095e-07,1.770104e-07,1.770112e-07,1.770120e-07,1.770129e-07,1.770137e-07,1.770145e-07,1.770154e-07,1.770162e-07,1.770170e-07,1.770179e-07,1.770187e-07,1.770195e-07,1.770204e-07,1.770212e-07,1.770220e-07,1.770229e-07,1.770237e-07,1.770246e-07,1.770254e-07,1.770262e-07,1.770271e-07,1.770279e-07,1.770287e-07,1.770296e-07,1.770304e-07,1.770312e-07,1.770321e-07,1.770329e-07,1.770337e-07,1.770346e-07,1.770354e-07,1.770362e-07,1.770371e-07,1.770379e-07,1.770387e-07,1.770396e-07,1.770404e-07,1.770412e-07,1.770421e-07,1.770429e-07,1.770437e-07,1.770446e-07,1.770454e-07,1.770462e-07,1.770471e-07,1.770479e-07,1.770487e-07,1.770496e-07,1.770504e-07,1.770512e-07,1.770521e-07,1.770529e-07,1.770537e-07,1.770546e-07,1.770554e-07,1.770562e-07,1.770571e-07,1.770579e-07,1.770587e-07,1.770596e-07,1.770604e-07,1.770612e-07,1.770620e-07,1.770629e-07,1.770637e-07,1.770645e-07,1.770654e-07,1.770662e-07,1.770670e-07,1.770679e-07,1.770687e-07,1.770695e-07,1.770704e-07,1.770712e-07,1.770720e-07,1.770729e-07,1.770737e-07,1.770745e-07,1.770753e-07,1.770762e-07,1.770770e-07,1.770778e-07,1.770787e-07,1.770795e-07,1.770803e-07,1.770812e-07,1.770820e-07,1.770828e-07,1.770837e-07,1.770845e-07,1.770853e-07,1.770861e-07,1.770870e-07,1.770878e-07,1.770886e-07,1.770895e-07,1.770903e-07,1.770911e-07,1.770920e-07,1.770928e-07,1.770936e-07,1.770944e-07,1.770953e-07,1.770961e-07,1.770969e-07,1.770978e-07,1.770986e-07,1.770994e-07,1.771002e-07,1.771011e-07,1.771019e-07,1.771027e-07,1.771036e-07,1.771044e-07,1.771052e-07,1.771061e-07,1.771069e-07,1.771077e-07,1.771085e-07,1.771094e-07,1.771102e-07,1.771110e-07,1.771119e-07,1.771127e-07,1.771135e-07,1.771143e-07,1.771152e-07,1.771160e-07,1.771168e-07,1.771176e-07,1.771185e-07,1.771193e-07,1.771201e-07,1.771210e-07,1.771218e-07,1.771226e-07,1.771234e-07,1.771243e-07,1.771251e-07,1.771259e-07,1.771267e-07,1.771276e-07,1.771284e-07,1.771292e-07,1.771301e-07,1.771309e-07,1.771317e-07,1.771325e-07,1.771334e-07,1.771342e-07,1.771350e-07,1.771358e-07,1.771367e-07,1.771375e-07,1.771383e-07,1.771392e-07,1.771400e-07,1.771408e-07,1.771416e-07,1.771425e-07,1.771433e-07,1.771441e-07,1.771449e-07,1.771458e-07,1.771466e-07,1.771474e-07,1.771482e-07,1.771491e-07,1.771499e-07,1.771507e-07,1.771515e-07,1.771524e-07,1.771532e-07,1.771540e-07,1.771548e-07,1.771557e-07,1.771565e-07,1.771573e-07,1.771581e-07,1.771590e-07,1.771598e-07,1.771606e-07,1.771614e-07,1.771623e-07,1.771631e-07,1.771639e-07,1.771647e-07,1.771656e-07,1.771664e-07,1.771672e-07,1.771680e-07,1.771689e-07,1.771697e-07,1.771705e-07,1.771713e-07,1.771722e-07,1.771730e-07,1.771738e-07,1.771746e-07,1.771755e-07,1.771763e-07,1.771771e-07,1.771779e-07,1.771787e-07,1.771796e-07,1.771804e-07,1.771812e-07,1.771820e-07,1.771829e-07,1.771837e-07,1.771845e-07,1.771853e-07,1.771862e-07,1.771870e-07,1.771878e-07,1.771886e-07,1.771894e-07,1.771903e-07,1.771911e-07,1.771919e-07,1.771927e-07,1.771936e-07,1.771944e-07,1.771952e-07,1.771960e-07,1.771969e-07,1.771977e-07,1.771985e-07,1.771993e-07,1.772001e-07,1.772010e-07,1.772018e-07,1.772026e-07,1.772034e-07,1.772043e-07,1.772051e-07,1.772059e-07,1.772067e-07,1.772075e-07,1.772084e-07,1.772092e-07,1.772100e-07,1.772108e-07,1.772116e-07,1.772125e-07,1.772133e-07,1.772141e-07,1.772149e-07,1.772157e-07,1.772166e-07,1.772174e-07,1.772182e-07,1.772190e-07,1.772199e-07,1.772207e-07,1.772215e-07,1.772223e-07,1.772231e-07,1.772240e-07,1.772248e-07,1.772256e-07,1.772264e-07,1.772272e-07,1.772281e-07,1.772289e-07,1.772297e-07,1.772305e-07,1.772313e-07,1.772322e-07,1.772330e-07,1.772338e-07,1.772346e-07,1.772354e-07,1.772363e-07,1.772371e-07,1.772379e-07,1.772387e-07,1.772395e-07,1.772404e-07,1.772412e-07,1.772420e-07,1.772428e-07,1.772436e-07,1.772444e-07,1.772453e-07,1.772461e-07,1.772469e-07,1.772477e-07,1.772485e-07,1.772494e-07,1.772502e-07,1.772510e-07,1.772518e-07,1.772526e-07,1.772535e-07,1.772543e-07,1.772551e-07,1.772559e-07,1.772567e-07,1.772575e-07,1.772584e-07,1.772592e-07,1.772600e-07,1.772608e-07,1.772616e-07,1.772624e-07,1.772633e-07,1.772641e-07,1.772649e-07,1.772657e-07,1.772665e-07,1.772674e-07,1.772682e-07,1.772690e-07,1.772698e-07,1.772706e-07,1.772714e-07,1.772723e-07,1.772731e-07,1.772739e-07,1.772747e-07,1.772755e-07,1.772763e-07,1.772772e-07,1.772780e-07,1.772788e-07,1.772796e-07,1.772804e-07,1.772812e-07,1.772821e-07,1.772829e-07,1.772837e-07,1.772845e-07,1.772853e-07,1.772861e-07,1.772870e-07,1.772878e-07,1.772886e-07,1.772894e-07,1.772902e-07,1.772910e-07,1.772918e-07,1.772927e-07,1.772935e-07,1.772943e-07,1.772951e-07,1.772959e-07,1.772967e-07,1.772976e-07,1.772984e-07,1.772992e-07,1.773000e-07,1.773008e-07,1.773016e-07,1.773024e-07,1.773033e-07,1.773041e-07,1.773049e-07,1.773057e-07,1.773065e-07,1.773073e-07,1.773081e-07,1.773090e-07,1.773098e-07,1.773106e-07,1.773114e-07,1.773122e-07,1.773130e-07,1.773138e-07,1.773147e-07,1.773155e-07,1.773163e-07,1.773171e-07,1.773179e-07,1.773187e-07,1.773195e-07,1.773204e-07,1.773212e-07,1.773220e-07,1.773228e-07,1.773236e-07,1.773244e-07,1.773252e-07,1.773261e-07,1.773269e-07,1.773277e-07,1.773285e-07,1.773293e-07,1.773301e-07,1.773309e-07,1.773317e-07,1.773326e-07,1.773334e-07,1.773342e-07,1.773350e-07,1.773358e-07,1.773366e-07,1.773374e-07,1.773382e-07,1.773391e-07,1.773399e-07,1.773407e-07,1.773415e-07,1.773423e-07,1.773431e-07,1.773439e-07,1.773447e-07,1.773456e-07,1.773464e-07,1.773472e-07,1.773480e-07,1.773488e-07,1.773496e-07,1.773504e-07,1.773512e-07,1.773520e-07,1.773529e-07,1.773537e-07,1.773545e-07,1.773553e-07,1.773561e-07,1.773569e-07,1.773577e-07,1.773585e-07,1.773593e-07,1.773602e-07,1.773610e-07,1.773618e-07,1.773626e-07,1.773634e-07,1.773642e-07,1.773650e-07,1.773658e-07,1.773666e-07,1.773674e-07,1.773683e-07,1.773691e-07,1.773699e-07,1.773707e-07,1.773715e-07,1.773723e-07,1.773731e-07,1.773739e-07,1.773747e-07,1.773756e-07,1.773764e-07,1.773772e-07,1.773780e-07,1.773788e-07,1.773796e-07,1.773804e-07,1.773812e-07,1.773820e-07,1.773828e-07,1.773836e-07,1.773845e-07,1.773853e-07,1.773861e-07,1.773869e-07,1.773877e-07,1.773885e-07,1.773893e-07,1.773901e-07,1.773909e-07,1.773917e-07,1.773925e-07,1.773934e-07,1.773942e-07,1.773950e-07,1.773958e-07,1.773966e-07,1.773974e-07,1.773982e-07,1.773990e-07,1.773998e-07,1.774006e-07,1.774014e-07,1.774022e-07,1.774030e-07,1.774039e-07,1.774047e-07,1.774055e-07,1.774063e-07,1.774071e-07,1.774079e-07,1.774087e-07,1.774095e-07,1.774103e-07,1.774111e-07,1.774119e-07,1.774127e-07,1.774135e-07,1.774144e-07,1.774152e-07,1.774160e-07,1.774168e-07,1.774176e-07,1.774184e-07,1.774192e-07,1.774200e-07,1.774208e-07,1.774216e-07,1.774224e-07,1.774232e-07,1.774240e-07,1.774248e-07,1.774256e-07,1.774265e-07,1.774273e-07,1.774281e-07,1.774289e-07,1.774297e-07,1.774305e-07,1.774313e-07,1.774321e-07,1.774329e-07,1.774337e-07,1.774345e-07,1.774353e-07,1.774361e-07,1.774369e-07,1.774377e-07,1.774385e-07,1.774393e-07,1.774401e-07,1.774410e-07,1.774418e-07,1.774426e-07,1.774434e-07,1.774442e-07,1.774450e-07,1.774458e-07,1.774466e-07,1.774474e-07,1.774482e-07,1.774490e-07,1.774498e-07,1.774506e-07,1.774514e-07,1.774522e-07,1.774530e-07,1.774538e-07,1.774546e-07,1.774554e-07,1.774562e-07,1.774570e-07,1.774579e-07,1.774587e-07,1.774595e-07,1.774603e-07,1.774611e-07,1.774619e-07,1.774627e-07,1.774635e-07,1.774643e-07,1.774651e-07,1.774659e-07,1.774667e-07,1.774675e-07,1.774683e-07,1.774691e-07,1.774699e-07,1.774707e-07,1.774715e-07,1.774723e-07,1.774731e-07,1.774739e-07,1.774747e-07,1.774755e-07,1.774763e-07,1.774771e-07,1.774779e-07,1.774787e-07,1.774795e-07,1.774803e-07,1.774811e-07,1.774819e-07,1.774828e-07,1.774836e-07,1.774844e-07,1.774852e-07,1.774860e-07,1.774868e-07,1.774876e-07,1.774884e-07,1.774892e-07,1.774900e-07,1.774908e-07,1.774916e-07,1.774924e-07,1.774932e-07,1.774940e-07,1.774948e-07,1.774956e-07,1.774964e-07,1.774972e-07,1.774980e-07,1.774988e-07,1.774996e-07,1.775004e-07,1.775012e-07,1.775020e-07,1.775028e-07,1.775036e-07,1.775044e-07,1.775052e-07,1.775060e-07,1.775068e-07,1.775076e-07,1.775084e-07,1.775092e-07,1.775100e-07,1.775108e-07,1.775116e-07,1.775124e-07,1.775132e-07,1.775140e-07,1.775148e-07,1.775156e-07,1.775164e-07,1.775172e-07,1.775180e-07,1.775188e-07,1.775196e-07,1.775204e-07,1.775212e-07,1.775220e-07,1.775228e-07,1.775236e-07,1.775244e-07,1.775252e-07,1.775260e-07,1.775268e-07,1.775276e-07,1.775284e-07,1.775292e-07,1.775300e-07,1.775308e-07,1.775316e-07,1.775324e-07,1.775332e-07,1.775340e-07,1.775348e-07,1.775356e-07,1.775364e-07,1.775372e-07,1.775380e-07,1.775388e-07,1.775396e-07,1.775404e-07,1.775412e-07,1.775420e-07,1.775428e-07,1.775436e-07,1.775444e-07,1.775452e-07,1.775460e-07,1.775468e-07,1.775476e-07,1.775484e-07,1.775492e-07,1.775500e-07,1.775507e-07,1.775515e-07,1.775523e-07,1.775531e-07,1.775539e-07,1.775547e-07,1.775555e-07,1.775563e-07,1.775571e-07,1.775579e-07,1.775587e-07,1.775595e-07,1.775603e-07,1.775611e-07,1.775619e-07,1.775627e-07,1.775635e-07,1.775643e-07,1.775651e-07,1.775659e-07,1.775667e-07,1.775675e-07,1.775683e-07,1.775691e-07,1.775699e-07,1.775707e-07,1.775715e-07,1.775723e-07,1.775731e-07,1.775739e-07,1.775747e-07,1.775755e-07,1.775762e-07,1.775770e-07,1.775778e-07,1.775786e-07,1.775794e-07,1.775802e-07,1.775810e-07,1.775818e-07,1.775826e-07,1.775834e-07,1.775842e-07,1.775850e-07,1.775858e-07,1.775866e-07,1.775874e-07,1.775882e-07,1.775890e-07,1.775898e-07,1.775906e-07,1.775914e-07,1.775922e-07,1.775929e-07,1.775937e-07,1.775945e-07,1.775953e-07,1.775961e-07,1.775969e-07,1.775977e-07,1.775985e-07,1.775993e-07,1.776001e-07,1.776009e-07,1.776017e-07,1.776025e-07,1.776033e-07,1.776041e-07,1.776049e-07,1.776057e-07,1.776065e-07,1.776072e-07,1.776080e-07,1.776088e-07,1.776096e-07,1.776104e-07,1.776112e-07,1.776120e-07,1.776128e-07,1.776136e-07,1.776144e-07,1.776152e-07,1.776160e-07,1.776168e-07,1.776176e-07,1.776184e-07,1.776191e-07,1.776199e-07,1.776207e-07,1.776215e-07,1.776223e-07,1.776231e-07,1.776239e-07,1.776247e-07,1.776255e-07,1.776263e-07,1.776271e-07,1.776279e-07,1.776287e-07,1.776295e-07,1.776302e-07,1.776310e-07,1.776318e-07,1.776326e-07,1.776334e-07,1.776342e-07,1.776350e-07,1.776358e-07,1.776366e-07,1.776374e-07,1.776382e-07,1.776390e-07,1.776397e-07,1.776405e-07,1.776413e-07,1.776421e-07,1.776429e-07,1.776437e-07,1.776445e-07,1.776453e-07,1.776461e-07,1.776469e-07,1.776477e-07,1.776485e-07,1.776492e-07,1.776500e-07,1.776508e-07,1.776516e-07,1.776524e-07,1.776532e-07,1.776540e-07,1.776548e-07,1.776556e-07,1.776564e-07,1.776571e-07,1.776579e-07,1.776587e-07,1.776595e-07,1.776603e-07,1.776611e-07,1.776619e-07,1.776627e-07,1.776635e-07,1.776643e-07,1.776650e-07,1.776658e-07,1.776666e-07,1.776674e-07,1.776682e-07,1.776690e-07,1.776698e-07,1.776706e-07,1.776714e-07,1.776722e-07,1.776729e-07,1.776737e-07,1.776745e-07,1.776753e-07,1.776761e-07,1.776769e-07,1.776777e-07,1.776785e-07,1.776793e-07,1.776800e-07,1.776808e-07,1.776816e-07,1.776824e-07,1.776832e-07,1.776840e-07,1.776848e-07,1.776856e-07,1.776864e-07,1.776871e-07,1.776879e-07,1.776887e-07,1.776895e-07,1.776903e-07,1.776911e-07,1.776919e-07,1.776927e-07,1.776934e-07,1.776942e-07,1.776950e-07,1.776958e-07,1.776966e-07,1.776974e-07,1.776982e-07,1.776990e-07,1.776998e-07,1.777005e-07,1.777013e-07,1.777021e-07,1.777029e-07,1.777037e-07,1.777045e-07,1.777053e-07,1.777060e-07,1.777068e-07,1.777076e-07,1.777084e-07,1.777092e-07,1.777100e-07,1.777108e-07,1.777116e-07,1.777123e-07,1.777131e-07,1.777139e-07,1.777147e-07,1.777155e-07,1.777163e-07,1.777171e-07,1.777179e-07,1.777186e-07,1.777194e-07,1.777202e-07,1.777210e-07,1.777218e-07,1.777226e-07,1.777234e-07,1.777241e-07,1.777249e-07,1.777257e-07,1.777265e-07,1.777273e-07,1.777281e-07,1.777289e-07,1.777296e-07,1.777304e-07,1.777312e-07,1.777320e-07,1.777328e-07,1.777336e-07,1.777344e-07,1.777351e-07,1.777359e-07,1.777367e-07,1.777375e-07,1.777383e-07,1.777391e-07,1.777398e-07,1.777406e-07,1.777414e-07,1.777422e-07,1.777430e-07,1.777438e-07,1.777446e-07,1.777453e-07,1.777461e-07,1.777469e-07,1.777477e-07,1.777485e-07,1.777493e-07,1.777500e-07,1.777508e-07,1.777516e-07,1.777524e-07,1.777532e-07,1.777540e-07,1.777547e-07,1.777555e-07,1.777563e-07,1.777571e-07,1.777579e-07,1.777587e-07,1.777594e-07,1.777602e-07,1.777610e-07,1.777618e-07,1.777626e-07,1.777634e-07,1.777641e-07,1.777649e-07,1.777657e-07,1.777665e-07,1.777673e-07,1.777681e-07,1.777688e-07,1.777696e-07,1.777704e-07,1.777712e-07,1.777720e-07,1.777728e-07,1.777735e-07,1.777743e-07,1.777751e-07,1.777759e-07,1.777767e-07,1.777775e-07,1.777782e-07,1.777790e-07,1.777798e-07,1.777806e-07,1.777814e-07,1.777821e-07,1.777829e-07,1.777837e-07,1.777845e-07,1.777853e-07,1.777861e-07,1.777868e-07,1.777876e-07,1.777884e-07,1.777892e-07,1.777900e-07,1.777907e-07,1.777915e-07,1.777923e-07,1.777931e-07,1.777939e-07,1.777947e-07,1.777954e-07,1.777962e-07,1.777970e-07,1.777978e-07,1.777986e-07,1.777993e-07,1.778001e-07,1.778009e-07,1.778017e-07,1.778025e-07,1.778032e-07,1.778040e-07,1.778048e-07,1.778056e-07,1.778064e-07,1.778071e-07,1.778079e-07,1.778087e-07,1.778095e-07,1.778103e-07,1.778110e-07,1.778118e-07,1.778126e-07,1.778134e-07,1.778142e-07,1.778149e-07,1.778157e-07,1.778165e-07,1.778173e-07,1.778181e-07,1.778188e-07,1.778196e-07,1.778204e-07,1.778212e-07,1.778220e-07,1.778227e-07,1.778235e-07,1.778243e-07,1.778251e-07,1.778259e-07,1.778266e-07,1.778274e-07,1.778282e-07,1.778290e-07,1.778298e-07,1.778305e-07,1.778313e-07,1.778321e-07,1.778329e-07,1.778336e-07,1.778344e-07,1.778352e-07,1.778360e-07,1.778368e-07,1.778375e-07,1.778383e-07,1.778391e-07,1.778399e-07,1.778406e-07,1.778414e-07,1.778422e-07,1.778430e-07,1.778438e-07,1.778445e-07,1.778453e-07,1.778461e-07,1.778469e-07,1.778476e-07,1.778484e-07,1.778492e-07,1.778500e-07,1.778508e-07,1.778515e-07,1.778523e-07,1.778531e-07,1.778539e-07,1.778546e-07,1.778554e-07,1.778562e-07,1.778570e-07,1.778578e-07,1.778585e-07,1.778593e-07,1.778601e-07,1.778609e-07,1.778616e-07,1.778624e-07,1.778632e-07,1.778640e-07,1.778647e-07,1.778655e-07,1.778663e-07,1.778671e-07,1.778678e-07,1.778686e-07,1.778694e-07,1.778702e-07,1.778710e-07,1.778717e-07,1.778725e-07,1.778733e-07,1.778741e-07,1.778748e-07,1.778756e-07,1.778764e-07,1.778772e-07,1.778779e-07,1.778787e-07,1.778795e-07,1.778803e-07,1.778810e-07,1.778818e-07,1.778826e-07,1.778834e-07,1.778841e-07,1.778849e-07,1.778857e-07,1.778865e-07,1.778872e-07,1.778880e-07,1.778888e-07,1.778896e-07,1.778903e-07,1.778911e-07,1.778919e-07,1.778927e-07,1.778934e-07,1.778942e-07,1.778950e-07,1.778958e-07,1.778965e-07,1.778973e-07,1.778981e-07,1.778989e-07,1.778996e-07,1.779004e-07,1.779012e-07,1.779020e-07,1.779027e-07,1.779035e-07,1.779043e-07,1.779050e-07,1.779058e-07,1.779066e-07,1.779074e-07,1.779081e-07,1.779089e-07,1.779097e-07,1.779105e-07,1.779112e-07,1.779120e-07,1.779128e-07,1.779136e-07,1.779143e-07,1.779151e-07,1.779159e-07,1.779166e-07,1.779174e-07,1.779182e-07,1.779190e-07,1.779197e-07,1.779205e-07,1.779213e-07,1.779221e-07,1.779228e-07,1.779236e-07,1.779244e-07,1.779251e-07,1.779259e-07,1.779267e-07,1.779275e-07,1.779282e-07,1.779290e-07,1.779298e-07,1.779306e-07,1.779313e-07,1.779321e-07,1.779329e-07,1.779336e-07,1.779344e-07,1.779352e-07,1.779360e-07,1.779367e-07,1.779375e-07,1.779383e-07,1.779390e-07,1.779398e-07,1.779406e-07,1.779414e-07,1.779421e-07,1.779429e-07,1.779437e-07,1.779444e-07,1.779452e-07,1.779460e-07,1.779468e-07,1.779475e-07,1.779483e-07,1.779491e-07,1.779498e-07,1.779506e-07,1.779514e-07,1.779522e-07,1.779529e-07,1.779537e-07,1.779545e-07,1.779552e-07,1.779560e-07,1.779568e-07,1.779575e-07,1.779583e-07,1.779591e-07,1.779599e-07,1.779606e-07,1.779614e-07,1.779622e-07,1.779629e-07,1.779637e-07,1.779645e-07,1.779652e-07,1.779660e-07,1.779668e-07,1.779676e-07,1.779683e-07,1.779691e-07,1.779699e-07,1.779706e-07,1.779714e-07,1.779722e-07,1.779729e-07,1.779737e-07,1.779745e-07,1.779752e-07,1.779760e-07,1.779768e-07,1.779776e-07,1.779783e-07,1.779791e-07,1.779799e-07,1.779806e-07,1.779814e-07,1.779822e-07,1.779829e-07,1.779837e-07,1.779845e-07,1.779852e-07,1.779860e-07,1.779868e-07,1.779875e-07,1.779883e-07,1.779891e-07,1.779899e-07,1.779906e-07,1.779914e-07,1.779922e-07,1.779929e-07,1.779937e-07,1.779945e-07,1.779952e-07,1.779960e-07,1.779968e-07,1.779975e-07,1.779983e-07,1.779991e-07,1.779998e-07,1.780006e-07,1.780014e-07,1.780021e-07,1.780029e-07,1.780037e-07,1.780044e-07,1.780052e-07,1.780060e-07,1.780067e-07,1.780075e-07,1.780083e-07,1.780090e-07,1.780098e-07,1.780106e-07,1.780113e-07,1.780121e-07,1.780129e-07,1.780136e-07,1.780144e-07,1.780152e-07,1.780159e-07,1.780167e-07,1.780175e-07,1.780182e-07,1.780190e-07,1.780198e-07,1.780205e-07,1.780213e-07,1.780221e-07,1.780228e-07,1.780236e-07,1.780244e-07,1.780251e-07,1.780259e-07,1.780267e-07,1.780274e-07,1.780282e-07,1.780290e-07,1.780297e-07,1.780305e-07,1.780313e-07,1.780320e-07,1.780328e-07,1.780336e-07,1.780343e-07,1.780351e-07,1.780358e-07,1.780366e-07,1.780374e-07,1.780381e-07,1.780389e-07,1.780397e-07,1.780404e-07,1.780412e-07,1.780420e-07,1.780427e-07,1.780435e-07,1.780443e-07,1.780450e-07,1.780458e-07,1.780466e-07,1.780473e-07,1.780481e-07,1.780488e-07,1.780496e-07,1.780504e-07,1.780511e-07,1.780519e-07,1.780527e-07,1.780534e-07,1.780542e-07,1.780550e-07,1.780557e-07,1.780565e-07,1.780573e-07,1.780580e-07,1.780588e-07,1.780595e-07,1.780603e-07,1.780611e-07,1.780618e-07,1.780626e-07,1.780634e-07,1.780641e-07,1.780649e-07,1.780657e-07,1.780664e-07,1.780672e-07,1.780679e-07,1.780687e-07,1.780695e-07,1.780702e-07,1.780710e-07,1.780718e-07,1.780725e-07,1.780733e-07,1.780740e-07,1.780748e-07,1.780756e-07,1.780763e-07,1.780771e-07,1.780779e-07,1.780786e-07,1.780794e-07,1.780801e-07,1.780809e-07,1.780817e-07,1.780824e-07,1.780832e-07,1.780840e-07,1.780847e-07,1.780855e-07,1.780862e-07,1.780870e-07,1.780878e-07,1.780885e-07,1.780893e-07,1.780900e-07,1.780908e-07,1.780916e-07,1.780923e-07,1.780931e-07,1.780939e-07,1.780946e-07,1.780954e-07,1.780961e-07,1.780969e-07,1.780977e-07,1.780984e-07,1.780992e-07,1.780999e-07,1.781007e-07,1.781015e-07,1.781022e-07,1.781030e-07,1.781037e-07,1.781045e-07,1.781053e-07,1.781060e-07,1.781068e-07,1.781075e-07,1.781083e-07,1.781091e-07,1.781098e-07,1.781106e-07,1.781114e-07,1.781121e-07,1.781129e-07,1.781136e-07,1.781144e-07,1.781152e-07,1.781159e-07,1.781167e-07,1.781174e-07,1.781182e-07,1.781189e-07,1.781197e-07,1.781205e-07,1.781212e-07,1.781220e-07,1.781227e-07,1.781235e-07,1.781243e-07,1.781250e-07,1.781258e-07,1.781265e-07,1.781273e-07,1.781281e-07,1.781288e-07,1.781296e-07,1.781303e-07,1.781311e-07,1.781319e-07,1.781326e-07,1.781334e-07,1.781341e-07,1.781349e-07,1.781357e-07,1.781364e-07,1.781372e-07,1.781379e-07,1.781387e-07,1.781394e-07,1.781402e-07,1.781410e-07,1.781417e-07,1.781425e-07,1.781432e-07,1.781440e-07,1.781448e-07,1.781455e-07,1.781463e-07,1.781470e-07,1.781478e-07,1.781485e-07,1.781493e-07,1.781501e-07,1.781508e-07,1.781516e-07,1.781523e-07,1.781531e-07,1.781538e-07,1.781546e-07,1.781554e-07,1.781561e-07,1.781569e-07,1.781576e-07,1.781584e-07,1.781591e-07,1.781599e-07,1.781607e-07,1.781614e-07,1.781622e-07,1.781629e-07,1.781637e-07,1.781644e-07,1.781652e-07,1.781660e-07,1.781667e-07,1.781675e-07,1.781682e-07,1.781690e-07,1.781697e-07,1.781705e-07,1.781713e-07,1.781720e-07,1.781728e-07,1.781735e-07,1.781743e-07,1.781750e-07,1.781758e-07,1.781765e-07,1.781773e-07,1.781781e-07,1.781788e-07,1.781796e-07,1.781803e-07,1.781811e-07,1.781818e-07,1.781826e-07,1.781833e-07,1.781841e-07,1.781849e-07,1.781856e-07,1.781864e-07,1.781871e-07,1.781879e-07,1.781886e-07,1.781894e-07,1.781901e-07,1.781909e-07,1.781917e-07,1.781924e-07,1.781932e-07,1.781939e-07,1.781947e-07,1.781954e-07,1.781962e-07,1.781969e-07,1.781977e-07,1.781984e-07,1.781992e-07,1.782000e-07,1.782007e-07,1.782015e-07,1.782022e-07,1.782030e-07,1.782037e-07,1.782045e-07,1.782052e-07,1.782060e-07,1.782067e-07,1.782075e-07,1.782082e-07,1.782090e-07,1.782098e-07,1.782105e-07,1.782113e-07,1.782120e-07,1.782128e-07,1.782135e-07,1.782143e-07,1.782150e-07,1.782158e-07,1.782165e-07,1.782173e-07,1.782180e-07,1.782188e-07,1.782196e-07,1.782203e-07,1.782211e-07,1.782218e-07,1.782226e-07,1.782233e-07,1.782241e-07,1.782248e-07,1.782256e-07,1.782263e-07,1.782271e-07,1.782278e-07,1.782286e-07,1.782293e-07,1.782301e-07,1.782308e-07,1.782316e-07,1.782323e-07,1.782331e-07,1.782339e-07,1.782346e-07,1.782354e-07,1.782361e-07,1.782369e-07,1.782376e-07,1.782384e-07,1.782391e-07,1.782399e-07,1.782406e-07,1.782414e-07,1.782421e-07,1.782429e-07,1.782436e-07,1.782444e-07,1.782451e-07,1.782459e-07,1.782466e-07,1.782474e-07,1.782481e-07,1.782489e-07,1.782496e-07,1.782504e-07,1.782511e-07,1.782519e-07,1.782526e-07,1.782534e-07,1.782541e-07,1.782549e-07,1.782556e-07,1.782564e-07,1.782571e-07,1.782579e-07,1.782586e-07,1.782594e-07,1.782602e-07,1.782609e-07,1.782617e-07,1.782624e-07,1.782632e-07,1.782639e-07,1.782647e-07,1.782654e-07,1.782662e-07,1.782669e-07,1.782677e-07,1.782684e-07,1.782692e-07,1.782699e-07,1.782707e-07,1.782714e-07,1.782722e-07,1.782729e-07,1.782737e-07,1.782744e-07,1.782752e-07,1.782759e-07,1.782767e-07,1.782774e-07,1.782781e-07,1.782789e-07,1.782796e-07,1.782804e-07,1.782811e-07,1.782819e-07,1.782826e-07,1.782834e-07,1.782841e-07,1.782849e-07,1.782856e-07,1.782864e-07,1.782871e-07,1.782879e-07,1.782886e-07,1.782894e-07,1.782901e-07,1.782909e-07,1.782916e-07,1.782924e-07,1.782931e-07,1.782939e-07,1.782946e-07,1.782954e-07,1.782961e-07,1.782969e-07,1.782976e-07,1.782984e-07,1.782991e-07,1.782999e-07,1.783006e-07,1.783014e-07,1.783021e-07,1.783029e-07,1.783036e-07,1.783043e-07,1.783051e-07,1.783058e-07,1.783066e-07,1.783073e-07,1.783081e-07,1.783088e-07,1.783096e-07,1.783103e-07,1.783111e-07,1.783118e-07,1.783126e-07,1.783133e-07,1.783141e-07,1.783148e-07,1.783156e-07,1.783163e-07,1.783171e-07,1.783178e-07,1.783185e-07,1.783193e-07,1.783200e-07,1.783208e-07,1.783215e-07,1.783223e-07,1.783230e-07,1.783238e-07,1.783245e-07,1.783253e-07,1.783260e-07,1.783268e-07,1.783275e-07,1.783282e-07,1.783290e-07,1.783297e-07,1.783305e-07,1.783312e-07,1.783320e-07,1.783327e-07,1.783335e-07,1.783342e-07,1.783350e-07,1.783357e-07,1.783365e-07,1.783372e-07,1.783379e-07,1.783387e-07,1.783394e-07,1.783402e-07,1.783409e-07,1.783417e-07,1.783424e-07,1.783432e-07,1.783439e-07,1.783447e-07,1.783454e-07,1.783461e-07,1.783469e-07,1.783476e-07,1.783484e-07,1.783491e-07,1.783499e-07,1.783506e-07,1.783514e-07,1.783521e-07,1.783528e-07,1.783536e-07,1.783543e-07,1.783551e-07,1.783558e-07,1.783566e-07,1.783573e-07,1.783581e-07,1.783588e-07,1.783595e-07,1.783603e-07,1.783610e-07,1.783618e-07,1.783625e-07,1.783633e-07,1.783640e-07,1.783648e-07,1.783655e-07,1.783662e-07,1.783670e-07,1.783677e-07,1.783685e-07,1.783692e-07,1.783700e-07,1.783707e-07,1.783714e-07,1.783722e-07,1.783729e-07,1.783737e-07,1.783744e-07,1.783752e-07,1.783759e-07,1.783766e-07,1.783774e-07,1.783781e-07,1.783789e-07,1.783796e-07,1.783804e-07,1.783811e-07,1.783818e-07,1.783826e-07,1.783833e-07,1.783841e-07,1.783848e-07,1.783856e-07,1.783863e-07,1.783870e-07,1.783878e-07,1.783885e-07,1.783893e-07,1.783900e-07,1.783908e-07,1.783915e-07,1.783922e-07,1.783930e-07,1.783937e-07,1.783945e-07,1.783952e-07,1.783960e-07,1.783967e-07,1.783974e-07,1.783982e-07,1.783989e-07,1.783997e-07,1.784004e-07,1.784011e-07,1.784019e-07,1.784026e-07,1.784034e-07,1.784041e-07,1.784049e-07,1.784056e-07,1.784063e-07,1.784071e-07,1.784078e-07,1.784086e-07,1.784093e-07,1.784100e-07,1.784108e-07,1.784115e-07,1.784123e-07,1.784130e-07,1.784137e-07,1.784145e-07,1.784152e-07,1.784160e-07,1.784167e-07,1.784174e-07,1.784182e-07,1.784189e-07,1.784197e-07,1.784204e-07,1.784211e-07,1.784219e-07,1.784226e-07,1.784234e-07,1.784241e-07,1.784248e-07,1.784256e-07,1.784263e-07,1.784271e-07,1.784278e-07,1.784285e-07,1.784293e-07,1.784300e-07,1.784308e-07,1.784315e-07,1.784322e-07,1.784330e-07,1.784337e-07,1.784345e-07,1.784352e-07,1.784359e-07,1.784367e-07,1.784374e-07,1.784382e-07,1.784389e-07,1.784396e-07,1.784404e-07,1.784411e-07,1.784419e-07,1.784426e-07,1.784433e-07,1.784441e-07,1.784448e-07,1.784455e-07,1.784463e-07,1.784470e-07,1.784478e-07,1.784485e-07,1.784492e-07,1.784500e-07,1.784507e-07,1.784515e-07,1.784522e-07,1.784529e-07,1.784537e-07,1.784544e-07,1.784551e-07,1.784559e-07,1.784566e-07,1.784574e-07,1.784581e-07,1.784588e-07,1.784596e-07,1.784603e-07,1.784611e-07,1.784618e-07,1.784625e-07,1.784633e-07,1.784640e-07,1.784647e-07,1.784655e-07,1.784662e-07,1.784670e-07,1.784677e-07,1.784684e-07,1.784692e-07,1.784699e-07,1.784706e-07,1.784714e-07,1.784721e-07,1.784728e-07,1.784736e-07,1.784743e-07,1.784751e-07,1.784758e-07,1.784765e-07,1.784773e-07,1.784780e-07,1.784787e-07,1.784795e-07,1.784802e-07,1.784810e-07,1.784817e-07,1.784824e-07,1.784832e-07,1.784839e-07,1.784846e-07,1.784854e-07,1.784861e-07,1.784868e-07,1.784876e-07,1.784883e-07,1.784890e-07,1.784898e-07,1.784905e-07,1.784913e-07,1.784920e-07,1.784927e-07,1.784935e-07,1.784942e-07,1.784949e-07,1.784957e-07,1.784964e-07,1.784971e-07,1.784979e-07,1.784986e-07,1.784993e-07,1.785001e-07,1.785008e-07,1.785016e-07,1.785023e-07,1.785030e-07,1.785038e-07,1.785045e-07,1.785052e-07,1.785060e-07,1.785067e-07,1.785074e-07,1.785082e-07,1.785089e-07,1.785096e-07,1.785104e-07,1.785111e-07,1.785118e-07,1.785126e-07,1.785133e-07,1.785140e-07,1.785148e-07,1.785155e-07,1.785162e-07,1.785170e-07,1.785177e-07,1.785184e-07,1.785192e-07,1.785199e-07,1.785207e-07,1.785214e-07,1.785221e-07,1.785229e-07,1.785236e-07,1.785243e-07,1.785251e-07,1.785258e-07,1.785265e-07,1.785273e-07,1.785280e-07,1.785287e-07,1.785295e-07,1.785302e-07,1.785309e-07,1.785317e-07,1.785324e-07,1.785331e-07,1.785339e-07,1.785346e-07,1.785353e-07,1.785361e-07,1.785368e-07,1.785375e-07,1.785383e-07,1.785390e-07,1.785397e-07,1.785405e-07,1.785412e-07,1.785419e-07,1.785426e-07,1.785434e-07,1.785441e-07,1.785448e-07,1.785456e-07,1.785463e-07,1.785470e-07,1.785478e-07,1.785485e-07,1.785492e-07,1.785500e-07,1.785507e-07,1.785514e-07,1.785522e-07,1.785529e-07,1.785536e-07,1.785544e-07,1.785551e-07,1.785558e-07,1.785566e-07,1.785573e-07,1.785580e-07,1.785588e-07,1.785595e-07,1.785602e-07,1.785609e-07,1.785617e-07,1.785624e-07,1.785631e-07,1.785639e-07,1.785646e-07,1.785653e-07,1.785661e-07,1.785668e-07,1.785675e-07,1.785683e-07,1.785690e-07,1.785697e-07,1.785705e-07,1.785712e-07,1.785719e-07,1.785726e-07,1.785734e-07,1.785741e-07,1.785748e-07,1.785756e-07,1.785763e-07,1.785770e-07,1.785778e-07,1.785785e-07,1.785792e-07,1.785799e-07,1.785807e-07,1.785814e-07,1.785821e-07,1.785829e-07,1.785836e-07,1.785843e-07,1.785851e-07,1.785858e-07,1.785865e-07,1.785872e-07,1.785880e-07,1.785887e-07,1.785894e-07,1.785902e-07,1.785909e-07,1.785916e-07,1.785924e-07,1.785931e-07,1.785938e-07,1.785945e-07,1.785953e-07,1.785960e-07,1.785967e-07,1.785975e-07,1.785982e-07,1.785989e-07,1.785996e-07,1.786004e-07,1.786011e-07,1.786018e-07,1.786026e-07,1.786033e-07,1.786040e-07,1.786047e-07,1.786055e-07,1.786062e-07,1.786069e-07,1.786077e-07,1.786084e-07,1.786091e-07,1.786098e-07,1.786106e-07,1.786113e-07,1.786120e-07,1.786128e-07,1.786135e-07,1.786142e-07,1.786149e-07,1.786157e-07,1.786164e-07,1.786171e-07,1.786179e-07,1.786186e-07,1.786193e-07,1.786200e-07,1.786208e-07,1.786215e-07,1.786222e-07,1.786230e-07,1.786237e-07,1.786244e-07,1.786251e-07,1.786259e-07,1.786266e-07,1.786273e-07,1.786280e-07,1.786288e-07,1.786295e-07,1.786302e-07,1.786310e-07,1.786317e-07,1.786324e-07,1.786331e-07,1.786339e-07,1.786346e-07,1.786353e-07,1.786360e-07,1.786368e-07,1.786375e-07,1.786382e-07,1.786389e-07,1.786397e-07,1.786404e-07,1.786411e-07,1.786419e-07,1.786426e-07,1.786433e-07,1.786440e-07,1.786448e-07,1.786455e-07,1.786462e-07,1.786469e-07,1.786477e-07,1.786484e-07,1.786491e-07,1.786498e-07,1.786506e-07,1.786513e-07,1.786520e-07,1.786527e-07,1.786535e-07,1.786542e-07,1.786549e-07,1.786556e-07,1.786564e-07,1.786571e-07,1.786578e-07,1.786585e-07,1.786593e-07,1.786600e-07,1.786607e-07,1.786614e-07,1.786622e-07,1.786629e-07,1.786636e-07,1.786643e-07,1.786651e-07,1.786658e-07,1.786665e-07,1.786672e-07,1.786680e-07,1.786687e-07,1.786694e-07,1.786701e-07,1.786709e-07,1.786716e-07,1.786723e-07,1.786730e-07,1.786738e-07,1.786745e-07,1.786752e-07,1.786759e-07,1.786767e-07,1.786774e-07,1.786781e-07,1.786788e-07,1.786796e-07,1.786803e-07,1.786810e-07,1.786817e-07,1.786825e-07,1.786832e-07,1.786839e-07,1.786846e-07,1.786854e-07,1.786861e-07,1.786868e-07,1.786875e-07,1.786882e-07,1.786890e-07,1.786897e-07,1.786904e-07,1.786911e-07,1.786919e-07,1.786926e-07,1.786933e-07,1.786940e-07,1.786948e-07,1.786955e-07,1.786962e-07,1.786969e-07,1.786976e-07,1.786984e-07,1.786991e-07,1.786998e-07,1.787005e-07,1.787013e-07,1.787020e-07,1.787027e-07,1.787034e-07,1.787041e-07,1.787049e-07,1.787056e-07,1.787063e-07,1.787070e-07,1.787078e-07,1.787085e-07,1.787092e-07,1.787099e-07,1.787107e-07,1.787114e-07,1.787121e-07,1.787128e-07,1.787135e-07,1.787143e-07,1.787150e-07,1.787157e-07,1.787164e-07,1.787171e-07,1.787179e-07,1.787186e-07,1.787193e-07,1.787200e-07,1.787208e-07,1.787215e-07,1.787222e-07,1.787229e-07,1.787236e-07,1.787244e-07,1.787251e-07,1.787258e-07,1.787265e-07,1.787272e-07,1.787280e-07,1.787287e-07,1.787294e-07,1.787301e-07,1.787309e-07,1.787316e-07,1.787323e-07,1.787330e-07,1.787337e-07,1.787345e-07,1.787352e-07,1.787359e-07,1.787366e-07,1.787373e-07,1.787381e-07,1.787388e-07,1.787395e-07,1.787402e-07,1.787409e-07,1.787417e-07,1.787424e-07,1.787431e-07,1.787438e-07,1.787445e-07,1.787453e-07,1.787460e-07,1.787467e-07,1.787474e-07,1.787481e-07,1.787489e-07,1.787496e-07,1.787503e-07,1.787510e-07,1.787517e-07,1.787525e-07,1.787532e-07,1.787539e-07,1.787546e-07,1.787553e-07,1.787561e-07,1.787568e-07,1.787575e-07,1.787582e-07,1.787589e-07,1.787596e-07,1.787604e-07,1.787611e-07,1.787618e-07,1.787625e-07,1.787632e-07,1.787640e-07,1.787647e-07,1.787654e-07,1.787661e-07,1.787668e-07,1.787676e-07,1.787683e-07,1.787690e-07,1.787697e-07,1.787704e-07,1.787711e-07,1.787719e-07,1.787726e-07,1.787733e-07,1.787740e-07,1.787747e-07,1.787755e-07,1.787762e-07,1.787769e-07,1.787776e-07,1.787783e-07,1.787790e-07,1.787798e-07,1.787805e-07,1.787812e-07,1.787819e-07,1.787826e-07,1.787834e-07,1.787841e-07,1.787848e-07,1.787855e-07,1.787862e-07,1.787869e-07,1.787877e-07,1.787884e-07,1.787891e-07,1.787898e-07,1.787905e-07,1.787912e-07,1.787920e-07,1.787927e-07,1.787934e-07,1.787941e-07,1.787948e-07,1.787955e-07,1.787963e-07,1.787970e-07,1.787977e-07,1.787984e-07,1.787991e-07,1.787998e-07,1.788006e-07,1.788013e-07,1.788020e-07,1.788027e-07,1.788034e-07,1.788041e-07,1.788049e-07,1.788056e-07,1.788063e-07,1.788070e-07,1.788077e-07,1.788084e-07,1.788092e-07,1.788099e-07,1.788106e-07,1.788113e-07,1.788120e-07,1.788127e-07,1.788135e-07,1.788142e-07,1.788149e-07,1.788156e-07,1.788163e-07,1.788170e-07,1.788177e-07,1.788185e-07,1.788192e-07,1.788199e-07,1.788206e-07,1.788213e-07,1.788220e-07,1.788228e-07,1.788235e-07,1.788242e-07,1.788249e-07,1.788256e-07,1.788263e-07,1.788270e-07,1.788278e-07,1.788285e-07,1.788292e-07,1.788299e-07,1.788306e-07,1.788313e-07,1.788320e-07,1.788328e-07,1.788335e-07,1.788342e-07,1.788349e-07,1.788356e-07,1.788363e-07,1.788370e-07,1.788378e-07,1.788385e-07,1.788392e-07,1.788399e-07,1.788406e-07,1.788413e-07,1.788420e-07,1.788428e-07,1.788435e-07,1.788442e-07,1.788449e-07,1.788456e-07,1.788463e-07,1.788470e-07,1.788478e-07,1.788485e-07,1.788492e-07,1.788499e-07,1.788506e-07,1.788513e-07,1.788520e-07,1.788527e-07,1.788535e-07,1.788542e-07,1.788549e-07,1.788556e-07,1.788563e-07,1.788570e-07,1.788577e-07,1.788585e-07,1.788592e-07,1.788599e-07,1.788606e-07,1.788613e-07,1.788620e-07,1.788627e-07,1.788634e-07,1.788642e-07,1.788649e-07,1.788656e-07,1.788663e-07,1.788670e-07,1.788677e-07,1.788684e-07,1.788691e-07,1.788699e-07,1.788706e-07,1.788713e-07,1.788720e-07,1.788727e-07,1.788734e-07,1.788741e-07,1.788748e-07,1.788756e-07,1.788763e-07,1.788770e-07,1.788777e-07,1.788784e-07,1.788791e-07,1.788798e-07,1.788805e-07,1.788812e-07,1.788820e-07,1.788827e-07,1.788834e-07,1.788841e-07,1.788848e-07,1.788855e-07,1.788862e-07,1.788869e-07,1.788876e-07,1.788884e-07,1.788891e-07,1.788898e-07,1.788905e-07,1.788912e-07,1.788919e-07,1.788926e-07,1.788933e-07,1.788940e-07,1.788948e-07,1.788955e-07,1.788962e-07,1.788969e-07,1.788976e-07,1.788983e-07,1.788990e-07,1.788997e-07,1.789004e-07,1.789012e-07,1.789019e-07,1.789026e-07,1.789033e-07,1.789040e-07,1.789047e-07,1.789054e-07,1.789061e-07,1.789068e-07,1.789075e-07,1.789083e-07,1.789090e-07,1.789097e-07,1.789104e-07,1.789111e-07,1.789118e-07,1.789125e-07,1.789132e-07,1.789139e-07,1.789146e-07,1.789154e-07,1.789161e-07,1.789168e-07,1.789175e-07,1.789182e-07,1.789189e-07,1.789196e-07,1.789203e-07,1.789210e-07,1.789217e-07,1.789224e-07,1.789232e-07,1.789239e-07,1.789246e-07,1.789253e-07,1.789260e-07,1.789267e-07,1.789274e-07,1.789281e-07,1.789288e-07,1.789295e-07,1.789302e-07,1.789309e-07,1.789317e-07,1.789324e-07,1.789331e-07,1.789338e-07,1.789345e-07,1.789352e-07,1.789359e-07,1.789366e-07,1.789373e-07,1.789380e-07,1.789387e-07,1.789394e-07,1.789402e-07,1.789409e-07,1.789416e-07,1.789423e-07,1.789430e-07,1.789437e-07,1.789444e-07,1.789451e-07,1.789458e-07,1.789465e-07,1.789472e-07,1.789479e-07,1.789486e-07,1.789494e-07,1.789501e-07,1.789508e-07,1.789515e-07,1.789522e-07,1.789529e-07,1.789536e-07,1.789543e-07,1.789550e-07,1.789557e-07,1.789564e-07,1.789571e-07,1.789578e-07,1.789585e-07,1.789593e-07,1.789600e-07,1.789607e-07,1.789614e-07,1.789621e-07,1.789628e-07,1.789635e-07,1.789642e-07,1.789649e-07,1.789656e-07,1.789663e-07,1.789670e-07,1.789677e-07,1.789684e-07,1.789691e-07,1.789699e-07,1.789706e-07,1.789713e-07,1.789720e-07,1.789727e-07,1.789734e-07,1.789741e-07,1.789748e-07,1.789755e-07,1.789762e-07,1.789769e-07,1.789776e-07,1.789783e-07,1.789790e-07,1.789797e-07,1.789804e-07,1.789811e-07,1.789819e-07,1.789826e-07,1.789833e-07,1.789840e-07,1.789847e-07,1.789854e-07,1.789861e-07,1.789868e-07,1.789875e-07,1.789882e-07,1.789889e-07,1.789896e-07,1.789903e-07,1.789910e-07,1.789917e-07,1.789924e-07,1.789931e-07,1.789938e-07,1.789945e-07,1.789952e-07,1.789960e-07,1.789967e-07,1.789974e-07,1.789981e-07,1.789988e-07,1.789995e-07,1.790002e-07,1.790009e-07,1.790016e-07,1.790023e-07,1.790030e-07,1.790037e-07,1.790044e-07,1.790051e-07,1.790058e-07,1.790065e-07,1.790072e-07,1.790079e-07,1.790086e-07,1.790093e-07,1.790100e-07,1.790107e-07,1.790114e-07,1.790121e-07,1.790129e-07,1.790136e-07,1.790143e-07,1.790150e-07,1.790157e-07,1.790164e-07,1.790171e-07,1.790178e-07,1.790185e-07,1.790192e-07,1.790199e-07,1.790206e-07,1.790213e-07,1.790220e-07,1.790227e-07,1.790234e-07,1.790241e-07,1.790248e-07,1.790255e-07,1.790262e-07,1.790269e-07,1.790276e-07,1.790283e-07,1.790290e-07,1.790297e-07,1.790304e-07,1.790311e-07,1.790318e-07,1.790325e-07,1.790332e-07,1.790339e-07,1.790346e-07,1.790353e-07,1.790360e-07,1.790367e-07,1.790375e-07,1.790382e-07,1.790389e-07,1.790396e-07,1.790403e-07,1.790410e-07,1.790417e-07,1.790424e-07,1.790431e-07,1.790438e-07,1.790445e-07,1.790452e-07,1.790459e-07,1.790466e-07,1.790473e-07,1.790480e-07,1.790487e-07,1.790494e-07,1.790501e-07,1.790508e-07,1.790515e-07,1.790522e-07,1.790529e-07,1.790536e-07,1.790543e-07,1.790550e-07,1.790557e-07,1.790564e-07,1.790571e-07,1.790578e-07,1.790585e-07,1.790592e-07,1.790599e-07,1.790606e-07,1.790613e-07,1.790620e-07,1.790627e-07,1.790634e-07,1.790641e-07,1.790648e-07,1.790655e-07,1.790662e-07,1.790669e-07,1.790676e-07,1.790683e-07,1.790690e-07,1.790697e-07,1.790704e-07,1.790711e-07,1.790718e-07,1.790725e-07,1.790732e-07,1.790739e-07,1.790746e-07,1.790753e-07,1.790760e-07,1.790767e-07,1.790774e-07,1.790781e-07,1.790788e-07,1.790795e-07,1.790802e-07,1.790809e-07,1.790816e-07,1.790823e-07,1.790830e-07,1.790837e-07,1.790844e-07,1.790851e-07,1.790858e-07,1.790865e-07,1.790872e-07,1.790879e-07,1.790886e-07,1.790893e-07,1.790900e-07,1.790907e-07,1.790914e-07,1.790921e-07,1.790928e-07,1.790935e-07,1.790942e-07,1.790949e-07,1.790956e-07,1.790963e-07,1.790970e-07,1.790977e-07,1.790984e-07,1.790991e-07,1.790998e-07,1.791005e-07,1.791012e-07,1.791019e-07,1.791026e-07,1.791033e-07,1.791040e-07,1.791047e-07,1.791054e-07,1.791061e-07,1.791068e-07,1.791074e-07,1.791081e-07,1.791088e-07,1.791095e-07,1.791102e-07,1.791109e-07,1.791116e-07,1.791123e-07,1.791130e-07,1.791137e-07,1.791144e-07,1.791151e-07,1.791158e-07,1.791165e-07,1.791172e-07,1.791179e-07,1.791186e-07,1.791193e-07,1.791200e-07,1.791207e-07,1.791214e-07,1.791221e-07,1.791228e-07,1.791235e-07,1.791242e-07,1.791249e-07,1.791256e-07,1.791263e-07,1.791270e-07,1.791277e-07,1.791284e-07,1.791291e-07,1.791298e-07,1.791305e-07,1.791312e-07,1.791318e-07,1.791325e-07,1.791332e-07,1.791339e-07,1.791346e-07,1.791353e-07,1.791360e-07,1.791367e-07,1.791374e-07,1.791381e-07,1.791388e-07,1.791395e-07,1.791402e-07,1.791409e-07,1.791416e-07,1.791423e-07,1.791430e-07,1.791437e-07,1.791444e-07,1.791451e-07,1.791458e-07,1.791465e-07,1.791472e-07,1.791479e-07,1.791486e-07,1.791492e-07,1.791499e-07,1.791506e-07,1.791513e-07,1.791520e-07,1.791527e-07,1.791534e-07,1.791541e-07,1.791548e-07,1.791555e-07,1.791562e-07,1.791569e-07,1.791576e-07,1.791583e-07,1.791590e-07,1.791597e-07,1.791604e-07,1.791611e-07,1.791618e-07,1.791625e-07,1.791631e-07,1.791638e-07,1.791645e-07,1.791652e-07,1.791659e-07,1.791666e-07,1.791673e-07,1.791680e-07,1.791687e-07,1.791694e-07,1.791701e-07,1.791708e-07,1.791715e-07,1.791722e-07,1.791729e-07,1.791736e-07,1.791743e-07,1.791749e-07,1.791756e-07,1.791763e-07,1.791770e-07,1.791777e-07,1.791784e-07,1.791791e-07,1.791798e-07,1.791805e-07,1.791812e-07,1.791819e-07,1.791826e-07,1.791833e-07,1.791840e-07,1.791847e-07,1.791854e-07,1.791860e-07,1.791867e-07,1.791874e-07,1.791881e-07,1.791888e-07,1.791895e-07,1.791902e-07,1.791909e-07,1.791916e-07,1.791923e-07,1.791930e-07,1.791937e-07,1.791944e-07,1.791951e-07,1.791957e-07,1.791964e-07,1.791971e-07,1.791978e-07,1.791985e-07,1.791992e-07,1.791999e-07,1.792006e-07,1.792013e-07,1.792020e-07,1.792027e-07,1.792034e-07,1.792041e-07,1.792047e-07,1.792054e-07,1.792061e-07,1.792068e-07,1.792075e-07,1.792082e-07,1.792089e-07,1.792096e-07,1.792103e-07,1.792110e-07,1.792117e-07,1.792124e-07,1.792130e-07,1.792137e-07,1.792144e-07,1.792151e-07,1.792158e-07,1.792165e-07,1.792172e-07,1.792179e-07,1.792186e-07,1.792193e-07,1.792200e-07,1.792207e-07,1.792213e-07,1.792220e-07,1.792227e-07,1.792234e-07,1.792241e-07,1.792248e-07,1.792255e-07,1.792262e-07,1.792269e-07,1.792276e-07,1.792283e-07,1.792289e-07,1.792296e-07,1.792303e-07,1.792310e-07,1.792317e-07,1.792324e-07,1.792331e-07,1.792338e-07,1.792345e-07,1.792352e-07,1.792358e-07,1.792365e-07,1.792372e-07,1.792379e-07,1.792386e-07,1.792393e-07,1.792400e-07,1.792407e-07,1.792414e-07,1.792421e-07,1.792427e-07,1.792434e-07,1.792441e-07,1.792448e-07,1.792455e-07,1.792462e-07,1.792469e-07,1.792476e-07,1.792483e-07,1.792490e-07,1.792496e-07,1.792503e-07,1.792510e-07,1.792517e-07,1.792524e-07,1.792531e-07,1.792538e-07,1.792545e-07,1.792552e-07,1.792558e-07,1.792565e-07,1.792572e-07,1.792579e-07,1.792586e-07,1.792593e-07,1.792600e-07,1.792607e-07,1.792614e-07,1.792620e-07,1.792627e-07,1.792634e-07,1.792641e-07,1.792648e-07,1.792655e-07,1.792662e-07,1.792669e-07,1.792676e-07,1.792682e-07,1.792689e-07,1.792696e-07,1.792703e-07,1.792710e-07,1.792717e-07,1.792724e-07,1.792731e-07,1.792737e-07,1.792744e-07,1.792751e-07,1.792758e-07,1.792765e-07,1.792772e-07,1.792779e-07,1.792786e-07,1.792793e-07,1.792799e-07,1.792806e-07,1.792813e-07,1.792820e-07,1.792827e-07,1.792834e-07,1.792841e-07,1.792848e-07,1.792854e-07,1.792861e-07,1.792868e-07,1.792875e-07,1.792882e-07,1.792889e-07,1.792896e-07,1.792902e-07,1.792909e-07,1.792916e-07,1.792923e-07,1.792930e-07,1.792937e-07,1.792944e-07,1.792951e-07,1.792957e-07,1.792964e-07,1.792971e-07,1.792978e-07,1.792985e-07,1.792992e-07,1.792999e-07,1.793006e-07,1.793012e-07,1.793019e-07,1.793026e-07,1.793033e-07,1.793040e-07,1.793047e-07,1.793054e-07,1.793060e-07,1.793067e-07,1.793074e-07,1.793081e-07,1.793088e-07,1.793095e-07,1.793102e-07,1.793108e-07,1.793115e-07,1.793122e-07,1.793129e-07,1.793136e-07,1.793143e-07,1.793150e-07,1.793156e-07,1.793163e-07,1.793170e-07,1.793177e-07,1.793184e-07,1.793191e-07,1.793198e-07,1.793204e-07,1.793211e-07,1.793218e-07,1.793225e-07,1.793232e-07,1.793239e-07,1.793246e-07,1.793252e-07,1.793259e-07,1.793266e-07,1.793273e-07,1.793280e-07,1.793287e-07,1.793293e-07,1.793300e-07,1.793307e-07,1.793314e-07,1.793321e-07,1.793328e-07,1.793335e-07,1.793341e-07,1.793348e-07,1.793355e-07,1.793362e-07,1.793369e-07,1.793376e-07,1.793382e-07,1.793389e-07,1.793396e-07,1.793403e-07,1.793410e-07,1.793417e-07,1.793423e-07,1.793430e-07,1.793437e-07,1.793444e-07,1.793451e-07,1.793458e-07,1.793465e-07,1.793471e-07,1.793478e-07,1.793485e-07,1.793492e-07,1.793499e-07,1.793506e-07,1.793512e-07,1.793519e-07,1.793526e-07,1.793533e-07,1.793540e-07,1.793547e-07,1.793553e-07,1.793560e-07,1.793567e-07,1.793574e-07,1.793581e-07,1.793588e-07,1.793594e-07,1.793601e-07,1.793608e-07,1.793615e-07,1.793622e-07,1.793628e-07,1.793635e-07,1.793642e-07,1.793649e-07,1.793656e-07,1.793663e-07,1.793669e-07,1.793676e-07,1.793683e-07,1.793690e-07,1.793697e-07,1.793704e-07,1.793710e-07,1.793717e-07,1.793724e-07,1.793731e-07,1.793738e-07,1.793744e-07,1.793751e-07,1.793758e-07,1.793765e-07,1.793772e-07,1.793779e-07,1.793785e-07,1.793792e-07,1.793799e-07,1.793806e-07,1.793813e-07,1.793819e-07,1.793826e-07,1.793833e-07,1.793840e-07,1.793847e-07,1.793854e-07,1.793860e-07,1.793867e-07,1.793874e-07,1.793881e-07,1.793888e-07,1.793894e-07,1.793901e-07,1.793908e-07,1.793915e-07,1.793922e-07,1.793929e-07,1.793935e-07,1.793942e-07,1.793949e-07,1.793956e-07,1.793963e-07,1.793969e-07,1.793976e-07,1.793983e-07,1.793990e-07,1.793997e-07,1.794003e-07,1.794010e-07,1.794017e-07,1.794024e-07,1.794031e-07,1.794037e-07,1.794044e-07,1.794051e-07,1.794058e-07,1.794065e-07,1.794071e-07,1.794078e-07,1.794085e-07,1.794092e-07,1.794099e-07,1.794105e-07,1.794112e-07,1.794119e-07,1.794126e-07,1.794133e-07,1.794139e-07,1.794146e-07,1.794153e-07,1.794160e-07,1.794167e-07,1.794173e-07,1.794180e-07,1.794187e-07,1.794194e-07,1.794201e-07,1.794207e-07,1.794214e-07,1.794221e-07,1.794228e-07,1.794235e-07,1.794241e-07,1.794248e-07,1.794255e-07,1.794262e-07,1.794269e-07,1.794275e-07,1.794282e-07,1.794289e-07,1.794296e-07,1.794302e-07,1.794309e-07,1.794316e-07,1.794323e-07,1.794330e-07,1.794336e-07,1.794343e-07,1.794350e-07,1.794357e-07,1.794364e-07,1.794370e-07,1.794377e-07,1.794384e-07,1.794391e-07,1.794397e-07,1.794404e-07,1.794411e-07,1.794418e-07,1.794425e-07,1.794431e-07,1.794438e-07,1.794445e-07,1.794452e-07,1.794458e-07,1.794465e-07,1.794472e-07,1.794479e-07,1.794486e-07,1.794492e-07,1.794499e-07,1.794506e-07,1.794513e-07,1.794519e-07,1.794526e-07,1.794533e-07,1.794540e-07,1.794547e-07,1.794553e-07,1.794560e-07,1.794567e-07,1.794574e-07,1.794580e-07,1.794587e-07,1.794594e-07,1.794601e-07,1.794608e-07,1.794614e-07,1.794621e-07,1.794628e-07,1.794635e-07,1.794641e-07,1.794648e-07,1.794655e-07,1.794662e-07,1.794668e-07,1.794675e-07,1.794682e-07,1.794689e-07,1.794696e-07,1.794702e-07,1.794709e-07,1.794716e-07,1.794723e-07,1.794729e-07,1.794736e-07,1.794743e-07,1.794750e-07,1.794756e-07,1.794763e-07,1.794770e-07,1.794777e-07,1.794783e-07,1.794790e-07,1.794797e-07,1.794804e-07,1.794810e-07,1.794817e-07,1.794824e-07,1.794831e-07,1.794837e-07,1.794844e-07,1.794851e-07,1.794858e-07,1.794865e-07,1.794871e-07,1.794878e-07,1.794885e-07,1.794892e-07,1.794898e-07,1.794905e-07,1.794912e-07,1.794919e-07,1.794925e-07,1.794932e-07,1.794939e-07,1.794946e-07,1.794952e-07,1.794959e-07,1.794966e-07,1.794973e-07,1.794979e-07,1.794986e-07,1.794993e-07,1.795000e-07,1.795006e-07,1.795013e-07,1.795020e-07,1.795027e-07,1.795033e-07,1.795040e-07,1.795047e-07,1.795054e-07,1.795060e-07,1.795067e-07,1.795074e-07,1.795080e-07,1.795087e-07,1.795094e-07,1.795101e-07,1.795107e-07,1.795114e-07,1.795121e-07,1.795128e-07,1.795134e-07,1.795141e-07,1.795148e-07,1.795155e-07,1.795161e-07,1.795168e-07,1.795175e-07,1.795182e-07,1.795188e-07,1.795195e-07,1.795202e-07,1.795209e-07,1.795215e-07,1.795222e-07,1.795229e-07,1.795235e-07,1.795242e-07,1.795249e-07,1.795256e-07,1.795262e-07,1.795269e-07,1.795276e-07,1.795283e-07,1.795289e-07,1.795296e-07,1.795303e-07,1.795310e-07,1.795316e-07,1.795323e-07,1.795330e-07,1.795336e-07,1.795343e-07,1.795350e-07,1.795357e-07,1.795363e-07,1.795370e-07,1.795377e-07,1.795384e-07,1.795390e-07,1.795397e-07,1.795404e-07,1.795410e-07,1.795417e-07,1.795424e-07,1.795431e-07,1.795437e-07,1.795444e-07,1.795451e-07,1.795457e-07,1.795464e-07,1.795471e-07,1.795478e-07,1.795484e-07,1.795491e-07,1.795498e-07,1.795505e-07,1.795511e-07,1.795518e-07,1.795525e-07,1.795531e-07,1.795538e-07,1.795545e-07,1.795552e-07,1.795558e-07,1.795565e-07,1.795572e-07,1.795578e-07,1.795585e-07,1.795592e-07,1.795599e-07,1.795605e-07,1.795612e-07,1.795619e-07,1.795625e-07,1.795632e-07,1.795639e-07,1.795646e-07,1.795652e-07,1.795659e-07,1.795666e-07,1.795672e-07,1.795679e-07,1.795686e-07,1.795693e-07,1.795699e-07,1.795706e-07,1.795713e-07,1.795719e-07,1.795726e-07,1.795733e-07,1.795739e-07,1.795746e-07,1.795753e-07,1.795760e-07,1.795766e-07,1.795773e-07,1.795780e-07,1.795786e-07,1.795793e-07,1.795800e-07,1.795806e-07,1.795813e-07,1.795820e-07,1.795827e-07,1.795833e-07,1.795840e-07,1.795847e-07,1.795853e-07,1.795860e-07,1.795867e-07,1.795873e-07,1.795880e-07,1.795887e-07,1.795894e-07,1.795900e-07,1.795907e-07,1.795914e-07,1.795920e-07,1.795927e-07,1.795934e-07,1.795940e-07,1.795947e-07,1.795954e-07,1.795961e-07,1.795967e-07,1.795974e-07,1.795981e-07,1.795987e-07,1.795994e-07,1.796001e-07,1.796007e-07,1.796014e-07,1.796021e-07,1.796027e-07,1.796034e-07,1.796041e-07,1.796047e-07,1.796054e-07,1.796061e-07,1.796068e-07,1.796074e-07,1.796081e-07,1.796088e-07,1.796094e-07,1.796101e-07,1.796108e-07,1.796114e-07,1.796121e-07,1.796128e-07,1.796134e-07,1.796141e-07,1.796148e-07,1.796154e-07,1.796161e-07,1.796168e-07,1.796174e-07,1.796181e-07,1.796188e-07,1.796195e-07,1.796201e-07,1.796208e-07,1.796215e-07,1.796221e-07,1.796228e-07,1.796235e-07,1.796241e-07,1.796248e-07,1.796255e-07,1.796261e-07,1.796268e-07,1.796275e-07,1.796281e-07,1.796288e-07,1.796295e-07,1.796301e-07,1.796308e-07,1.796315e-07,1.796321e-07,1.796328e-07,1.796335e-07,1.796341e-07,1.796348e-07,1.796355e-07,1.796361e-07,1.796368e-07,1.796375e-07,1.796381e-07,1.796388e-07,1.796395e-07,1.796401e-07,1.796408e-07,1.796415e-07,1.796421e-07,1.796428e-07,1.796435e-07,1.796441e-07,1.796448e-07,1.796455e-07,1.796461e-07,1.796468e-07,1.796475e-07,1.796481e-07,1.796488e-07,1.796495e-07,1.796501e-07,1.796508e-07,1.796515e-07,1.796521e-07,1.796528e-07,1.796535e-07,1.796541e-07,1.796548e-07,1.796555e-07,1.796561e-07,1.796568e-07,1.796575e-07,1.796581e-07,1.796588e-07,1.796595e-07,1.796601e-07,1.796608e-07,1.796615e-07,1.796621e-07,1.796628e-07,1.796634e-07,1.796641e-07,1.796648e-07,1.796654e-07,1.796661e-07,1.796668e-07,1.796674e-07,1.796681e-07,1.796688e-07,1.796694e-07,1.796701e-07,1.796708e-07,1.796714e-07,1.796721e-07,1.796728e-07,1.796734e-07,1.796741e-07,1.796748e-07,1.796754e-07,1.796761e-07,1.796767e-07,1.796774e-07,1.796781e-07,1.796787e-07,1.796794e-07,1.796801e-07,1.796807e-07,1.796814e-07,1.796821e-07,1.796827e-07,1.796834e-07,1.796841e-07,1.796847e-07,1.796854e-07,1.796860e-07,1.796867e-07,1.796874e-07,1.796880e-07,1.796887e-07,1.796894e-07,1.796900e-07,1.796907e-07,1.796914e-07,1.796920e-07,1.796927e-07,1.796934e-07,1.796940e-07,1.796947e-07,1.796953e-07,1.796960e-07,1.796967e-07,1.796973e-07,1.796980e-07,1.796987e-07,1.796993e-07,1.797000e-07,1.797006e-07,1.797013e-07,1.797020e-07,1.797026e-07,1.797033e-07,1.797040e-07,1.797046e-07,1.797053e-07,1.797060e-07,1.797066e-07,1.797073e-07,1.797079e-07,1.797086e-07,1.797093e-07,1.797099e-07,1.797106e-07,1.797113e-07,1.797119e-07,1.797126e-07,1.797132e-07,1.797139e-07,1.797146e-07,1.797152e-07,1.797159e-07,1.797166e-07,1.797172e-07,1.797179e-07,1.797185e-07,1.797192e-07,1.797199e-07,1.797205e-07,1.797212e-07,1.797219e-07,1.797225e-07,1.797232e-07,1.797238e-07,1.797245e-07,1.797252e-07,1.797258e-07,1.797265e-07,1.797271e-07,1.797278e-07,1.797285e-07,1.797291e-07,1.797298e-07,1.797305e-07,1.797311e-07,1.797318e-07,1.797324e-07,1.797331e-07,1.797338e-07,1.797344e-07,1.797351e-07,1.797357e-07,1.797364e-07,1.797371e-07,1.797377e-07,1.797384e-07,1.797391e-07,1.797397e-07,1.797404e-07,1.797410e-07,1.797417e-07,1.797424e-07,1.797430e-07,1.797437e-07,1.797443e-07,1.797450e-07,1.797457e-07,1.797463e-07,1.797470e-07,1.797476e-07,1.797483e-07,1.797490e-07,1.797496e-07,1.797503e-07,1.797509e-07,1.797516e-07,1.797523e-07,1.797529e-07,1.797536e-07,1.797542e-07,1.797549e-07,1.797556e-07,1.797562e-07,1.797569e-07,1.797576e-07,1.797582e-07,1.797589e-07,1.797595e-07,1.797602e-07,1.797609e-07,1.797615e-07,1.797622e-07,1.797628e-07,1.797635e-07,1.797641e-07,1.797648e-07,1.797655e-07,1.797661e-07,1.797668e-07,1.797674e-07,1.797681e-07,1.797688e-07,1.797694e-07,1.797701e-07,1.797707e-07,1.797714e-07,1.797721e-07,1.797727e-07,1.797734e-07,1.797740e-07,1.797747e-07,1.797754e-07,1.797760e-07,1.797767e-07,1.797773e-07,1.797780e-07,1.797787e-07,1.797793e-07,1.797800e-07,1.797806e-07,1.797813e-07,1.797819e-07,1.797826e-07,1.797833e-07,1.797839e-07,1.797846e-07,1.797852e-07,1.797859e-07,1.797866e-07,1.797872e-07,1.797879e-07,1.797885e-07,1.797892e-07,1.797898e-07,1.797905e-07,1.797912e-07,1.797918e-07,1.797925e-07,1.797931e-07,1.797938e-07,1.797945e-07,1.797951e-07,1.797958e-07,1.797964e-07,1.797971e-07,1.797977e-07,1.797984e-07,1.797991e-07,1.797997e-07,1.798004e-07,1.798010e-07,1.798017e-07,1.798023e-07,1.798030e-07,1.798037e-07,1.798043e-07,1.798050e-07,1.798056e-07,1.798063e-07,1.798069e-07,1.798076e-07,1.798083e-07,1.798089e-07,1.798096e-07,1.798102e-07,1.798109e-07,1.798115e-07,1.798122e-07,1.798129e-07,1.798135e-07,1.798142e-07,1.798148e-07,1.798155e-07,1.798161e-07,1.798168e-07,1.798175e-07,1.798181e-07,1.798188e-07,1.798194e-07,1.798201e-07,1.798207e-07,1.798214e-07,1.798221e-07,1.798227e-07,1.798234e-07,1.798240e-07,1.798247e-07,1.798253e-07,1.798260e-07,1.798266e-07,1.798273e-07,1.798280e-07,1.798286e-07,1.798293e-07,1.798299e-07,1.798306e-07,1.798312e-07,1.798319e-07,1.798326e-07,1.798332e-07,1.798339e-07,1.798345e-07,1.798352e-07,1.798358e-07,1.798365e-07,1.798371e-07,1.798378e-07,1.798385e-07,1.798391e-07,1.798398e-07,1.798404e-07,1.798411e-07,1.798417e-07,1.798424e-07,1.798430e-07,1.798437e-07,1.798443e-07,1.798450e-07,1.798457e-07,1.798463e-07,1.798470e-07,1.798476e-07,1.798483e-07,1.798489e-07,1.798496e-07,1.798502e-07,1.798509e-07,1.798516e-07,1.798522e-07,1.798529e-07,1.798535e-07,1.798542e-07,1.798548e-07,1.798555e-07,1.798561e-07,1.798568e-07,1.798574e-07,1.798581e-07,1.798588e-07,1.798594e-07,1.798601e-07,1.798607e-07,1.798614e-07,1.798620e-07,1.798627e-07,1.798633e-07,1.798640e-07,1.798646e-07,1.798653e-07,1.798659e-07,1.798666e-07,1.798673e-07,1.798679e-07,1.798686e-07,1.798692e-07,1.798699e-07,1.798705e-07,1.798712e-07,1.798718e-07,1.798725e-07,1.798731e-07,1.798738e-07,1.798744e-07,1.798751e-07,1.798758e-07,1.798764e-07,1.798771e-07,1.798777e-07,1.798784e-07,1.798790e-07,1.798797e-07,1.798803e-07,1.798810e-07,1.798816e-07,1.798823e-07,1.798829e-07,1.798836e-07,1.798842e-07,1.798849e-07,1.798855e-07,1.798862e-07,1.798869e-07,1.798875e-07,1.798882e-07,1.798888e-07,1.798895e-07,1.798901e-07,1.798908e-07,1.798914e-07,1.798921e-07,1.798927e-07,1.798934e-07,1.798940e-07,1.798947e-07,1.798953e-07,1.798960e-07,1.798966e-07,1.798973e-07,1.798979e-07,1.798986e-07,1.798993e-07,1.798999e-07,1.799006e-07,1.799012e-07,1.799019e-07,1.799025e-07,1.799032e-07,1.799038e-07,1.799045e-07,1.799051e-07,1.799058e-07,1.799064e-07,1.799071e-07,1.799077e-07,1.799084e-07,1.799090e-07,1.799097e-07,1.799103e-07,1.799110e-07,1.799116e-07,1.799123e-07,1.799129e-07,1.799136e-07,1.799142e-07,1.799149e-07,1.799155e-07,1.799162e-07,1.799168e-07,1.799175e-07,1.799181e-07,1.799188e-07,1.799194e-07,1.799201e-07,1.799207e-07,1.799214e-07,1.799221e-07,1.799227e-07,1.799234e-07,1.799240e-07,1.799247e-07,1.799253e-07,1.799260e-07,1.799266e-07,1.799273e-07,1.799279e-07,1.799286e-07,1.799292e-07,1.799299e-07,1.799305e-07,1.799312e-07,1.799318e-07,1.799325e-07,1.799331e-07,1.799338e-07,1.799344e-07,1.799351e-07,1.799357e-07,1.799364e-07,1.799370e-07,1.799377e-07,1.799383e-07,1.799390e-07,1.799396e-07,1.799403e-07,1.799409e-07,1.799416e-07,1.799422e-07,1.799429e-07,1.799435e-07,1.799442e-07,1.799448e-07,1.799455e-07,1.799461e-07,1.799468e-07,1.799474e-07,1.799481e-07,1.799487e-07,1.799494e-07,1.799500e-07,1.799506e-07,1.799513e-07,1.799519e-07,1.799526e-07,1.799532e-07,1.799539e-07,1.799545e-07,1.799552e-07,1.799558e-07,1.799565e-07,1.799571e-07,1.799578e-07,1.799584e-07,1.799591e-07,1.799597e-07,1.799604e-07,1.799610e-07,1.799617e-07,1.799623e-07,1.799630e-07,1.799636e-07,1.799643e-07,1.799649e-07,1.799656e-07,1.799662e-07,1.799669e-07,1.799675e-07,1.799682e-07,1.799688e-07,1.799695e-07,1.799701e-07,1.799708e-07,1.799714e-07,1.799721e-07,1.799727e-07,1.799733e-07,1.799740e-07,1.799746e-07,1.799753e-07,1.799759e-07,1.799766e-07,1.799772e-07,1.799779e-07,1.799785e-07,1.799792e-07,1.799798e-07,1.799805e-07,1.799811e-07,1.799818e-07,1.799824e-07,1.799831e-07,1.799837e-07,1.799844e-07,1.799850e-07,1.799857e-07,1.799863e-07,1.799869e-07,1.799876e-07,1.799882e-07,1.799889e-07,1.799895e-07,1.799902e-07,1.799908e-07,1.799915e-07,1.799921e-07,1.799928e-07,1.799934e-07,1.799941e-07,1.799947e-07,1.799954e-07,1.799960e-07,1.799967e-07,1.799973e-07,1.799979e-07,1.799986e-07,1.799992e-07,1.799999e-07,1.800005e-07,1.800012e-07,1.800018e-07,1.800025e-07,1.800031e-07,1.800038e-07,1.800044e-07,1.800051e-07,1.800057e-07,1.800063e-07,1.800070e-07,1.800076e-07,1.800083e-07,1.800089e-07,1.800096e-07,1.800102e-07,1.800109e-07,1.800115e-07,1.800122e-07,1.800128e-07,1.800135e-07,1.800141e-07,1.800147e-07,1.800154e-07,1.800160e-07,1.800167e-07,1.800173e-07,1.800180e-07,1.800186e-07,1.800193e-07,1.800199e-07,1.800206e-07,1.800212e-07,1.800218e-07,1.800225e-07,1.800231e-07,1.800238e-07,1.800244e-07,1.800251e-07,1.800257e-07,1.800264e-07,1.800270e-07,1.800276e-07,1.800283e-07,1.800289e-07,1.800296e-07,1.800302e-07,1.800309e-07,1.800315e-07,1.800322e-07,1.800328e-07,1.800334e-07,1.800341e-07,1.800347e-07,1.800354e-07,1.800360e-07,1.800367e-07,1.800373e-07,1.800380e-07,1.800386e-07,1.800392e-07,1.800399e-07,1.800405e-07,1.800412e-07,1.800418e-07,1.800425e-07,1.800431e-07,1.800438e-07,1.800444e-07,1.800450e-07,1.800457e-07,1.800463e-07,1.800470e-07,1.800476e-07,1.800483e-07,1.800489e-07,1.800496e-07,1.800502e-07,1.800508e-07,1.800515e-07,1.800521e-07,1.800528e-07,1.800534e-07,1.800541e-07,1.800547e-07,1.800553e-07,1.800560e-07,1.800566e-07,1.800573e-07,1.800579e-07,1.800586e-07,1.800592e-07,1.800598e-07,1.800605e-07,1.800611e-07,1.800618e-07,1.800624e-07,1.800631e-07,1.800637e-07,1.800643e-07,1.800650e-07,1.800656e-07,1.800663e-07,1.800669e-07,1.800676e-07,1.800682e-07,1.800688e-07,1.800695e-07,1.800701e-07,1.800708e-07,1.800714e-07,1.800721e-07,1.800727e-07,1.800733e-07,1.800740e-07,1.800746e-07,1.800753e-07,1.800759e-07,1.800766e-07,1.800772e-07,1.800778e-07,1.800785e-07,1.800791e-07,1.800798e-07,1.800804e-07,1.800811e-07,1.800817e-07,1.800823e-07,1.800830e-07,1.800836e-07,1.800843e-07,1.800849e-07,1.800855e-07,1.800862e-07,1.800868e-07,1.800875e-07,1.800881e-07,1.800888e-07,1.800894e-07,1.800900e-07,1.800907e-07,1.800913e-07,1.800920e-07,1.800926e-07,1.800932e-07,1.800939e-07,1.800945e-07,1.800952e-07,1.800958e-07,1.800964e-07,1.800971e-07,1.800977e-07,1.800984e-07,1.800990e-07,1.800997e-07,1.801003e-07,1.801009e-07,1.801016e-07,1.801022e-07,1.801029e-07,1.801035e-07,1.801041e-07,1.801048e-07,1.801054e-07,1.801061e-07,1.801067e-07,1.801073e-07,1.801080e-07,1.801086e-07,1.801093e-07,1.801099e-07,1.801105e-07,1.801112e-07,1.801118e-07,1.801125e-07,1.801131e-07,1.801137e-07,1.801144e-07,1.801150e-07,1.801157e-07,1.801163e-07,1.801169e-07,1.801176e-07,1.801182e-07,1.801189e-07,1.801195e-07,1.801201e-07,1.801208e-07,1.801214e-07,1.801221e-07,1.801227e-07,1.801233e-07,1.801240e-07,1.801246e-07,1.801253e-07,1.801259e-07,1.801265e-07,1.801272e-07,1.801278e-07,1.801285e-07,1.801291e-07,1.801297e-07,1.801304e-07,1.801310e-07,1.801317e-07,1.801323e-07,1.801329e-07,1.801336e-07,1.801342e-07,1.801349e-07,1.801355e-07,1.801361e-07,1.801368e-07,1.801374e-07,1.801380e-07,1.801387e-07,1.801393e-07,1.801400e-07,1.801406e-07,1.801412e-07,1.801419e-07,1.801425e-07,1.801432e-07,1.801438e-07,1.801444e-07,1.801451e-07,1.801457e-07,1.801463e-07,1.801470e-07,1.801476e-07,1.801483e-07,1.801489e-07,1.801495e-07,1.801502e-07,1.801508e-07,1.801515e-07,1.801521e-07,1.801527e-07,1.801534e-07,1.801540e-07,1.801546e-07,1.801553e-07,1.801559e-07,1.801566e-07,1.801572e-07,1.801578e-07,1.801585e-07,1.801591e-07,1.801597e-07,1.801604e-07,1.801610e-07,1.801617e-07,1.801623e-07,1.801629e-07,1.801636e-07,1.801642e-07,1.801648e-07,1.801655e-07,1.801661e-07,1.801668e-07,1.801674e-07,1.801680e-07,1.801687e-07,1.801693e-07,1.801699e-07,1.801706e-07,1.801712e-07,1.801719e-07,1.801725e-07,1.801731e-07,1.801738e-07,1.801744e-07,1.801750e-07,1.801757e-07,1.801763e-07,1.801769e-07,1.801776e-07,1.801782e-07,1.801789e-07,1.801795e-07,1.801801e-07,1.801808e-07,1.801814e-07,1.801820e-07,1.801827e-07,1.801833e-07,1.801840e-07,1.801846e-07,1.801852e-07,1.801859e-07,1.801865e-07,1.801871e-07,1.801878e-07,1.801884e-07,1.801890e-07,1.801897e-07,1.801903e-07,1.801909e-07,1.801916e-07,1.801922e-07,1.801929e-07,1.801935e-07,1.801941e-07,1.801948e-07,1.801954e-07,1.801960e-07,1.801967e-07,1.801973e-07,1.801979e-07,1.801986e-07,1.801992e-07,1.801998e-07,1.802005e-07,1.802011e-07,1.802018e-07,1.802024e-07,1.802030e-07,1.802037e-07,1.802043e-07,1.802049e-07,1.802056e-07,1.802062e-07,1.802068e-07,1.802075e-07,1.802081e-07,1.802087e-07,1.802094e-07,1.802100e-07,1.802106e-07,1.802113e-07,1.802119e-07,1.802126e-07,1.802132e-07,1.802138e-07,1.802145e-07,1.802151e-07,1.802157e-07,1.802164e-07,1.802170e-07,1.802176e-07,1.802183e-07,1.802189e-07,1.802195e-07,1.802202e-07,1.802208e-07,1.802214e-07,1.802221e-07,1.802227e-07,1.802233e-07,1.802240e-07,1.802246e-07,1.802252e-07,1.802259e-07,1.802265e-07,1.802271e-07,1.802278e-07,1.802284e-07,1.802290e-07,1.802297e-07,1.802303e-07,1.802309e-07,1.802316e-07,1.802322e-07,1.802328e-07,1.802335e-07,1.802341e-07,1.802347e-07,1.802354e-07,1.802360e-07,1.802366e-07,1.802373e-07,1.802379e-07,1.802385e-07,1.802392e-07,1.802398e-07,1.802404e-07,1.802411e-07,1.802417e-07,1.802423e-07,1.802430e-07,1.802436e-07,1.802442e-07,1.802449e-07,1.802455e-07,1.802461e-07,1.802468e-07,1.802474e-07,1.802480e-07,1.802487e-07,1.802493e-07,1.802499e-07,1.802506e-07,1.802512e-07,1.802518e-07,1.802525e-07,1.802531e-07,1.802537e-07,1.802544e-07,1.802550e-07,1.802556e-07,1.802563e-07,1.802569e-07,1.802575e-07,1.802582e-07,1.802588e-07,1.802594e-07,1.802601e-07,1.802607e-07,1.802613e-07,1.802620e-07,1.802626e-07,1.802632e-07,1.802639e-07,1.802645e-07,1.802651e-07,1.802657e-07,1.802664e-07,1.802670e-07,1.802676e-07,1.802683e-07,1.802689e-07,1.802695e-07,1.802702e-07,1.802708e-07,1.802714e-07,1.802721e-07,1.802727e-07,1.802733e-07,1.802740e-07,1.802746e-07,1.802752e-07,1.802759e-07,1.802765e-07,1.802771e-07,1.802777e-07,1.802784e-07,1.802790e-07,1.802796e-07,1.802803e-07,1.802809e-07,1.802815e-07,1.802822e-07,1.802828e-07,1.802834e-07,1.802841e-07,1.802847e-07,1.802853e-07,1.802860e-07,1.802866e-07,1.802872e-07,1.802878e-07,1.802885e-07,1.802891e-07,1.802897e-07,1.802904e-07,1.802910e-07,1.802916e-07,1.802923e-07,1.802929e-07,1.802935e-07,1.802941e-07,1.802948e-07,1.802954e-07,1.802960e-07,1.802967e-07,1.802973e-07,1.802979e-07,1.802986e-07,1.802992e-07,1.802998e-07,1.803004e-07,1.803011e-07,1.803017e-07,1.803023e-07,1.803030e-07,1.803036e-07,1.803042e-07,1.803049e-07,1.803055e-07,1.803061e-07,1.803067e-07,1.803074e-07,1.803080e-07,1.803086e-07,1.803093e-07,1.803099e-07,1.803105e-07,1.803112e-07,1.803118e-07,1.803124e-07,1.803130e-07,1.803137e-07,1.803143e-07,1.803149e-07,1.803156e-07,1.803162e-07,1.803168e-07,1.803174e-07,1.803181e-07,1.803187e-07,1.803193e-07,1.803200e-07,1.803206e-07,1.803212e-07,1.803218e-07,1.803225e-07,1.803231e-07,1.803237e-07,1.803244e-07,1.803250e-07,1.803256e-07,1.803263e-07,1.803269e-07,1.803275e-07,1.803281e-07,1.803288e-07,1.803294e-07,1.803300e-07,1.803306e-07,1.803313e-07,1.803319e-07,1.803325e-07,1.803332e-07,1.803338e-07,1.803344e-07,1.803350e-07,1.803357e-07,1.803363e-07,1.803369e-07,1.803376e-07,1.803382e-07,1.803388e-07,1.803394e-07,1.803401e-07,1.803407e-07,1.803413e-07,1.803420e-07,1.803426e-07,1.803432e-07,1.803438e-07,1.803445e-07,1.803451e-07,1.803457e-07,1.803463e-07,1.803470e-07,1.803476e-07,1.803482e-07,1.803489e-07,1.803495e-07,1.803501e-07,1.803507e-07,1.803514e-07,1.803520e-07,1.803526e-07,1.803532e-07,1.803539e-07,1.803545e-07,1.803551e-07,1.803558e-07,1.803564e-07,1.803570e-07,1.803576e-07,1.803583e-07,1.803589e-07,1.803595e-07,1.803601e-07,1.803608e-07,1.803614e-07,1.803620e-07,1.803627e-07,1.803633e-07,1.803639e-07,1.803645e-07,1.803652e-07,1.803658e-07,1.803664e-07,1.803670e-07,1.803677e-07,1.803683e-07,1.803689e-07,1.803695e-07,1.803702e-07,1.803708e-07,1.803714e-07,1.803720e-07,1.803727e-07,1.803733e-07,1.803739e-07,1.803746e-07,1.803752e-07,1.803758e-07,1.803764e-07,1.803771e-07,1.803777e-07,1.803783e-07,1.803789e-07,1.803796e-07,1.803802e-07,1.803808e-07,1.803814e-07,1.803821e-07,1.803827e-07,1.803833e-07,1.803839e-07,1.803846e-07,1.803852e-07,1.803858e-07,1.803864e-07,1.803871e-07,1.803877e-07,1.803883e-07,1.803889e-07,1.803896e-07,1.803902e-07,1.803908e-07,1.803914e-07,1.803921e-07,1.803927e-07,1.803933e-07,1.803939e-07,1.803946e-07,1.803952e-07,1.803958e-07,1.803964e-07,1.803971e-07,1.803977e-07,1.803983e-07,1.803989e-07,1.803996e-07,1.804002e-07,1.804008e-07,1.804014e-07,1.804021e-07,1.804027e-07,1.804033e-07,1.804039e-07,1.804046e-07,1.804052e-07,1.804058e-07,1.804064e-07,1.804071e-07,1.804077e-07,1.804083e-07,1.804089e-07,1.804096e-07,1.804102e-07,1.804108e-07,1.804114e-07,1.804121e-07,1.804127e-07,1.804133e-07,1.804139e-07,1.804145e-07,1.804152e-07,1.804158e-07,1.804164e-07,1.804170e-07,1.804177e-07,1.804183e-07,1.804189e-07,1.804195e-07,1.804202e-07,1.804208e-07,1.804214e-07,1.804220e-07,1.804227e-07,1.804233e-07,1.804239e-07,1.804245e-07,1.804251e-07,1.804258e-07,1.804264e-07,1.804270e-07,1.804276e-07,1.804283e-07,1.804289e-07,1.804295e-07,1.804301e-07,1.804308e-07,1.804314e-07,1.804320e-07,1.804326e-07,1.804332e-07,1.804339e-07,1.804345e-07,1.804351e-07,1.804357e-07,1.804364e-07,1.804370e-07,1.804376e-07,1.804382e-07,1.804389e-07,1.804395e-07,1.804401e-07,1.804407e-07,1.804413e-07,1.804420e-07,1.804426e-07,1.804432e-07,1.804438e-07,1.804445e-07,1.804451e-07,1.804457e-07,1.804463e-07,1.804469e-07,1.804476e-07,1.804482e-07,1.804488e-07,1.804494e-07,1.804501e-07,1.804507e-07,1.804513e-07,1.804519e-07,1.804525e-07,1.804532e-07,1.804538e-07,1.804544e-07,1.804550e-07,1.804556e-07,1.804563e-07,1.804569e-07,1.804575e-07,1.804581e-07,1.804588e-07,1.804594e-07,1.804600e-07,1.804606e-07,1.804612e-07,1.804619e-07,1.804625e-07,1.804631e-07,1.804637e-07,1.804643e-07,1.804650e-07,1.804656e-07,1.804662e-07,1.804668e-07,1.804675e-07,1.804681e-07,1.804687e-07,1.804693e-07,1.804699e-07,1.804706e-07,1.804712e-07,1.804718e-07,1.804724e-07,1.804730e-07,1.804737e-07,1.804743e-07,1.804749e-07,1.804755e-07,1.804761e-07,1.804768e-07,1.804774e-07,1.804780e-07,1.804786e-07,1.804792e-07,1.804799e-07,1.804805e-07,1.804811e-07,1.804817e-07,1.804823e-07,1.804830e-07,1.804836e-07,1.804842e-07,1.804848e-07,1.804855e-07,1.804861e-07,1.804867e-07,1.804873e-07,1.804879e-07,1.804886e-07,1.804892e-07,1.804898e-07,1.804904e-07,1.804910e-07,1.804916e-07,1.804923e-07,1.804929e-07,1.804935e-07,1.804941e-07,1.804947e-07,1.804954e-07,1.804960e-07,1.804966e-07,1.804972e-07,1.804978e-07,1.804985e-07,1.804991e-07,1.804997e-07,1.805003e-07,1.805009e-07,1.805016e-07,1.805022e-07,1.805028e-07,1.805034e-07,1.805040e-07,1.805047e-07,1.805053e-07,1.805059e-07,1.805065e-07,1.805071e-07,1.805078e-07,1.805084e-07,1.805090e-07,1.805096e-07,1.805102e-07,1.805108e-07,1.805115e-07,1.805121e-07,1.805127e-07,1.805133e-07,1.805139e-07,1.805146e-07,1.805152e-07,1.805158e-07,1.805164e-07,1.805170e-07,1.805176e-07,1.805183e-07,1.805189e-07,1.805195e-07,1.805201e-07,1.805207e-07,1.805214e-07,1.805220e-07,1.805226e-07,1.805232e-07,1.805238e-07,1.805244e-07,1.805251e-07,1.805257e-07,1.805263e-07,1.805269e-07,1.805275e-07,1.805282e-07,1.805288e-07,1.805294e-07,1.805300e-07,1.805306e-07,1.805312e-07,1.805319e-07,1.805325e-07,1.805331e-07,1.805337e-07,1.805343e-07,1.805350e-07,1.805356e-07,1.805362e-07,1.805368e-07,1.805374e-07,1.805380e-07,1.805387e-07,1.805393e-07,1.805399e-07,1.805405e-07,1.805411e-07,1.805417e-07,1.805424e-07,1.805430e-07,1.805436e-07,1.805442e-07,1.805448e-07,1.805454e-07,1.805461e-07,1.805467e-07,1.805473e-07,1.805479e-07,1.805485e-07,1.805491e-07,1.805498e-07,1.805504e-07,1.805510e-07,1.805516e-07,1.805522e-07,1.805528e-07,1.805535e-07,1.805541e-07,1.805547e-07,1.805553e-07,1.805559e-07,1.805565e-07,1.805572e-07,1.805578e-07,1.805584e-07,1.805590e-07,1.805596e-07,1.805602e-07,1.805609e-07,1.805615e-07,1.805621e-07,1.805627e-07,1.805633e-07,1.805639e-07,1.805646e-07,1.805652e-07,1.805658e-07,1.805664e-07,1.805670e-07,1.805676e-07,1.805682e-07,1.805689e-07,1.805695e-07,1.805701e-07,1.805707e-07,1.805713e-07,1.805719e-07,1.805726e-07,1.805732e-07,1.805738e-07,1.805744e-07,1.805750e-07,1.805756e-07,1.805762e-07,1.805769e-07,1.805775e-07,1.805781e-07,1.805787e-07,1.805793e-07,1.805799e-07,1.805806e-07,1.805812e-07,1.805818e-07,1.805824e-07,1.805830e-07,1.805836e-07,1.805842e-07,1.805849e-07,1.805855e-07,1.805861e-07,1.805867e-07,1.805873e-07,1.805879e-07,1.805885e-07,1.805892e-07,1.805898e-07,1.805904e-07,1.805910e-07,1.805916e-07,1.805922e-07,1.805928e-07,1.805935e-07,1.805941e-07,1.805947e-07,1.805953e-07,1.805959e-07,1.805965e-07,1.805971e-07,1.805978e-07,1.805984e-07,1.805990e-07,1.805996e-07,1.806002e-07,1.806008e-07,1.806014e-07,1.806021e-07,1.806027e-07,1.806033e-07,1.806039e-07,1.806045e-07,1.806051e-07,1.806057e-07,1.806064e-07,1.806070e-07,1.806076e-07,1.806082e-07,1.806088e-07,1.806094e-07,1.806100e-07,1.806107e-07,1.806113e-07,1.806119e-07,1.806125e-07,1.806131e-07,1.806137e-07,1.806143e-07,1.806149e-07,1.806156e-07,1.806162e-07,1.806168e-07,1.806174e-07,1.806180e-07,1.806186e-07,1.806192e-07,1.806198e-07,1.806205e-07,1.806211e-07,1.806217e-07,1.806223e-07,1.806229e-07,1.806235e-07,1.806241e-07,1.806248e-07,1.806254e-07,1.806260e-07,1.806266e-07,1.806272e-07,1.806278e-07,1.806284e-07,1.806290e-07,1.806297e-07,1.806303e-07,1.806309e-07,1.806315e-07,1.806321e-07,1.806327e-07,1.806333e-07,1.806339e-07,1.806346e-07,1.806352e-07,1.806358e-07,1.806364e-07,1.806370e-07,1.806376e-07,1.806382e-07,1.806388e-07,1.806394e-07,1.806401e-07,1.806407e-07,1.806413e-07,1.806419e-07,1.806425e-07,1.806431e-07,1.806437e-07,1.806443e-07,1.806450e-07,1.806456e-07,1.806462e-07,1.806468e-07,1.806474e-07,1.806480e-07,1.806486e-07,1.806492e-07,1.806498e-07,1.806505e-07,1.806511e-07,1.806517e-07,1.806523e-07,1.806529e-07,1.806535e-07,1.806541e-07,1.806547e-07,1.806553e-07,1.806560e-07,1.806566e-07,1.806572e-07,1.806578e-07,1.806584e-07,1.806590e-07,1.806596e-07,1.806602e-07,1.806608e-07,1.806615e-07,1.806621e-07,1.806627e-07,1.806633e-07,1.806639e-07,1.806645e-07,1.806651e-07,1.806657e-07,1.806663e-07,1.806670e-07,1.806676e-07,1.806682e-07,1.806688e-07,1.806694e-07,1.806700e-07,1.806706e-07,1.806712e-07,1.806718e-07,1.806724e-07,1.806731e-07,1.806737e-07,1.806743e-07,1.806749e-07,1.806755e-07,1.806761e-07,1.806767e-07,1.806773e-07,1.806779e-07,1.806785e-07,1.806792e-07,1.806798e-07,1.806804e-07,1.806810e-07,1.806816e-07,1.806822e-07,1.806828e-07,1.806834e-07,1.806840e-07,1.806846e-07,1.806853e-07,1.806859e-07,1.806865e-07,1.806871e-07,1.806877e-07,1.806883e-07,1.806889e-07,1.806895e-07,1.806901e-07,1.806907e-07,1.806913e-07,1.806920e-07,1.806926e-07,1.806932e-07,1.806938e-07,1.806944e-07,1.806950e-07,1.806956e-07,1.806962e-07,1.806968e-07,1.806974e-07,1.806980e-07,1.806987e-07,1.806993e-07,1.806999e-07,1.807005e-07,1.807011e-07,1.807017e-07,1.807023e-07,1.807029e-07,1.807035e-07,1.807041e-07,1.807047e-07,1.807053e-07,1.807060e-07,1.807066e-07,1.807072e-07,1.807078e-07,1.807084e-07,1.807090e-07,1.807096e-07,1.807102e-07,1.807108e-07,1.807114e-07,1.807120e-07,1.807126e-07,1.807133e-07,1.807139e-07,1.807145e-07,1.807151e-07,1.807157e-07,1.807163e-07,1.807169e-07,1.807175e-07,1.807181e-07,1.807187e-07,1.807193e-07,1.807199e-07,1.807206e-07,1.807212e-07,1.807218e-07,1.807224e-07,1.807230e-07,1.807236e-07,1.807242e-07,1.807248e-07,1.807254e-07,1.807260e-07,1.807266e-07,1.807272e-07,1.807278e-07,1.807284e-07,1.807291e-07,1.807297e-07,1.807303e-07,1.807309e-07,1.807315e-07,1.807321e-07,1.807327e-07,1.807333e-07,1.807339e-07,1.807345e-07,1.807351e-07,1.807357e-07,1.807363e-07,1.807369e-07,1.807376e-07,1.807382e-07,1.807388e-07,1.807394e-07,1.807400e-07,1.807406e-07,1.807412e-07,1.807418e-07,1.807424e-07,1.807430e-07,1.807436e-07,1.807442e-07,1.807448e-07,1.807454e-07,1.807460e-07,1.807467e-07,1.807473e-07,1.807479e-07,1.807485e-07,1.807491e-07,1.807497e-07,1.807503e-07,1.807509e-07,1.807515e-07,1.807521e-07,1.807527e-07,1.807533e-07,1.807539e-07,1.807545e-07,1.807551e-07,1.807557e-07,1.807564e-07,1.807570e-07,1.807576e-07,1.807582e-07,1.807588e-07,1.807594e-07,1.807600e-07,1.807606e-07,1.807612e-07,1.807618e-07,1.807624e-07,1.807630e-07,1.807636e-07,1.807642e-07,1.807648e-07,1.807654e-07,1.807660e-07,1.807666e-07,1.807673e-07,1.807679e-07,1.807685e-07,1.807691e-07,1.807697e-07,1.807703e-07,1.807709e-07,1.807715e-07,1.807721e-07,1.807727e-07,1.807733e-07,1.807739e-07,1.807745e-07,1.807751e-07,1.807757e-07,1.807763e-07,1.807769e-07,1.807775e-07,1.807781e-07,1.807787e-07,1.807793e-07,1.807800e-07,1.807806e-07,1.807812e-07,1.807818e-07,1.807824e-07,1.807830e-07,1.807836e-07,1.807842e-07,1.807848e-07,1.807854e-07,1.807860e-07,1.807866e-07,1.807872e-07,1.807878e-07,1.807884e-07,1.807890e-07,1.807896e-07,1.807902e-07,1.807908e-07,1.807914e-07,1.807920e-07,1.807926e-07,1.807932e-07,1.807939e-07,1.807945e-07,1.807951e-07,1.807957e-07,1.807963e-07,1.807969e-07,1.807975e-07,1.807981e-07,1.807987e-07,1.807993e-07,1.807999e-07,1.808005e-07,1.808011e-07,1.808017e-07,1.808023e-07,1.808029e-07,1.808035e-07,1.808041e-07,1.808047e-07,1.808053e-07,1.808059e-07,1.808065e-07,1.808071e-07,1.808077e-07,1.808083e-07,1.808089e-07,1.808095e-07,1.808101e-07,1.808107e-07,1.808114e-07,1.808120e-07,1.808126e-07,1.808132e-07,1.808138e-07,1.808144e-07,1.808150e-07,1.808156e-07,1.808162e-07,1.808168e-07,1.808174e-07,1.808180e-07,1.808186e-07,1.808192e-07,1.808198e-07,1.808204e-07,1.808210e-07,1.808216e-07,1.808222e-07,1.808228e-07,1.808234e-07,1.808240e-07,1.808246e-07,1.808252e-07,1.808258e-07,1.808264e-07,1.808270e-07,1.808276e-07,1.808282e-07,1.808288e-07,1.808294e-07,1.808300e-07,1.808306e-07,1.808312e-07,1.808318e-07,1.808324e-07,1.808330e-07,1.808336e-07,1.808342e-07,1.808348e-07,1.808354e-07,1.808360e-07,1.808366e-07,1.808373e-07,1.808379e-07,1.808385e-07,1.808391e-07,1.808397e-07,1.808403e-07,1.808409e-07,1.808415e-07,1.808421e-07,1.808427e-07,1.808433e-07,1.808439e-07,1.808445e-07,1.808451e-07,1.808457e-07,1.808463e-07,1.808469e-07,1.808475e-07,1.808481e-07,1.808487e-07,1.808493e-07,1.808499e-07,1.808505e-07,1.808511e-07,1.808517e-07,1.808523e-07,1.808529e-07,1.808535e-07,1.808541e-07,1.808547e-07,1.808553e-07,1.808559e-07,1.808565e-07,1.808571e-07,1.808577e-07,1.808583e-07,1.808589e-07,1.808595e-07,1.808601e-07,1.808607e-07,1.808613e-07,1.808619e-07,1.808625e-07,1.808631e-07,1.808637e-07,1.808643e-07,1.808649e-07,1.808655e-07,1.808661e-07,1.808667e-07,1.808673e-07,1.808679e-07,1.808685e-07,1.808691e-07,1.808697e-07,1.808703e-07,1.808709e-07,1.808715e-07,1.808721e-07,1.808727e-07,1.808733e-07,1.808739e-07,1.808745e-07,1.808751e-07,1.808757e-07,1.808763e-07,1.808769e-07,1.808775e-07,1.808781e-07,1.808787e-07,1.808793e-07,1.808799e-07,1.808805e-07,1.808811e-07,1.808817e-07,1.808823e-07,1.808829e-07,1.808835e-07,1.808841e-07,1.808847e-07,1.808853e-07,1.808859e-07,1.808865e-07,1.808871e-07,1.808877e-07,1.808883e-07,1.808889e-07,1.808895e-07,1.808901e-07,1.808907e-07,1.808913e-07,1.808919e-07,1.808925e-07,1.808931e-07,1.808937e-07,1.808943e-07,1.808949e-07,1.808955e-07,1.808961e-07,1.808967e-07,1.808973e-07,1.808979e-07,1.808985e-07,1.808991e-07,1.808997e-07,1.809003e-07,1.809009e-07,1.809014e-07,1.809020e-07,1.809026e-07,1.809032e-07,1.809038e-07,1.809044e-07,1.809050e-07,1.809056e-07,1.809062e-07,1.809068e-07,1.809074e-07,1.809080e-07,1.809086e-07,1.809092e-07,1.809098e-07,1.809104e-07,1.809110e-07,1.809116e-07,1.809122e-07,1.809128e-07,1.809134e-07,1.809140e-07,1.809146e-07,1.809152e-07,1.809158e-07,1.809164e-07,1.809170e-07,1.809176e-07,1.809182e-07,1.809188e-07,1.809194e-07,1.809200e-07,1.809206e-07,1.809212e-07,1.809218e-07,1.809224e-07,1.809230e-07,1.809236e-07,1.809242e-07,1.809248e-07,1.809254e-07,1.809260e-07,1.809266e-07,1.809271e-07,1.809277e-07,1.809283e-07,1.809289e-07,1.809295e-07,1.809301e-07,1.809307e-07,1.809313e-07,1.809319e-07,1.809325e-07,1.809331e-07,1.809337e-07,1.809343e-07,1.809349e-07,1.809355e-07,1.809361e-07,1.809367e-07,1.809373e-07,1.809379e-07,1.809385e-07,1.809391e-07,1.809397e-07,1.809403e-07,1.809409e-07,1.809415e-07,1.809421e-07,1.809427e-07,1.809433e-07,1.809439e-07,1.809444e-07,1.809450e-07,1.809456e-07,1.809462e-07,1.809468e-07,1.809474e-07,1.809480e-07,1.809486e-07,1.809492e-07,1.809498e-07,1.809504e-07,1.809510e-07,1.809516e-07,1.809522e-07,1.809528e-07,1.809534e-07,1.809540e-07,1.809546e-07,1.809552e-07,1.809558e-07,1.809564e-07,1.809570e-07,1.809576e-07,1.809582e-07,1.809587e-07,1.809593e-07,1.809599e-07,1.809605e-07,1.809611e-07,1.809617e-07,1.809623e-07,1.809629e-07,1.809635e-07,1.809641e-07,1.809647e-07,1.809653e-07,1.809659e-07,1.809665e-07,1.809671e-07,1.809677e-07,1.809683e-07,1.809689e-07,1.809695e-07,1.809701e-07,1.809706e-07,1.809712e-07,1.809718e-07,1.809724e-07,1.809730e-07,1.809736e-07,1.809742e-07,1.809748e-07,1.809754e-07,1.809760e-07,1.809766e-07,1.809772e-07,1.809778e-07,1.809784e-07,1.809790e-07,1.809796e-07,1.809802e-07,1.809808e-07,1.809814e-07,1.809819e-07,1.809825e-07,1.809831e-07,1.809837e-07,1.809843e-07,1.809849e-07,1.809855e-07,1.809861e-07,1.809867e-07,1.809873e-07,1.809879e-07,1.809885e-07,1.809891e-07,1.809897e-07,1.809903e-07,1.809909e-07,1.809914e-07,1.809920e-07,1.809926e-07,1.809932e-07,1.809938e-07,1.809944e-07,1.809950e-07,1.809956e-07,1.809962e-07,1.809968e-07,1.809974e-07,1.809980e-07,1.809986e-07,1.809992e-07,1.809998e-07,1.810004e-07,1.810009e-07,1.810015e-07,1.810021e-07,1.810027e-07,1.810033e-07,1.810039e-07,1.810045e-07,1.810051e-07,1.810057e-07,1.810063e-07,1.810069e-07,1.810075e-07,1.810081e-07,1.810087e-07,1.810092e-07,1.810098e-07,1.810104e-07,1.810110e-07,1.810116e-07,1.810122e-07,1.810128e-07,1.810134e-07,1.810140e-07,1.810146e-07,1.810152e-07,1.810158e-07,1.810164e-07,1.810170e-07,1.810175e-07,1.810181e-07,1.810187e-07,1.810193e-07,1.810199e-07,1.810205e-07,1.810211e-07,1.810217e-07,1.810223e-07,1.810229e-07,1.810235e-07,1.810241e-07,1.810247e-07,1.810252e-07,1.810258e-07,1.810264e-07,1.810270e-07,1.810276e-07,1.810282e-07,1.810288e-07,1.810294e-07,1.810300e-07,1.810306e-07,1.810312e-07,1.810318e-07,1.810323e-07,1.810329e-07,1.810335e-07,1.810341e-07,1.810347e-07,1.810353e-07,1.810359e-07,1.810365e-07,1.810371e-07,1.810377e-07,1.810383e-07,1.810389e-07,1.810394e-07,1.810400e-07,1.810406e-07,1.810412e-07,1.810418e-07,1.810424e-07,1.810430e-07,1.810436e-07,1.810442e-07,1.810448e-07,1.810454e-07,1.810459e-07,1.810465e-07,1.810471e-07,1.810477e-07,1.810483e-07,1.810489e-07,1.810495e-07,1.810501e-07,1.810507e-07,1.810513e-07,1.810519e-07,1.810524e-07,1.810530e-07,1.810536e-07,1.810542e-07,1.810548e-07,1.810554e-07,1.810560e-07,1.810566e-07,1.810572e-07,1.810578e-07,1.810583e-07,1.810589e-07,1.810595e-07,1.810601e-07,1.810607e-07,1.810613e-07,1.810619e-07,1.810625e-07,1.810631e-07,1.810637e-07,1.810643e-07,1.810648e-07,1.810654e-07,1.810660e-07,1.810666e-07,1.810672e-07,1.810678e-07,1.810684e-07,1.810690e-07,1.810696e-07,1.810701e-07,1.810707e-07,1.810713e-07,1.810719e-07,1.810725e-07,1.810731e-07,1.810737e-07,1.810743e-07,1.810749e-07,1.810755e-07,1.810760e-07,1.810766e-07,1.810772e-07,1.810778e-07,1.810784e-07,1.810790e-07,1.810796e-07,1.810802e-07,1.810808e-07,1.810813e-07,1.810819e-07,1.810825e-07,1.810831e-07,1.810837e-07,1.810843e-07,1.810849e-07,1.810855e-07,1.810861e-07,1.810867e-07,1.810872e-07,1.810878e-07,1.810884e-07,1.810890e-07,1.810896e-07,1.810902e-07,1.810908e-07,1.810914e-07,1.810920e-07,1.810925e-07,1.810931e-07,1.810937e-07,1.810943e-07,1.810949e-07,1.810955e-07,1.810961e-07,1.810967e-07,1.810972e-07,1.810978e-07,1.810984e-07,1.810990e-07,1.810996e-07,1.811002e-07,1.811008e-07,1.811014e-07,1.811020e-07,1.811025e-07,1.811031e-07,1.811037e-07,1.811043e-07,1.811049e-07,1.811055e-07,1.811061e-07,1.811067e-07,1.811072e-07,1.811078e-07,1.811084e-07,1.811090e-07,1.811096e-07,1.811102e-07,1.811108e-07,1.811114e-07,1.811119e-07,1.811125e-07,1.811131e-07,1.811137e-07,1.811143e-07,1.811149e-07,1.811155e-07,1.811161e-07,1.811166e-07,1.811172e-07,1.811178e-07,1.811184e-07,1.811190e-07,1.811196e-07,1.811202e-07,1.811208e-07,1.811213e-07,1.811219e-07,1.811225e-07,1.811231e-07,1.811237e-07,1.811243e-07,1.811249e-07,1.811255e-07,1.811260e-07,1.811266e-07,1.811272e-07,1.811278e-07,1.811284e-07,1.811290e-07,1.811296e-07,1.811301e-07,1.811307e-07,1.811313e-07,1.811319e-07,1.811325e-07,1.811331e-07,1.811337e-07,1.811343e-07,1.811348e-07,1.811354e-07,1.811360e-07,1.811366e-07,1.811372e-07,1.811378e-07,1.811384e-07,1.811389e-07,1.811395e-07,1.811401e-07,1.811407e-07,1.811413e-07,1.811419e-07,1.811425e-07,1.811430e-07,1.811436e-07,1.811442e-07,1.811448e-07,1.811454e-07,1.811460e-07,1.811466e-07,1.811472e-07,1.811477e-07,1.811483e-07,1.811489e-07,1.811495e-07,1.811501e-07,1.811507e-07,1.811513e-07,1.811518e-07,1.811524e-07,1.811530e-07,1.811536e-07,1.811542e-07,1.811548e-07,1.811554e-07,1.811559e-07,1.811565e-07,1.811571e-07,1.811577e-07,1.811583e-07,1.811589e-07,1.811594e-07,1.811600e-07,1.811606e-07,1.811612e-07,1.811618e-07,1.811624e-07,1.811630e-07,1.811635e-07,1.811641e-07,1.811647e-07,1.811653e-07,1.811659e-07,1.811665e-07,1.811671e-07,1.811676e-07,1.811682e-07,1.811688e-07,1.811694e-07,1.811700e-07,1.811706e-07,1.811711e-07,1.811717e-07,1.811723e-07,1.811729e-07,1.811735e-07,1.811741e-07,1.811747e-07,1.811752e-07,1.811758e-07,1.811764e-07,1.811770e-07,1.811776e-07,1.811782e-07,1.811787e-07,1.811793e-07,1.811799e-07,1.811805e-07,1.811811e-07,1.811817e-07,1.811823e-07,1.811828e-07,1.811834e-07,1.811840e-07,1.811846e-07,1.811852e-07,1.811858e-07,1.811863e-07,1.811869e-07,1.811875e-07,1.811881e-07,1.811887e-07,1.811893e-07,1.811898e-07,1.811904e-07,1.811910e-07,1.811916e-07,1.811922e-07,1.811928e-07,1.811933e-07,1.811939e-07,1.811945e-07,1.811951e-07,1.811957e-07,1.811963e-07,1.811968e-07,1.811974e-07,1.811980e-07,1.811986e-07,1.811992e-07,1.811998e-07,1.812003e-07,1.812009e-07,1.812015e-07,1.812021e-07,1.812027e-07,1.812033e-07,1.812038e-07,1.812044e-07,1.812050e-07,1.812056e-07,1.812062e-07,1.812068e-07,1.812073e-07,1.812079e-07,1.812085e-07,1.812091e-07,1.812097e-07,1.812103e-07,1.812108e-07,1.812114e-07,1.812120e-07,1.812126e-07,1.812132e-07,1.812137e-07,1.812143e-07,1.812149e-07,1.812155e-07,1.812161e-07,1.812167e-07,1.812172e-07,1.812178e-07,1.812184e-07,1.812190e-07,1.812196e-07,1.812202e-07,1.812207e-07,1.812213e-07,1.812219e-07,1.812225e-07,1.812231e-07,1.812236e-07,1.812242e-07,1.812248e-07,1.812254e-07,1.812260e-07,1.812266e-07,1.812271e-07,1.812277e-07,1.812283e-07,1.812289e-07,1.812295e-07,1.812300e-07,1.812306e-07,1.812312e-07,1.812318e-07,1.812324e-07,1.812330e-07,1.812335e-07,1.812341e-07,1.812347e-07,1.812353e-07,1.812359e-07,1.812364e-07,1.812370e-07,1.812376e-07,1.812382e-07,1.812388e-07,1.812394e-07,1.812399e-07,1.812405e-07,1.812411e-07,1.812417e-07,1.812423e-07,1.812428e-07,1.812434e-07,1.812440e-07,1.812446e-07,1.812452e-07,1.812457e-07,1.812463e-07,1.812469e-07,1.812475e-07,1.812481e-07,1.812486e-07,1.812492e-07,1.812498e-07,1.812504e-07,1.812510e-07,1.812516e-07,1.812521e-07,1.812527e-07,1.812533e-07,1.812539e-07,1.812545e-07,1.812550e-07,1.812556e-07,1.812562e-07,1.812568e-07,1.812574e-07,1.812579e-07,1.812585e-07,1.812591e-07,1.812597e-07,1.812603e-07,1.812608e-07,1.812614e-07,1.812620e-07,1.812626e-07,1.812632e-07,1.812637e-07,1.812643e-07,1.812649e-07,1.812655e-07,1.812661e-07,1.812666e-07,1.812672e-07,1.812678e-07,1.812684e-07,1.812690e-07,1.812695e-07,1.812701e-07,1.812707e-07,1.812713e-07,1.812719e-07,1.812724e-07,1.812730e-07,1.812736e-07,1.812742e-07,1.812748e-07,1.812753e-07,1.812759e-07,1.812765e-07,1.812771e-07,1.812777e-07,1.812782e-07,1.812788e-07,1.812794e-07,1.812800e-07,1.812805e-07,1.812811e-07,1.812817e-07,1.812823e-07,1.812829e-07,1.812834e-07,1.812840e-07,1.812846e-07,1.812852e-07,1.812858e-07,1.812863e-07,1.812869e-07,1.812875e-07,1.812881e-07,1.812887e-07,1.812892e-07,1.812898e-07,1.812904e-07,1.812910e-07,1.812915e-07,1.812921e-07,1.812927e-07,1.812933e-07,1.812939e-07,1.812944e-07,1.812950e-07,1.812956e-07,1.812962e-07,1.812968e-07,1.812973e-07,1.812979e-07,1.812985e-07,1.812991e-07,1.812996e-07,1.813002e-07,1.813008e-07,1.813014e-07,1.813020e-07,1.813025e-07,1.813031e-07,1.813037e-07,1.813043e-07,1.813048e-07,1.813054e-07,1.813060e-07,1.813066e-07,1.813072e-07,1.813077e-07,1.813083e-07,1.813089e-07,1.813095e-07,1.813100e-07,1.813106e-07,1.813112e-07,1.813118e-07,1.813124e-07,1.813129e-07,1.813135e-07,1.813141e-07,1.813147e-07,1.813152e-07,1.813158e-07,1.813164e-07,1.813170e-07,1.813176e-07,1.813181e-07,1.813187e-07,1.813193e-07,1.813199e-07,1.813204e-07,1.813210e-07,1.813216e-07,1.813222e-07,1.813228e-07,1.813233e-07,1.813239e-07,1.813245e-07,1.813251e-07,1.813256e-07,1.813262e-07,1.813268e-07,1.813274e-07,1.813279e-07,1.813285e-07,1.813291e-07,1.813297e-07,1.813303e-07,1.813308e-07,1.813314e-07,1.813320e-07,1.813326e-07,1.813331e-07,1.813337e-07,1.813343e-07,1.813349e-07,1.813354e-07,1.813360e-07,1.813366e-07,1.813372e-07,1.813377e-07,1.813383e-07,1.813389e-07,1.813395e-07,1.813401e-07,1.813406e-07,1.813412e-07,1.813418e-07,1.813424e-07,1.813429e-07,1.813435e-07,1.813441e-07,1.813447e-07,1.813452e-07,1.813458e-07,1.813464e-07,1.813470e-07,1.813475e-07,1.813481e-07,1.813487e-07,1.813493e-07,1.813498e-07,1.813504e-07,1.813510e-07,1.813516e-07,1.813521e-07,1.813527e-07,1.813533e-07,1.813539e-07,1.813545e-07,1.813550e-07,1.813556e-07,1.813562e-07,1.813568e-07,1.813573e-07,1.813579e-07,1.813585e-07,1.813591e-07,1.813596e-07,1.813602e-07,1.813608e-07,1.813614e-07,1.813619e-07,1.813625e-07,1.813631e-07,1.813637e-07,1.813642e-07,1.813648e-07,1.813654e-07,1.813660e-07,1.813665e-07,1.813671e-07,1.813677e-07,1.813683e-07,1.813688e-07,1.813694e-07,1.813700e-07,1.813706e-07,1.813711e-07,1.813717e-07,1.813723e-07,1.813729e-07,1.813734e-07,1.813740e-07,1.813746e-07,1.813752e-07,1.813757e-07,1.813763e-07,1.813769e-07,1.813774e-07,1.813780e-07,1.813786e-07,1.813792e-07,1.813797e-07,1.813803e-07,1.813809e-07,1.813815e-07,1.813820e-07,1.813826e-07,1.813832e-07,1.813838e-07,1.813843e-07,1.813849e-07,1.813855e-07,1.813861e-07,1.813866e-07,1.813872e-07,1.813878e-07,1.813884e-07,1.813889e-07,1.813895e-07,1.813901e-07,1.813907e-07,1.813912e-07,1.813918e-07,1.813924e-07,1.813929e-07,1.813935e-07,1.813941e-07,1.813947e-07,1.813952e-07,1.813958e-07,1.813964e-07,1.813970e-07,1.813975e-07,1.813981e-07,1.813987e-07,1.813993e-07,1.813998e-07,1.814004e-07,1.814010e-07,1.814015e-07,1.814021e-07,1.814027e-07,1.814033e-07,1.814038e-07,1.814044e-07,1.814050e-07,1.814056e-07,1.814061e-07,1.814067e-07,1.814073e-07,1.814079e-07,1.814084e-07,1.814090e-07,1.814096e-07,1.814101e-07,1.814107e-07,1.814113e-07,1.814119e-07,1.814124e-07,1.814130e-07,1.814136e-07,1.814142e-07,1.814147e-07,1.814153e-07,1.814159e-07,1.814164e-07,1.814170e-07,1.814176e-07,1.814182e-07,1.814187e-07,1.814193e-07,1.814199e-07,1.814205e-07,1.814210e-07,1.814216e-07,1.814222e-07,1.814227e-07,1.814233e-07,1.814239e-07,1.814245e-07,1.814250e-07,1.814256e-07,1.814262e-07,1.814267e-07,1.814273e-07,1.814279e-07,1.814285e-07,1.814290e-07,1.814296e-07,1.814302e-07,1.814307e-07,1.814313e-07,1.814319e-07,1.814325e-07,1.814330e-07,1.814336e-07,1.814342e-07,1.814347e-07,1.814353e-07,1.814359e-07,1.814365e-07,1.814370e-07,1.814376e-07,1.814382e-07,1.814387e-07,1.814393e-07,1.814399e-07,1.814405e-07,1.814410e-07,1.814416e-07,1.814422e-07,1.814427e-07,1.814433e-07,1.814439e-07,1.814445e-07,1.814450e-07,1.814456e-07,1.814462e-07,1.814467e-07,1.814473e-07,1.814479e-07,1.814485e-07,1.814490e-07,1.814496e-07,1.814502e-07,1.814507e-07,1.814513e-07,1.814519e-07,1.814525e-07,1.814530e-07,1.814536e-07,1.814542e-07,1.814547e-07,1.814553e-07,1.814559e-07,1.814564e-07,1.814570e-07,1.814576e-07,1.814582e-07,1.814587e-07,1.814593e-07,1.814599e-07,1.814604e-07,1.814610e-07,1.814616e-07,1.814622e-07,1.814627e-07,1.814633e-07,1.814639e-07,1.814644e-07,1.814650e-07,1.814656e-07,1.814661e-07,1.814667e-07,1.814673e-07,1.814679e-07,1.814684e-07,1.814690e-07,1.814696e-07,1.814701e-07,1.814707e-07,1.814713e-07,1.814718e-07,1.814724e-07,1.814730e-07,1.814736e-07,1.814741e-07,1.814747e-07,1.814753e-07,1.814758e-07,1.814764e-07,1.814770e-07,1.814775e-07,1.814781e-07,1.814787e-07,1.814792e-07,1.814798e-07,1.814804e-07,1.814810e-07,1.814815e-07,1.814821e-07,1.814827e-07,1.814832e-07,1.814838e-07,1.814844e-07,1.814849e-07,1.814855e-07,1.814861e-07,1.814866e-07,1.814872e-07,1.814878e-07,1.814884e-07,1.814889e-07,1.814895e-07,1.814901e-07,1.814906e-07,1.814912e-07,1.814918e-07,1.814923e-07,1.814929e-07,1.814935e-07,1.814940e-07,1.814946e-07,1.814952e-07,1.814957e-07,1.814963e-07,1.814969e-07,1.814975e-07,1.814980e-07,1.814986e-07,1.814992e-07,1.814997e-07,1.815003e-07,1.815009e-07,1.815014e-07,1.815020e-07,1.815026e-07,1.815031e-07,1.815037e-07,1.815043e-07,1.815048e-07,1.815054e-07,1.815060e-07,1.815065e-07,1.815071e-07,1.815077e-07,1.815083e-07,1.815088e-07,1.815094e-07,1.815100e-07,1.815105e-07,1.815111e-07,1.815117e-07,1.815122e-07,1.815128e-07,1.815134e-07,1.815139e-07,1.815145e-07,1.815151e-07,1.815156e-07,1.815162e-07,1.815168e-07,1.815173e-07,1.815179e-07,1.815185e-07,1.815190e-07,1.815196e-07,1.815202e-07,1.815207e-07,1.815213e-07,1.815219e-07,1.815224e-07,1.815230e-07,1.815236e-07,1.815241e-07,1.815247e-07,1.815253e-07,1.815258e-07,1.815264e-07,1.815270e-07,1.815275e-07,1.815281e-07,1.815287e-07,1.815292e-07,1.815298e-07,1.815304e-07,1.815309e-07,1.815315e-07,1.815321e-07,1.815326e-07,1.815332e-07,1.815338e-07,1.815344e-07,1.815349e-07,1.815355e-07,1.815361e-07,1.815366e-07,1.815372e-07,1.815378e-07,1.815383e-07,1.815389e-07,1.815394e-07,1.815400e-07,1.815406e-07,1.815411e-07,1.815417e-07,1.815423e-07,1.815428e-07,1.815434e-07,1.815440e-07,1.815445e-07,1.815451e-07,1.815457e-07,1.815462e-07,1.815468e-07,1.815474e-07,1.815479e-07,1.815485e-07,1.815491e-07,1.815496e-07,1.815502e-07,1.815508e-07,1.815513e-07,1.815519e-07,1.815525e-07,1.815530e-07,1.815536e-07,1.815542e-07,1.815547e-07,1.815553e-07,1.815559e-07,1.815564e-07,1.815570e-07,1.815576e-07,1.815581e-07,1.815587e-07,1.815593e-07,1.815598e-07,1.815604e-07,1.815610e-07,1.815615e-07,1.815621e-07,1.815627e-07,1.815632e-07,1.815638e-07,1.815643e-07,1.815649e-07,1.815655e-07,1.815660e-07,1.815666e-07,1.815672e-07,1.815677e-07,1.815683e-07,1.815689e-07,1.815694e-07,1.815700e-07,1.815706e-07,1.815711e-07,1.815717e-07,1.815723e-07,1.815728e-07,1.815734e-07,1.815740e-07,1.815745e-07,1.815751e-07,1.815756e-07,1.815762e-07,1.815768e-07,1.815773e-07,1.815779e-07,1.815785e-07,1.815790e-07,1.815796e-07,1.815802e-07,1.815807e-07,1.815813e-07,1.815819e-07,1.815824e-07,1.815830e-07,1.815836e-07,1.815841e-07,1.815847e-07,1.815852e-07,1.815858e-07,1.815864e-07,1.815869e-07,1.815875e-07,1.815881e-07,1.815886e-07,1.815892e-07,1.815898e-07,1.815903e-07,1.815909e-07,1.815914e-07,1.815920e-07,1.815926e-07,1.815931e-07,1.815937e-07,1.815943e-07,1.815948e-07,1.815954e-07,1.815960e-07,1.815965e-07,1.815971e-07,1.815977e-07,1.815982e-07,1.815988e-07,1.815993e-07,1.815999e-07,1.816005e-07,1.816010e-07,1.816016e-07,1.816022e-07,1.816027e-07,1.816033e-07,1.816039e-07,1.816044e-07,1.816050e-07,1.816055e-07,1.816061e-07,1.816067e-07,1.816072e-07,1.816078e-07,1.816084e-07,1.816089e-07,1.816095e-07,1.816100e-07,1.816106e-07,1.816112e-07,1.816117e-07,1.816123e-07,1.816129e-07,1.816134e-07,1.816140e-07,1.816145e-07,1.816151e-07,1.816157e-07,1.816162e-07,1.816168e-07,1.816174e-07,1.816179e-07,1.816185e-07,1.816191e-07,1.816196e-07,1.816202e-07,1.816207e-07,1.816213e-07,1.816219e-07,1.816224e-07,1.816230e-07,1.816236e-07,1.816241e-07,1.816247e-07,1.816252e-07,1.816258e-07,1.816264e-07,1.816269e-07,1.816275e-07,1.816280e-07,1.816286e-07,1.816292e-07,1.816297e-07,1.816303e-07,1.816309e-07,1.816314e-07,1.816320e-07,1.816325e-07,1.816331e-07,1.816337e-07,1.816342e-07,1.816348e-07,1.816354e-07,1.816359e-07,1.816365e-07,1.816370e-07,1.816376e-07,1.816382e-07,1.816387e-07,1.816393e-07,1.816398e-07,1.816404e-07,1.816410e-07,1.816415e-07,1.816421e-07,1.816427e-07,1.816432e-07,1.816438e-07,1.816443e-07,1.816449e-07,1.816455e-07,1.816460e-07,1.816466e-07,1.816471e-07,1.816477e-07,1.816483e-07,1.816488e-07,1.816494e-07,1.816500e-07,1.816505e-07,1.816511e-07,1.816516e-07,1.816522e-07,1.816528e-07,1.816533e-07,1.816539e-07,1.816544e-07,1.816550e-07,1.816556e-07,1.816561e-07,1.816567e-07,1.816572e-07,1.816578e-07,1.816584e-07,1.816589e-07,1.816595e-07,1.816601e-07,1.816606e-07,1.816612e-07,1.816617e-07,1.816623e-07,1.816629e-07,1.816634e-07,1.816640e-07,1.816645e-07,1.816651e-07,1.816657e-07,1.816662e-07,1.816668e-07,1.816673e-07,1.816679e-07,1.816685e-07,1.816690e-07,1.816696e-07,1.816701e-07,1.816707e-07,1.816713e-07,1.816718e-07,1.816724e-07,1.816729e-07,1.816735e-07,1.816741e-07,1.816746e-07,1.816752e-07,1.816757e-07,1.816763e-07,1.816769e-07,1.816774e-07,1.816780e-07,1.816785e-07,1.816791e-07,1.816797e-07,1.816802e-07,1.816808e-07,1.816813e-07,1.816819e-07,1.816825e-07,1.816830e-07,1.816836e-07,1.816841e-07,1.816847e-07,1.816853e-07,1.816858e-07,1.816864e-07,1.816869e-07,1.816875e-07,1.816880e-07,1.816886e-07,1.816892e-07,1.816897e-07,1.816903e-07,1.816908e-07,1.816914e-07,1.816920e-07,1.816925e-07,1.816931e-07,1.816936e-07,1.816942e-07,1.816948e-07,1.816953e-07,1.816959e-07,1.816964e-07,1.816970e-07,1.816976e-07,1.816981e-07,1.816987e-07,1.816992e-07,1.816998e-07,1.817003e-07,1.817009e-07,1.817015e-07,1.817020e-07,1.817026e-07,1.817031e-07,1.817037e-07,1.817043e-07,1.817048e-07,1.817054e-07,1.817059e-07,1.817065e-07,1.817071e-07,1.817076e-07,1.817082e-07,1.817087e-07,1.817093e-07,1.817098e-07,1.817104e-07,1.817110e-07,1.817115e-07,1.817121e-07,1.817126e-07,1.817132e-07,1.817137e-07,1.817143e-07,1.817149e-07,1.817154e-07,1.817160e-07,1.817165e-07,1.817171e-07,1.817177e-07,1.817182e-07,1.817188e-07,1.817193e-07,1.817199e-07,1.817204e-07,1.817210e-07,1.817216e-07,1.817221e-07,1.817227e-07,1.817232e-07,1.817238e-07,1.817243e-07,1.817249e-07,1.817255e-07,1.817260e-07,1.817266e-07,1.817271e-07,1.817277e-07,1.817283e-07,1.817288e-07,1.817294e-07,1.817299e-07,1.817305e-07,1.817310e-07,1.817316e-07,1.817322e-07,1.817327e-07,1.817333e-07,1.817338e-07,1.817344e-07,1.817349e-07,1.817355e-07,1.817361e-07,1.817366e-07,1.817372e-07,1.817377e-07,1.817383e-07,1.817388e-07,1.817394e-07,1.817399e-07,1.817405e-07,1.817411e-07,1.817416e-07,1.817422e-07,1.817427e-07,1.817433e-07,1.817438e-07,1.817444e-07,1.817450e-07,1.817455e-07,1.817461e-07,1.817466e-07,1.817472e-07,1.817477e-07,1.817483e-07,1.817489e-07,1.817494e-07,1.817500e-07,1.817505e-07,1.817511e-07,1.817516e-07,1.817522e-07,1.817527e-07,1.817533e-07,1.817539e-07,1.817544e-07,1.817550e-07,1.817555e-07,1.817561e-07,1.817566e-07,1.817572e-07,1.817578e-07,1.817583e-07,1.817589e-07,1.817594e-07,1.817600e-07,1.817605e-07,1.817611e-07,1.817616e-07,1.817622e-07,1.817628e-07,1.817633e-07,1.817639e-07,1.817644e-07,1.817650e-07,1.817655e-07,1.817661e-07,1.817666e-07,1.817672e-07,1.817678e-07,1.817683e-07,1.817689e-07,1.817694e-07,1.817700e-07,1.817705e-07,1.817711e-07,1.817716e-07,1.817722e-07,1.817728e-07,1.817733e-07,1.817739e-07,1.817744e-07,1.817750e-07,1.817755e-07,1.817761e-07,1.817766e-07,1.817772e-07,1.817778e-07,1.817783e-07,1.817789e-07,1.817794e-07,1.817800e-07,1.817805e-07,1.817811e-07,1.817816e-07,1.817822e-07,1.817827e-07,1.817833e-07,1.817839e-07,1.817844e-07,1.817850e-07,1.817855e-07,1.817861e-07,1.817866e-07,1.817872e-07,1.817877e-07,1.817883e-07,1.817888e-07,1.817894e-07,1.817900e-07,1.817905e-07,1.817911e-07,1.817916e-07,1.817922e-07,1.817927e-07,1.817933e-07,1.817938e-07,1.817944e-07,1.817949e-07,1.817955e-07,1.817961e-07,1.817966e-07,1.817972e-07,1.817977e-07,1.817983e-07,1.817988e-07,1.817994e-07,1.817999e-07,1.818005e-07,1.818010e-07,1.818016e-07,1.818021e-07,1.818027e-07,1.818033e-07,1.818038e-07,1.818044e-07,1.818049e-07,1.818055e-07,1.818060e-07,1.818066e-07,1.818071e-07,1.818077e-07,1.818082e-07,1.818088e-07,1.818093e-07,1.818099e-07,1.818105e-07,1.818110e-07,1.818116e-07,1.818121e-07,1.818127e-07,1.818132e-07,1.818138e-07,1.818143e-07,1.818149e-07,1.818154e-07,1.818160e-07,1.818165e-07,1.818171e-07,1.818176e-07,1.818182e-07,1.818188e-07,1.818193e-07,1.818199e-07,1.818204e-07,1.818210e-07,1.818215e-07,1.818221e-07,1.818226e-07,1.818232e-07,1.818237e-07,1.818243e-07,1.818248e-07,1.818254e-07,1.818259e-07,1.818265e-07,1.818270e-07,1.818276e-07,1.818282e-07,1.818287e-07,1.818293e-07,1.818298e-07,1.818304e-07,1.818309e-07,1.818315e-07,1.818320e-07,1.818326e-07,1.818331e-07,1.818337e-07,1.818342e-07,1.818348e-07,1.818353e-07,1.818359e-07,1.818364e-07,1.818370e-07,1.818375e-07,1.818381e-07,1.818386e-07,1.818392e-07,1.818397e-07,1.818403e-07,1.818409e-07,1.818414e-07,1.818420e-07,1.818425e-07,1.818431e-07,1.818436e-07,1.818442e-07,1.818447e-07,1.818453e-07,1.818458e-07,1.818464e-07,1.818469e-07,1.818475e-07,1.818480e-07,1.818486e-07,1.818491e-07,1.818497e-07,1.818502e-07,1.818508e-07,1.818513e-07,1.818519e-07,1.818524e-07,1.818530e-07,1.818535e-07,1.818541e-07,1.818546e-07,1.818552e-07,1.818557e-07,1.818563e-07,1.818569e-07,1.818574e-07,1.818580e-07,1.818585e-07,1.818591e-07,1.818596e-07,1.818602e-07,1.818607e-07,1.818613e-07,1.818618e-07,1.818624e-07,1.818629e-07,1.818635e-07,1.818640e-07,1.818646e-07,1.818651e-07,1.818657e-07,1.818662e-07,1.818668e-07,1.818673e-07,1.818679e-07,1.818684e-07,1.818690e-07,1.818695e-07,1.818701e-07,1.818706e-07,1.818712e-07,1.818717e-07,1.818723e-07,1.818728e-07,1.818734e-07,1.818739e-07,1.818745e-07,1.818750e-07,1.818756e-07,1.818761e-07,1.818767e-07,1.818772e-07,1.818778e-07,1.818783e-07,1.818789e-07,1.818794e-07,1.818800e-07,1.818805e-07,1.818811e-07,1.818816e-07,1.818822e-07,1.818827e-07,1.818833e-07,1.818838e-07,1.818844e-07,1.818849e-07,1.818855e-07,1.818860e-07,1.818866e-07,1.818871e-07,1.818877e-07,1.818882e-07,1.818888e-07,1.818893e-07,1.818899e-07,1.818904e-07,1.818910e-07,1.818915e-07,1.818921e-07,1.818926e-07,1.818932e-07,1.818937e-07,1.818943e-07,1.818948e-07,1.818954e-07,1.818959e-07,1.818965e-07,1.818970e-07,1.818976e-07,1.818981e-07,1.818987e-07,1.818992e-07,1.818998e-07,1.819003e-07,1.819009e-07,1.819014e-07,1.819020e-07,1.819025e-07,1.819031e-07,1.819036e-07,1.819042e-07,1.819047e-07,1.819053e-07,1.819058e-07,1.819064e-07,1.819069e-07,1.819075e-07,1.819080e-07,1.819086e-07,1.819091e-07,1.819097e-07,1.819102e-07,1.819108e-07,1.819113e-07,1.819118e-07,1.819124e-07,1.819129e-07,1.819135e-07,1.819140e-07,1.819146e-07,1.819151e-07,1.819157e-07,1.819162e-07,1.819168e-07,1.819173e-07,1.819179e-07,1.819184e-07,1.819190e-07,1.819195e-07,1.819201e-07,1.819206e-07,1.819212e-07,1.819217e-07,1.819223e-07,1.819228e-07,1.819234e-07,1.819239e-07,1.819245e-07,1.819250e-07,1.819256e-07,1.819261e-07,1.819267e-07,1.819272e-07,1.819278e-07,1.819283e-07,1.819288e-07,1.819294e-07,1.819299e-07,1.819305e-07,1.819310e-07,1.819316e-07,1.819321e-07,1.819327e-07,1.819332e-07,1.819338e-07,1.819343e-07,1.819349e-07,1.819354e-07,1.819360e-07,1.819365e-07,1.819371e-07,1.819376e-07,1.819382e-07,1.819387e-07,1.819393e-07,1.819398e-07,1.819403e-07,1.819409e-07,1.819414e-07,1.819420e-07,1.819425e-07,1.819431e-07,1.819436e-07,1.819442e-07,1.819447e-07,1.819453e-07,1.819458e-07,1.819464e-07,1.819469e-07,1.819475e-07,1.819480e-07,1.819486e-07,1.819491e-07,1.819496e-07,1.819502e-07,1.819507e-07,1.819513e-07,1.819518e-07,1.819524e-07,1.819529e-07,1.819535e-07,1.819540e-07,1.819546e-07,1.819551e-07,1.819557e-07,1.819562e-07,1.819568e-07,1.819573e-07,1.819578e-07,1.819584e-07,1.819589e-07,1.819595e-07,1.819600e-07,1.819606e-07,1.819611e-07,1.819617e-07,1.819622e-07,1.819628e-07,1.819633e-07,1.819639e-07,1.819644e-07,1.819649e-07,1.819655e-07,1.819660e-07,1.819666e-07,1.819671e-07,1.819677e-07,1.819682e-07,1.819688e-07,1.819693e-07,1.819699e-07,1.819704e-07,1.819710e-07,1.819715e-07,1.819720e-07,1.819726e-07,1.819731e-07,1.819737e-07,1.819742e-07,1.819748e-07,1.819753e-07,1.819759e-07,1.819764e-07,1.819770e-07,1.819775e-07,1.819781e-07,1.819786e-07,1.819791e-07,1.819797e-07,1.819802e-07,1.819808e-07,1.819813e-07,1.819819e-07,1.819824e-07,1.819830e-07,1.819835e-07,1.819841e-07,1.819846e-07,1.819851e-07,1.819857e-07,1.819862e-07,1.819868e-07,1.819873e-07,1.819879e-07,1.819884e-07,1.819890e-07,1.819895e-07,1.819900e-07,1.819906e-07,1.819911e-07,1.819917e-07,1.819922e-07,1.819928e-07,1.819933e-07,1.819939e-07,1.819944e-07,1.819950e-07,1.819955e-07,1.819960e-07,1.819966e-07,1.819971e-07,1.819977e-07,1.819982e-07,1.819988e-07,1.819993e-07,1.819999e-07,1.820004e-07,1.820009e-07,1.820015e-07,1.820020e-07,1.820026e-07,1.820031e-07,1.820037e-07,1.820042e-07,1.820048e-07,1.820053e-07,1.820058e-07,1.820064e-07,1.820069e-07,1.820075e-07,1.820080e-07,1.820086e-07,1.820091e-07,1.820097e-07,1.820102e-07,1.820107e-07,1.820113e-07,1.820118e-07,1.820124e-07,1.820129e-07,1.820135e-07,1.820140e-07,1.820145e-07,1.820151e-07,1.820156e-07,1.820162e-07,1.820167e-07,1.820173e-07,1.820178e-07,1.820184e-07,1.820189e-07,1.820194e-07,1.820200e-07,1.820205e-07,1.820211e-07,1.820216e-07,1.820222e-07,1.820227e-07,1.820232e-07,1.820238e-07,1.820243e-07,1.820249e-07,1.820254e-07,1.820260e-07,1.820265e-07,1.820270e-07,1.820276e-07,1.820281e-07,1.820287e-07,1.820292e-07,1.820298e-07,1.820303e-07,1.820309e-07,1.820314e-07,1.820319e-07,1.820325e-07,1.820330e-07,1.820336e-07,1.820341e-07,1.820347e-07,1.820352e-07,1.820357e-07,1.820363e-07,1.820368e-07,1.820374e-07,1.820379e-07,1.820385e-07,1.820390e-07,1.820395e-07,1.820401e-07,1.820406e-07,1.820412e-07,1.820417e-07,1.820423e-07,1.820428e-07,1.820433e-07,1.820439e-07,1.820444e-07,1.820450e-07,1.820455e-07,1.820460e-07,1.820466e-07,1.820471e-07,1.820477e-07,1.820482e-07,1.820488e-07,1.820493e-07,1.820498e-07,1.820504e-07,1.820509e-07,1.820515e-07,1.820520e-07,1.820526e-07,1.820531e-07,1.820536e-07,1.820542e-07,1.820547e-07,1.820553e-07,1.820558e-07,1.820564e-07,1.820569e-07,1.820574e-07,1.820580e-07,1.820585e-07,1.820591e-07,1.820596e-07,1.820601e-07,1.820607e-07,1.820612e-07,1.820618e-07,1.820623e-07,1.820629e-07,1.820634e-07,1.820639e-07,1.820645e-07,1.820650e-07,1.820656e-07,1.820661e-07,1.820666e-07,1.820672e-07,1.820677e-07,1.820683e-07,1.820688e-07,1.820693e-07,1.820699e-07,1.820704e-07,1.820710e-07,1.820715e-07,1.820721e-07,1.820726e-07,1.820731e-07,1.820737e-07,1.820742e-07,1.820748e-07,1.820753e-07,1.820758e-07,1.820764e-07,1.820769e-07,1.820775e-07,1.820780e-07,1.820785e-07,1.820791e-07,1.820796e-07,1.820802e-07,1.820807e-07,1.820813e-07,1.820818e-07,1.820823e-07,1.820829e-07,1.820834e-07,1.820840e-07,1.820845e-07,1.820850e-07,1.820856e-07,1.820861e-07,1.820867e-07,1.820872e-07,1.820877e-07,1.820883e-07,1.820888e-07,1.820894e-07,1.820899e-07,1.820904e-07,1.820910e-07,1.820915e-07,1.820921e-07,1.820926e-07,1.820931e-07,1.820937e-07,1.820942e-07,1.820948e-07,1.820953e-07,1.820958e-07,1.820964e-07,1.820969e-07,1.820975e-07,1.820980e-07,1.820985e-07,1.820991e-07,1.820996e-07,1.821002e-07,1.821007e-07,1.821012e-07,1.821018e-07,1.821023e-07,1.821029e-07,1.821034e-07,1.821039e-07,1.821045e-07,1.821050e-07,1.821056e-07,1.821061e-07,1.821066e-07,1.821072e-07,1.821077e-07,1.821083e-07,1.821088e-07,1.821093e-07,1.821099e-07,1.821104e-07,1.821110e-07,1.821115e-07,1.821120e-07,1.821126e-07,1.821131e-07,1.821137e-07,1.821142e-07,1.821147e-07,1.821153e-07,1.821158e-07,1.821163e-07,1.821169e-07,1.821174e-07,1.821180e-07,1.821185e-07,1.821190e-07,1.821196e-07,1.821201e-07,1.821207e-07,1.821212e-07,1.821217e-07,1.821223e-07,1.821228e-07,1.821234e-07,1.821239e-07,1.821244e-07,1.821250e-07,1.821255e-07,1.821260e-07,1.821266e-07,1.821271e-07,1.821277e-07,1.821282e-07,1.821287e-07,1.821293e-07,1.821298e-07,1.821304e-07,1.821309e-07,1.821314e-07,1.821320e-07,1.821325e-07,1.821331e-07,1.821336e-07,1.821341e-07,1.821347e-07,1.821352e-07,1.821357e-07,1.821363e-07,1.821368e-07,1.821374e-07,1.821379e-07,1.821384e-07,1.821390e-07,1.821395e-07,1.821400e-07,1.821406e-07,1.821411e-07,1.821417e-07,1.821422e-07,1.821427e-07,1.821433e-07,1.821438e-07,1.821444e-07,1.821449e-07,1.821454e-07,1.821460e-07,1.821465e-07,1.821470e-07,1.821476e-07,1.821481e-07,1.821487e-07,1.821492e-07,1.821497e-07,1.821503e-07,1.821508e-07,1.821513e-07,1.821519e-07,1.821524e-07,1.821530e-07,1.821535e-07,1.821540e-07,1.821546e-07,1.821551e-07,1.821556e-07,1.821562e-07,1.821567e-07,1.821573e-07,1.821578e-07,1.821583e-07,1.821589e-07,1.821594e-07,1.821599e-07,1.821605e-07,1.821610e-07,1.821615e-07,1.821621e-07,1.821626e-07,1.821632e-07,1.821637e-07,1.821642e-07,1.821648e-07,1.821653e-07,1.821658e-07,1.821664e-07,1.821669e-07,1.821675e-07,1.821680e-07,1.821685e-07,1.821691e-07,1.821696e-07,1.821701e-07,1.821707e-07,1.821712e-07,1.821717e-07,1.821723e-07,1.821728e-07,1.821734e-07,1.821739e-07,1.821744e-07,1.821750e-07,1.821755e-07,1.821760e-07,1.821766e-07,1.821771e-07,1.821776e-07,1.821782e-07,1.821787e-07,1.821793e-07,1.821798e-07,1.821803e-07,1.821809e-07,1.821814e-07,1.821819e-07,1.821825e-07,1.821830e-07,1.821835e-07,1.821841e-07,1.821846e-07,1.821852e-07,1.821857e-07,1.821862e-07,1.821868e-07,1.821873e-07,1.821878e-07,1.821884e-07,1.821889e-07,1.821894e-07,1.821900e-07,1.821905e-07,1.821911e-07,1.821916e-07,1.821921e-07,1.821927e-07,1.821932e-07,1.821937e-07,1.821943e-07,1.821948e-07,1.821953e-07,1.821959e-07,1.821964e-07,1.821969e-07,1.821975e-07,1.821980e-07,1.821985e-07,1.821991e-07,1.821996e-07,1.822002e-07,1.822007e-07,1.822012e-07,1.822018e-07,1.822023e-07,1.822028e-07,1.822034e-07,1.822039e-07,1.822044e-07,1.822050e-07,1.822055e-07,1.822060e-07,1.822066e-07,1.822071e-07,1.822076e-07,1.822082e-07,1.822087e-07,1.822092e-07,1.822098e-07,1.822103e-07,1.822109e-07,1.822114e-07,1.822119e-07,1.822125e-07,1.822130e-07,1.822135e-07,1.822141e-07,1.822146e-07,1.822151e-07,1.822157e-07,1.822162e-07,1.822167e-07,1.822173e-07,1.822178e-07,1.822183e-07,1.822189e-07,1.822194e-07,1.822199e-07,1.822205e-07,1.822210e-07,1.822215e-07,1.822221e-07,1.822226e-07,1.822231e-07,1.822237e-07,1.822242e-07,1.822248e-07,1.822253e-07,1.822258e-07,1.822264e-07,1.822269e-07,1.822274e-07,1.822280e-07,1.822285e-07,1.822290e-07,1.822296e-07,1.822301e-07,1.822306e-07,1.822312e-07,1.822317e-07,1.822322e-07,1.822328e-07,1.822333e-07,1.822338e-07,1.822344e-07,1.822349e-07,1.822354e-07,1.822360e-07,1.822365e-07,1.822370e-07,1.822376e-07,1.822381e-07,1.822386e-07,1.822392e-07,1.822397e-07,1.822402e-07,1.822408e-07,1.822413e-07,1.822418e-07,1.822424e-07,1.822429e-07,1.822434e-07,1.822440e-07,1.822445e-07,1.822450e-07,1.822456e-07,1.822461e-07,1.822466e-07,1.822472e-07,1.822477e-07,1.822482e-07,1.822488e-07,1.822493e-07,1.822498e-07,1.822504e-07,1.822509e-07,1.822514e-07,1.822520e-07,1.822525e-07,1.822530e-07,1.822536e-07,1.822541e-07,1.822546e-07,1.822552e-07,1.822557e-07,1.822562e-07,1.822568e-07,1.822573e-07,1.822578e-07,1.822584e-07,1.822589e-07,1.822594e-07,1.822600e-07,1.822605e-07,1.822610e-07,1.822615e-07,1.822621e-07,1.822626e-07,1.822631e-07,1.822637e-07,1.822642e-07,1.822647e-07,1.822653e-07,1.822658e-07,1.822663e-07,1.822669e-07,1.822674e-07,1.822679e-07,1.822685e-07,1.822690e-07,1.822695e-07,1.822701e-07,1.822706e-07,1.822711e-07,1.822717e-07,1.822722e-07,1.822727e-07,1.822733e-07,1.822738e-07,1.822743e-07,1.822749e-07,1.822754e-07,1.822759e-07,1.822764e-07,1.822770e-07,1.822775e-07,1.822780e-07,1.822786e-07,1.822791e-07,1.822796e-07,1.822802e-07,1.822807e-07,1.822812e-07,1.822818e-07,1.822823e-07,1.822828e-07,1.822834e-07,1.822839e-07,1.822844e-07,1.822850e-07,1.822855e-07,1.822860e-07,1.822865e-07,1.822871e-07,1.822876e-07,1.822881e-07,1.822887e-07,1.822892e-07,1.822897e-07,1.822903e-07,1.822908e-07,1.822913e-07,1.822919e-07,1.822924e-07,1.822929e-07,1.822935e-07,1.822940e-07,1.822945e-07,1.822950e-07,1.822956e-07,1.822961e-07,1.822966e-07,1.822972e-07,1.822977e-07,1.822982e-07,1.822988e-07,1.822993e-07,1.822998e-07,1.823004e-07,1.823009e-07,1.823014e-07,1.823019e-07,1.823025e-07,1.823030e-07,1.823035e-07,1.823041e-07,1.823046e-07,1.823051e-07,1.823057e-07,1.823062e-07,1.823067e-07,1.823073e-07,1.823078e-07,1.823083e-07,1.823088e-07,1.823094e-07,1.823099e-07,1.823104e-07,1.823110e-07,1.823115e-07,1.823120e-07,1.823126e-07,1.823131e-07,1.823136e-07,1.823141e-07,1.823147e-07,1.823152e-07,1.823157e-07,1.823163e-07,1.823168e-07,1.823173e-07,1.823179e-07,1.823184e-07,1.823189e-07,1.823194e-07,1.823200e-07,1.823205e-07,1.823210e-07,1.823216e-07,1.823221e-07,1.823226e-07,1.823232e-07,1.823237e-07,1.823242e-07,1.823247e-07,1.823253e-07,1.823258e-07,1.823263e-07,1.823269e-07,1.823274e-07,1.823279e-07,1.823284e-07,1.823290e-07,1.823295e-07,1.823300e-07,1.823306e-07,1.823311e-07,1.823316e-07,1.823322e-07,1.823327e-07,1.823332e-07,1.823337e-07,1.823343e-07,1.823348e-07,1.823353e-07,1.823359e-07,1.823364e-07,1.823369e-07,1.823374e-07,1.823380e-07,1.823385e-07,1.823390e-07,1.823396e-07,1.823401e-07,1.823406e-07,1.823411e-07,1.823417e-07,1.823422e-07,1.823427e-07,1.823433e-07,1.823438e-07,1.823443e-07,1.823448e-07,1.823454e-07,1.823459e-07,1.823464e-07,1.823470e-07,1.823475e-07,1.823480e-07,1.823485e-07,1.823491e-07,1.823496e-07,1.823501e-07,1.823507e-07,1.823512e-07,1.823517e-07,1.823522e-07,1.823528e-07,1.823533e-07,1.823538e-07,1.823544e-07,1.823549e-07,1.823554e-07,1.823559e-07,1.823565e-07,1.823570e-07,1.823575e-07,1.823581e-07,1.823586e-07,1.823591e-07,1.823596e-07,1.823602e-07,1.823607e-07,1.823612e-07,1.823618e-07,1.823623e-07,1.823628e-07,1.823633e-07,1.823639e-07,1.823644e-07,1.823649e-07,1.823654e-07,1.823660e-07,1.823665e-07,1.823670e-07,1.823676e-07,1.823681e-07,1.823686e-07,1.823691e-07,1.823697e-07,1.823702e-07,1.823707e-07,1.823713e-07,1.823718e-07,1.823723e-07,1.823728e-07,1.823734e-07,1.823739e-07,1.823744e-07,1.823749e-07,1.823755e-07,1.823760e-07,1.823765e-07,1.823771e-07,1.823776e-07,1.823781e-07,1.823786e-07,1.823792e-07,1.823797e-07,1.823802e-07,1.823807e-07,1.823813e-07,1.823818e-07,1.823823e-07,1.823829e-07,1.823834e-07,1.823839e-07,1.823844e-07,1.823850e-07,1.823855e-07,1.823860e-07,1.823865e-07,1.823871e-07,1.823876e-07,1.823881e-07,1.823886e-07,1.823892e-07,1.823897e-07,1.823902e-07,1.823908e-07,1.823913e-07,1.823918e-07,1.823923e-07,1.823929e-07,1.823934e-07,1.823939e-07,1.823944e-07,1.823950e-07,1.823955e-07,1.823960e-07,1.823965e-07,1.823971e-07,1.823976e-07,1.823981e-07,1.823987e-07,1.823992e-07,1.823997e-07,1.824002e-07,1.824008e-07,1.824013e-07,1.824018e-07,1.824023e-07,1.824029e-07,1.824034e-07,1.824039e-07,1.824044e-07,1.824050e-07,1.824055e-07,1.824060e-07,1.824065e-07,1.824071e-07,1.824076e-07,1.824081e-07,1.824086e-07,1.824092e-07,1.824097e-07,1.824102e-07,1.824107e-07,1.824113e-07,1.824118e-07,1.824123e-07,1.824129e-07,1.824134e-07,1.824139e-07,1.824144e-07,1.824150e-07,1.824155e-07,1.824160e-07,1.824165e-07,1.824171e-07,1.824176e-07,1.824181e-07,1.824186e-07,1.824192e-07,1.824197e-07,1.824202e-07,1.824207e-07,1.824213e-07,1.824218e-07,1.824223e-07,1.824228e-07,1.824234e-07,1.824239e-07,1.824244e-07,1.824249e-07,1.824255e-07,1.824260e-07,1.824265e-07,1.824270e-07,1.824276e-07,1.824281e-07,1.824286e-07,1.824291e-07,1.824297e-07,1.824302e-07,1.824307e-07,1.824312e-07,1.824318e-07,1.824323e-07,1.824328e-07,1.824333e-07,1.824339e-07,1.824344e-07,1.824349e-07,1.824354e-07,1.824360e-07,1.824365e-07,1.824370e-07,1.824375e-07,1.824381e-07,1.824386e-07,1.824391e-07,1.824396e-07,1.824402e-07,1.824407e-07,1.824412e-07,1.824417e-07,1.824422e-07,1.824428e-07,1.824433e-07,1.824438e-07,1.824443e-07,1.824449e-07,1.824454e-07,1.824459e-07,1.824464e-07,1.824470e-07,1.824475e-07,1.824480e-07,1.824485e-07,1.824491e-07,1.824496e-07,1.824501e-07,1.824506e-07,1.824512e-07,1.824517e-07,1.824522e-07,1.824527e-07,1.824533e-07,1.824538e-07,1.824543e-07,1.824548e-07,1.824553e-07,1.824559e-07,1.824564e-07,1.824569e-07,1.824574e-07,1.824580e-07,1.824585e-07,1.824590e-07,1.824595e-07,1.824601e-07,1.824606e-07,1.824611e-07,1.824616e-07,1.824622e-07,1.824627e-07,1.824632e-07,1.824637e-07,1.824642e-07,1.824648e-07,1.824653e-07,1.824658e-07,1.824663e-07,1.824669e-07,1.824674e-07,1.824679e-07,1.824684e-07,1.824690e-07,1.824695e-07,1.824700e-07,1.824705e-07,1.824710e-07,1.824716e-07,1.824721e-07,1.824726e-07,1.824731e-07,1.824737e-07,1.824742e-07,1.824747e-07,1.824752e-07,1.824758e-07,1.824763e-07,1.824768e-07,1.824773e-07,1.824778e-07,1.824784e-07,1.824789e-07,1.824794e-07,1.824799e-07,1.824805e-07,1.824810e-07,1.824815e-07,1.824820e-07,1.824825e-07,1.824831e-07,1.824836e-07,1.824841e-07,1.824846e-07,1.824852e-07,1.824857e-07,1.824862e-07,1.824867e-07,1.824872e-07,1.824878e-07,1.824883e-07,1.824888e-07,1.824893e-07,1.824899e-07,1.824904e-07,1.824909e-07,1.824914e-07,1.824919e-07,1.824925e-07,1.824930e-07,1.824935e-07,1.824940e-07,1.824946e-07,1.824951e-07,1.824956e-07,1.824961e-07,1.824966e-07,1.824972e-07,1.824977e-07,1.824982e-07,1.824987e-07,1.824993e-07,1.824998e-07,1.825003e-07,1.825008e-07,1.825013e-07,1.825019e-07,1.825024e-07,1.825029e-07,1.825034e-07,1.825040e-07,1.825045e-07,1.825050e-07,1.825055e-07,1.825060e-07,1.825066e-07,1.825071e-07,1.825076e-07,1.825081e-07,1.825086e-07,1.825092e-07,1.825097e-07,1.825102e-07,1.825107e-07,1.825112e-07,1.825118e-07,1.825123e-07,1.825128e-07,1.825133e-07,1.825139e-07,1.825144e-07,1.825149e-07,1.825154e-07,1.825159e-07,1.825165e-07,1.825170e-07,1.825175e-07,1.825180e-07,1.825185e-07,1.825191e-07,1.825196e-07,1.825201e-07,1.825206e-07,1.825211e-07,1.825217e-07,1.825222e-07,1.825227e-07,1.825232e-07,1.825238e-07,1.825243e-07,1.825248e-07,1.825253e-07,1.825258e-07,1.825264e-07,1.825269e-07,1.825274e-07,1.825279e-07,1.825284e-07,1.825290e-07,1.825295e-07,1.825300e-07,1.825305e-07,1.825310e-07,1.825316e-07,1.825321e-07,1.825326e-07,1.825331e-07,1.825336e-07,1.825342e-07,1.825347e-07,1.825352e-07,1.825357e-07,1.825362e-07,1.825368e-07,1.825373e-07,1.825378e-07,1.825383e-07,1.825388e-07,1.825394e-07,1.825399e-07,1.825404e-07,1.825409e-07,1.825414e-07,1.825420e-07,1.825425e-07,1.825430e-07,1.825435e-07,1.825440e-07,1.825446e-07,1.825451e-07,1.825456e-07,1.825461e-07,1.825466e-07,1.825472e-07,1.825477e-07,1.825482e-07,1.825487e-07,1.825492e-07,1.825498e-07,1.825503e-07,1.825508e-07,1.825513e-07,1.825518e-07,1.825524e-07,1.825529e-07,1.825534e-07,1.825539e-07,1.825544e-07,1.825549e-07,1.825555e-07,1.825560e-07,1.825565e-07,1.825570e-07,1.825575e-07,1.825581e-07,1.825586e-07,1.825591e-07,1.825596e-07,1.825601e-07,1.825607e-07,1.825612e-07,1.825617e-07,1.825622e-07,1.825627e-07,1.825633e-07,1.825638e-07,1.825643e-07,1.825648e-07,1.825653e-07,1.825658e-07,1.825664e-07,1.825669e-07,1.825674e-07,1.825679e-07,1.825684e-07,1.825690e-07,1.825695e-07,1.825700e-07,1.825705e-07,1.825710e-07,1.825716e-07,1.825721e-07,1.825726e-07,1.825731e-07,1.825736e-07,1.825741e-07,1.825747e-07,1.825752e-07,1.825757e-07,1.825762e-07,1.825767e-07,1.825773e-07,1.825778e-07,1.825783e-07,1.825788e-07,1.825793e-07,1.825798e-07,1.825804e-07,1.825809e-07,1.825814e-07,1.825819e-07,1.825824e-07,1.825830e-07,1.825835e-07,1.825840e-07,1.825845e-07,1.825850e-07,1.825855e-07,1.825861e-07,1.825866e-07,1.825871e-07,1.825876e-07,1.825881e-07,1.825887e-07,1.825892e-07,1.825897e-07,1.825902e-07,1.825907e-07,1.825912e-07,1.825918e-07,1.825923e-07,1.825928e-07,1.825933e-07,1.825938e-07,1.825943e-07,1.825949e-07,1.825954e-07,1.825959e-07,1.825964e-07,1.825969e-07,1.825974e-07,1.825980e-07,1.825985e-07,1.825990e-07,1.825995e-07,1.826000e-07,1.826006e-07,1.826011e-07,1.826016e-07,1.826021e-07,1.826026e-07,1.826031e-07,1.826037e-07,1.826042e-07,1.826047e-07,1.826052e-07,1.826057e-07,1.826062e-07,1.826068e-07,1.826073e-07,1.826078e-07,1.826083e-07,1.826088e-07,1.826093e-07,1.826099e-07,1.826104e-07,1.826109e-07,1.826114e-07,1.826119e-07,1.826124e-07,1.826130e-07,1.826135e-07,1.826140e-07,1.826145e-07,1.826150e-07,1.826155e-07,1.826161e-07,1.826166e-07,1.826171e-07,1.826176e-07,1.826181e-07,1.826186e-07,1.826192e-07,1.826197e-07,1.826202e-07,1.826207e-07,1.826212e-07,1.826217e-07,1.826223e-07,1.826228e-07,1.826233e-07,1.826238e-07,1.826243e-07,1.826248e-07,1.826254e-07,1.826259e-07,1.826264e-07,1.826269e-07,1.826274e-07,1.826279e-07,1.826284e-07,1.826290e-07,1.826295e-07,1.826300e-07,1.826305e-07,1.826310e-07,1.826315e-07,1.826321e-07,1.826326e-07,1.826331e-07,1.826336e-07,1.826341e-07,1.826346e-07,1.826352e-07,1.826357e-07,1.826362e-07,1.826367e-07,1.826372e-07,1.826377e-07,1.826382e-07,1.826388e-07,1.826393e-07,1.826398e-07,1.826403e-07,1.826408e-07,1.826413e-07,1.826419e-07,1.826424e-07,1.826429e-07,1.826434e-07,1.826439e-07,1.826444e-07,1.826449e-07,1.826455e-07,1.826460e-07,1.826465e-07,1.826470e-07,1.826475e-07,1.826480e-07,1.826486e-07,1.826491e-07,1.826496e-07,1.826501e-07,1.826506e-07,1.826511e-07,1.826516e-07,1.826522e-07,1.826527e-07,1.826532e-07,1.826537e-07,1.826542e-07,1.826547e-07,1.826552e-07,1.826558e-07,1.826563e-07,1.826568e-07,1.826573e-07,1.826578e-07,1.826583e-07,1.826589e-07,1.826594e-07,1.826599e-07,1.826604e-07,1.826609e-07,1.826614e-07,1.826619e-07,1.826625e-07,1.826630e-07,1.826635e-07,1.826640e-07,1.826645e-07,1.826650e-07,1.826655e-07,1.826661e-07,1.826666e-07,1.826671e-07,1.826676e-07,1.826681e-07,1.826686e-07,1.826691e-07,1.826697e-07,1.826702e-07,1.826707e-07,1.826712e-07,1.826717e-07,1.826722e-07,1.826727e-07,1.826733e-07,1.826738e-07,1.826743e-07,1.826748e-07,1.826753e-07,1.826758e-07,1.826763e-07,1.826769e-07,1.826774e-07,1.826779e-07,1.826784e-07,1.826789e-07,1.826794e-07,1.826799e-07,1.826804e-07,1.826810e-07,1.826815e-07,1.826820e-07,1.826825e-07,1.826830e-07,1.826835e-07,1.826840e-07,1.826846e-07,1.826851e-07,1.826856e-07,1.826861e-07,1.826866e-07,1.826871e-07,1.826876e-07,1.826882e-07,1.826887e-07,1.826892e-07,1.826897e-07,1.826902e-07,1.826907e-07,1.826912e-07,1.826917e-07,1.826923e-07,1.826928e-07,1.826933e-07,1.826938e-07,1.826943e-07,1.826948e-07,1.826953e-07,1.826958e-07,1.826964e-07,1.826969e-07,1.826974e-07,1.826979e-07,1.826984e-07,1.826989e-07,1.826994e-07,1.827000e-07,1.827005e-07,1.827010e-07,1.827015e-07,1.827020e-07,1.827025e-07,1.827030e-07,1.827035e-07,1.827041e-07,1.827046e-07,1.827051e-07,1.827056e-07,1.827061e-07,1.827066e-07,1.827071e-07,1.827076e-07,1.827082e-07,1.827087e-07,1.827092e-07,1.827097e-07,1.827102e-07,1.827107e-07,1.827112e-07,1.827117e-07,1.827123e-07,1.827128e-07,1.827133e-07,1.827138e-07,1.827143e-07,1.827148e-07,1.827153e-07,1.827158e-07,1.827164e-07,1.827169e-07,1.827174e-07,1.827179e-07,1.827184e-07,1.827189e-07,1.827194e-07,1.827199e-07,1.827204e-07,1.827210e-07,1.827215e-07,1.827220e-07,1.827225e-07,1.827230e-07,1.827235e-07,1.827240e-07,1.827245e-07,1.827251e-07,1.827256e-07,1.827261e-07,1.827266e-07,1.827271e-07,1.827276e-07,1.827281e-07,1.827286e-07,1.827291e-07,1.827297e-07,1.827302e-07,1.827307e-07,1.827312e-07,1.827317e-07,1.827322e-07,1.827327e-07,1.827332e-07,1.827337e-07,1.827343e-07,1.827348e-07,1.827353e-07,1.827358e-07,1.827363e-07,1.827368e-07,1.827373e-07,1.827378e-07,1.827384e-07,1.827389e-07,1.827394e-07,1.827399e-07,1.827404e-07,1.827409e-07,1.827414e-07,1.827419e-07,1.827424e-07,1.827430e-07,1.827435e-07,1.827440e-07,1.827445e-07,1.827450e-07,1.827455e-07,1.827460e-07,1.827465e-07,1.827470e-07,1.827475e-07,1.827481e-07,1.827486e-07,1.827491e-07,1.827496e-07,1.827501e-07,1.827506e-07,1.827511e-07,1.827516e-07,1.827521e-07,1.827527e-07,1.827532e-07,1.827537e-07,1.827542e-07,1.827547e-07,1.827552e-07,1.827557e-07,1.827562e-07,1.827567e-07,1.827572e-07,1.827578e-07,1.827583e-07,1.827588e-07,1.827593e-07,1.827598e-07,1.827603e-07,1.827608e-07,1.827613e-07,1.827618e-07,1.827624e-07,1.827629e-07,1.827634e-07,1.827639e-07,1.827644e-07,1.827649e-07,1.827654e-07,1.827659e-07,1.827664e-07,1.827669e-07,1.827675e-07,1.827680e-07,1.827685e-07,1.827690e-07,1.827695e-07,1.827700e-07,1.827705e-07,1.827710e-07,1.827715e-07,1.827720e-07,1.827725e-07,1.827731e-07,1.827736e-07,1.827741e-07,1.827746e-07,1.827751e-07,1.827756e-07,1.827761e-07,1.827766e-07,1.827771e-07,1.827776e-07,1.827782e-07,1.827787e-07,1.827792e-07,1.827797e-07,1.827802e-07,1.827807e-07,1.827812e-07,1.827817e-07,1.827822e-07,1.827827e-07,1.827832e-07,1.827838e-07,1.827843e-07,1.827848e-07,1.827853e-07,1.827858e-07,1.827863e-07,1.827868e-07,1.827873e-07,1.827878e-07,1.827883e-07,1.827888e-07,1.827894e-07,1.827899e-07,1.827904e-07,1.827909e-07,1.827914e-07,1.827919e-07,1.827924e-07,1.827929e-07,1.827934e-07,1.827939e-07,1.827944e-07,1.827950e-07,1.827955e-07,1.827960e-07,1.827965e-07,1.827970e-07,1.827975e-07,1.827980e-07,1.827985e-07,1.827990e-07,1.827995e-07,1.828000e-07,1.828005e-07,1.828011e-07,1.828016e-07,1.828021e-07,1.828026e-07,1.828031e-07,1.828036e-07,1.828041e-07,1.828046e-07,1.828051e-07,1.828056e-07,1.828061e-07,1.828066e-07,1.828072e-07,1.828077e-07,1.828082e-07,1.828087e-07,1.828092e-07,1.828097e-07,1.828102e-07,1.828107e-07,1.828112e-07,1.828117e-07,1.828122e-07,1.828127e-07,1.828132e-07,1.828138e-07,1.828143e-07,1.828148e-07,1.828153e-07,1.828158e-07,1.828163e-07,1.828168e-07,1.828173e-07,1.828178e-07,1.828183e-07,1.828188e-07,1.828193e-07,1.828198e-07,1.828204e-07,1.828209e-07,1.828214e-07,1.828219e-07,1.828224e-07,1.828229e-07,1.828234e-07,1.828239e-07,1.828244e-07,1.828249e-07,1.828254e-07,1.828259e-07,1.828264e-07,1.828270e-07,1.828275e-07,1.828280e-07,1.828285e-07,1.828290e-07,1.828295e-07,1.828300e-07,1.828305e-07,1.828310e-07,1.828315e-07,1.828320e-07,1.828325e-07,1.828330e-07,1.828335e-07,1.828341e-07,1.828346e-07,1.828351e-07,1.828356e-07,1.828361e-07,1.828366e-07,1.828371e-07,1.828376e-07,1.828381e-07,1.828386e-07,1.828391e-07,1.828396e-07,1.828401e-07,1.828406e-07,1.828411e-07,1.828417e-07,1.828422e-07,1.828427e-07,1.828432e-07,1.828437e-07,1.828442e-07,1.828447e-07,1.828452e-07,1.828457e-07,1.828462e-07,1.828467e-07,1.828472e-07,1.828477e-07,1.828482e-07,1.828487e-07,1.828493e-07,1.828498e-07,1.828503e-07,1.828508e-07,1.828513e-07,1.828518e-07,1.828523e-07,1.828528e-07,1.828533e-07,1.828538e-07,1.828543e-07,1.828548e-07,1.828553e-07,1.828558e-07,1.828563e-07,1.828568e-07,1.828574e-07,1.828579e-07,1.828584e-07,1.828589e-07,1.828594e-07,1.828599e-07,1.828604e-07,1.828609e-07,1.828614e-07,1.828619e-07,1.828624e-07,1.828629e-07,1.828634e-07,1.828639e-07,1.828644e-07,1.828649e-07,1.828654e-07,1.828659e-07,1.828665e-07,1.828670e-07,1.828675e-07,1.828680e-07,1.828685e-07,1.828690e-07,1.828695e-07,1.828700e-07,1.828705e-07,1.828710e-07,1.828715e-07,1.828720e-07,1.828725e-07,1.828730e-07,1.828735e-07,1.828740e-07,1.828745e-07,1.828750e-07,1.828756e-07,1.828761e-07,1.828766e-07,1.828771e-07,1.828776e-07,1.828781e-07,1.828786e-07,1.828791e-07,1.828796e-07,1.828801e-07,1.828806e-07,1.828811e-07,1.828816e-07,1.828821e-07,1.828826e-07,1.828831e-07,1.828836e-07,1.828841e-07,1.828846e-07,1.828851e-07,1.828857e-07,1.828862e-07,1.828867e-07,1.828872e-07,1.828877e-07,1.828882e-07,1.828887e-07,1.828892e-07,1.828897e-07,1.828902e-07,1.828907e-07,1.828912e-07,1.828917e-07,1.828922e-07,1.828927e-07,1.828932e-07,1.828937e-07,1.828942e-07,1.828947e-07,1.828952e-07,1.828957e-07,1.828962e-07,1.828967e-07,1.828973e-07,1.828978e-07,1.828983e-07,1.828988e-07,1.828993e-07,1.828998e-07,1.829003e-07,1.829008e-07,1.829013e-07,1.829018e-07,1.829023e-07,1.829028e-07,1.829033e-07,1.829038e-07,1.829043e-07,1.829048e-07,1.829053e-07,1.829058e-07,1.829063e-07,1.829068e-07,1.829073e-07,1.829078e-07,1.829083e-07,1.829088e-07,1.829093e-07,1.829099e-07,1.829104e-07,1.829109e-07,1.829114e-07,1.829119e-07,1.829124e-07,1.829129e-07,1.829134e-07,1.829139e-07,1.829144e-07,1.829149e-07,1.829154e-07,1.829159e-07,1.829164e-07,1.829169e-07,1.829174e-07,1.829179e-07,1.829184e-07,1.829189e-07,1.829194e-07,1.829199e-07,1.829204e-07,1.829209e-07,1.829214e-07,1.829219e-07,1.829224e-07,1.829229e-07,1.829234e-07,1.829239e-07,1.829245e-07,1.829250e-07,1.829255e-07,1.829260e-07,1.829265e-07,1.829270e-07,1.829275e-07,1.829280e-07,1.829285e-07,1.829290e-07,1.829295e-07,1.829300e-07,1.829305e-07,1.829310e-07,1.829315e-07,1.829320e-07,1.829325e-07,1.829330e-07,1.829335e-07,1.829340e-07,1.829345e-07,1.829350e-07,1.829355e-07,1.829360e-07,1.829365e-07,1.829370e-07,1.829375e-07,1.829380e-07,1.829385e-07,1.829390e-07,1.829395e-07,1.829400e-07,1.829405e-07,1.829410e-07,1.829415e-07,1.829420e-07,1.829425e-07,1.829430e-07,1.829436e-07,1.829441e-07,1.829446e-07,1.829451e-07,1.829456e-07,1.829461e-07,1.829466e-07,1.829471e-07,1.829476e-07,1.829481e-07,1.829486e-07,1.829491e-07,1.829496e-07,1.829501e-07,1.829506e-07,1.829511e-07,1.829516e-07,1.829521e-07,1.829526e-07,1.829531e-07,1.829536e-07,1.829541e-07,1.829546e-07,1.829551e-07,1.829556e-07,1.829561e-07,1.829566e-07,1.829571e-07,1.829576e-07,1.829581e-07,1.829586e-07,1.829591e-07,1.829596e-07,1.829601e-07,1.829606e-07,1.829611e-07,1.829616e-07,1.829621e-07,1.829626e-07,1.829631e-07,1.829636e-07,1.829641e-07,1.829646e-07,1.829651e-07,1.829656e-07,1.829661e-07,1.829666e-07,1.829671e-07,1.829676e-07,1.829681e-07,1.829686e-07,1.829691e-07,1.829696e-07,1.829701e-07,1.829706e-07,1.829711e-07,1.829716e-07,1.829721e-07,1.829726e-07,1.829731e-07,1.829736e-07,1.829741e-07,1.829746e-07,1.829751e-07,1.829756e-07,1.829762e-07,1.829767e-07,1.829772e-07,1.829777e-07,1.829782e-07,1.829787e-07,1.829792e-07,1.829797e-07,1.829802e-07,1.829807e-07,1.829812e-07,1.829817e-07,1.829822e-07,1.829827e-07,1.829832e-07,1.829837e-07,1.829842e-07,1.829847e-07,1.829852e-07,1.829857e-07,1.829862e-07,1.829867e-07,1.829872e-07,1.829877e-07,1.829882e-07,1.829887e-07,1.829892e-07,1.829897e-07,1.829902e-07,1.829907e-07,1.829912e-07,1.829917e-07,1.829922e-07,1.829927e-07,1.829932e-07,1.829937e-07,1.829942e-07,1.829947e-07,1.829952e-07,1.829957e-07,1.829962e-07,1.829967e-07,1.829972e-07,1.829977e-07,1.829982e-07,1.829987e-07,1.829992e-07,1.829997e-07,1.830002e-07,1.830007e-07,1.830012e-07,1.830017e-07,1.830022e-07,1.830027e-07,1.830032e-07,1.830037e-07,1.830042e-07,1.830047e-07,1.830052e-07,1.830057e-07,1.830062e-07,1.830067e-07,1.830072e-07,1.830077e-07,1.830082e-07,1.830087e-07,1.830092e-07,1.830097e-07,1.830102e-07,1.830107e-07,1.830112e-07,1.830117e-07,1.830122e-07,1.830127e-07,1.830132e-07,1.830137e-07,1.830142e-07,1.830147e-07,1.830152e-07,1.830156e-07,1.830161e-07,1.830166e-07,1.830171e-07,1.830176e-07,1.830181e-07,1.830186e-07,1.830191e-07,1.830196e-07,1.830201e-07,1.830206e-07,1.830211e-07,1.830216e-07,1.830221e-07,1.830226e-07,1.830231e-07,1.830236e-07,1.830241e-07,1.830246e-07,1.830251e-07,1.830256e-07,1.830261e-07,1.830266e-07,1.830271e-07,1.830276e-07,1.830281e-07,1.830286e-07,1.830291e-07,1.830296e-07,1.830301e-07,1.830306e-07,1.830311e-07,1.830316e-07,1.830321e-07,1.830326e-07,1.830331e-07,1.830336e-07,1.830341e-07,1.830346e-07,1.830351e-07,1.830356e-07,1.830361e-07,1.830366e-07,1.830371e-07,1.830376e-07,1.830381e-07,1.830386e-07,1.830391e-07,1.830396e-07,1.830401e-07,1.830406e-07,1.830411e-07,1.830416e-07,1.830421e-07,1.830426e-07,1.830431e-07,1.830436e-07,1.830441e-07,1.830446e-07,1.830451e-07,1.830456e-07,1.830461e-07,1.830466e-07,1.830471e-07,1.830476e-07,1.830480e-07,1.830485e-07,1.830490e-07,1.830495e-07,1.830500e-07,1.830505e-07,1.830510e-07,1.830515e-07,1.830520e-07,1.830525e-07,1.830530e-07,1.830535e-07,1.830540e-07,1.830545e-07,1.830550e-07,1.830555e-07,1.830560e-07,1.830565e-07,1.830570e-07,1.830575e-07,1.830580e-07,1.830585e-07,1.830590e-07,1.830595e-07,1.830600e-07,1.830605e-07,1.830610e-07,1.830615e-07,1.830620e-07,1.830625e-07,1.830630e-07,1.830635e-07,1.830640e-07,1.830645e-07,1.830650e-07,1.830655e-07,1.830660e-07,1.830665e-07,1.830669e-07,1.830674e-07,1.830679e-07,1.830684e-07,1.830689e-07,1.830694e-07,1.830699e-07,1.830704e-07,1.830709e-07,1.830714e-07,1.830719e-07,1.830724e-07,1.830729e-07,1.830734e-07,1.830739e-07,1.830744e-07,1.830749e-07,1.830754e-07,1.830759e-07,1.830764e-07,1.830769e-07,1.830774e-07,1.830779e-07,1.830784e-07,1.830789e-07,1.830794e-07,1.830799e-07,1.830804e-07,1.830809e-07,1.830814e-07,1.830818e-07,1.830823e-07,1.830828e-07,1.830833e-07,1.830838e-07,1.830843e-07,1.830848e-07,1.830853e-07,1.830858e-07,1.830863e-07,1.830868e-07,1.830873e-07,1.830878e-07,1.830883e-07,1.830888e-07,1.830893e-07,1.830898e-07,1.830903e-07,1.830908e-07,1.830913e-07,1.830918e-07,1.830923e-07,1.830928e-07,1.830933e-07,1.830938e-07,1.830942e-07,1.830947e-07,1.830952e-07,1.830957e-07,1.830962e-07,1.830967e-07,1.830972e-07,1.830977e-07,1.830982e-07,1.830987e-07,1.830992e-07,1.830997e-07,1.831002e-07,1.831007e-07,1.831012e-07,1.831017e-07,1.831022e-07,1.831027e-07,1.831032e-07,1.831037e-07,1.831042e-07,1.831047e-07,1.831052e-07,1.831056e-07,1.831061e-07,1.831066e-07,1.831071e-07,1.831076e-07,1.831081e-07,1.831086e-07,1.831091e-07,1.831096e-07,1.831101e-07,1.831106e-07,1.831111e-07,1.831116e-07,1.831121e-07,1.831126e-07,1.831131e-07,1.831136e-07,1.831141e-07,1.831146e-07,1.831151e-07,1.831155e-07,1.831160e-07,1.831165e-07,1.831170e-07,1.831175e-07,1.831180e-07,1.831185e-07,1.831190e-07,1.831195e-07,1.831200e-07,1.831205e-07,1.831210e-07,1.831215e-07,1.831220e-07,1.831225e-07,1.831230e-07,1.831235e-07,1.831240e-07,1.831245e-07,1.831249e-07,1.831254e-07,1.831259e-07,1.831264e-07,1.831269e-07,1.831274e-07,1.831279e-07,1.831284e-07,1.831289e-07,1.831294e-07,1.831299e-07,1.831304e-07,1.831309e-07,1.831314e-07,1.831319e-07,1.831324e-07,1.831329e-07,1.831334e-07,1.831338e-07,1.831343e-07,1.831348e-07,1.831353e-07,1.831358e-07,1.831363e-07,1.831368e-07,1.831373e-07,1.831378e-07,1.831383e-07,1.831388e-07,1.831393e-07,1.831398e-07,1.831403e-07,1.831408e-07,1.831413e-07,1.831417e-07,1.831422e-07,1.831427e-07,1.831432e-07,1.831437e-07,1.831442e-07,1.831447e-07,1.831452e-07,1.831457e-07,1.831462e-07,1.831467e-07,1.831472e-07,1.831477e-07,1.831482e-07,1.831487e-07,1.831492e-07,1.831496e-07,1.831501e-07,1.831506e-07,1.831511e-07,1.831516e-07,1.831521e-07,1.831526e-07,1.831531e-07,1.831536e-07,1.831541e-07,1.831546e-07,1.831551e-07,1.831556e-07,1.831561e-07,1.831566e-07,1.831570e-07,1.831575e-07,1.831580e-07,1.831585e-07,1.831590e-07,1.831595e-07,1.831600e-07,1.831605e-07,1.831610e-07,1.831615e-07,1.831620e-07,1.831625e-07,1.831630e-07,1.831635e-07,1.831639e-07,1.831644e-07,1.831649e-07,1.831654e-07,1.831659e-07,1.831664e-07,1.831669e-07,1.831674e-07,1.831679e-07,1.831684e-07,1.831689e-07,1.831694e-07,1.831699e-07,1.831704e-07,1.831708e-07,1.831713e-07,1.831718e-07,1.831723e-07,1.831728e-07,1.831733e-07,1.831738e-07,1.831743e-07,1.831748e-07,1.831753e-07,1.831758e-07,1.831763e-07,1.831768e-07,1.831772e-07,1.831777e-07,1.831782e-07,1.831787e-07,1.831792e-07,1.831797e-07,1.831802e-07,1.831807e-07,1.831812e-07,1.831817e-07,1.831822e-07,1.831827e-07,1.831832e-07,1.831836e-07,1.831841e-07,1.831846e-07,1.831851e-07,1.831856e-07,1.831861e-07,1.831866e-07,1.831871e-07,1.831876e-07,1.831881e-07,1.831886e-07,1.831891e-07,1.831895e-07,1.831900e-07,1.831905e-07,1.831910e-07,1.831915e-07,1.831920e-07,1.831925e-07,1.831930e-07,1.831935e-07,1.831940e-07,1.831945e-07,1.831950e-07,1.831954e-07,1.831959e-07,1.831964e-07,1.831969e-07,1.831974e-07,1.831979e-07,1.831984e-07,1.831989e-07,1.831994e-07,1.831999e-07,1.832004e-07,1.832009e-07,1.832013e-07,1.832018e-07,1.832023e-07,1.832028e-07,1.832033e-07,1.832038e-07,1.832043e-07,1.832048e-07,1.832053e-07,1.832058e-07,1.832063e-07,1.832067e-07,1.832072e-07,1.832077e-07,1.832082e-07,1.832087e-07,1.832092e-07,1.832097e-07,1.832102e-07,1.832107e-07,1.832112e-07,1.832117e-07,1.832121e-07,1.832126e-07,1.832131e-07,1.832136e-07,1.832141e-07,1.832146e-07,1.832151e-07,1.832156e-07,1.832161e-07,1.832166e-07,1.832171e-07,1.832175e-07,1.832180e-07,1.832185e-07,1.832190e-07,1.832195e-07,1.832200e-07,1.832205e-07,1.832210e-07,1.832215e-07,1.832220e-07,1.832224e-07,1.832229e-07,1.832234e-07,1.832239e-07,1.832244e-07,1.832249e-07,1.832254e-07,1.832259e-07,1.832264e-07,1.832269e-07,1.832274e-07,1.832278e-07,1.832283e-07,1.832288e-07,1.832293e-07,1.832298e-07,1.832303e-07,1.832308e-07,1.832313e-07,1.832318e-07,1.832323e-07,1.832327e-07,1.832332e-07,1.832337e-07,1.832342e-07,1.832347e-07,1.832352e-07,1.832357e-07,1.832362e-07,1.832367e-07,1.832371e-07,1.832376e-07,1.832381e-07,1.832386e-07,1.832391e-07,1.832396e-07,1.832401e-07,1.832406e-07,1.832411e-07,1.832416e-07,1.832420e-07,1.832425e-07,1.832430e-07,1.832435e-07,1.832440e-07,1.832445e-07,1.832450e-07,1.832455e-07,1.832460e-07,1.832465e-07,1.832469e-07,1.832474e-07,1.832479e-07,1.832484e-07,1.832489e-07,1.832494e-07,1.832499e-07,1.832504e-07,1.832509e-07,1.832513e-07,1.832518e-07,1.832523e-07,1.832528e-07,1.832533e-07,1.832538e-07,1.832543e-07,1.832548e-07,1.832553e-07,1.832557e-07,1.832562e-07,1.832567e-07,1.832572e-07,1.832577e-07,1.832582e-07,1.832587e-07,1.832592e-07,1.832597e-07,1.832601e-07,1.832606e-07,1.832611e-07,1.832616e-07,1.832621e-07,1.832626e-07,1.832631e-07,1.832636e-07,1.832641e-07,1.832645e-07,1.832650e-07,1.832655e-07,1.832660e-07,1.832665e-07,1.832670e-07,1.832675e-07,1.832680e-07,1.832685e-07,1.832689e-07,1.832694e-07,1.832699e-07,1.832704e-07,1.832709e-07,1.832714e-07,1.832719e-07,1.832724e-07,1.832728e-07,1.832733e-07,1.832738e-07,1.832743e-07,1.832748e-07,1.832753e-07,1.832758e-07,1.832763e-07,1.832768e-07,1.832772e-07,1.832777e-07,1.832782e-07,1.832787e-07,1.832792e-07,1.832797e-07,1.832802e-07,1.832807e-07,1.832811e-07,1.832816e-07,1.832821e-07,1.832826e-07,1.832831e-07,1.832836e-07,1.832841e-07,1.832846e-07,1.832850e-07,1.832855e-07,1.832860e-07,1.832865e-07,1.832870e-07,1.832875e-07,1.832880e-07,1.832885e-07,1.832889e-07,1.832894e-07,1.832899e-07,1.832904e-07,1.832909e-07,1.832914e-07,1.832919e-07,1.832924e-07,1.832928e-07,1.832933e-07,1.832938e-07,1.832943e-07,1.832948e-07,1.832953e-07,1.832958e-07,1.832963e-07,1.832967e-07,1.832972e-07,1.832977e-07,1.832982e-07,1.832987e-07,1.832992e-07,1.832997e-07,1.833002e-07,1.833006e-07,1.833011e-07,1.833016e-07,1.833021e-07,1.833026e-07,1.833031e-07,1.833036e-07,1.833041e-07,1.833045e-07,1.833050e-07,1.833055e-07,1.833060e-07,1.833065e-07,1.833070e-07,1.833075e-07,1.833079e-07,1.833084e-07,1.833089e-07,1.833094e-07,1.833099e-07,1.833104e-07,1.833109e-07,1.833114e-07,1.833118e-07,1.833123e-07,1.833128e-07,1.833133e-07,1.833138e-07,1.833143e-07,1.833148e-07,1.833152e-07,1.833157e-07,1.833162e-07,1.833167e-07,1.833172e-07,1.833177e-07,1.833182e-07,1.833187e-07,1.833191e-07,1.833196e-07,1.833201e-07,1.833206e-07,1.833211e-07,1.833216e-07,1.833221e-07,1.833225e-07,1.833230e-07,1.833235e-07,1.833240e-07,1.833245e-07,1.833250e-07,1.833255e-07,1.833259e-07,1.833264e-07,1.833269e-07,1.833274e-07,1.833279e-07,1.833284e-07,1.833289e-07,1.833293e-07,1.833298e-07,1.833303e-07,1.833308e-07,1.833313e-07,1.833318e-07,1.833323e-07,1.833327e-07,1.833332e-07,1.833337e-07,1.833342e-07,1.833347e-07,1.833352e-07,1.833357e-07,1.833361e-07,1.833366e-07,1.833371e-07,1.833376e-07,1.833381e-07,1.833386e-07,1.833391e-07,1.833395e-07,1.833400e-07,1.833405e-07,1.833410e-07,1.833415e-07,1.833420e-07,1.833425e-07,1.833429e-07,1.833434e-07,1.833439e-07,1.833444e-07,1.833449e-07,1.833454e-07,1.833459e-07,1.833463e-07,1.833468e-07,1.833473e-07,1.833478e-07,1.833483e-07,1.833488e-07,1.833493e-07,1.833497e-07,1.833502e-07,1.833507e-07,1.833512e-07,1.833517e-07,1.833522e-07,1.833526e-07,1.833531e-07,1.833536e-07,1.833541e-07,1.833546e-07,1.833551e-07,1.833556e-07,1.833560e-07,1.833565e-07,1.833570e-07,1.833575e-07,1.833580e-07,1.833585e-07,1.833590e-07,1.833594e-07,1.833599e-07,1.833604e-07,1.833609e-07,1.833614e-07,1.833619e-07,1.833623e-07,1.833628e-07,1.833633e-07,1.833638e-07,1.833643e-07,1.833648e-07,1.833653e-07,1.833657e-07,1.833662e-07,1.833667e-07,1.833672e-07,1.833677e-07,1.833682e-07,1.833686e-07,1.833691e-07,1.833696e-07,1.833701e-07,1.833706e-07,1.833711e-07,1.833715e-07,1.833720e-07,1.833725e-07,1.833730e-07,1.833735e-07,1.833740e-07,1.833745e-07,1.833749e-07,1.833754e-07,1.833759e-07,1.833764e-07,1.833769e-07,1.833774e-07,1.833778e-07,1.833783e-07,1.833788e-07,1.833793e-07,1.833798e-07,1.833803e-07,1.833807e-07,1.833812e-07,1.833817e-07,1.833822e-07,1.833827e-07,1.833832e-07,1.833836e-07,1.833841e-07,1.833846e-07,1.833851e-07,1.833856e-07,1.833861e-07,1.833865e-07,1.833870e-07,1.833875e-07,1.833880e-07,1.833885e-07,1.833890e-07,1.833894e-07,1.833899e-07,1.833904e-07,1.833909e-07,1.833914e-07,1.833919e-07,1.833923e-07,1.833928e-07,1.833933e-07,1.833938e-07,1.833943e-07,1.833948e-07,1.833952e-07,1.833957e-07,1.833962e-07,1.833967e-07,1.833972e-07,1.833977e-07,1.833981e-07,1.833986e-07,1.833991e-07,1.833996e-07,1.834001e-07,1.834006e-07,1.834010e-07,1.834015e-07,1.834020e-07,1.834025e-07,1.834030e-07,1.834035e-07,1.834039e-07,1.834044e-07,1.834049e-07,1.834054e-07,1.834059e-07,1.834064e-07,1.834068e-07,1.834073e-07,1.834078e-07,1.834083e-07,1.834088e-07,1.834092e-07,1.834097e-07,1.834102e-07,1.834107e-07,1.834112e-07,1.834117e-07,1.834121e-07,1.834126e-07,1.834131e-07,1.834136e-07,1.834141e-07,1.834146e-07,1.834150e-07,1.834155e-07,1.834160e-07,1.834165e-07,1.834170e-07,1.834174e-07,1.834179e-07,1.834184e-07,1.834189e-07,1.834194e-07,1.834199e-07,1.834203e-07,1.834208e-07,1.834213e-07,1.834218e-07,1.834223e-07,1.834228e-07,1.834232e-07,1.834237e-07,1.834242e-07,1.834247e-07,1.834252e-07,1.834256e-07,1.834261e-07,1.834266e-07,1.834271e-07,1.834276e-07,1.834281e-07,1.834285e-07,1.834290e-07,1.834295e-07,1.834300e-07,1.834305e-07,1.834309e-07,1.834314e-07,1.834319e-07,1.834324e-07,1.834329e-07,1.834334e-07,1.834338e-07,1.834343e-07,1.834348e-07,1.834353e-07,1.834358e-07,1.834362e-07,1.834367e-07,1.834372e-07,1.834377e-07,1.834382e-07,1.834386e-07,1.834391e-07,1.834396e-07,1.834401e-07,1.834406e-07,1.834411e-07,1.834415e-07,1.834420e-07,1.834425e-07,1.834430e-07,1.834435e-07,1.834439e-07,1.834444e-07,1.834449e-07,1.834454e-07,1.834459e-07,1.834463e-07,1.834468e-07,1.834473e-07,1.834478e-07,1.834483e-07,1.834488e-07,1.834492e-07,1.834497e-07,1.834502e-07,1.834507e-07,1.834512e-07,1.834516e-07,1.834521e-07,1.834526e-07,1.834531e-07,1.834536e-07,1.834540e-07,1.834545e-07,1.834550e-07,1.834555e-07,1.834560e-07,1.834564e-07,1.834569e-07,1.834574e-07,1.834579e-07,1.834584e-07,1.834588e-07,1.834593e-07,1.834598e-07,1.834603e-07,1.834608e-07,1.834613e-07,1.834617e-07,1.834622e-07,1.834627e-07,1.834632e-07,1.834637e-07,1.834641e-07,1.834646e-07,1.834651e-07,1.834656e-07,1.834661e-07,1.834665e-07,1.834670e-07,1.834675e-07,1.834680e-07,1.834685e-07,1.834689e-07,1.834694e-07,1.834699e-07,1.834704e-07,1.834709e-07,1.834713e-07,1.834718e-07,1.834723e-07,1.834728e-07,1.834733e-07,1.834737e-07,1.834742e-07,1.834747e-07,1.834752e-07,1.834757e-07,1.834761e-07,1.834766e-07,1.834771e-07,1.834776e-07,1.834781e-07,1.834785e-07,1.834790e-07,1.834795e-07,1.834800e-07,1.834805e-07,1.834809e-07,1.834814e-07,1.834819e-07,1.834824e-07,1.834829e-07,1.834833e-07,1.834838e-07,1.834843e-07,1.834848e-07,1.834852e-07,1.834857e-07,1.834862e-07,1.834867e-07,1.834872e-07,1.834876e-07,1.834881e-07,1.834886e-07,1.834891e-07,1.834896e-07,1.834900e-07,1.834905e-07,1.834910e-07,1.834915e-07,1.834920e-07,1.834924e-07,1.834929e-07,1.834934e-07,1.834939e-07,1.834944e-07,1.834948e-07,1.834953e-07,1.834958e-07,1.834963e-07,1.834968e-07,1.834972e-07,1.834977e-07,1.834982e-07,1.834987e-07,1.834991e-07,1.834996e-07,1.835001e-07,1.835006e-07,1.835011e-07,1.835015e-07,1.835020e-07,1.835025e-07,1.835030e-07,1.835035e-07,1.835039e-07,1.835044e-07,1.835049e-07,1.835054e-07,1.835058e-07,1.835063e-07,1.835068e-07,1.835073e-07,1.835078e-07,1.835082e-07,1.835087e-07,1.835092e-07,1.835097e-07,1.835102e-07,1.835106e-07,1.835111e-07,1.835116e-07,1.835121e-07,1.835125e-07,1.835130e-07,1.835135e-07,1.835140e-07,1.835145e-07,1.835149e-07,1.835154e-07,1.835159e-07,1.835164e-07,1.835169e-07,1.835173e-07,1.835178e-07,1.835183e-07,1.835188e-07,1.835192e-07,1.835197e-07,1.835202e-07,1.835207e-07,1.835212e-07,1.835216e-07,1.835221e-07,1.835226e-07,1.835231e-07,1.835235e-07,1.835240e-07,1.835245e-07,1.835250e-07,1.835255e-07,1.835259e-07,1.835264e-07,1.835269e-07,1.835274e-07,1.835278e-07,1.835283e-07,1.835288e-07,1.835293e-07,1.835298e-07,1.835302e-07,1.835307e-07,1.835312e-07,1.835317e-07,1.835321e-07,1.835326e-07,1.835331e-07,1.835336e-07,1.835341e-07,1.835345e-07,1.835350e-07,1.835355e-07,1.835360e-07,1.835364e-07,1.835369e-07,1.835374e-07,1.835379e-07,1.835383e-07,1.835388e-07,1.835393e-07,1.835398e-07,1.835403e-07,1.835407e-07,1.835412e-07,1.835417e-07,1.835422e-07,1.835426e-07,1.835431e-07,1.835436e-07,1.835441e-07,1.835446e-07,1.835450e-07,1.835455e-07,1.835460e-07,1.835465e-07,1.835469e-07,1.835474e-07,1.835479e-07,1.835484e-07,1.835488e-07,1.835493e-07,1.835498e-07,1.835503e-07,1.835507e-07,1.835512e-07,1.835517e-07,1.835522e-07,1.835527e-07,1.835531e-07,1.835536e-07,1.835541e-07,1.835546e-07,1.835550e-07,1.835555e-07,1.835560e-07,1.835565e-07,1.835569e-07,1.835574e-07,1.835579e-07,1.835584e-07,1.835589e-07,1.835593e-07,1.835598e-07,1.835603e-07,1.835608e-07,1.835612e-07,1.835617e-07,1.835622e-07,1.835627e-07,1.835631e-07,1.835636e-07,1.835641e-07,1.835646e-07,1.835650e-07,1.835655e-07,1.835660e-07,1.835665e-07,1.835669e-07,1.835674e-07,1.835679e-07,1.835684e-07,1.835689e-07,1.835693e-07,1.835698e-07,1.835703e-07,1.835708e-07,1.835712e-07,1.835717e-07,1.835722e-07,1.835727e-07,1.835731e-07,1.835736e-07,1.835741e-07,1.835746e-07,1.835750e-07,1.835755e-07,1.835760e-07,1.835765e-07,1.835769e-07,1.835774e-07,1.835779e-07,1.835784e-07,1.835788e-07,1.835793e-07,1.835798e-07,1.835803e-07,1.835807e-07,1.835812e-07,1.835817e-07,1.835822e-07,1.835826e-07,1.835831e-07,1.835836e-07,1.835841e-07,1.835846e-07,1.835850e-07,1.835855e-07,1.835860e-07,1.835865e-07,1.835869e-07,1.835874e-07,1.835879e-07,1.835884e-07,1.835888e-07,1.835893e-07,1.835898e-07,1.835903e-07,1.835907e-07,1.835912e-07,1.835917e-07,1.835922e-07,1.835926e-07,1.835931e-07,1.835936e-07,1.835941e-07,1.835945e-07,1.835950e-07,1.835955e-07,1.835960e-07,1.835964e-07,1.835969e-07,1.835974e-07,1.835979e-07,1.835983e-07,1.835988e-07,1.835993e-07,1.835998e-07,1.836002e-07,1.836007e-07,1.836012e-07,1.836017e-07,1.836021e-07,1.836026e-07,1.836031e-07,1.836036e-07,1.836040e-07,1.836045e-07,1.836050e-07,1.836055e-07,1.836059e-07,1.836064e-07,1.836069e-07,1.836073e-07,1.836078e-07,1.836083e-07,1.836088e-07,1.836092e-07,1.836097e-07,1.836102e-07,1.836107e-07,1.836111e-07,1.836116e-07,1.836121e-07,1.836126e-07,1.836130e-07,1.836135e-07,1.836140e-07,1.836145e-07,1.836149e-07,1.836154e-07,1.836159e-07,1.836164e-07,1.836168e-07,1.836173e-07,1.836178e-07,1.836183e-07,1.836187e-07,1.836192e-07,1.836197e-07,1.836202e-07,1.836206e-07,1.836211e-07,1.836216e-07,1.836220e-07,1.836225e-07,1.836230e-07,1.836235e-07,1.836239e-07,1.836244e-07,1.836249e-07,1.836254e-07,1.836258e-07,1.836263e-07,1.836268e-07,1.836273e-07,1.836277e-07,1.836282e-07,1.836287e-07,1.836292e-07,1.836296e-07,1.836301e-07,1.836306e-07,1.836310e-07,1.836315e-07,1.836320e-07,1.836325e-07,1.836329e-07,1.836334e-07,1.836339e-07,1.836344e-07,1.836348e-07,1.836353e-07,1.836358e-07,1.836363e-07,1.836367e-07,1.836372e-07,1.836377e-07,1.836381e-07,1.836386e-07,1.836391e-07,1.836396e-07,1.836400e-07,1.836405e-07,1.836410e-07,1.836415e-07,1.836419e-07,1.836424e-07,1.836429e-07,1.836434e-07,1.836438e-07,1.836443e-07,1.836448e-07,1.836452e-07,1.836457e-07,1.836462e-07,1.836467e-07,1.836471e-07,1.836476e-07,1.836481e-07,1.836486e-07,1.836490e-07,1.836495e-07,1.836500e-07,1.836504e-07,1.836509e-07,1.836514e-07,1.836519e-07,1.836523e-07,1.836528e-07,1.836533e-07,1.836538e-07,1.836542e-07,1.836547e-07,1.836552e-07,1.836556e-07,1.836561e-07,1.836566e-07,1.836571e-07,1.836575e-07,1.836580e-07,1.836585e-07,1.836590e-07,1.836594e-07,1.836599e-07,1.836604e-07,1.836608e-07,1.836613e-07,1.836618e-07,1.836623e-07,1.836627e-07,1.836632e-07,1.836637e-07,1.836641e-07,1.836646e-07,1.836651e-07,1.836656e-07,1.836660e-07,1.836665e-07,1.836670e-07,1.836674e-07,1.836679e-07,1.836684e-07,1.836689e-07,1.836693e-07,1.836698e-07,1.836703e-07,1.836708e-07,1.836712e-07,1.836717e-07,1.836722e-07,1.836726e-07,1.836731e-07,1.836736e-07,1.836741e-07,1.836745e-07,1.836750e-07,1.836755e-07,1.836759e-07,1.836764e-07,1.836769e-07,1.836774e-07,1.836778e-07,1.836783e-07,1.836788e-07,1.836792e-07,1.836797e-07,1.836802e-07,1.836807e-07,1.836811e-07,1.836816e-07,1.836821e-07,1.836825e-07,1.836830e-07,1.836835e-07,1.836840e-07,1.836844e-07,1.836849e-07,1.836854e-07,1.836858e-07,1.836863e-07,1.836868e-07,1.836873e-07,1.836877e-07,1.836882e-07,1.836887e-07,1.836891e-07,1.836896e-07,1.836901e-07,1.836906e-07,1.836910e-07,1.836915e-07,1.836920e-07,1.836924e-07,1.836929e-07,1.836934e-07,1.836939e-07,1.836943e-07,1.836948e-07,1.836953e-07,1.836957e-07,1.836962e-07,1.836967e-07,1.836971e-07,1.836976e-07,1.836981e-07,1.836986e-07,1.836990e-07,1.836995e-07,1.837000e-07,1.837004e-07,1.837009e-07,1.837014e-07,1.837019e-07,1.837023e-07,1.837028e-07,1.837033e-07,1.837037e-07,1.837042e-07,1.837047e-07,1.837052e-07,1.837056e-07,1.837061e-07,1.837066e-07,1.837070e-07,1.837075e-07,1.837080e-07,1.837084e-07,1.837089e-07,1.837094e-07,1.837099e-07,1.837103e-07,1.837108e-07,1.837113e-07,1.837117e-07,1.837122e-07,1.837127e-07,1.837131e-07,1.837136e-07,1.837141e-07,1.837146e-07,1.837150e-07,1.837155e-07,1.837160e-07,1.837164e-07,1.837169e-07,1.837174e-07,1.837178e-07,1.837183e-07,1.837188e-07,1.837193e-07,1.837197e-07,1.837202e-07,1.837207e-07,1.837211e-07,1.837216e-07,1.837221e-07,1.837225e-07,1.837230e-07,1.837235e-07,1.837240e-07,1.837244e-07,1.837249e-07,1.837254e-07,1.837258e-07,1.837263e-07,1.837268e-07,1.837272e-07,1.837277e-07,1.837282e-07,1.837287e-07,1.837291e-07,1.837296e-07,1.837301e-07,1.837305e-07,1.837310e-07,1.837315e-07,1.837319e-07,1.837324e-07,1.837329e-07,1.837333e-07,1.837338e-07,1.837343e-07,1.837348e-07,1.837352e-07,1.837357e-07,1.837362e-07,1.837366e-07,1.837371e-07,1.837376e-07,1.837380e-07,1.837385e-07,1.837390e-07,1.837394e-07,1.837399e-07,1.837404e-07,1.837409e-07,1.837413e-07,1.837418e-07,1.837423e-07,1.837427e-07,1.837432e-07,1.837437e-07,1.837441e-07,1.837446e-07,1.837451e-07,1.837455e-07,1.837460e-07,1.837465e-07,1.837470e-07,1.837474e-07,1.837479e-07,1.837484e-07,1.837488e-07,1.837493e-07,1.837498e-07,1.837502e-07,1.837507e-07,1.837512e-07,1.837516e-07,1.837521e-07,1.837526e-07,1.837530e-07,1.837535e-07,1.837540e-07,1.837544e-07,1.837549e-07,1.837554e-07,1.837559e-07,1.837563e-07,1.837568e-07,1.837573e-07,1.837577e-07,1.837582e-07,1.837587e-07,1.837591e-07,1.837596e-07,1.837601e-07,1.837605e-07,1.837610e-07,1.837615e-07,1.837619e-07,1.837624e-07,1.837629e-07,1.837633e-07,1.837638e-07,1.837643e-07,1.837648e-07,1.837652e-07,1.837657e-07,1.837662e-07,1.837666e-07,1.837671e-07,1.837676e-07,1.837680e-07,1.837685e-07,1.837690e-07,1.837694e-07,1.837699e-07,1.837704e-07,1.837708e-07,1.837713e-07,1.837718e-07,1.837722e-07,1.837727e-07,1.837732e-07,1.837736e-07,1.837741e-07,1.837746e-07,1.837750e-07,1.837755e-07,1.837760e-07,1.837764e-07,1.837769e-07,1.837774e-07,1.837779e-07,1.837783e-07,1.837788e-07,1.837793e-07,1.837797e-07,1.837802e-07,1.837807e-07,1.837811e-07,1.837816e-07,1.837821e-07,1.837825e-07,1.837830e-07,1.837835e-07,1.837839e-07,1.837844e-07,1.837849e-07,1.837853e-07,1.837858e-07,1.837863e-07,1.837867e-07,1.837872e-07,1.837877e-07,1.837881e-07,1.837886e-07,1.837891e-07,1.837895e-07,1.837900e-07,1.837905e-07,1.837909e-07,1.837914e-07,1.837919e-07,1.837923e-07,1.837928e-07,1.837933e-07,1.837937e-07,1.837942e-07,1.837947e-07,1.837951e-07,1.837956e-07,1.837961e-07,1.837965e-07,1.837970e-07,1.837975e-07,1.837979e-07,1.837984e-07,1.837989e-07,1.837993e-07,1.837998e-07,1.838003e-07,1.838007e-07,1.838012e-07,1.838017e-07,1.838021e-07,1.838026e-07,1.838031e-07,1.838035e-07,1.838040e-07,1.838045e-07,1.838049e-07,1.838054e-07,1.838059e-07,1.838063e-07,1.838068e-07,1.838073e-07,1.838077e-07,1.838082e-07,1.838087e-07,1.838091e-07,1.838096e-07,1.838101e-07,1.838105e-07,1.838110e-07,1.838115e-07,1.838119e-07,1.838124e-07,1.838129e-07,1.838133e-07,1.838138e-07,1.838143e-07,1.838147e-07,1.838152e-07,1.838157e-07,1.838161e-07,1.838166e-07,1.838171e-07,1.838175e-07,1.838180e-07,1.838185e-07,1.838189e-07,1.838194e-07,1.838199e-07,1.838203e-07,1.838208e-07,1.838213e-07,1.838217e-07,1.838222e-07,1.838227e-07,1.838231e-07,1.838236e-07,1.838241e-07,1.838245e-07,1.838250e-07,1.838254e-07,1.838259e-07,1.838264e-07,1.838268e-07,1.838273e-07,1.838278e-07,1.838282e-07,1.838287e-07,1.838292e-07,1.838296e-07,1.838301e-07,1.838306e-07,1.838310e-07,1.838315e-07,1.838320e-07,1.838324e-07,1.838329e-07,1.838334e-07,1.838338e-07,1.838343e-07,1.838348e-07,1.838352e-07,1.838357e-07,1.838362e-07,1.838366e-07,1.838371e-07,1.838375e-07,1.838380e-07,1.838385e-07,1.838389e-07,1.838394e-07,1.838399e-07,1.838403e-07,1.838408e-07,1.838413e-07,1.838417e-07,1.838422e-07,1.838427e-07,1.838431e-07,1.838436e-07,1.838441e-07,1.838445e-07,1.838450e-07,1.838455e-07,1.838459e-07,1.838464e-07,1.838468e-07,1.838473e-07,1.838478e-07,1.838482e-07,1.838487e-07,1.838492e-07,1.838496e-07,1.838501e-07,1.838506e-07,1.838510e-07,1.838515e-07,1.838520e-07,1.838524e-07,1.838529e-07,1.838534e-07,1.838538e-07,1.838543e-07,1.838547e-07,1.838552e-07,1.838557e-07,1.838561e-07,1.838566e-07,1.838571e-07,1.838575e-07,1.838580e-07,1.838585e-07,1.838589e-07,1.838594e-07,1.838599e-07,1.838603e-07,1.838608e-07,1.838613e-07,1.838617e-07,1.838622e-07,1.838626e-07,1.838631e-07,1.838636e-07,1.838640e-07,1.838645e-07,1.838650e-07,1.838654e-07,1.838659e-07,1.838664e-07,1.838668e-07,1.838673e-07,1.838677e-07,1.838682e-07,1.838687e-07,1.838691e-07,1.838696e-07,1.838701e-07,1.838705e-07,1.838710e-07,1.838715e-07,1.838719e-07,1.838724e-07,1.838729e-07,1.838733e-07,1.838738e-07,1.838742e-07,1.838747e-07,1.838752e-07,1.838756e-07,1.838761e-07,1.838766e-07,1.838770e-07,1.838775e-07,1.838780e-07,1.838784e-07,1.838789e-07,1.838793e-07,1.838798e-07,1.838803e-07,1.838807e-07,1.838812e-07,1.838817e-07,1.838821e-07,1.838826e-07,1.838830e-07,1.838835e-07,1.838840e-07,1.838844e-07,1.838849e-07,1.838854e-07,1.838858e-07,1.838863e-07,1.838868e-07,1.838872e-07,1.838877e-07,1.838881e-07,1.838886e-07,1.838891e-07,1.838895e-07,1.838900e-07,1.838905e-07,1.838909e-07,1.838914e-07,1.838919e-07,1.838923e-07,1.838928e-07,1.838932e-07,1.838937e-07,1.838942e-07,1.838946e-07,1.838951e-07,1.838956e-07,1.838960e-07,1.838965e-07,1.838969e-07,1.838974e-07,1.838979e-07,1.838983e-07,1.838988e-07,1.838993e-07,1.838997e-07,1.839002e-07,1.839006e-07,1.839011e-07,1.839016e-07,1.839020e-07,1.839025e-07,1.839030e-07,1.839034e-07,1.839039e-07,1.839043e-07,1.839048e-07,1.839053e-07,1.839057e-07,1.839062e-07,1.839067e-07,1.839071e-07,1.839076e-07,1.839080e-07,1.839085e-07,1.839090e-07,1.839094e-07,1.839099e-07,1.839104e-07,1.839108e-07,1.839113e-07,1.839117e-07,1.839122e-07,1.839127e-07,1.839131e-07,1.839136e-07,1.839141e-07,1.839145e-07,1.839150e-07,1.839154e-07,1.839159e-07,1.839164e-07,1.839168e-07,1.839173e-07,1.839178e-07,1.839182e-07,1.839187e-07,1.839191e-07,1.839196e-07,1.839201e-07,1.839205e-07,1.839210e-07,1.839214e-07,1.839219e-07,1.839224e-07,1.839228e-07,1.839233e-07,1.839238e-07,1.839242e-07,1.839247e-07,1.839251e-07,1.839256e-07,1.839261e-07,1.839265e-07,1.839270e-07,1.839275e-07,1.839279e-07,1.839284e-07,1.839288e-07,1.839293e-07,1.839298e-07,1.839302e-07,1.839307e-07,1.839311e-07,1.839316e-07,1.839321e-07,1.839325e-07,1.839330e-07,1.839334e-07,1.839339e-07,1.839344e-07,1.839348e-07,1.839353e-07,1.839358e-07,1.839362e-07,1.839367e-07,1.839371e-07,1.839376e-07,1.839381e-07,1.839385e-07,1.839390e-07,1.839394e-07,1.839399e-07,1.839404e-07,1.839408e-07,1.839413e-07,1.839418e-07,1.839422e-07,1.839427e-07,1.839431e-07,1.839436e-07,1.839441e-07,1.839445e-07,1.839450e-07,1.839454e-07,1.839459e-07,1.839464e-07,1.839468e-07,1.839473e-07,1.839477e-07,1.839482e-07,1.839487e-07,1.839491e-07,1.839496e-07,1.839500e-07,1.839505e-07,1.839510e-07,1.839514e-07,1.839519e-07,1.839524e-07,1.839528e-07,1.839533e-07,1.839537e-07,1.839542e-07,1.839547e-07,1.839551e-07,1.839556e-07,1.839560e-07,1.839565e-07,1.839570e-07,1.839574e-07,1.839579e-07,1.839583e-07,1.839588e-07,1.839593e-07,1.839597e-07,1.839602e-07,1.839606e-07,1.839611e-07,1.839616e-07,1.839620e-07,1.839625e-07,1.839629e-07,1.839634e-07,1.839639e-07,1.839643e-07,1.839648e-07,1.839652e-07,1.839657e-07,1.839662e-07,1.839666e-07,1.839671e-07,1.839675e-07,1.839680e-07,1.839685e-07,1.839689e-07,1.839694e-07,1.839698e-07,1.839703e-07,1.839708e-07,1.839712e-07,1.839717e-07,1.839721e-07,1.839726e-07,1.839731e-07,1.839735e-07,1.839740e-07,1.839744e-07,1.839749e-07,1.839754e-07,1.839758e-07,1.839763e-07,1.839767e-07,1.839772e-07,1.839777e-07,1.839781e-07,1.839786e-07,1.839790e-07,1.839795e-07,1.839800e-07,1.839804e-07,1.839809e-07,1.839813e-07,1.839818e-07,1.839823e-07,1.839827e-07,1.839832e-07,1.839836e-07,1.839841e-07,1.839846e-07,1.839850e-07,1.839855e-07,1.839859e-07,1.839864e-07,1.839868e-07,1.839873e-07,1.839878e-07,1.839882e-07,1.839887e-07,1.839891e-07,1.839896e-07,1.839901e-07,1.839905e-07,1.839910e-07,1.839914e-07,1.839919e-07,1.839924e-07,1.839928e-07,1.839933e-07,1.839937e-07,1.839942e-07,1.839947e-07,1.839951e-07,1.839956e-07,1.839960e-07,1.839965e-07,1.839969e-07,1.839974e-07,1.839979e-07,1.839983e-07,1.839988e-07,1.839992e-07,1.839997e-07,1.840002e-07,1.840006e-07,1.840011e-07,1.840015e-07,1.840020e-07,1.840025e-07,1.840029e-07,1.840034e-07,1.840038e-07,1.840043e-07,1.840047e-07,1.840052e-07,1.840057e-07,1.840061e-07,1.840066e-07,1.840070e-07,1.840075e-07,1.840080e-07,1.840084e-07,1.840089e-07,1.840093e-07,1.840098e-07,1.840102e-07,1.840107e-07,1.840112e-07,1.840116e-07,1.840121e-07,1.840125e-07,1.840130e-07,1.840135e-07,1.840139e-07,1.840144e-07,1.840148e-07,1.840153e-07,1.840157e-07,1.840162e-07,1.840167e-07,1.840171e-07,1.840176e-07,1.840180e-07,1.840185e-07,1.840190e-07,1.840194e-07,1.840199e-07,1.840203e-07,1.840208e-07,1.840212e-07,1.840217e-07,1.840222e-07,1.840226e-07,1.840231e-07,1.840235e-07,1.840240e-07,1.840244e-07,1.840249e-07,1.840254e-07,1.840258e-07,1.840263e-07,1.840267e-07,1.840272e-07,1.840277e-07,1.840281e-07,1.840286e-07,1.840290e-07,1.840295e-07,1.840299e-07,1.840304e-07,1.840309e-07,1.840313e-07,1.840318e-07,1.840322e-07,1.840327e-07,1.840331e-07,1.840336e-07,1.840341e-07,1.840345e-07,1.840350e-07,1.840354e-07,1.840359e-07,1.840363e-07,1.840368e-07,1.840373e-07,1.840377e-07,1.840382e-07,1.840386e-07,1.840391e-07,1.840395e-07,1.840400e-07,1.840405e-07,1.840409e-07,1.840414e-07,1.840418e-07,1.840423e-07,1.840427e-07,1.840432e-07,1.840437e-07,1.840441e-07,1.840446e-07,1.840450e-07,1.840455e-07,1.840459e-07,1.840464e-07,1.840469e-07,1.840473e-07,1.840478e-07,1.840482e-07,1.840487e-07,1.840491e-07,1.840496e-07,1.840501e-07,1.840505e-07,1.840510e-07,1.840514e-07,1.840519e-07,1.840523e-07,1.840528e-07,1.840533e-07,1.840537e-07,1.840542e-07,1.840546e-07,1.840551e-07,1.840555e-07,1.840560e-07,1.840565e-07,1.840569e-07,1.840574e-07,1.840578e-07,1.840583e-07,1.840587e-07,1.840592e-07,1.840596e-07,1.840601e-07,1.840606e-07,1.840610e-07,1.840615e-07,1.840619e-07,1.840624e-07,1.840628e-07,1.840633e-07,1.840638e-07,1.840642e-07,1.840647e-07,1.840651e-07,1.840656e-07,1.840660e-07,1.840665e-07,1.840669e-07,1.840674e-07,1.840679e-07,1.840683e-07,1.840688e-07,1.840692e-07,1.840697e-07,1.840701e-07,1.840706e-07,1.840711e-07,1.840715e-07,1.840720e-07,1.840724e-07,1.840729e-07,1.840733e-07,1.840738e-07,1.840742e-07,1.840747e-07,1.840752e-07,1.840756e-07,1.840761e-07,1.840765e-07,1.840770e-07,1.840774e-07,1.840779e-07,1.840783e-07,1.840788e-07,1.840793e-07,1.840797e-07,1.840802e-07,1.840806e-07,1.840811e-07,1.840815e-07,1.840820e-07,1.840824e-07,1.840829e-07,1.840834e-07,1.840838e-07,1.840843e-07,1.840847e-07,1.840852e-07,1.840856e-07,1.840861e-07,1.840865e-07,1.840870e-07,1.840875e-07,1.840879e-07,1.840884e-07,1.840888e-07,1.840893e-07,1.840897e-07,1.840902e-07,1.840906e-07,1.840911e-07,1.840916e-07,1.840920e-07,1.840925e-07,1.840929e-07,1.840934e-07,1.840938e-07,1.840943e-07,1.840947e-07,1.840952e-07,1.840956e-07,1.840961e-07,1.840966e-07,1.840970e-07,1.840975e-07,1.840979e-07,1.840984e-07,1.840988e-07,1.840993e-07,1.840997e-07,1.841002e-07,1.841007e-07,1.841011e-07,1.841016e-07,1.841020e-07,1.841025e-07,1.841029e-07,1.841034e-07,1.841038e-07,1.841043e-07,1.841047e-07,1.841052e-07,1.841057e-07,1.841061e-07,1.841066e-07,1.841070e-07,1.841075e-07,1.841079e-07,1.841084e-07,1.841088e-07,1.841093e-07,1.841097e-07,1.841102e-07,1.841107e-07,1.841111e-07,1.841116e-07,1.841120e-07,1.841125e-07,1.841129e-07,1.841134e-07,1.841138e-07,1.841143e-07,1.841147e-07,1.841152e-07,1.841157e-07,1.841161e-07,1.841166e-07,1.841170e-07,1.841175e-07,1.841179e-07,1.841184e-07,1.841188e-07,1.841193e-07,1.841197e-07,1.841202e-07,1.841206e-07,1.841211e-07,1.841216e-07,1.841220e-07,1.841225e-07,1.841229e-07,1.841234e-07,1.841238e-07,1.841243e-07,1.841247e-07,1.841252e-07,1.841256e-07,1.841261e-07,1.841265e-07,1.841270e-07,1.841275e-07,1.841279e-07,1.841284e-07,1.841288e-07,1.841293e-07,1.841297e-07,1.841302e-07,1.841306e-07,1.841311e-07,1.841315e-07,1.841320e-07,1.841324e-07,1.841329e-07,1.841334e-07,1.841338e-07,1.841343e-07,1.841347e-07,1.841352e-07,1.841356e-07,1.841361e-07,1.841365e-07,1.841370e-07,1.841374e-07,1.841379e-07,1.841383e-07,1.841388e-07,1.841392e-07,1.841397e-07,1.841402e-07,1.841406e-07,1.841411e-07,1.841415e-07,1.841420e-07,1.841424e-07,1.841429e-07,1.841433e-07,1.841438e-07,1.841442e-07,1.841447e-07,1.841451e-07,1.841456e-07,1.841460e-07,1.841465e-07,1.841470e-07,1.841474e-07,1.841479e-07,1.841483e-07,1.841488e-07,1.841492e-07,1.841497e-07,1.841501e-07,1.841506e-07,1.841510e-07,1.841515e-07,1.841519e-07,1.841524e-07,1.841528e-07,1.841533e-07,1.841537e-07,1.841542e-07,1.841547e-07,1.841551e-07,1.841556e-07,1.841560e-07,1.841565e-07,1.841569e-07,1.841574e-07,1.841578e-07,1.841583e-07,1.841587e-07,1.841592e-07,1.841596e-07,1.841601e-07,1.841605e-07,1.841610e-07,1.841614e-07,1.841619e-07,1.841623e-07,1.841628e-07,1.841633e-07,1.841637e-07,1.841642e-07,1.841646e-07,1.841651e-07,1.841655e-07,1.841660e-07,1.841664e-07,1.841669e-07,1.841673e-07,1.841678e-07,1.841682e-07,1.841687e-07,1.841691e-07,1.841696e-07,1.841700e-07,1.841705e-07,1.841709e-07,1.841714e-07,1.841718e-07,1.841723e-07,1.841727e-07,1.841732e-07,1.841737e-07,1.841741e-07,1.841746e-07,1.841750e-07,1.841755e-07,1.841759e-07,1.841764e-07,1.841768e-07,1.841773e-07,1.841777e-07,1.841782e-07,1.841786e-07,1.841791e-07,1.841795e-07,1.841800e-07,1.841804e-07,1.841809e-07,1.841813e-07,1.841818e-07,1.841822e-07,1.841827e-07,1.841831e-07,1.841836e-07,1.841840e-07,1.841845e-07,1.841849e-07,1.841854e-07,1.841858e-07,1.841863e-07,1.841868e-07,1.841872e-07,1.841877e-07,1.841881e-07,1.841886e-07,1.841890e-07,1.841895e-07,1.841899e-07,1.841904e-07,1.841908e-07,1.841913e-07,1.841917e-07,1.841922e-07,1.841926e-07,1.841931e-07,1.841935e-07,1.841940e-07,1.841944e-07,1.841949e-07,1.841953e-07,1.841958e-07,1.841962e-07,1.841967e-07,1.841971e-07,1.841976e-07,1.841980e-07,1.841985e-07,1.841989e-07,1.841994e-07,1.841998e-07,1.842003e-07,1.842007e-07,1.842012e-07,1.842016e-07,1.842021e-07,1.842025e-07,1.842030e-07,1.842034e-07,1.842039e-07,1.842043e-07,1.842048e-07,1.842052e-07,1.842057e-07,1.842061e-07,1.842066e-07,1.842071e-07,1.842075e-07,1.842080e-07,1.842084e-07,1.842089e-07,1.842093e-07,1.842098e-07,1.842102e-07,1.842107e-07,1.842111e-07,1.842116e-07,1.842120e-07,1.842125e-07,1.842129e-07,1.842134e-07,1.842138e-07,1.842143e-07,1.842147e-07,1.842152e-07,1.842156e-07,1.842161e-07,1.842165e-07,1.842170e-07,1.842174e-07,1.842179e-07,1.842183e-07,1.842188e-07,1.842192e-07,1.842197e-07,1.842201e-07,1.842206e-07,1.842210e-07,1.842215e-07,1.842219e-07,1.842224e-07,1.842228e-07,1.842233e-07,1.842237e-07,1.842242e-07,1.842246e-07,1.842251e-07,1.842255e-07,1.842260e-07,1.842264e-07,1.842269e-07,1.842273e-07,1.842278e-07,1.842282e-07,1.842287e-07,1.842291e-07,1.842296e-07,1.842300e-07,1.842305e-07,1.842309e-07,1.842314e-07,1.842318e-07,1.842323e-07,1.842327e-07,1.842332e-07,1.842336e-07,1.842341e-07,1.842345e-07,1.842350e-07,1.842354e-07,1.842359e-07,1.842363e-07,1.842368e-07,1.842372e-07,1.842377e-07,1.842381e-07,1.842386e-07,1.842390e-07,1.842395e-07,1.842399e-07,1.842404e-07,1.842408e-07,1.842413e-07,1.842417e-07,1.842422e-07,1.842426e-07,1.842431e-07,1.842435e-07,1.842439e-07,1.842444e-07,1.842448e-07,1.842453e-07,1.842457e-07,1.842462e-07,1.842466e-07,1.842471e-07,1.842475e-07,1.842480e-07,1.842484e-07,1.842489e-07,1.842493e-07,1.842498e-07,1.842502e-07,1.842507e-07,1.842511e-07,1.842516e-07,1.842520e-07,1.842525e-07,1.842529e-07,1.842534e-07,1.842538e-07,1.842543e-07,1.842547e-07,1.842552e-07,1.842556e-07,1.842561e-07,1.842565e-07,1.842570e-07,1.842574e-07,1.842579e-07,1.842583e-07,1.842588e-07,1.842592e-07,1.842597e-07,1.842601e-07,1.842606e-07,1.842610e-07,1.842615e-07,1.842619e-07,1.842624e-07,1.842628e-07,1.842633e-07,1.842637e-07,1.842641e-07,1.842646e-07,1.842650e-07,1.842655e-07,1.842659e-07,1.842664e-07,1.842668e-07,1.842673e-07,1.842677e-07,1.842682e-07,1.842686e-07,1.842691e-07,1.842695e-07,1.842700e-07,1.842704e-07,1.842709e-07,1.842713e-07,1.842718e-07,1.842722e-07,1.842727e-07,1.842731e-07,1.842736e-07,1.842740e-07,1.842745e-07,1.842749e-07,1.842754e-07,1.842758e-07,1.842763e-07,1.842767e-07,1.842771e-07,1.842776e-07,1.842780e-07,1.842785e-07,1.842789e-07,1.842794e-07,1.842798e-07,1.842803e-07,1.842807e-07,1.842812e-07,1.842816e-07,1.842821e-07,1.842825e-07,1.842830e-07,1.842834e-07,1.842839e-07,1.842843e-07,1.842848e-07,1.842852e-07,1.842857e-07,1.842861e-07,1.842866e-07,1.842870e-07,1.842874e-07,1.842879e-07,1.842883e-07,1.842888e-07,1.842892e-07,1.842897e-07,1.842901e-07,1.842906e-07,1.842910e-07,1.842915e-07,1.842919e-07,1.842924e-07,1.842928e-07,1.842933e-07,1.842937e-07,1.842942e-07,1.842946e-07,1.842951e-07,1.842955e-07,1.842959e-07,1.842964e-07,1.842968e-07,1.842973e-07,1.842977e-07,1.842982e-07,1.842986e-07,1.842991e-07,1.842995e-07,1.843000e-07,1.843004e-07,1.843009e-07,1.843013e-07,1.843018e-07,1.843022e-07,1.843027e-07,1.843031e-07,1.843036e-07,1.843040e-07,1.843044e-07,1.843049e-07,1.843053e-07,1.843058e-07,1.843062e-07,1.843067e-07,1.843071e-07,1.843076e-07,1.843080e-07,1.843085e-07,1.843089e-07,1.843094e-07,1.843098e-07,1.843103e-07,1.843107e-07,1.843111e-07,1.843116e-07,1.843120e-07,1.843125e-07,1.843129e-07,1.843134e-07,1.843138e-07,1.843143e-07,1.843147e-07,1.843152e-07,1.843156e-07,1.843161e-07,1.843165e-07,1.843170e-07,1.843174e-07,1.843178e-07,1.843183e-07,1.843187e-07,1.843192e-07,1.843196e-07,1.843201e-07,1.843205e-07,1.843210e-07,1.843214e-07,1.843219e-07,1.843223e-07,1.843228e-07,1.843232e-07,1.843236e-07,1.843241e-07,1.843245e-07,1.843250e-07,1.843254e-07,1.843259e-07,1.843263e-07,1.843268e-07,1.843272e-07,1.843277e-07,1.843281e-07,1.843286e-07,1.843290e-07,1.843294e-07,1.843299e-07,1.843303e-07,1.843308e-07,1.843312e-07,1.843317e-07,1.843321e-07,1.843326e-07,1.843330e-07,1.843335e-07,1.843339e-07,1.843344e-07,1.843348e-07,1.843352e-07,1.843357e-07,1.843361e-07,1.843366e-07,1.843370e-07,1.843375e-07,1.843379e-07,1.843384e-07,1.843388e-07,1.843393e-07,1.843397e-07,1.843401e-07,1.843406e-07,1.843410e-07,1.843415e-07,1.843419e-07,1.843424e-07,1.843428e-07,1.843433e-07,1.843437e-07,1.843442e-07,1.843446e-07,1.843450e-07,1.843455e-07,1.843459e-07,1.843464e-07,1.843468e-07,1.843473e-07,1.843477e-07,1.843482e-07,1.843486e-07,1.843491e-07,1.843495e-07,1.843499e-07,1.843504e-07,1.843508e-07,1.843513e-07,1.843517e-07,1.843522e-07,1.843526e-07,1.843531e-07,1.843535e-07,1.843540e-07,1.843544e-07,1.843548e-07,1.843553e-07,1.843557e-07,1.843562e-07,1.843566e-07,1.843571e-07,1.843575e-07,1.843580e-07,1.843584e-07,1.843588e-07,1.843593e-07,1.843597e-07,1.843602e-07,1.843606e-07,1.843611e-07,1.843615e-07,1.843620e-07,1.843624e-07,1.843628e-07,1.843633e-07,1.843637e-07,1.843642e-07,1.843646e-07,1.843651e-07,1.843655e-07,1.843660e-07,1.843664e-07,1.843669e-07,1.843673e-07,1.843677e-07,1.843682e-07,1.843686e-07,1.843691e-07,1.843695e-07,1.843700e-07,1.843704e-07,1.843709e-07,1.843713e-07,1.843717e-07,1.843722e-07,1.843726e-07,1.843731e-07,1.843735e-07,1.843740e-07,1.843744e-07,1.843749e-07,1.843753e-07,1.843757e-07,1.843762e-07,1.843766e-07,1.843771e-07,1.843775e-07,1.843780e-07,1.843784e-07,1.843788e-07,1.843793e-07,1.843797e-07,1.843802e-07,1.843806e-07,1.843811e-07,1.843815e-07,1.843820e-07,1.843824e-07,1.843828e-07,1.843833e-07,1.843837e-07,1.843842e-07,1.843846e-07,1.843851e-07,1.843855e-07,1.843860e-07,1.843864e-07,1.843868e-07,1.843873e-07,1.843877e-07,1.843882e-07,1.843886e-07,1.843891e-07,1.843895e-07,1.843899e-07,1.843904e-07,1.843908e-07,1.843913e-07,1.843917e-07,1.843922e-07,1.843926e-07,1.843931e-07,1.843935e-07,1.843939e-07,1.843944e-07,1.843948e-07,1.843953e-07,1.843957e-07,1.843962e-07,1.843966e-07,1.843970e-07,1.843975e-07,1.843979e-07,1.843984e-07,1.843988e-07,1.843993e-07,1.843997e-07,1.844001e-07,1.844006e-07,1.844010e-07,1.844015e-07,1.844019e-07,1.844024e-07,1.844028e-07,1.844032e-07,1.844037e-07,1.844041e-07,1.844046e-07,1.844050e-07,1.844055e-07,1.844059e-07,1.844064e-07,1.844068e-07,1.844072e-07,1.844077e-07,1.844081e-07,1.844086e-07,1.844090e-07,1.844095e-07,1.844099e-07,1.844103e-07,1.844108e-07,1.844112e-07,1.844117e-07,1.844121e-07,1.844126e-07,1.844130e-07,1.844134e-07,1.844139e-07,1.844143e-07,1.844148e-07,1.844152e-07,1.844157e-07,1.844161e-07,1.844165e-07,1.844170e-07,1.844174e-07,1.844179e-07,1.844183e-07,1.844188e-07,1.844192e-07,1.844196e-07,1.844201e-07,1.844205e-07,1.844210e-07,1.844214e-07,1.844218e-07,1.844223e-07,1.844227e-07,1.844232e-07,1.844236e-07,1.844241e-07,1.844245e-07,1.844249e-07,1.844254e-07,1.844258e-07,1.844263e-07,1.844267e-07,1.844272e-07,1.844276e-07,1.844280e-07,1.844285e-07,1.844289e-07,1.844294e-07,1.844298e-07,1.844303e-07,1.844307e-07,1.844311e-07,1.844316e-07,1.844320e-07,1.844325e-07,1.844329e-07,1.844333e-07,1.844338e-07,1.844342e-07,1.844347e-07,1.844351e-07,1.844356e-07,1.844360e-07,1.844364e-07,1.844369e-07,1.844373e-07,1.844378e-07,1.844382e-07,1.844387e-07,1.844391e-07,1.844395e-07,1.844400e-07,1.844404e-07,1.844409e-07,1.844413e-07,1.844417e-07,1.844422e-07,1.844426e-07,1.844431e-07,1.844435e-07,1.844440e-07,1.844444e-07,1.844448e-07,1.844453e-07,1.844457e-07,1.844462e-07,1.844466e-07,1.844470e-07,1.844475e-07,1.844479e-07,1.844484e-07,1.844488e-07,1.844492e-07,1.844497e-07,1.844501e-07,1.844506e-07,1.844510e-07,1.844515e-07,1.844519e-07,1.844523e-07,1.844528e-07,1.844532e-07,1.844537e-07,1.844541e-07,1.844545e-07,1.844550e-07,1.844554e-07,1.844559e-07,1.844563e-07,1.844568e-07,1.844572e-07,1.844576e-07,1.844581e-07,1.844585e-07,1.844590e-07,1.844594e-07,1.844598e-07,1.844603e-07,1.844607e-07,1.844612e-07,1.844616e-07,1.844620e-07,1.844625e-07,1.844629e-07,1.844634e-07,1.844638e-07,1.844642e-07,1.844647e-07,1.844651e-07,1.844656e-07,1.844660e-07,1.844665e-07,1.844669e-07,1.844673e-07,1.844678e-07,1.844682e-07,1.844687e-07,1.844691e-07,1.844695e-07,1.844700e-07,1.844704e-07,1.844709e-07,1.844713e-07,1.844717e-07,1.844722e-07,1.844726e-07,1.844731e-07,1.844735e-07,1.844739e-07,1.844744e-07,1.844748e-07,1.844753e-07,1.844757e-07,1.844761e-07,1.844766e-07,1.844770e-07,1.844775e-07,1.844779e-07,1.844783e-07,1.844788e-07,1.844792e-07,1.844797e-07,1.844801e-07,1.844806e-07,1.844810e-07,1.844814e-07,1.844819e-07,1.844823e-07,1.844828e-07,1.844832e-07,1.844836e-07,1.844841e-07,1.844845e-07,1.844850e-07,1.844854e-07,1.844858e-07,1.844863e-07,1.844867e-07,1.844872e-07,1.844876e-07,1.844880e-07,1.844885e-07,1.844889e-07,1.844894e-07,1.844898e-07,1.844902e-07,1.844907e-07,1.844911e-07,1.844916e-07,1.844920e-07,1.844924e-07,1.844929e-07,1.844933e-07,1.844938e-07,1.844942e-07,1.844946e-07,1.844951e-07,1.844955e-07,1.844959e-07,1.844964e-07,1.844968e-07,1.844973e-07,1.844977e-07,1.844981e-07,1.844986e-07,1.844990e-07,1.844995e-07,1.844999e-07,1.845003e-07,1.845008e-07,1.845012e-07,1.845017e-07,1.845021e-07,1.845025e-07,1.845030e-07,1.845034e-07,1.845039e-07,1.845043e-07,1.845047e-07,1.845052e-07,1.845056e-07,1.845061e-07,1.845065e-07,1.845069e-07,1.845074e-07,1.845078e-07,1.845083e-07,1.845087e-07,1.845091e-07,1.845096e-07,1.845100e-07,1.845104e-07,1.845109e-07,1.845113e-07,1.845118e-07,1.845122e-07,1.845126e-07,1.845131e-07,1.845135e-07,1.845140e-07,1.845144e-07,1.845148e-07,1.845153e-07,1.845157e-07,1.845162e-07,1.845166e-07,1.845170e-07,1.845175e-07,1.845179e-07,1.845184e-07,1.845188e-07,1.845192e-07,1.845197e-07,1.845201e-07,1.845205e-07,1.845210e-07,1.845214e-07,1.845219e-07,1.845223e-07,1.845227e-07,1.845232e-07,1.845236e-07,1.845241e-07,1.845245e-07,1.845249e-07,1.845254e-07,1.845258e-07,1.845262e-07,1.845267e-07,1.845271e-07,1.845276e-07,1.845280e-07,1.845284e-07,1.845289e-07,1.845293e-07,1.845298e-07,1.845302e-07,1.845306e-07,1.845311e-07,1.845315e-07,1.845319e-07,1.845324e-07,1.845328e-07,1.845333e-07,1.845337e-07,1.845341e-07,1.845346e-07,1.845350e-07,1.845355e-07,1.845359e-07,1.845363e-07,1.845368e-07,1.845372e-07,1.845376e-07,1.845381e-07,1.845385e-07,1.845390e-07,1.845394e-07,1.845398e-07,1.845403e-07,1.845407e-07,1.845411e-07,1.845416e-07,1.845420e-07,1.845425e-07,1.845429e-07,1.845433e-07,1.845438e-07,1.845442e-07,1.845447e-07,1.845451e-07,1.845455e-07,1.845460e-07,1.845464e-07,1.845468e-07,1.845473e-07,1.845477e-07,1.845482e-07,1.845486e-07,1.845490e-07,1.845495e-07,1.845499e-07,1.845503e-07,1.845508e-07,1.845512e-07,1.845517e-07,1.845521e-07,1.845525e-07,1.845530e-07,1.845534e-07,1.845538e-07,1.845543e-07,1.845547e-07,1.845552e-07,1.845556e-07,1.845560e-07,1.845565e-07,1.845569e-07,1.845573e-07,1.845578e-07,1.845582e-07,1.845587e-07,1.845591e-07,1.845595e-07,1.845600e-07,1.845604e-07,1.845608e-07,1.845613e-07,1.845617e-07,1.845622e-07,1.845626e-07,1.845630e-07,1.845635e-07,1.845639e-07,1.845643e-07,1.845648e-07,1.845652e-07,1.845657e-07,1.845661e-07,1.845665e-07,1.845670e-07,1.845674e-07,1.845678e-07,1.845683e-07,1.845687e-07,1.845691e-07,1.845696e-07,1.845700e-07,1.845705e-07,1.845709e-07,1.845713e-07,1.845718e-07,1.845722e-07,1.845726e-07,1.845731e-07,1.845735e-07,1.845740e-07,1.845744e-07,1.845748e-07,1.845753e-07,1.845757e-07,1.845761e-07,1.845766e-07,1.845770e-07,1.845774e-07,1.845779e-07,1.845783e-07,1.845788e-07,1.845792e-07,1.845796e-07,1.845801e-07,1.845805e-07,1.845809e-07,1.845814e-07,1.845818e-07,1.845822e-07,1.845827e-07,1.845831e-07,1.845836e-07,1.845840e-07,1.845844e-07,1.845849e-07,1.845853e-07,1.845857e-07,1.845862e-07,1.845866e-07,1.845870e-07,1.845875e-07,1.845879e-07,1.845884e-07,1.845888e-07,1.845892e-07,1.845897e-07,1.845901e-07,1.845905e-07,1.845910e-07,1.845914e-07,1.845918e-07,1.845923e-07,1.845927e-07,1.845932e-07,1.845936e-07,1.845940e-07,1.845945e-07,1.845949e-07,1.845953e-07,1.845958e-07,1.845962e-07,1.845966e-07,1.845971e-07,1.845975e-07,1.845979e-07,1.845984e-07,1.845988e-07,1.845993e-07,1.845997e-07,1.846001e-07,1.846006e-07,1.846010e-07,1.846014e-07,1.846019e-07,1.846023e-07,1.846027e-07,1.846032e-07,1.846036e-07,1.846040e-07,1.846045e-07,1.846049e-07,1.846054e-07,1.846058e-07,1.846062e-07,1.846067e-07,1.846071e-07,1.846075e-07,1.846080e-07,1.846084e-07,1.846088e-07,1.846093e-07,1.846097e-07,1.846101e-07,1.846106e-07,1.846110e-07,1.846115e-07,1.846119e-07,1.846123e-07,1.846128e-07,1.846132e-07,1.846136e-07,1.846141e-07,1.846145e-07,1.846149e-07,1.846154e-07,1.846158e-07,1.846162e-07,1.846167e-07,1.846171e-07,1.846175e-07,1.846180e-07,1.846184e-07,1.846189e-07,1.846193e-07,1.846197e-07,1.846202e-07,1.846206e-07,1.846210e-07,1.846215e-07,1.846219e-07,1.846223e-07,1.846228e-07,1.846232e-07,1.846236e-07,1.846241e-07,1.846245e-07,1.846249e-07,1.846254e-07,1.846258e-07,1.846262e-07,1.846267e-07,1.846271e-07,1.846275e-07,1.846280e-07,1.846284e-07,1.846289e-07,1.846293e-07,1.846297e-07,1.846302e-07,1.846306e-07,1.846310e-07,1.846315e-07,1.846319e-07,1.846323e-07,1.846328e-07,1.846332e-07,1.846336e-07,1.846341e-07,1.846345e-07,1.846349e-07,1.846354e-07,1.846358e-07,1.846362e-07,1.846367e-07,1.846371e-07,1.846375e-07,1.846380e-07,1.846384e-07,1.846388e-07,1.846393e-07,1.846397e-07,1.846401e-07,1.846406e-07,1.846410e-07,1.846415e-07,1.846419e-07,1.846423e-07,1.846428e-07,1.846432e-07,1.846436e-07,1.846441e-07,1.846445e-07,1.846449e-07,1.846454e-07,1.846458e-07,1.846462e-07,1.846467e-07,1.846471e-07,1.846475e-07,1.846480e-07,1.846484e-07,1.846488e-07,1.846493e-07,1.846497e-07,1.846501e-07,1.846506e-07,1.846510e-07,1.846514e-07,1.846519e-07,1.846523e-07,1.846527e-07,1.846532e-07,1.846536e-07,1.846540e-07,1.846545e-07,1.846549e-07,1.846553e-07,1.846558e-07,1.846562e-07,1.846566e-07,1.846571e-07,1.846575e-07,1.846579e-07,1.846584e-07,1.846588e-07,1.846592e-07,1.846597e-07,1.846601e-07,1.846605e-07,1.846610e-07,1.846614e-07,1.846618e-07,1.846623e-07,1.846627e-07,1.846631e-07,1.846636e-07,1.846640e-07,1.846644e-07,1.846649e-07,1.846653e-07,1.846657e-07,1.846662e-07,1.846666e-07,1.846670e-07,1.846675e-07,1.846679e-07,1.846683e-07,1.846688e-07,1.846692e-07,1.846696e-07,1.846701e-07,1.846705e-07,1.846709e-07,1.846714e-07,1.846718e-07,1.846722e-07,1.846727e-07,1.846731e-07,1.846735e-07,1.846740e-07,1.846744e-07,1.846748e-07,1.846753e-07,1.846757e-07,1.846761e-07,1.846766e-07,1.846770e-07,1.846774e-07,1.846779e-07,1.846783e-07,1.846787e-07,1.846792e-07,1.846796e-07,1.846800e-07,1.846805e-07,1.846809e-07,1.846813e-07,1.846818e-07,1.846822e-07,1.846826e-07,1.846831e-07,1.846835e-07,1.846839e-07,1.846844e-07,1.846848e-07,1.846852e-07,1.846857e-07,1.846861e-07,1.846865e-07,1.846870e-07,1.846874e-07,1.846878e-07,1.846883e-07,1.846887e-07,1.846891e-07,1.846896e-07,1.846900e-07,1.846904e-07,1.846909e-07,1.846913e-07,1.846917e-07,1.846921e-07,1.846926e-07,1.846930e-07,1.846934e-07,1.846939e-07,1.846943e-07,1.846947e-07,1.846952e-07,1.846956e-07,1.846960e-07,1.846965e-07,1.846969e-07,1.846973e-07,1.846978e-07,1.846982e-07,1.846986e-07,1.846991e-07,1.846995e-07,1.846999e-07,1.847004e-07,1.847008e-07,1.847012e-07,1.847017e-07,1.847021e-07,1.847025e-07,1.847030e-07,1.847034e-07,1.847038e-07,1.847042e-07,1.847047e-07,1.847051e-07,1.847055e-07,1.847060e-07,1.847064e-07,1.847068e-07,1.847073e-07,1.847077e-07,1.847081e-07,1.847086e-07,1.847090e-07,1.847094e-07,1.847099e-07,1.847103e-07,1.847107e-07,1.847112e-07,1.847116e-07,1.847120e-07,1.847125e-07,1.847129e-07,1.847133e-07,1.847137e-07,1.847142e-07,1.847146e-07,1.847150e-07,1.847155e-07,1.847159e-07,1.847163e-07,1.847168e-07,1.847172e-07,1.847176e-07,1.847181e-07,1.847185e-07,1.847189e-07,1.847194e-07,1.847198e-07,1.847202e-07,1.847206e-07,1.847211e-07,1.847215e-07,1.847219e-07,1.847224e-07,1.847228e-07,1.847232e-07,1.847237e-07,1.847241e-07,1.847245e-07,1.847250e-07,1.847254e-07,1.847258e-07,1.847263e-07,1.847267e-07,1.847271e-07,1.847275e-07,1.847280e-07,1.847284e-07,1.847288e-07,1.847293e-07,1.847297e-07,1.847301e-07,1.847306e-07,1.847310e-07,1.847314e-07,1.847319e-07,1.847323e-07,1.847327e-07,1.847331e-07,1.847336e-07,1.847340e-07,1.847344e-07,1.847349e-07,1.847353e-07,1.847357e-07,1.847362e-07,1.847366e-07,1.847370e-07,1.847375e-07,1.847379e-07,1.847383e-07,1.847387e-07,1.847392e-07,1.847396e-07,1.847400e-07,1.847405e-07,1.847409e-07,1.847413e-07,1.847418e-07,1.847422e-07,1.847426e-07,1.847431e-07,1.847435e-07,1.847439e-07,1.847443e-07,1.847448e-07,1.847452e-07,1.847456e-07,1.847461e-07,1.847465e-07,1.847469e-07,1.847474e-07,1.847478e-07,1.847482e-07,1.847486e-07,1.847491e-07,1.847495e-07,1.847499e-07,1.847504e-07,1.847508e-07,1.847512e-07,1.847517e-07,1.847521e-07,1.847525e-07,1.847530e-07,1.847534e-07,1.847538e-07,1.847542e-07,1.847547e-07,1.847551e-07,1.847555e-07,1.847560e-07,1.847564e-07,1.847568e-07,1.847573e-07,1.847577e-07,1.847581e-07,1.847585e-07,1.847590e-07,1.847594e-07,1.847598e-07,1.847603e-07,1.847607e-07,1.847611e-07,1.847615e-07,1.847620e-07,1.847624e-07,1.847628e-07,1.847633e-07,1.847637e-07,1.847641e-07,1.847646e-07,1.847650e-07,1.847654e-07,1.847658e-07,1.847663e-07,1.847667e-07,1.847671e-07,1.847676e-07,1.847680e-07,1.847684e-07,1.847689e-07,1.847693e-07,1.847697e-07,1.847701e-07,1.847706e-07,1.847710e-07,1.847714e-07,1.847719e-07,1.847723e-07,1.847727e-07,1.847731e-07,1.847736e-07,1.847740e-07,1.847744e-07,1.847749e-07,1.847753e-07,1.847757e-07,1.847762e-07,1.847766e-07,1.847770e-07,1.847774e-07,1.847779e-07,1.847783e-07,1.847787e-07,1.847792e-07,1.847796e-07,1.847800e-07,1.847804e-07,1.847809e-07,1.847813e-07,1.847817e-07,1.847822e-07,1.847826e-07,1.847830e-07,1.847834e-07,1.847839e-07,1.847843e-07,1.847847e-07,1.847852e-07,1.847856e-07,1.847860e-07,1.847865e-07,1.847869e-07,1.847873e-07,1.847877e-07,1.847882e-07,1.847886e-07,1.847890e-07,1.847895e-07,1.847899e-07,1.847903e-07,1.847907e-07,1.847912e-07,1.847916e-07,1.847920e-07,1.847925e-07,1.847929e-07,1.847933e-07,1.847937e-07,1.847942e-07,1.847946e-07,1.847950e-07,1.847955e-07,1.847959e-07,1.847963e-07,1.847967e-07,1.847972e-07,1.847976e-07,1.847980e-07,1.847985e-07,1.847989e-07,1.847993e-07,1.847997e-07,1.848002e-07,1.848006e-07,1.848010e-07,1.848015e-07,1.848019e-07,1.848023e-07,1.848027e-07,1.848032e-07,1.848036e-07,1.848040e-07,1.848044e-07,1.848049e-07,1.848053e-07,1.848057e-07,1.848062e-07,1.848066e-07,1.848070e-07,1.848074e-07,1.848079e-07,1.848083e-07,1.848087e-07,1.848092e-07,1.848096e-07,1.848100e-07,1.848104e-07,1.848109e-07,1.848113e-07,1.848117e-07,1.848122e-07,1.848126e-07,1.848130e-07,1.848134e-07,1.848139e-07,1.848143e-07,1.848147e-07,1.848151e-07,1.848156e-07,1.848160e-07,1.848164e-07,1.848169e-07,1.848173e-07,1.848177e-07,1.848181e-07,1.848186e-07,1.848190e-07,1.848194e-07,1.848199e-07,1.848203e-07,1.848207e-07,1.848211e-07,1.848216e-07,1.848220e-07,1.848224e-07,1.848228e-07,1.848233e-07,1.848237e-07,1.848241e-07,1.848246e-07,1.848250e-07,1.848254e-07,1.848258e-07,1.848263e-07,1.848267e-07,1.848271e-07,1.848276e-07,1.848280e-07,1.848284e-07,1.848288e-07,1.848293e-07,1.848297e-07,1.848301e-07,1.848305e-07,1.848310e-07,1.848314e-07,1.848318e-07,1.848323e-07,1.848327e-07,1.848331e-07,1.848335e-07,1.848340e-07,1.848344e-07,1.848348e-07,1.848352e-07,1.848357e-07,1.848361e-07,1.848365e-07,1.848369e-07,1.848374e-07,1.848378e-07,1.848382e-07,1.848387e-07,1.848391e-07,1.848395e-07,1.848399e-07,1.848404e-07,1.848408e-07,1.848412e-07,1.848416e-07,1.848421e-07,1.848425e-07,1.848429e-07,1.848434e-07,1.848438e-07,1.848442e-07,1.848446e-07,1.848451e-07,1.848455e-07,1.848459e-07,1.848463e-07,1.848468e-07,1.848472e-07,1.848476e-07,1.848480e-07,1.848485e-07,1.848489e-07,1.848493e-07,1.848498e-07,1.848502e-07,1.848506e-07,1.848510e-07,1.848515e-07,1.848519e-07,1.848523e-07,1.848527e-07,1.848532e-07,1.848536e-07,1.848540e-07,1.848544e-07,1.848549e-07,1.848553e-07,1.848557e-07,1.848561e-07,1.848566e-07,1.848570e-07,1.848574e-07,1.848579e-07,1.848583e-07,1.848587e-07,1.848591e-07,1.848596e-07,1.848600e-07,1.848604e-07,1.848608e-07,1.848613e-07,1.848617e-07,1.848621e-07,1.848625e-07,1.848630e-07,1.848634e-07,1.848638e-07,1.848642e-07,1.848647e-07,1.848651e-07,1.848655e-07,1.848659e-07,1.848664e-07,1.848668e-07,1.848672e-07,1.848677e-07,1.848681e-07,1.848685e-07,1.848689e-07,1.848694e-07,1.848698e-07,1.848702e-07,1.848706e-07,1.848711e-07,1.848715e-07,1.848719e-07,1.848723e-07,1.848728e-07,1.848732e-07,1.848736e-07,1.848740e-07,1.848745e-07,1.848749e-07,1.848753e-07,1.848757e-07,1.848762e-07,1.848766e-07,1.848770e-07,1.848774e-07,1.848779e-07,1.848783e-07,1.848787e-07,1.848791e-07,1.848796e-07,1.848800e-07,1.848804e-07,1.848808e-07,1.848813e-07,1.848817e-07,1.848821e-07,1.848826e-07,1.848830e-07,1.848834e-07,1.848838e-07,1.848843e-07,1.848847e-07,1.848851e-07,1.848855e-07,1.848860e-07,1.848864e-07,1.848868e-07,1.848872e-07,1.848877e-07,1.848881e-07,1.848885e-07,1.848889e-07,1.848894e-07,1.848898e-07,1.848902e-07,1.848906e-07,1.848911e-07,1.848915e-07,1.848919e-07,1.848923e-07,1.848928e-07,1.848932e-07,1.848936e-07,1.848940e-07,1.848945e-07,1.848949e-07,1.848953e-07,1.848957e-07,1.848962e-07,1.848966e-07,1.848970e-07,1.848974e-07,1.848979e-07,1.848983e-07,1.848987e-07,1.848991e-07,1.848996e-07,1.849000e-07,1.849004e-07,1.849008e-07,1.849013e-07,1.849017e-07,1.849021e-07,1.849025e-07,1.849029e-07,1.849034e-07,1.849038e-07,1.849042e-07,1.849046e-07,1.849051e-07,1.849055e-07,1.849059e-07,1.849063e-07,1.849068e-07,1.849072e-07,1.849076e-07,1.849080e-07,1.849085e-07,1.849089e-07,1.849093e-07,1.849097e-07,1.849102e-07,1.849106e-07,1.849110e-07,1.849114e-07,1.849119e-07,1.849123e-07,1.849127e-07,1.849131e-07,1.849136e-07,1.849140e-07,1.849144e-07,1.849148e-07,1.849153e-07,1.849157e-07,1.849161e-07,1.849165e-07,1.849170e-07,1.849174e-07,1.849178e-07,1.849182e-07,1.849187e-07,1.849191e-07,1.849195e-07,1.849199e-07,1.849203e-07,1.849208e-07,1.849212e-07,1.849216e-07,1.849220e-07,1.849225e-07,1.849229e-07,1.849233e-07,1.849237e-07,1.849242e-07,1.849246e-07,1.849250e-07,1.849254e-07,1.849259e-07,1.849263e-07,1.849267e-07,1.849271e-07,1.849276e-07,1.849280e-07,1.849284e-07,1.849288e-07,1.849292e-07,1.849297e-07,1.849301e-07,1.849305e-07,1.849309e-07,1.849314e-07,1.849318e-07,1.849322e-07,1.849326e-07,1.849331e-07,1.849335e-07,1.849339e-07,1.849343e-07,1.849348e-07,1.849352e-07,1.849356e-07,1.849360e-07,1.849364e-07,1.849369e-07,1.849373e-07,1.849377e-07,1.849381e-07,1.849386e-07,1.849390e-07,1.849394e-07,1.849398e-07,1.849403e-07,1.849407e-07,1.849411e-07,1.849415e-07,1.849419e-07,1.849424e-07,1.849428e-07,1.849432e-07,1.849436e-07,1.849441e-07,1.849445e-07,1.849449e-07,1.849453e-07,1.849458e-07,1.849462e-07,1.849466e-07,1.849470e-07,1.849474e-07,1.849479e-07,1.849483e-07,1.849487e-07,1.849491e-07,1.849496e-07,1.849500e-07,1.849504e-07,1.849508e-07,1.849513e-07,1.849517e-07,1.849521e-07,1.849525e-07,1.849529e-07,1.849534e-07,1.849538e-07,1.849542e-07,1.849546e-07,1.849551e-07,1.849555e-07,1.849559e-07,1.849563e-07,1.849568e-07,1.849572e-07,1.849576e-07,1.849580e-07,1.849584e-07,1.849589e-07,1.849593e-07,1.849597e-07,1.849601e-07,1.849606e-07,1.849610e-07,1.849614e-07,1.849618e-07,1.849622e-07,1.849627e-07,1.849631e-07,1.849635e-07,1.849639e-07,1.849644e-07,1.849648e-07,1.849652e-07,1.849656e-07,1.849660e-07,1.849665e-07,1.849669e-07,1.849673e-07,1.849677e-07,1.849682e-07,1.849686e-07,1.849690e-07,1.849694e-07,1.849698e-07,1.849703e-07,1.849707e-07,1.849711e-07,1.849715e-07,1.849720e-07,1.849724e-07,1.849728e-07,1.849732e-07,1.849736e-07,1.849741e-07,1.849745e-07,1.849749e-07,1.849753e-07,1.849758e-07,1.849762e-07,1.849766e-07,1.849770e-07,1.849774e-07,1.849779e-07,1.849783e-07,1.849787e-07,1.849791e-07,1.849796e-07,1.849800e-07,1.849804e-07,1.849808e-07,1.849812e-07,1.849817e-07,1.849821e-07,1.849825e-07,1.849829e-07,1.849833e-07,1.849838e-07,1.849842e-07,1.849846e-07,1.849850e-07,1.849855e-07,1.849859e-07,1.849863e-07,1.849867e-07,1.849871e-07,1.849876e-07,1.849880e-07,1.849884e-07,1.849888e-07,1.849893e-07,1.849897e-07,1.849901e-07,1.849905e-07,1.849909e-07,1.849914e-07,1.849918e-07,1.849922e-07,1.849926e-07,1.849930e-07,1.849935e-07,1.849939e-07,1.849943e-07,1.849947e-07,1.849952e-07,1.849956e-07,1.849960e-07,1.849964e-07,1.849968e-07,1.849973e-07,1.849977e-07,1.849981e-07,1.849985e-07,1.849989e-07,1.849994e-07,1.849998e-07,1.850002e-07,1.850006e-07,1.850010e-07,1.850015e-07,1.850019e-07,1.850023e-07,1.850027e-07,1.850032e-07,1.850036e-07,1.850040e-07,1.850044e-07,1.850048e-07,1.850053e-07,1.850057e-07,1.850061e-07,1.850065e-07,1.850069e-07,1.850074e-07,1.850078e-07,1.850082e-07,1.850086e-07,1.850090e-07,1.850095e-07,1.850099e-07,1.850103e-07,1.850107e-07,1.850111e-07,1.850116e-07,1.850120e-07,1.850124e-07,1.850128e-07,1.850133e-07,1.850137e-07,1.850141e-07,1.850145e-07,1.850149e-07,1.850154e-07,1.850158e-07,1.850162e-07,1.850166e-07,1.850170e-07,1.850175e-07,1.850179e-07,1.850183e-07,1.850187e-07,1.850191e-07,1.850196e-07,1.850200e-07,1.850204e-07,1.850208e-07,1.850212e-07,1.850217e-07,1.850221e-07,1.850225e-07,1.850229e-07,1.850233e-07,1.850238e-07,1.850242e-07,1.850246e-07,1.850250e-07,1.850254e-07,1.850259e-07,1.850263e-07,1.850267e-07,1.850271e-07,1.850275e-07,1.850280e-07,1.850284e-07,1.850288e-07,1.850292e-07,1.850296e-07,1.850301e-07,1.850305e-07,1.850309e-07,1.850313e-07,1.850317e-07,1.850322e-07,1.850326e-07,1.850330e-07,1.850334e-07,1.850338e-07,1.850343e-07,1.850347e-07,1.850351e-07,1.850355e-07,1.850359e-07,1.850364e-07,1.850368e-07,1.850372e-07,1.850376e-07,1.850380e-07,1.850385e-07,1.850389e-07,1.850393e-07,1.850397e-07,1.850401e-07,1.850406e-07,1.850410e-07,1.850414e-07,1.850418e-07,1.850422e-07,1.850427e-07,1.850431e-07,1.850435e-07,1.850439e-07,1.850443e-07,1.850448e-07,1.850452e-07,1.850456e-07,1.850460e-07,1.850464e-07,1.850469e-07,1.850473e-07,1.850477e-07,1.850481e-07,1.850485e-07,1.850489e-07,1.850494e-07,1.850498e-07,1.850502e-07,1.850506e-07,1.850510e-07,1.850515e-07,1.850519e-07,1.850523e-07,1.850527e-07,1.850531e-07,1.850536e-07,1.850540e-07,1.850544e-07,1.850548e-07,1.850552e-07,1.850557e-07,1.850561e-07,1.850565e-07,1.850569e-07,1.850573e-07,1.850578e-07,1.850582e-07,1.850586e-07,1.850590e-07,1.850594e-07,1.850598e-07,1.850603e-07,1.850607e-07,1.850611e-07,1.850615e-07,1.850619e-07,1.850624e-07,1.850628e-07,1.850632e-07,1.850636e-07,1.850640e-07,1.850645e-07,1.850649e-07,1.850653e-07,1.850657e-07,1.850661e-07,1.850665e-07,1.850670e-07,1.850674e-07,1.850678e-07,1.850682e-07,1.850686e-07,1.850691e-07,1.850695e-07,1.850699e-07,1.850703e-07,1.850707e-07,1.850712e-07,1.850716e-07,1.850720e-07,1.850724e-07,1.850728e-07,1.850732e-07,1.850737e-07,1.850741e-07,1.850745e-07,1.850749e-07,1.850753e-07,1.850758e-07,1.850762e-07,1.850766e-07,1.850770e-07,1.850774e-07,1.850778e-07,1.850783e-07,1.850787e-07,1.850791e-07,1.850795e-07,1.850799e-07,1.850804e-07,1.850808e-07,1.850812e-07,1.850816e-07,1.850820e-07,1.850824e-07,1.850829e-07,1.850833e-07,1.850837e-07,1.850841e-07,1.850845e-07,1.850850e-07,1.850854e-07,1.850858e-07,1.850862e-07,1.850866e-07,1.850870e-07,1.850875e-07,1.850879e-07,1.850883e-07,1.850887e-07,1.850891e-07,1.850896e-07,1.850900e-07,1.850904e-07,1.850908e-07,1.850912e-07,1.850916e-07,1.850921e-07,1.850925e-07,1.850929e-07,1.850933e-07,1.850937e-07,1.850942e-07,1.850946e-07,1.850950e-07,1.850954e-07,1.850958e-07,1.850962e-07,1.850967e-07,1.850971e-07,1.850975e-07,1.850979e-07,1.850983e-07,1.850987e-07,1.850992e-07,1.850996e-07,1.851000e-07,1.851004e-07,1.851008e-07,1.851012e-07,1.851017e-07,1.851021e-07,1.851025e-07,1.851029e-07,1.851033e-07,1.851038e-07,1.851042e-07,1.851046e-07,1.851050e-07,1.851054e-07,1.851058e-07,1.851063e-07,1.851067e-07,1.851071e-07,1.851075e-07,1.851079e-07,1.851083e-07,1.851088e-07,1.851092e-07,1.851096e-07,1.851100e-07,1.851104e-07,1.851108e-07,1.851113e-07,1.851117e-07,1.851121e-07,1.851125e-07,1.851129e-07,1.851133e-07,1.851138e-07,1.851142e-07,1.851146e-07,1.851150e-07,1.851154e-07,1.851159e-07,1.851163e-07,1.851167e-07,1.851171e-07,1.851175e-07,1.851179e-07,1.851184e-07,1.851188e-07,1.851192e-07,1.851196e-07,1.851200e-07,1.851204e-07,1.851209e-07,1.851213e-07,1.851217e-07,1.851221e-07,1.851225e-07,1.851229e-07,1.851234e-07,1.851238e-07,1.851242e-07,1.851246e-07,1.851250e-07,1.851254e-07,1.851259e-07,1.851263e-07,1.851267e-07,1.851271e-07,1.851275e-07,1.851279e-07,1.851284e-07,1.851288e-07,1.851292e-07,1.851296e-07,1.851300e-07,1.851304e-07,1.851309e-07,1.851313e-07,1.851317e-07,1.851321e-07,1.851325e-07,1.851329e-07,1.851334e-07,1.851338e-07,1.851342e-07,1.851346e-07,1.851350e-07,1.851354e-07,1.851358e-07,1.851363e-07,1.851367e-07,1.851371e-07,1.851375e-07,1.851379e-07,1.851383e-07,1.851388e-07,1.851392e-07,1.851396e-07,1.851400e-07,1.851404e-07,1.851408e-07,1.851413e-07,1.851417e-07,1.851421e-07,1.851425e-07,1.851429e-07,1.851433e-07,1.851438e-07,1.851442e-07,1.851446e-07,1.851450e-07,1.851454e-07,1.851458e-07,1.851462e-07,1.851467e-07,1.851471e-07,1.851475e-07,1.851479e-07,1.851483e-07,1.851487e-07,1.851492e-07,1.851496e-07,1.851500e-07,1.851504e-07,1.851508e-07,1.851512e-07,1.851517e-07,1.851521e-07,1.851525e-07,1.851529e-07,1.851533e-07,1.851537e-07,1.851541e-07,1.851546e-07,1.851550e-07,1.851554e-07,1.851558e-07,1.851562e-07,1.851566e-07,1.851571e-07,1.851575e-07,1.851579e-07,1.851583e-07,1.851587e-07,1.851591e-07,1.851595e-07,1.851600e-07,1.851604e-07,1.851608e-07,1.851612e-07,1.851616e-07,1.851620e-07,1.851625e-07,1.851629e-07,1.851633e-07,1.851637e-07,1.851641e-07,1.851645e-07,1.851649e-07,1.851654e-07,1.851658e-07,1.851662e-07,1.851666e-07,1.851670e-07,1.851674e-07,1.851679e-07,1.851683e-07,1.851687e-07,1.851691e-07,1.851695e-07,1.851699e-07,1.851703e-07,1.851708e-07,1.851712e-07,1.851716e-07,1.851720e-07,1.851724e-07,1.851728e-07,1.851732e-07,1.851737e-07,1.851741e-07,1.851745e-07,1.851749e-07,1.851753e-07,1.851757e-07,1.851762e-07,1.851766e-07,1.851770e-07,1.851774e-07,1.851778e-07,1.851782e-07,1.851786e-07,1.851791e-07,1.851795e-07,1.851799e-07,1.851803e-07,1.851807e-07,1.851811e-07,1.851815e-07,1.851820e-07,1.851824e-07,1.851828e-07,1.851832e-07,1.851836e-07,1.851840e-07,1.851844e-07,1.851849e-07,1.851853e-07,1.851857e-07,1.851861e-07,1.851865e-07,1.851869e-07,1.851873e-07,1.851878e-07,1.851882e-07,1.851886e-07,1.851890e-07,1.851894e-07,1.851898e-07,1.851902e-07,1.851907e-07,1.851911e-07,1.851915e-07,1.851919e-07,1.851923e-07,1.851927e-07,1.851931e-07,1.851936e-07,1.851940e-07,1.851944e-07,1.851948e-07,1.851952e-07,1.851956e-07,1.851960e-07,1.851965e-07,1.851969e-07,1.851973e-07,1.851977e-07,1.851981e-07,1.851985e-07,1.851989e-07,1.851994e-07,1.851998e-07,1.852002e-07,1.852006e-07,1.852010e-07,1.852014e-07,1.852018e-07,1.852023e-07,1.852027e-07,1.852031e-07,1.852035e-07,1.852039e-07,1.852043e-07,1.852047e-07,1.852052e-07,1.852056e-07,1.852060e-07,1.852064e-07,1.852068e-07,1.852072e-07,1.852076e-07,1.852080e-07,1.852085e-07,1.852089e-07,1.852093e-07,1.852097e-07,1.852101e-07,1.852105e-07,1.852109e-07,1.852114e-07,1.852118e-07,1.852122e-07,1.852126e-07,1.852130e-07,1.852134e-07,1.852138e-07,1.852143e-07,1.852147e-07,1.852151e-07,1.852155e-07,1.852159e-07,1.852163e-07,1.852167e-07,1.852171e-07,1.852176e-07,1.852180e-07,1.852184e-07,1.852188e-07,1.852192e-07,1.852196e-07,1.852200e-07,1.852205e-07,1.852209e-07,1.852213e-07,1.852217e-07,1.852221e-07,1.852225e-07,1.852229e-07,1.852233e-07,1.852238e-07,1.852242e-07,1.852246e-07,1.852250e-07,1.852254e-07,1.852258e-07,1.852262e-07,1.852266e-07,1.852271e-07,1.852275e-07,1.852279e-07,1.852283e-07,1.852287e-07,1.852291e-07,1.852295e-07,1.852300e-07,1.852304e-07,1.852308e-07,1.852312e-07,1.852316e-07,1.852320e-07,1.852324e-07,1.852328e-07,1.852333e-07,1.852337e-07,1.852341e-07,1.852345e-07,1.852349e-07,1.852353e-07,1.852357e-07,1.852361e-07,1.852366e-07,1.852370e-07,1.852374e-07,1.852378e-07,1.852382e-07,1.852386e-07,1.852390e-07,1.852394e-07,1.852399e-07,1.852403e-07,1.852407e-07,1.852411e-07,1.852415e-07,1.852419e-07,1.852423e-07,1.852427e-07,1.852432e-07,1.852436e-07,1.852440e-07,1.852444e-07,1.852448e-07,1.852452e-07,1.852456e-07,1.852460e-07,1.852465e-07,1.852469e-07,1.852473e-07,1.852477e-07,1.852481e-07,1.852485e-07,1.852489e-07,1.852493e-07,1.852498e-07,1.852502e-07,1.852506e-07,1.852510e-07,1.852514e-07,1.852518e-07,1.852522e-07,1.852526e-07,1.852531e-07,1.852535e-07,1.852539e-07,1.852543e-07,1.852547e-07,1.852551e-07,1.852555e-07,1.852559e-07,1.852563e-07,1.852568e-07,1.852572e-07,1.852576e-07,1.852580e-07,1.852584e-07,1.852588e-07,1.852592e-07,1.852596e-07,1.852601e-07,1.852605e-07,1.852609e-07,1.852613e-07,1.852617e-07,1.852621e-07,1.852625e-07,1.852629e-07,1.852633e-07,1.852638e-07,1.852642e-07,1.852646e-07,1.852650e-07,1.852654e-07,1.852658e-07,1.852662e-07,1.852666e-07,1.852671e-07,1.852675e-07,1.852679e-07,1.852683e-07,1.852687e-07,1.852691e-07,1.852695e-07,1.852699e-07,1.852703e-07,1.852708e-07,1.852712e-07,1.852716e-07,1.852720e-07,1.852724e-07,1.852728e-07,1.852732e-07,1.852736e-07,1.852740e-07,1.852745e-07,1.852749e-07,1.852753e-07,1.852757e-07,1.852761e-07,1.852765e-07,1.852769e-07,1.852773e-07,1.852777e-07,1.852782e-07,1.852786e-07,1.852790e-07,1.852794e-07,1.852798e-07,1.852802e-07,1.852806e-07,1.852810e-07,1.852814e-07,1.852819e-07,1.852823e-07,1.852827e-07,1.852831e-07,1.852835e-07,1.852839e-07,1.852843e-07,1.852847e-07,1.852851e-07,1.852856e-07,1.852860e-07,1.852864e-07,1.852868e-07,1.852872e-07,1.852876e-07,1.852880e-07,1.852884e-07,1.852888e-07,1.852893e-07,1.852897e-07,1.852901e-07,1.852905e-07,1.852909e-07,1.852913e-07,1.852917e-07,1.852921e-07,1.852925e-07,1.852930e-07,1.852934e-07,1.852938e-07,1.852942e-07,1.852946e-07,1.852950e-07,1.852954e-07,1.852958e-07,1.852962e-07,1.852966e-07,1.852971e-07,1.852975e-07,1.852979e-07,1.852983e-07,1.852987e-07,1.852991e-07,1.852995e-07,1.852999e-07,1.853003e-07,1.853008e-07,1.853012e-07,1.853016e-07,1.853020e-07,1.853024e-07,1.853028e-07,1.853032e-07,1.853036e-07,1.853040e-07,1.853044e-07,1.853049e-07,1.853053e-07,1.853057e-07,1.853061e-07,1.853065e-07,1.853069e-07,1.853073e-07,1.853077e-07,1.853081e-07,1.853085e-07,1.853090e-07,1.853094e-07,1.853098e-07,1.853102e-07,1.853106e-07,1.853110e-07,1.853114e-07,1.853118e-07,1.853122e-07,1.853126e-07,1.853131e-07,1.853135e-07,1.853139e-07,1.853143e-07,1.853147e-07,1.853151e-07,1.853155e-07,1.853159e-07,1.853163e-07,1.853167e-07,1.853172e-07,1.853176e-07,1.853180e-07,1.853184e-07,1.853188e-07,1.853192e-07,1.853196e-07,1.853200e-07,1.853204e-07,1.853208e-07,1.853213e-07,1.853217e-07,1.853221e-07,1.853225e-07,1.853229e-07,1.853233e-07,1.853237e-07,1.853241e-07,1.853245e-07,1.853249e-07,1.853254e-07,1.853258e-07,1.853262e-07,1.853266e-07,1.853270e-07,1.853274e-07,1.853278e-07,1.853282e-07,1.853286e-07,1.853290e-07,1.853294e-07,1.853299e-07,1.853303e-07,1.853307e-07,1.853311e-07,1.853315e-07,1.853319e-07,1.853323e-07,1.853327e-07,1.853331e-07,1.853335e-07,1.853339e-07,1.853344e-07,1.853348e-07,1.853352e-07,1.853356e-07,1.853360e-07,1.853364e-07,1.853368e-07,1.853372e-07,1.853376e-07,1.853380e-07,1.853384e-07,1.853389e-07,1.853393e-07,1.853397e-07,1.853401e-07,1.853405e-07,1.853409e-07,1.853413e-07,1.853417e-07,1.853421e-07,1.853425e-07,1.853429e-07,1.853434e-07,1.853438e-07,1.853442e-07,1.853446e-07,1.853450e-07,1.853454e-07,1.853458e-07,1.853462e-07,1.853466e-07,1.853470e-07,1.853474e-07,1.853479e-07,1.853483e-07,1.853487e-07,1.853491e-07,1.853495e-07,1.853499e-07,1.853503e-07,1.853507e-07,1.853511e-07,1.853515e-07,1.853519e-07,1.853523e-07,1.853528e-07,1.853532e-07,1.853536e-07,1.853540e-07,1.853544e-07,1.853548e-07,1.853552e-07,1.853556e-07,1.853560e-07,1.853564e-07,1.853568e-07,1.853572e-07,1.853577e-07,1.853581e-07,1.853585e-07,1.853589e-07,1.853593e-07,1.853597e-07,1.853601e-07,1.853605e-07,1.853609e-07,1.853613e-07,1.853617e-07,1.853621e-07,1.853626e-07,1.853630e-07,1.853634e-07,1.853638e-07,1.853642e-07,1.853646e-07,1.853650e-07,1.853654e-07,1.853658e-07,1.853662e-07,1.853666e-07,1.853670e-07,1.853675e-07,1.853679e-07,1.853683e-07,1.853687e-07,1.853691e-07,1.853695e-07,1.853699e-07,1.853703e-07,1.853707e-07,1.853711e-07,1.853715e-07,1.853719e-07,1.853724e-07,1.853728e-07,1.853732e-07,1.853736e-07,1.853740e-07,1.853744e-07,1.853748e-07,1.853752e-07,1.853756e-07,1.853760e-07,1.853764e-07,1.853768e-07,1.853772e-07,1.853777e-07,1.853781e-07,1.853785e-07,1.853789e-07,1.853793e-07,1.853797e-07,1.853801e-07,1.853805e-07,1.853809e-07,1.853813e-07,1.853817e-07,1.853821e-07,1.853825e-07,1.853830e-07,1.853834e-07,1.853838e-07,1.853842e-07,1.853846e-07,1.853850e-07,1.853854e-07,1.853858e-07,1.853862e-07,1.853866e-07,1.853870e-07,1.853874e-07,1.853878e-07,1.853882e-07,1.853887e-07,1.853891e-07,1.853895e-07,1.853899e-07,1.853903e-07,1.853907e-07,1.853911e-07,1.853915e-07,1.853919e-07,1.853923e-07,1.853927e-07,1.853931e-07,1.853935e-07,1.853939e-07,1.853944e-07,1.853948e-07,1.853952e-07,1.853956e-07,1.853960e-07,1.853964e-07,1.853968e-07,1.853972e-07,1.853976e-07,1.853980e-07,1.853984e-07,1.853988e-07,1.853992e-07,1.853996e-07,1.854001e-07,1.854005e-07,1.854009e-07,1.854013e-07,1.854017e-07,1.854021e-07,1.854025e-07,1.854029e-07,1.854033e-07,1.854037e-07,1.854041e-07,1.854045e-07,1.854049e-07,1.854053e-07,1.854057e-07,1.854062e-07,1.854066e-07,1.854070e-07,1.854074e-07,1.854078e-07,1.854082e-07,1.854086e-07,1.854090e-07,1.854094e-07,1.854098e-07,1.854102e-07,1.854106e-07,1.854110e-07,1.854114e-07,1.854118e-07,1.854123e-07,1.854127e-07,1.854131e-07,1.854135e-07,1.854139e-07,1.854143e-07,1.854147e-07,1.854151e-07,1.854155e-07,1.854159e-07,1.854163e-07,1.854167e-07,1.854171e-07,1.854175e-07,1.854179e-07,1.854184e-07,1.854188e-07,1.854192e-07,1.854196e-07,1.854200e-07,1.854204e-07,1.854208e-07,1.854212e-07,1.854216e-07,1.854220e-07,1.854224e-07,1.854228e-07,1.854232e-07,1.854236e-07,1.854240e-07,1.854244e-07,1.854248e-07,1.854253e-07,1.854257e-07,1.854261e-07,1.854265e-07,1.854269e-07,1.854273e-07,1.854277e-07,1.854281e-07,1.854285e-07,1.854289e-07,1.854293e-07,1.854297e-07,1.854301e-07,1.854305e-07,1.854309e-07,1.854313e-07,1.854318e-07,1.854322e-07,1.854326e-07,1.854330e-07,1.854334e-07,1.854338e-07,1.854342e-07,1.854346e-07,1.854350e-07,1.854354e-07,1.854358e-07,1.854362e-07,1.854366e-07,1.854370e-07,1.854374e-07,1.854378e-07,1.854382e-07,1.854386e-07,1.854391e-07,1.854395e-07,1.854399e-07,1.854403e-07,1.854407e-07,1.854411e-07,1.854415e-07,1.854419e-07,1.854423e-07,1.854427e-07,1.854431e-07,1.854435e-07,1.854439e-07,1.854443e-07,1.854447e-07,1.854451e-07,1.854455e-07,1.854459e-07,1.854464e-07,1.854468e-07,1.854472e-07,1.854476e-07,1.854480e-07,1.854484e-07,1.854488e-07,1.854492e-07,1.854496e-07,1.854500e-07,1.854504e-07,1.854508e-07,1.854512e-07,1.854516e-07,1.854520e-07,1.854524e-07,1.854528e-07,1.854532e-07,1.854536e-07,1.854540e-07,1.854545e-07,1.854549e-07,1.854553e-07,1.854557e-07,1.854561e-07,1.854565e-07,1.854569e-07,1.854573e-07,1.854577e-07,1.854581e-07,1.854585e-07,1.854589e-07,1.854593e-07,1.854597e-07,1.854601e-07,1.854605e-07,1.854609e-07,1.854613e-07,1.854617e-07,1.854621e-07,1.854626e-07,1.854630e-07,1.854634e-07,1.854638e-07,1.854642e-07,1.854646e-07,1.854650e-07,1.854654e-07,1.854658e-07,1.854662e-07,1.854666e-07,1.854670e-07,1.854674e-07,1.854678e-07,1.854682e-07,1.854686e-07,1.854690e-07,1.854694e-07,1.854698e-07,1.854702e-07,1.854706e-07,1.854710e-07,1.854715e-07,1.854719e-07,1.854723e-07,1.854727e-07,1.854731e-07,1.854735e-07,1.854739e-07,1.854743e-07,1.854747e-07,1.854751e-07,1.854755e-07,1.854759e-07,1.854763e-07,1.854767e-07,1.854771e-07,1.854775e-07,1.854779e-07,1.854783e-07,1.854787e-07,1.854791e-07,1.854795e-07,1.854799e-07,1.854803e-07,1.854808e-07,1.854812e-07,1.854816e-07,1.854820e-07,1.854824e-07,1.854828e-07,1.854832e-07,1.854836e-07,1.854840e-07,1.854844e-07,1.854848e-07,1.854852e-07,1.854856e-07,1.854860e-07,1.854864e-07,1.854868e-07,1.854872e-07,1.854876e-07,1.854880e-07,1.854884e-07,1.854888e-07,1.854892e-07,1.854896e-07,1.854900e-07,1.854904e-07,1.854908e-07,1.854913e-07,1.854917e-07,1.854921e-07,1.854925e-07,1.854929e-07,1.854933e-07,1.854937e-07,1.854941e-07,1.854945e-07,1.854949e-07,1.854953e-07,1.854957e-07,1.854961e-07,1.854965e-07,1.854969e-07,1.854973e-07,1.854977e-07,1.854981e-07,1.854985e-07,1.854989e-07,1.854993e-07,1.854997e-07,1.855001e-07,1.855005e-07,1.855009e-07,1.855013e-07,1.855017e-07,1.855021e-07,1.855026e-07,1.855030e-07,1.855034e-07,1.855038e-07,1.855042e-07,1.855046e-07,1.855050e-07,1.855054e-07,1.855058e-07,1.855062e-07,1.855066e-07,1.855070e-07,1.855074e-07,1.855078e-07,1.855082e-07,1.855086e-07,1.855090e-07,1.855094e-07,1.855098e-07,1.855102e-07,1.855106e-07,1.855110e-07,1.855114e-07,1.855118e-07,1.855122e-07,1.855126e-07,1.855130e-07,1.855134e-07,1.855138e-07,1.855142e-07,1.855146e-07,1.855151e-07,1.855155e-07,1.855159e-07,1.855163e-07,1.855167e-07,1.855171e-07,1.855175e-07,1.855179e-07,1.855183e-07,1.855187e-07,1.855191e-07,1.855195e-07,1.855199e-07,1.855203e-07,1.855207e-07,1.855211e-07,1.855215e-07,1.855219e-07,1.855223e-07,1.855227e-07,1.855231e-07,1.855235e-07,1.855239e-07,1.855243e-07,1.855247e-07,1.855251e-07,1.855255e-07,1.855259e-07,1.855263e-07,1.855267e-07,1.855271e-07,1.855275e-07,1.855279e-07,1.855283e-07,1.855287e-07,1.855291e-07,1.855295e-07,1.855299e-07,1.855304e-07,1.855308e-07,1.855312e-07,1.855316e-07,1.855320e-07,1.855324e-07,1.855328e-07,1.855332e-07,1.855336e-07,1.855340e-07,1.855344e-07,1.855348e-07,1.855352e-07,1.855356e-07,1.855360e-07,1.855364e-07,1.855368e-07,1.855372e-07,1.855376e-07,1.855380e-07,1.855384e-07,1.855388e-07,1.855392e-07,1.855396e-07,1.855400e-07,1.855404e-07,1.855408e-07,1.855412e-07,1.855416e-07,1.855420e-07,1.855424e-07,1.855428e-07,1.855432e-07,1.855436e-07,1.855440e-07,1.855444e-07,1.855448e-07,1.855452e-07,1.855456e-07,1.855460e-07,1.855464e-07,1.855468e-07,1.855472e-07,1.855476e-07,1.855480e-07,1.855484e-07,1.855488e-07,1.855492e-07,1.855497e-07,1.855501e-07,1.855505e-07,1.855509e-07,1.855513e-07,1.855517e-07,1.855521e-07,1.855525e-07,1.855529e-07,1.855533e-07,1.855537e-07,1.855541e-07,1.855545e-07,1.855549e-07,1.855553e-07,1.855557e-07,1.855561e-07,1.855565e-07,1.855569e-07,1.855573e-07,1.855577e-07,1.855581e-07,1.855585e-07,1.855589e-07,1.855593e-07,1.855597e-07,1.855601e-07,1.855605e-07,1.855609e-07,1.855613e-07,1.855617e-07,1.855621e-07,1.855625e-07,1.855629e-07,1.855633e-07,1.855637e-07,1.855641e-07,1.855645e-07,1.855649e-07,1.855653e-07,1.855657e-07,1.855661e-07,1.855665e-07,1.855669e-07,1.855673e-07,1.855677e-07,1.855681e-07,1.855685e-07,1.855689e-07,1.855693e-07,1.855697e-07,1.855701e-07,1.855705e-07,1.855709e-07,1.855713e-07,1.855717e-07,1.855721e-07,1.855725e-07,1.855729e-07,1.855733e-07,1.855737e-07,1.855741e-07,1.855745e-07,1.855749e-07,1.855753e-07,1.855757e-07,1.855761e-07,1.855765e-07,1.855769e-07,1.855773e-07,1.855777e-07,1.855781e-07,1.855785e-07,1.855789e-07,1.855793e-07,1.855797e-07,1.855801e-07,1.855805e-07,1.855809e-07,1.855813e-07,1.855817e-07,1.855821e-07,1.855825e-07,1.855829e-07,1.855833e-07,1.855837e-07,1.855841e-07,1.855845e-07,1.855849e-07,1.855854e-07,1.855858e-07,1.855862e-07,1.855866e-07,1.855870e-07,1.855874e-07,1.855878e-07,1.855882e-07,1.855886e-07,1.855890e-07,1.855894e-07,1.855898e-07,1.855902e-07,1.855906e-07,1.855910e-07,1.855914e-07,1.855918e-07,1.855922e-07,1.855926e-07,1.855930e-07,1.855934e-07,1.855938e-07,1.855942e-07,1.855946e-07,1.855950e-07,1.855954e-07,1.855958e-07,1.855962e-07,1.855966e-07,1.855970e-07,1.855974e-07,1.855978e-07,1.855982e-07,1.855986e-07,1.855990e-07,1.855994e-07,1.855998e-07,1.856002e-07,1.856006e-07,1.856010e-07,1.856014e-07,1.856018e-07,1.856022e-07,1.856026e-07,1.856030e-07,1.856034e-07,1.856038e-07,1.856042e-07,1.856046e-07,1.856050e-07,1.856054e-07,1.856058e-07,1.856062e-07,1.856066e-07,1.856070e-07,1.856074e-07,1.856078e-07,1.856082e-07,1.856086e-07,1.856090e-07,1.856094e-07,1.856098e-07,1.856102e-07,1.856106e-07,1.856110e-07,1.856114e-07,1.856118e-07,1.856122e-07,1.856126e-07,1.856130e-07,1.856134e-07,1.856138e-07,1.856142e-07,1.856146e-07,1.856150e-07,1.856153e-07,1.856157e-07,1.856161e-07,1.856165e-07,1.856169e-07,1.856173e-07,1.856177e-07,1.856181e-07,1.856185e-07,1.856189e-07,1.856193e-07,1.856197e-07,1.856201e-07,1.856205e-07,1.856209e-07,1.856213e-07,1.856217e-07,1.856221e-07,1.856225e-07,1.856229e-07,1.856233e-07,1.856237e-07,1.856241e-07,1.856245e-07,1.856249e-07,1.856253e-07,1.856257e-07,1.856261e-07,1.856265e-07,1.856269e-07,1.856273e-07,1.856277e-07,1.856281e-07,1.856285e-07,1.856289e-07,1.856293e-07,1.856297e-07,1.856301e-07,1.856305e-07,1.856309e-07,1.856313e-07,1.856317e-07,1.856321e-07,1.856325e-07,1.856329e-07,1.856333e-07,1.856337e-07,1.856341e-07,1.856345e-07,1.856349e-07,1.856353e-07,1.856357e-07,1.856361e-07,1.856365e-07,1.856369e-07,1.856373e-07,1.856377e-07,1.856381e-07,1.856385e-07,1.856389e-07,1.856393e-07,1.856397e-07,1.856401e-07,1.856405e-07,1.856409e-07,1.856413e-07,1.856417e-07,1.856421e-07,1.856425e-07,1.856429e-07,1.856433e-07,1.856437e-07,1.856441e-07,1.856445e-07,1.856449e-07,1.856453e-07,1.856457e-07,1.856461e-07,1.856465e-07,1.856469e-07,1.856473e-07,1.856477e-07,1.856481e-07,1.856485e-07,1.856489e-07,1.856493e-07,1.856497e-07,1.856501e-07,1.856505e-07,1.856508e-07,1.856512e-07,1.856516e-07,1.856520e-07,1.856524e-07,1.856528e-07,1.856532e-07,1.856536e-07,1.856540e-07,1.856544e-07,1.856548e-07,1.856552e-07,1.856556e-07,1.856560e-07,1.856564e-07,1.856568e-07,1.856572e-07,1.856576e-07,1.856580e-07,1.856584e-07,1.856588e-07,1.856592e-07,1.856596e-07,1.856600e-07,1.856604e-07,1.856608e-07,1.856612e-07,1.856616e-07,1.856620e-07,1.856624e-07,1.856628e-07,1.856632e-07,1.856636e-07,1.856640e-07,1.856644e-07,1.856648e-07,1.856652e-07,1.856656e-07,1.856660e-07,1.856664e-07,1.856668e-07,1.856672e-07,1.856676e-07,1.856680e-07,1.856684e-07,1.856688e-07,1.856692e-07,1.856696e-07,1.856700e-07,1.856703e-07,1.856707e-07,1.856711e-07,1.856715e-07,1.856719e-07,1.856723e-07,1.856727e-07,1.856731e-07,1.856735e-07,1.856739e-07,1.856743e-07,1.856747e-07,1.856751e-07,1.856755e-07,1.856759e-07,1.856763e-07,1.856767e-07,1.856771e-07,1.856775e-07,1.856779e-07,1.856783e-07,1.856787e-07,1.856791e-07,1.856795e-07,1.856799e-07,1.856803e-07,1.856807e-07,1.856811e-07,1.856815e-07,1.856819e-07,1.856823e-07,1.856827e-07,1.856831e-07,1.856835e-07,1.856839e-07,1.856843e-07,1.856847e-07,1.856851e-07,1.856854e-07,1.856858e-07,1.856862e-07,1.856866e-07,1.856870e-07,1.856874e-07,1.856878e-07,1.856882e-07,1.856886e-07,1.856890e-07,1.856894e-07,1.856898e-07,1.856902e-07,1.856906e-07,1.856910e-07,1.856914e-07,1.856918e-07,1.856922e-07,1.856926e-07,1.856930e-07,1.856934e-07,1.856938e-07,1.856942e-07,1.856946e-07,1.856950e-07,1.856954e-07,1.856958e-07,1.856962e-07,1.856966e-07,1.856970e-07,1.856974e-07,1.856978e-07,1.856981e-07,1.856985e-07,1.856989e-07,1.856993e-07,1.856997e-07,1.857001e-07,1.857005e-07,1.857009e-07,1.857013e-07,1.857017e-07,1.857021e-07,1.857025e-07,1.857029e-07,1.857033e-07,1.857037e-07,1.857041e-07,1.857045e-07,1.857049e-07,1.857053e-07,1.857057e-07,1.857061e-07,1.857065e-07,1.857069e-07,1.857073e-07,1.857077e-07,1.857081e-07,1.857085e-07,1.857089e-07,1.857092e-07,1.857096e-07,1.857100e-07,1.857104e-07,1.857108e-07,1.857112e-07,1.857116e-07,1.857120e-07,1.857124e-07,1.857128e-07,1.857132e-07,1.857136e-07,1.857140e-07,1.857144e-07,1.857148e-07,1.857152e-07,1.857156e-07,1.857160e-07,1.857164e-07,1.857168e-07,1.857172e-07,1.857176e-07,1.857180e-07,1.857184e-07,1.857188e-07,1.857192e-07,1.857195e-07,1.857199e-07,1.857203e-07,1.857207e-07,1.857211e-07,1.857215e-07,1.857219e-07,1.857223e-07,1.857227e-07,1.857231e-07,1.857235e-07,1.857239e-07,1.857243e-07,1.857247e-07,1.857251e-07,1.857255e-07,1.857259e-07,1.857263e-07,1.857267e-07,1.857271e-07,1.857275e-07,1.857279e-07,1.857283e-07,1.857287e-07,1.857290e-07,1.857294e-07,1.857298e-07,1.857302e-07,1.857306e-07,1.857310e-07,1.857314e-07,1.857318e-07,1.857322e-07,1.857326e-07,1.857330e-07,1.857334e-07,1.857338e-07,1.857342e-07,1.857346e-07,1.857350e-07,1.857354e-07,1.857358e-07,1.857362e-07,1.857366e-07,1.857370e-07,1.857374e-07,1.857377e-07,1.857381e-07,1.857385e-07,1.857389e-07,1.857393e-07,1.857397e-07,1.857401e-07,1.857405e-07,1.857409e-07,1.857413e-07,1.857417e-07,1.857421e-07,1.857425e-07,1.857429e-07,1.857433e-07,1.857437e-07,1.857441e-07,1.857445e-07,1.857449e-07,1.857453e-07,1.857456e-07,1.857460e-07,1.857464e-07,1.857468e-07,1.857472e-07,1.857476e-07,1.857480e-07,1.857484e-07,1.857488e-07,1.857492e-07,1.857496e-07,1.857500e-07,1.857504e-07,1.857508e-07,1.857512e-07,1.857516e-07,1.857520e-07,1.857524e-07,1.857528e-07,1.857532e-07,1.857535e-07,1.857539e-07,1.857543e-07,1.857547e-07,1.857551e-07,1.857555e-07,1.857559e-07,1.857563e-07,1.857567e-07,1.857571e-07,1.857575e-07,1.857579e-07,1.857583e-07,1.857587e-07,1.857591e-07,1.857595e-07,1.857599e-07,1.857603e-07,1.857607e-07,1.857610e-07,1.857614e-07,1.857618e-07,1.857622e-07,1.857626e-07,1.857630e-07,1.857634e-07,1.857638e-07,1.857642e-07,1.857646e-07,1.857650e-07,1.857654e-07,1.857658e-07,1.857662e-07,1.857666e-07,1.857670e-07,1.857674e-07,1.857678e-07,1.857681e-07,1.857685e-07,1.857689e-07,1.857693e-07,1.857697e-07,1.857701e-07,1.857705e-07,1.857709e-07,1.857713e-07,1.857717e-07,1.857721e-07,1.857725e-07,1.857729e-07,1.857733e-07,1.857737e-07,1.857741e-07,1.857745e-07,1.857748e-07,1.857752e-07,1.857756e-07,1.857760e-07,1.857764e-07,1.857768e-07,1.857772e-07,1.857776e-07,1.857780e-07,1.857784e-07,1.857788e-07,1.857792e-07,1.857796e-07,1.857800e-07,1.857804e-07,1.857808e-07,1.857812e-07,1.857815e-07,1.857819e-07,1.857823e-07,1.857827e-07,1.857831e-07,1.857835e-07,1.857839e-07,1.857843e-07,1.857847e-07,1.857851e-07,1.857855e-07,1.857859e-07,1.857863e-07,1.857867e-07,1.857871e-07,1.857875e-07,1.857878e-07,1.857882e-07,1.857886e-07,1.857890e-07,1.857894e-07,1.857898e-07,1.857902e-07,1.857906e-07,1.857910e-07,1.857914e-07,1.857918e-07,1.857922e-07,1.857926e-07,1.857930e-07,1.857934e-07,1.857937e-07,1.857941e-07,1.857945e-07,1.857949e-07,1.857953e-07,1.857957e-07,1.857961e-07,1.857965e-07,1.857969e-07,1.857973e-07,1.857977e-07,1.857981e-07,1.857985e-07,1.857989e-07,1.857993e-07,1.857996e-07,1.858000e-07,1.858004e-07,1.858008e-07,1.858012e-07,1.858016e-07,1.858020e-07,1.858024e-07,1.858028e-07,1.858032e-07,1.858036e-07,1.858040e-07,1.858044e-07,1.858048e-07,1.858052e-07,1.858055e-07,1.858059e-07,1.858063e-07,1.858067e-07,1.858071e-07,1.858075e-07,1.858079e-07,1.858083e-07,1.858087e-07,1.858091e-07,1.858095e-07,1.858099e-07,1.858103e-07,1.858107e-07,1.858110e-07,1.858114e-07,1.858118e-07,1.858122e-07,1.858126e-07,1.858130e-07,1.858134e-07,1.858138e-07,1.858142e-07,1.858146e-07,1.858150e-07,1.858154e-07,1.858158e-07,1.858162e-07,1.858165e-07,1.858169e-07,1.858173e-07,1.858177e-07,1.858181e-07,1.858185e-07,1.858189e-07,1.858193e-07,1.858197e-07,1.858201e-07,1.858205e-07,1.858209e-07,1.858213e-07,1.858216e-07,1.858220e-07,1.858224e-07,1.858228e-07,1.858232e-07,1.858236e-07,1.858240e-07,1.858244e-07,1.858248e-07,1.858252e-07,1.858256e-07,1.858260e-07,1.858264e-07,1.858267e-07,1.858271e-07,1.858275e-07,1.858279e-07,1.858283e-07,1.858287e-07,1.858291e-07,1.858295e-07,1.858299e-07,1.858303e-07,1.858307e-07,1.858311e-07,1.858315e-07,1.858318e-07,1.858322e-07,1.858326e-07,1.858330e-07,1.858334e-07,1.858338e-07,1.858342e-07,1.858346e-07,1.858350e-07,1.858354e-07,1.858358e-07,1.858362e-07,1.858366e-07,1.858369e-07,1.858373e-07,1.858377e-07,1.858381e-07,1.858385e-07,1.858389e-07,1.858393e-07,1.858397e-07,1.858401e-07,1.858405e-07,1.858409e-07,1.858413e-07,1.858416e-07,1.858420e-07,1.858424e-07,1.858428e-07,1.858432e-07,1.858436e-07,1.858440e-07,1.858444e-07,1.858448e-07,1.858452e-07,1.858456e-07,1.858460e-07,1.858463e-07,1.858467e-07,1.858471e-07,1.858475e-07,1.858479e-07,1.858483e-07,1.858487e-07,1.858491e-07,1.858495e-07,1.858499e-07,1.858503e-07,1.858507e-07,1.858510e-07,1.858514e-07,1.858518e-07,1.858522e-07,1.858526e-07,1.858530e-07,1.858534e-07,1.858538e-07,1.858542e-07,1.858546e-07,1.858550e-07,1.858554e-07,1.858557e-07,1.858561e-07,1.858565e-07,1.858569e-07,1.858573e-07,1.858577e-07,1.858581e-07,1.858585e-07,1.858589e-07,1.858593e-07,1.858597e-07,1.858600e-07,1.858604e-07,1.858608e-07,1.858612e-07,1.858616e-07,1.858620e-07,1.858624e-07,1.858628e-07,1.858632e-07,1.858636e-07,1.858640e-07,1.858643e-07,1.858647e-07,1.858651e-07,1.858655e-07,1.858659e-07,1.858663e-07,1.858667e-07,1.858671e-07,1.858675e-07,1.858679e-07,1.858683e-07,1.858686e-07,1.858690e-07,1.858694e-07,1.858698e-07,1.858702e-07,1.858706e-07,1.858710e-07,1.858714e-07,1.858718e-07,1.858722e-07,1.858726e-07,1.858729e-07,1.858733e-07,1.858737e-07,1.858741e-07,1.858745e-07,1.858749e-07,1.858753e-07,1.858757e-07,1.858761e-07,1.858765e-07,1.858769e-07,1.858772e-07,1.858776e-07,1.858780e-07,1.858784e-07,1.858788e-07,1.858792e-07,1.858796e-07,1.858800e-07,1.858804e-07,1.858808e-07,1.858812e-07,1.858815e-07,1.858819e-07,1.858823e-07,1.858827e-07,1.858831e-07,1.858835e-07,1.858839e-07,1.858843e-07,1.858847e-07,1.858851e-07,1.858854e-07,1.858858e-07,1.858862e-07,1.858866e-07,1.858870e-07,1.858874e-07,1.858878e-07,1.858882e-07,1.858886e-07,1.858890e-07,1.858893e-07,1.858897e-07,1.858901e-07,1.858905e-07,1.858909e-07,1.858913e-07,1.858917e-07,1.858921e-07,1.858925e-07,1.858929e-07,1.858933e-07,1.858936e-07,1.858940e-07,1.858944e-07,1.858948e-07,1.858952e-07,1.858956e-07,1.858960e-07,1.858964e-07,1.858968e-07,1.858972e-07,1.858975e-07,1.858979e-07,1.858983e-07,1.858987e-07,1.858991e-07,1.858995e-07,1.858999e-07,1.859003e-07,1.859007e-07,1.859011e-07,1.859014e-07,1.859018e-07,1.859022e-07,1.859026e-07,1.859030e-07,1.859034e-07,1.859038e-07,1.859042e-07,1.859046e-07,1.859049e-07,1.859053e-07,1.859057e-07,1.859061e-07,1.859065e-07,1.859069e-07,1.859073e-07,1.859077e-07,1.859081e-07,1.859085e-07,1.859088e-07,1.859092e-07,1.859096e-07,1.859100e-07,1.859104e-07,1.859108e-07,1.859112e-07,1.859116e-07,1.859120e-07,1.859123e-07,1.859127e-07,1.859131e-07,1.859135e-07,1.859139e-07,1.859143e-07,1.859147e-07,1.859151e-07,1.859155e-07,1.859159e-07,1.859162e-07,1.859166e-07,1.859170e-07,1.859174e-07,1.859178e-07,1.859182e-07,1.859186e-07,1.859190e-07,1.859194e-07,1.859197e-07,1.859201e-07,1.859205e-07,1.859209e-07,1.859213e-07,1.859217e-07,1.859221e-07,1.859225e-07,1.859229e-07,1.859232e-07,1.859236e-07,1.859240e-07,1.859244e-07,1.859248e-07,1.859252e-07,1.859256e-07,1.859260e-07,1.859264e-07,1.859268e-07,1.859271e-07,1.859275e-07,1.859279e-07,1.859283e-07,1.859287e-07,1.859291e-07,1.859295e-07,1.859299e-07,1.859303e-07,1.859306e-07,1.859310e-07,1.859314e-07,1.859318e-07,1.859322e-07,1.859326e-07,1.859330e-07,1.859334e-07,1.859337e-07,1.859341e-07,1.859345e-07,1.859349e-07,1.859353e-07,1.859357e-07,1.859361e-07,1.859365e-07,1.859369e-07,1.859372e-07,1.859376e-07,1.859380e-07,1.859384e-07,1.859388e-07,1.859392e-07,1.859396e-07,1.859400e-07,1.859404e-07,1.859407e-07,1.859411e-07,1.859415e-07,1.859419e-07,1.859423e-07,1.859427e-07,1.859431e-07,1.859435e-07,1.859439e-07,1.859442e-07,1.859446e-07,1.859450e-07,1.859454e-07,1.859458e-07,1.859462e-07,1.859466e-07,1.859470e-07,1.859473e-07,1.859477e-07,1.859481e-07,1.859485e-07,1.859489e-07,1.859493e-07,1.859497e-07,1.859501e-07,1.859505e-07,1.859508e-07,1.859512e-07,1.859516e-07,1.859520e-07,1.859524e-07,1.859528e-07,1.859532e-07,1.859536e-07,1.859539e-07,1.859543e-07,1.859547e-07,1.859551e-07,1.859555e-07,1.859559e-07,1.859563e-07,1.859567e-07,1.859571e-07,1.859574e-07,1.859578e-07,1.859582e-07,1.859586e-07,1.859590e-07,1.859594e-07,1.859598e-07,1.859602e-07,1.859605e-07,1.859609e-07,1.859613e-07,1.859617e-07,1.859621e-07,1.859625e-07,1.859629e-07,1.859633e-07,1.859636e-07,1.859640e-07,1.859644e-07,1.859648e-07,1.859652e-07,1.859656e-07,1.859660e-07,1.859664e-07,1.859667e-07,1.859671e-07,1.859675e-07,1.859679e-07,1.859683e-07,1.859687e-07,1.859691e-07,1.859695e-07,1.859698e-07,1.859702e-07,1.859706e-07,1.859710e-07,1.859714e-07,1.859718e-07,1.859722e-07,1.859726e-07,1.859729e-07,1.859733e-07,1.859737e-07,1.859741e-07,1.859745e-07,1.859749e-07,1.859753e-07,1.859757e-07,1.859760e-07,1.859764e-07,1.859768e-07,1.859772e-07,1.859776e-07,1.859780e-07,1.859784e-07,1.859788e-07,1.859791e-07,1.859795e-07,1.859799e-07,1.859803e-07,1.859807e-07,1.859811e-07,1.859815e-07,1.859819e-07,1.859822e-07,1.859826e-07,1.859830e-07,1.859834e-07,1.859838e-07,1.859842e-07,1.859846e-07,1.859850e-07,1.859853e-07,1.859857e-07,1.859861e-07,1.859865e-07,1.859869e-07,1.859873e-07,1.859877e-07,1.859880e-07,1.859884e-07,1.859888e-07,1.859892e-07,1.859896e-07,1.859900e-07,1.859904e-07,1.859908e-07,1.859911e-07,1.859915e-07,1.859919e-07,1.859923e-07,1.859927e-07,1.859931e-07,1.859935e-07,1.859938e-07,1.859942e-07,1.859946e-07,1.859950e-07,1.859954e-07,1.859958e-07,1.859962e-07,1.859966e-07,1.859969e-07,1.859973e-07,1.859977e-07,1.859981e-07,1.859985e-07,1.859989e-07,1.859993e-07,1.859996e-07,1.860000e-07,1.860004e-07,1.860008e-07,1.860012e-07,1.860016e-07,1.860020e-07,1.860024e-07,1.860027e-07,1.860031e-07,1.860035e-07,1.860039e-07,1.860043e-07,1.860047e-07,1.860051e-07,1.860054e-07,1.860058e-07,1.860062e-07,1.860066e-07,1.860070e-07,1.860074e-07,1.860078e-07,1.860081e-07,1.860085e-07,1.860089e-07,1.860093e-07,1.860097e-07,1.860101e-07,1.860105e-07,1.860109e-07,1.860112e-07,1.860116e-07,1.860120e-07,1.860124e-07,1.860128e-07,1.860132e-07,1.860136e-07,1.860139e-07,1.860143e-07,1.860147e-07,1.860151e-07,1.860155e-07,1.860159e-07,1.860163e-07,1.860166e-07,1.860170e-07,1.860174e-07,1.860178e-07,1.860182e-07,1.860186e-07,1.860190e-07,1.860193e-07,1.860197e-07,1.860201e-07,1.860205e-07,1.860209e-07,1.860213e-07,1.860217e-07,1.860220e-07,1.860224e-07,1.860228e-07,1.860232e-07,1.860236e-07,1.860240e-07,1.860244e-07,1.860247e-07,1.860251e-07,1.860255e-07,1.860259e-07,1.860263e-07,1.860267e-07,1.860271e-07,1.860274e-07,1.860278e-07,1.860282e-07,1.860286e-07,1.860290e-07,1.860294e-07,1.860298e-07,1.860301e-07,1.860305e-07,1.860309e-07,1.860313e-07,1.860317e-07,1.860321e-07,1.860325e-07,1.860328e-07,1.860332e-07,1.860336e-07,1.860340e-07,1.860344e-07,1.860348e-07,1.860352e-07,1.860355e-07,1.860359e-07,1.860363e-07,1.860367e-07,1.860371e-07,1.860375e-07,1.860379e-07,1.860382e-07,1.860386e-07,1.860390e-07,1.860394e-07,1.860398e-07,1.860402e-07,1.860406e-07,1.860409e-07,1.860413e-07,1.860417e-07,1.860421e-07,1.860425e-07,1.860429e-07,1.860432e-07,1.860436e-07,1.860440e-07,1.860444e-07,1.860448e-07,1.860452e-07,1.860456e-07,1.860459e-07,1.860463e-07,1.860467e-07,1.860471e-07,1.860475e-07,1.860479e-07,1.860483e-07,1.860486e-07,1.860490e-07,1.860494e-07,1.860498e-07,1.860502e-07,1.860506e-07,1.860509e-07,1.860513e-07,1.860517e-07,1.860521e-07,1.860525e-07,1.860529e-07,1.860533e-07,1.860536e-07,1.860540e-07,1.860544e-07,1.860548e-07,1.860552e-07,1.860556e-07,1.860559e-07,1.860563e-07,1.860567e-07,1.860571e-07,1.860575e-07,1.860579e-07,1.860583e-07,1.860586e-07,1.860590e-07,1.860594e-07,1.860598e-07,1.860602e-07,1.860606e-07,1.860609e-07,1.860613e-07,1.860617e-07,1.860621e-07,1.860625e-07,1.860629e-07,1.860633e-07,1.860636e-07,1.860640e-07,1.860644e-07,1.860648e-07,1.860652e-07,1.860656e-07,1.860659e-07,1.860663e-07,1.860667e-07,1.860671e-07,1.860675e-07,1.860679e-07,1.860683e-07,1.860686e-07,1.860690e-07,1.860694e-07,1.860698e-07,1.860702e-07,1.860706e-07,1.860709e-07,1.860713e-07,1.860717e-07,1.860721e-07,1.860725e-07,1.860729e-07,1.860732e-07,1.860736e-07,1.860740e-07,1.860744e-07,1.860748e-07,1.860752e-07,1.860756e-07,1.860759e-07,1.860763e-07,1.860767e-07,1.860771e-07,1.860775e-07,1.860779e-07,1.860782e-07,1.860786e-07,1.860790e-07,1.860794e-07,1.860798e-07,1.860802e-07,1.860805e-07,1.860809e-07,1.860813e-07,1.860817e-07,1.860821e-07,1.860825e-07,1.860828e-07,1.860832e-07,1.860836e-07,1.860840e-07,1.860844e-07,1.860848e-07,1.860851e-07,1.860855e-07,1.860859e-07,1.860863e-07,1.860867e-07,1.860871e-07,1.860875e-07,1.860878e-07,1.860882e-07,1.860886e-07,1.860890e-07,1.860894e-07,1.860898e-07,1.860901e-07,1.860905e-07,1.860909e-07,1.860913e-07,1.860917e-07,1.860921e-07,1.860924e-07,1.860928e-07,1.860932e-07,1.860936e-07,1.860940e-07,1.860944e-07,1.860947e-07,1.860951e-07,1.860955e-07,1.860959e-07,1.860963e-07,1.860967e-07,1.860970e-07,1.860974e-07,1.860978e-07,1.860982e-07,1.860986e-07,1.860990e-07,1.860993e-07,1.860997e-07,1.861001e-07,1.861005e-07,1.861009e-07,1.861013e-07,1.861016e-07,1.861020e-07,1.861024e-07,1.861028e-07,1.861032e-07,1.861036e-07,1.861039e-07,1.861043e-07,1.861047e-07,1.861051e-07,1.861055e-07,1.861059e-07,1.861062e-07,1.861066e-07,1.861070e-07,1.861074e-07,1.861078e-07,1.861081e-07,1.861085e-07,1.861089e-07,1.861093e-07,1.861097e-07,1.861101e-07,1.861104e-07,1.861108e-07,1.861112e-07,1.861116e-07,1.861120e-07,1.861124e-07,1.861127e-07,1.861131e-07,1.861135e-07,1.861139e-07,1.861143e-07,1.861147e-07,1.861150e-07,1.861154e-07,1.861158e-07,1.861162e-07,1.861166e-07,1.861170e-07,1.861173e-07,1.861177e-07,1.861181e-07,1.861185e-07,1.861189e-07,1.861193e-07,1.861196e-07,1.861200e-07,1.861204e-07,1.861208e-07,1.861212e-07,1.861215e-07,1.861219e-07,1.861223e-07,1.861227e-07,1.861231e-07,1.861235e-07,1.861238e-07,1.861242e-07,1.861246e-07,1.861250e-07,1.861254e-07,1.861258e-07,1.861261e-07,1.861265e-07,1.861269e-07,1.861273e-07,1.861277e-07,1.861280e-07,1.861284e-07,1.861288e-07,1.861292e-07,1.861296e-07,1.861300e-07,1.861303e-07,1.861307e-07,1.861311e-07,1.861315e-07,1.861319e-07,1.861323e-07,1.861326e-07,1.861330e-07,1.861334e-07,1.861338e-07,1.861342e-07,1.861345e-07,1.861349e-07,1.861353e-07,1.861357e-07,1.861361e-07,1.861365e-07,1.861368e-07,1.861372e-07,1.861376e-07,1.861380e-07,1.861384e-07,1.861387e-07,1.861391e-07,1.861395e-07,1.861399e-07,1.861403e-07,1.861407e-07,1.861410e-07,1.861414e-07,1.861418e-07,1.861422e-07,1.861426e-07,1.861429e-07,1.861433e-07,1.861437e-07,1.861441e-07,1.861445e-07,1.861449e-07,1.861452e-07,1.861456e-07,1.861460e-07,1.861464e-07,1.861468e-07,1.861471e-07,1.861475e-07,1.861479e-07,1.861483e-07,1.861487e-07,1.861491e-07,1.861494e-07,1.861498e-07,1.861502e-07,1.861506e-07,1.861510e-07,1.861513e-07,1.861517e-07,1.861521e-07,1.861525e-07,1.861529e-07,1.861533e-07,1.861536e-07,1.861540e-07,1.861544e-07,1.861548e-07,1.861552e-07,1.861555e-07,1.861559e-07,1.861563e-07,1.861567e-07,1.861571e-07,1.861574e-07,1.861578e-07,1.861582e-07,1.861586e-07,1.861590e-07,1.861594e-07,1.861597e-07,1.861601e-07,1.861605e-07,1.861609e-07,1.861613e-07,1.861616e-07,1.861620e-07,1.861624e-07,1.861628e-07,1.861632e-07,1.861635e-07,1.861639e-07,1.861643e-07,1.861647e-07,1.861651e-07,1.861655e-07,1.861658e-07,1.861662e-07,1.861666e-07,1.861670e-07,1.861674e-07,1.861677e-07,1.861681e-07,1.861685e-07,1.861689e-07,1.861693e-07,1.861696e-07,1.861700e-07,1.861704e-07,1.861708e-07,1.861712e-07,1.861716e-07,1.861719e-07,1.861723e-07,1.861727e-07,1.861731e-07,1.861735e-07,1.861738e-07,1.861742e-07,1.861746e-07,1.861750e-07,1.861754e-07,1.861757e-07,1.861761e-07,1.861765e-07,1.861769e-07,1.861773e-07,1.861776e-07,1.861780e-07,1.861784e-07,1.861788e-07,1.861792e-07,1.861795e-07,1.861799e-07,1.861803e-07,1.861807e-07,1.861811e-07,1.861814e-07,1.861818e-07,1.861822e-07,1.861826e-07,1.861830e-07,1.861834e-07,1.861837e-07,1.861841e-07,1.861845e-07,1.861849e-07,1.861853e-07,1.861856e-07,1.861860e-07,1.861864e-07,1.861868e-07,1.861872e-07,1.861875e-07,1.861879e-07,1.861883e-07,1.861887e-07,1.861891e-07,1.861894e-07,1.861898e-07,1.861902e-07,1.861906e-07,1.861910e-07,1.861913e-07,1.861917e-07,1.861921e-07,1.861925e-07,1.861929e-07,1.861932e-07,1.861936e-07,1.861940e-07,1.861944e-07,1.861948e-07,1.861951e-07,1.861955e-07,1.861959e-07,1.861963e-07,1.861967e-07,1.861970e-07,1.861974e-07,1.861978e-07,1.861982e-07,1.861986e-07,1.861989e-07,1.861993e-07,1.861997e-07,1.862001e-07,1.862005e-07,1.862008e-07,1.862012e-07,1.862016e-07,1.862020e-07,1.862024e-07,1.862027e-07,1.862031e-07,1.862035e-07,1.862039e-07,1.862043e-07,1.862046e-07,1.862050e-07,1.862054e-07,1.862058e-07,1.862062e-07,1.862065e-07,1.862069e-07,1.862073e-07,1.862077e-07,1.862081e-07,1.862084e-07,1.862088e-07,1.862092e-07,1.862096e-07,1.862100e-07,1.862103e-07,1.862107e-07,1.862111e-07,1.862115e-07,1.862119e-07,1.862122e-07,1.862126e-07,1.862130e-07,1.862134e-07,1.862138e-07,1.862141e-07,1.862145e-07,1.862149e-07,1.862153e-07,1.862157e-07,1.862160e-07,1.862164e-07,1.862168e-07,1.862172e-07,1.862175e-07,1.862179e-07,1.862183e-07,1.862187e-07,1.862191e-07,1.862194e-07,1.862198e-07,1.862202e-07,1.862206e-07,1.862210e-07,1.862213e-07,1.862217e-07,1.862221e-07,1.862225e-07,1.862229e-07,1.862232e-07,1.862236e-07,1.862240e-07,1.862244e-07,1.862248e-07,1.862251e-07,1.862255e-07,1.862259e-07,1.862263e-07,1.862267e-07,1.862270e-07,1.862274e-07,1.862278e-07,1.862282e-07,1.862285e-07,1.862289e-07,1.862293e-07,1.862297e-07,1.862301e-07,1.862304e-07,1.862308e-07,1.862312e-07,1.862316e-07,1.862320e-07,1.862323e-07,1.862327e-07,1.862331e-07,1.862335e-07,1.862339e-07,1.862342e-07,1.862346e-07,1.862350e-07,1.862354e-07,1.862357e-07,1.862361e-07,1.862365e-07,1.862369e-07,1.862373e-07,1.862376e-07,1.862380e-07,1.862384e-07,1.862388e-07,1.862392e-07,1.862395e-07,1.862399e-07,1.862403e-07,1.862407e-07,1.862410e-07,1.862414e-07,1.862418e-07,1.862422e-07,1.862426e-07,1.862429e-07,1.862433e-07,1.862437e-07,1.862441e-07,1.862445e-07,1.862448e-07,1.862452e-07,1.862456e-07,1.862460e-07,1.862463e-07,1.862467e-07,1.862471e-07,1.862475e-07,1.862479e-07,1.862482e-07,1.862486e-07,1.862490e-07,1.862494e-07,1.862498e-07,1.862501e-07,1.862505e-07,1.862509e-07,1.862513e-07,1.862516e-07,1.862520e-07,1.862524e-07,1.862528e-07,1.862532e-07,1.862535e-07,1.862539e-07,1.862543e-07,1.862547e-07,1.862550e-07,1.862554e-07,1.862558e-07,1.862562e-07,1.862566e-07,1.862569e-07,1.862573e-07,1.862577e-07,1.862581e-07,1.862585e-07,1.862588e-07,1.862592e-07,1.862596e-07,1.862600e-07,1.862603e-07,1.862607e-07,1.862611e-07,1.862615e-07,1.862619e-07,1.862622e-07,1.862626e-07,1.862630e-07,1.862634e-07,1.862637e-07,1.862641e-07,1.862645e-07,1.862649e-07,1.862653e-07,1.862656e-07,1.862660e-07,1.862664e-07,1.862668e-07,1.862671e-07,1.862675e-07,1.862679e-07,1.862683e-07,1.862687e-07,1.862690e-07,1.862694e-07,1.862698e-07,1.862702e-07,1.862705e-07,1.862709e-07,1.862713e-07,1.862717e-07,1.862721e-07,1.862724e-07,1.862728e-07,1.862732e-07,1.862736e-07,1.862739e-07,1.862743e-07,1.862747e-07,1.862751e-07,1.862755e-07,1.862758e-07,1.862762e-07,1.862766e-07,1.862770e-07,1.862773e-07,1.862777e-07,1.862781e-07,1.862785e-07,1.862789e-07,1.862792e-07,1.862796e-07,1.862800e-07,1.862804e-07,1.862807e-07,1.862811e-07,1.862815e-07,1.862819e-07,1.862822e-07,1.862826e-07,1.862830e-07,1.862834e-07,1.862838e-07,1.862841e-07,1.862845e-07,1.862849e-07,1.862853e-07,1.862856e-07,1.862860e-07,1.862864e-07,1.862868e-07,1.862872e-07,1.862875e-07,1.862879e-07,1.862883e-07,1.862887e-07,1.862890e-07,1.862894e-07,1.862898e-07,1.862902e-07,1.862905e-07,1.862909e-07,1.862913e-07,1.862917e-07,1.862921e-07,1.862924e-07,1.862928e-07,1.862932e-07,1.862936e-07,1.862939e-07,1.862943e-07,1.862947e-07,1.862951e-07,1.862954e-07,1.862958e-07,1.862962e-07,1.862966e-07,1.862970e-07,1.862973e-07,1.862977e-07,1.862981e-07,1.862985e-07,1.862988e-07,1.862992e-07,1.862996e-07,1.863000e-07,1.863003e-07,1.863007e-07,1.863011e-07,1.863015e-07,1.863019e-07,1.863022e-07,1.863026e-07,1.863030e-07,1.863034e-07,1.863037e-07,1.863041e-07,1.863045e-07,1.863049e-07,1.863052e-07,1.863056e-07,1.863060e-07,1.863064e-07,1.863067e-07,1.863071e-07,1.863075e-07,1.863079e-07,1.863083e-07,1.863086e-07,1.863090e-07,1.863094e-07,1.863098e-07,1.863101e-07,1.863105e-07,1.863109e-07,1.863113e-07,1.863116e-07,1.863120e-07,1.863124e-07,1.863128e-07,1.863131e-07,1.863135e-07,1.863139e-07,1.863143e-07,1.863147e-07,1.863150e-07,1.863154e-07,1.863158e-07,1.863162e-07,1.863165e-07,1.863169e-07,1.863173e-07,1.863177e-07,1.863180e-07,1.863184e-07,1.863188e-07,1.863192e-07,1.863195e-07,1.863199e-07,1.863203e-07,1.863207e-07,1.863210e-07,1.863214e-07,1.863218e-07,1.863222e-07,1.863225e-07,1.863229e-07,1.863233e-07,1.863237e-07,1.863241e-07,1.863244e-07,1.863248e-07,1.863252e-07,1.863256e-07,1.863259e-07,1.863263e-07,1.863267e-07,1.863271e-07,1.863274e-07,1.863278e-07,1.863282e-07,1.863286e-07,1.863289e-07,1.863293e-07,1.863297e-07,1.863301e-07,1.863304e-07,1.863308e-07,1.863312e-07,1.863316e-07,1.863319e-07,1.863323e-07,1.863327e-07,1.863331e-07,1.863334e-07,1.863338e-07,1.863342e-07,1.863346e-07,1.863350e-07,1.863353e-07,1.863357e-07,1.863361e-07,1.863365e-07,1.863368e-07,1.863372e-07,1.863376e-07,1.863380e-07,1.863383e-07,1.863387e-07,1.863391e-07,1.863395e-07,1.863398e-07,1.863402e-07,1.863406e-07,1.863410e-07,1.863413e-07,1.863417e-07,1.863421e-07,1.863425e-07,1.863428e-07,1.863432e-07,1.863436e-07,1.863440e-07,1.863443e-07,1.863447e-07,1.863451e-07,1.863455e-07,1.863458e-07,1.863462e-07,1.863466e-07,1.863470e-07,1.863473e-07,1.863477e-07,1.863481e-07,1.863485e-07,1.863488e-07,1.863492e-07,1.863496e-07,1.863500e-07,1.863503e-07,1.863507e-07,1.863511e-07,1.863515e-07,1.863518e-07,1.863522e-07,1.863526e-07,1.863530e-07,1.863533e-07,1.863537e-07,1.863541e-07,1.863545e-07,1.863548e-07,1.863552e-07,1.863556e-07,1.863560e-07,1.863563e-07,1.863567e-07,1.863571e-07,1.863575e-07,1.863578e-07,1.863582e-07,1.863586e-07,1.863590e-07,1.863593e-07,1.863597e-07,1.863601e-07,1.863605e-07,1.863608e-07,1.863612e-07,1.863616e-07,1.863620e-07,1.863623e-07,1.863627e-07,1.863631e-07,1.863635e-07,1.863638e-07,1.863642e-07,1.863646e-07,1.863650e-07,1.863653e-07,1.863657e-07,1.863661e-07,1.863665e-07,1.863668e-07,1.863672e-07,1.863676e-07,1.863680e-07,1.863683e-07,1.863687e-07,1.863691e-07,1.863695e-07,1.863698e-07,1.863702e-07,1.863706e-07,1.863710e-07,1.863713e-07,1.863717e-07,1.863721e-07,1.863725e-07,1.863728e-07,1.863732e-07,1.863736e-07,1.863739e-07,1.863743e-07,1.863747e-07,1.863751e-07,1.863754e-07,1.863758e-07,1.863762e-07,1.863766e-07,1.863769e-07,1.863773e-07,1.863777e-07,1.863781e-07,1.863784e-07,1.863788e-07,1.863792e-07,1.863796e-07,1.863799e-07,1.863803e-07,1.863807e-07,1.863811e-07,1.863814e-07,1.863818e-07,1.863822e-07,1.863826e-07,1.863829e-07,1.863833e-07,1.863837e-07,1.863841e-07,1.863844e-07,1.863848e-07,1.863852e-07,1.863855e-07,1.863859e-07,1.863863e-07,1.863867e-07,1.863870e-07,1.863874e-07,1.863878e-07,1.863882e-07,1.863885e-07,1.863889e-07,1.863893e-07,1.863897e-07,1.863900e-07,1.863904e-07,1.863908e-07,1.863912e-07,1.863915e-07,1.863919e-07,1.863923e-07,1.863927e-07,1.863930e-07,1.863934e-07,1.863938e-07,1.863941e-07,1.863945e-07,1.863949e-07,1.863953e-07,1.863956e-07,1.863960e-07,1.863964e-07,1.863968e-07,1.863971e-07,1.863975e-07,1.863979e-07,1.863983e-07,1.863986e-07,1.863990e-07,1.863994e-07,1.863998e-07,1.864001e-07,1.864005e-07,1.864009e-07,1.864012e-07,1.864016e-07,1.864020e-07,1.864024e-07,1.864027e-07,1.864031e-07,1.864035e-07,1.864039e-07,1.864042e-07,1.864046e-07,1.864050e-07,1.864054e-07,1.864057e-07,1.864061e-07,1.864065e-07,1.864068e-07,1.864072e-07,1.864076e-07,1.864080e-07,1.864083e-07,1.864087e-07,1.864091e-07,1.864095e-07,1.864098e-07,1.864102e-07,1.864106e-07,1.864110e-07,1.864113e-07,1.864117e-07,1.864121e-07,1.864124e-07,1.864128e-07,1.864132e-07,1.864136e-07,1.864139e-07,1.864143e-07,1.864147e-07,1.864151e-07,1.864154e-07,1.864158e-07,1.864162e-07,1.864165e-07,1.864169e-07,1.864173e-07,1.864177e-07,1.864180e-07,1.864184e-07,1.864188e-07,1.864192e-07,1.864195e-07,1.864199e-07,1.864203e-07,1.864207e-07,1.864210e-07,1.864214e-07,1.864218e-07,1.864221e-07,1.864225e-07,1.864229e-07,1.864233e-07,1.864236e-07,1.864240e-07,1.864244e-07,1.864248e-07,1.864251e-07,1.864255e-07,1.864259e-07,1.864262e-07,1.864266e-07,1.864270e-07,1.864274e-07,1.864277e-07,1.864281e-07,1.864285e-07,1.864289e-07,1.864292e-07,1.864296e-07,1.864300e-07,1.864303e-07,1.864307e-07,1.864311e-07,1.864315e-07,1.864318e-07,1.864322e-07,1.864326e-07,1.864329e-07,1.864333e-07,1.864337e-07,1.864341e-07,1.864344e-07,1.864348e-07,1.864352e-07,1.864356e-07,1.864359e-07,1.864363e-07,1.864367e-07,1.864370e-07,1.864374e-07,1.864378e-07,1.864382e-07,1.864385e-07,1.864389e-07,1.864393e-07,1.864397e-07,1.864400e-07,1.864404e-07,1.864408e-07,1.864411e-07,1.864415e-07,1.864419e-07,1.864423e-07,1.864426e-07,1.864430e-07,1.864434e-07,1.864437e-07,1.864441e-07,1.864445e-07,1.864449e-07,1.864452e-07,1.864456e-07,1.864460e-07,1.864463e-07,1.864467e-07,1.864471e-07,1.864475e-07,1.864478e-07,1.864482e-07,1.864486e-07,1.864490e-07,1.864493e-07,1.864497e-07,1.864501e-07,1.864504e-07,1.864508e-07,1.864512e-07,1.864516e-07,1.864519e-07,1.864523e-07,1.864527e-07,1.864530e-07,1.864534e-07,1.864538e-07,1.864542e-07,1.864545e-07,1.864549e-07,1.864553e-07,1.864556e-07,1.864560e-07,1.864564e-07,1.864568e-07,1.864571e-07,1.864575e-07,1.864579e-07,1.864582e-07,1.864586e-07,1.864590e-07,1.864594e-07,1.864597e-07,1.864601e-07,1.864605e-07,1.864608e-07,1.864612e-07,1.864616e-07,1.864620e-07,1.864623e-07,1.864627e-07,1.864631e-07,1.864635e-07,1.864638e-07,1.864642e-07,1.864646e-07,1.864649e-07,1.864653e-07,1.864657e-07,1.864661e-07,1.864664e-07,1.864668e-07,1.864672e-07,1.864675e-07,1.864679e-07,1.864683e-07,1.864687e-07,1.864690e-07,1.864694e-07,1.864698e-07,1.864701e-07,1.864705e-07,1.864709e-07,1.864712e-07,1.864716e-07,1.864720e-07,1.864724e-07,1.864727e-07,1.864731e-07,1.864735e-07,1.864738e-07,1.864742e-07,1.864746e-07,1.864750e-07,1.864753e-07,1.864757e-07,1.864761e-07,1.864764e-07,1.864768e-07,1.864772e-07,1.864776e-07,1.864779e-07,1.864783e-07,1.864787e-07,1.864790e-07,1.864794e-07,1.864798e-07,1.864802e-07,1.864805e-07,1.864809e-07,1.864813e-07,1.864816e-07,1.864820e-07,1.864824e-07,1.864828e-07,1.864831e-07,1.864835e-07,1.864839e-07,1.864842e-07,1.864846e-07,1.864850e-07,1.864853e-07,1.864857e-07,1.864861e-07,1.864865e-07,1.864868e-07,1.864872e-07,1.864876e-07,1.864879e-07,1.864883e-07,1.864887e-07,1.864891e-07,1.864894e-07,1.864898e-07,1.864902e-07,1.864905e-07,1.864909e-07,1.864913e-07,1.864917e-07,1.864920e-07,1.864924e-07,1.864928e-07,1.864931e-07,1.864935e-07,1.864939e-07,1.864942e-07,1.864946e-07,1.864950e-07,1.864954e-07,1.864957e-07,1.864961e-07,1.864965e-07,1.864968e-07,1.864972e-07,1.864976e-07,1.864979e-07,1.864983e-07,1.864987e-07,1.864991e-07,1.864994e-07,1.864998e-07,1.865002e-07,1.865005e-07,1.865009e-07,1.865013e-07,1.865017e-07,1.865020e-07,1.865024e-07,1.865028e-07,1.865031e-07,1.865035e-07,1.865039e-07,1.865042e-07,1.865046e-07,1.865050e-07,1.865054e-07,1.865057e-07,1.865061e-07,1.865065e-07,1.865068e-07,1.865072e-07,1.865076e-07,1.865079e-07,1.865083e-07,1.865087e-07,1.865091e-07,1.865094e-07,1.865098e-07,1.865102e-07,1.865105e-07,1.865109e-07,1.865113e-07,1.865116e-07,1.865120e-07,1.865124e-07,1.865128e-07,1.865131e-07,1.865135e-07,1.865139e-07,1.865142e-07,1.865146e-07,1.865150e-07,1.865153e-07,1.865157e-07,1.865161e-07,1.865165e-07,1.865168e-07,1.865172e-07,1.865176e-07,1.865179e-07,1.865183e-07,1.865187e-07,1.865190e-07,1.865194e-07,1.865198e-07,1.865202e-07,1.865205e-07,1.865209e-07,1.865213e-07,1.865216e-07,1.865220e-07,1.865224e-07,1.865227e-07,1.865231e-07,1.865235e-07,1.865238e-07,1.865242e-07,1.865246e-07,1.865250e-07,1.865253e-07,1.865257e-07,1.865261e-07,1.865264e-07,1.865268e-07,1.865272e-07,1.865275e-07,1.865279e-07,1.865283e-07,1.865287e-07,1.865290e-07,1.865294e-07,1.865298e-07,1.865301e-07,1.865305e-07,1.865309e-07,1.865312e-07,1.865316e-07,1.865320e-07,1.865323e-07,1.865327e-07,1.865331e-07,1.865335e-07,1.865338e-07,1.865342e-07,1.865346e-07,1.865349e-07,1.865353e-07,1.865357e-07,1.865360e-07,1.865364e-07,1.865368e-07,1.865371e-07,1.865375e-07,1.865379e-07,1.865383e-07,1.865386e-07,1.865390e-07,1.865394e-07,1.865397e-07,1.865401e-07,1.865405e-07,1.865408e-07,1.865412e-07,1.865416e-07,1.865419e-07,1.865423e-07,1.865427e-07,1.865431e-07,1.865434e-07,1.865438e-07,1.865442e-07,1.865445e-07,1.865449e-07,1.865453e-07,1.865456e-07,1.865460e-07,1.865464e-07,1.865467e-07,1.865471e-07,1.865475e-07,1.865478e-07,1.865482e-07,1.865486e-07,1.865490e-07,1.865493e-07,1.865497e-07,1.865501e-07,1.865504e-07,1.865508e-07,1.865512e-07,1.865515e-07,1.865519e-07,1.865523e-07,1.865526e-07,1.865530e-07,1.865534e-07,1.865537e-07,1.865541e-07,1.865545e-07,1.865549e-07,1.865552e-07,1.865556e-07,1.865560e-07,1.865563e-07,1.865567e-07,1.865571e-07,1.865574e-07,1.865578e-07,1.865582e-07,1.865585e-07,1.865589e-07,1.865593e-07,1.865596e-07,1.865600e-07,1.865604e-07,1.865607e-07,1.865611e-07,1.865615e-07,1.865619e-07,1.865622e-07,1.865626e-07,1.865630e-07,1.865633e-07,1.865637e-07,1.865641e-07,1.865644e-07,1.865648e-07,1.865652e-07,1.865655e-07,1.865659e-07,1.865663e-07,1.865666e-07,1.865670e-07,1.865674e-07,1.865677e-07,1.865681e-07,1.865685e-07,1.865689e-07,1.865692e-07,1.865696e-07,1.865700e-07,1.865703e-07,1.865707e-07,1.865711e-07,1.865714e-07,1.865718e-07,1.865722e-07,1.865725e-07,1.865729e-07,1.865733e-07,1.865736e-07,1.865740e-07,1.865744e-07,1.865747e-07,1.865751e-07,1.865755e-07,1.865758e-07,1.865762e-07,1.865766e-07,1.865769e-07,1.865773e-07,1.865777e-07,1.865781e-07,1.865784e-07,1.865788e-07,1.865792e-07,1.865795e-07,1.865799e-07,1.865803e-07,1.865806e-07,1.865810e-07,1.865814e-07,1.865817e-07,1.865821e-07,1.865825e-07,1.865828e-07,1.865832e-07,1.865836e-07,1.865839e-07,1.865843e-07,1.865847e-07,1.865850e-07,1.865854e-07,1.865858e-07,1.865861e-07,1.865865e-07,1.865869e-07,1.865872e-07,1.865876e-07,1.865880e-07,1.865883e-07,1.865887e-07,1.865891e-07,1.865894e-07,1.865898e-07,1.865902e-07,1.865906e-07,1.865909e-07,1.865913e-07,1.865917e-07,1.865920e-07,1.865924e-07,1.865928e-07,1.865931e-07,1.865935e-07,1.865939e-07,1.865942e-07,1.865946e-07,1.865950e-07,1.865953e-07,1.865957e-07,1.865961e-07,1.865964e-07,1.865968e-07,1.865972e-07,1.865975e-07,1.865979e-07,1.865983e-07,1.865986e-07,1.865990e-07,1.865994e-07,1.865997e-07,1.866001e-07,1.866005e-07,1.866008e-07,1.866012e-07,1.866016e-07,1.866019e-07,1.866023e-07,1.866027e-07,1.866030e-07,1.866034e-07,1.866038e-07,1.866041e-07,1.866045e-07,1.866049e-07,1.866052e-07,1.866056e-07,1.866060e-07,1.866063e-07,1.866067e-07,1.866071e-07,1.866074e-07,1.866078e-07,1.866082e-07,1.866085e-07,1.866089e-07,1.866093e-07,1.866096e-07,1.866100e-07,1.866104e-07,1.866107e-07,1.866111e-07,1.866115e-07,1.866118e-07,1.866122e-07,1.866126e-07,1.866129e-07,1.866133e-07,1.866137e-07,1.866140e-07,1.866144e-07,1.866148e-07,1.866151e-07,1.866155e-07,1.866159e-07,1.866162e-07,1.866166e-07,1.866170e-07,1.866173e-07,1.866177e-07,1.866181e-07,1.866184e-07,1.866188e-07,1.866192e-07,1.866195e-07,1.866199e-07,1.866203e-07,1.866206e-07,1.866210e-07,1.866214e-07,1.866217e-07,1.866221e-07,1.866225e-07,1.866228e-07,1.866232e-07,1.866236e-07,1.866239e-07,1.866243e-07,1.866247e-07,1.866250e-07,1.866254e-07,1.866258e-07,1.866261e-07,1.866265e-07,1.866269e-07,1.866272e-07,1.866276e-07,1.866280e-07,1.866283e-07,1.866287e-07,1.866291e-07,1.866294e-07,1.866298e-07,1.866302e-07,1.866305e-07,1.866309e-07,1.866313e-07,1.866316e-07,1.866320e-07,1.866324e-07,1.866327e-07,1.866331e-07,1.866335e-07,1.866338e-07,1.866342e-07,1.866346e-07,1.866349e-07,1.866353e-07,1.866357e-07,1.866360e-07,1.866364e-07,1.866368e-07,1.866371e-07,1.866375e-07,1.866379e-07,1.866382e-07,1.866386e-07,1.866390e-07,1.866393e-07,1.866397e-07,1.866401e-07,1.866404e-07,1.866408e-07,1.866412e-07,1.866415e-07,1.866419e-07,1.866423e-07,1.866426e-07,1.866430e-07,1.866433e-07,1.866437e-07,1.866441e-07,1.866444e-07,1.866448e-07,1.866452e-07,1.866455e-07,1.866459e-07,1.866463e-07,1.866466e-07,1.866470e-07,1.866474e-07,1.866477e-07,1.866481e-07,1.866485e-07,1.866488e-07,1.866492e-07,1.866496e-07,1.866499e-07,1.866503e-07,1.866507e-07,1.866510e-07,1.866514e-07,1.866518e-07,1.866521e-07,1.866525e-07,1.866529e-07,1.866532e-07,1.866536e-07,1.866540e-07,1.866543e-07,1.866547e-07,1.866550e-07,1.866554e-07,1.866558e-07,1.866561e-07,1.866565e-07,1.866569e-07,1.866572e-07,1.866576e-07,1.866580e-07,1.866583e-07,1.866587e-07,1.866591e-07,1.866594e-07,1.866598e-07,1.866602e-07,1.866605e-07,1.866609e-07,1.866613e-07,1.866616e-07,1.866620e-07,1.866624e-07,1.866627e-07,1.866631e-07,1.866635e-07,1.866638e-07,1.866642e-07,1.866645e-07,1.866649e-07,1.866653e-07,1.866656e-07,1.866660e-07,1.866664e-07,1.866667e-07,1.866671e-07,1.866675e-07,1.866678e-07,1.866682e-07,1.866686e-07,1.866689e-07,1.866693e-07,1.866697e-07,1.866700e-07,1.866704e-07,1.866708e-07,1.866711e-07,1.866715e-07,1.866718e-07,1.866722e-07,1.866726e-07,1.866729e-07,1.866733e-07,1.866737e-07,1.866740e-07,1.866744e-07,1.866748e-07,1.866751e-07,1.866755e-07,1.866759e-07,1.866762e-07,1.866766e-07,1.866770e-07,1.866773e-07,1.866777e-07,1.866781e-07,1.866784e-07,1.866788e-07,1.866791e-07,1.866795e-07,1.866799e-07,1.866802e-07,1.866806e-07,1.866810e-07,1.866813e-07,1.866817e-07,1.866821e-07,1.866824e-07,1.866828e-07,1.866832e-07,1.866835e-07,1.866839e-07,1.866842e-07,1.866846e-07,1.866850e-07,1.866853e-07,1.866857e-07,1.866861e-07,1.866864e-07,1.866868e-07,1.866872e-07,1.866875e-07,1.866879e-07,1.866883e-07,1.866886e-07,1.866890e-07,1.866894e-07,1.866897e-07,1.866901e-07,1.866904e-07,1.866908e-07,1.866912e-07,1.866915e-07,1.866919e-07,1.866923e-07,1.866926e-07,1.866930e-07,1.866934e-07,1.866937e-07,1.866941e-07,1.866945e-07,1.866948e-07,1.866952e-07,1.866955e-07,1.866959e-07,1.866963e-07,1.866966e-07,1.866970e-07,1.866974e-07,1.866977e-07,1.866981e-07,1.866985e-07,1.866988e-07,1.866992e-07,1.866995e-07,1.866999e-07,1.867003e-07,1.867006e-07,1.867010e-07,1.867014e-07,1.867017e-07,1.867021e-07,1.867025e-07,1.867028e-07,1.867032e-07,1.867036e-07,1.867039e-07,1.867043e-07,1.867046e-07,1.867050e-07,1.867054e-07,1.867057e-07,1.867061e-07,1.867065e-07,1.867068e-07,1.867072e-07,1.867076e-07,1.867079e-07,1.867083e-07,1.867086e-07,1.867090e-07,1.867094e-07,1.867097e-07,1.867101e-07,1.867105e-07,1.867108e-07,1.867112e-07,1.867116e-07,1.867119e-07,1.867123e-07,1.867126e-07,1.867130e-07,1.867134e-07,1.867137e-07,1.867141e-07,1.867145e-07,1.867148e-07,1.867152e-07,1.867156e-07,1.867159e-07,1.867163e-07,1.867166e-07,1.867170e-07,1.867174e-07,1.867177e-07,1.867181e-07,1.867185e-07,1.867188e-07,1.867192e-07,1.867196e-07,1.867199e-07,1.867203e-07,1.867206e-07,1.867210e-07,1.867214e-07,1.867217e-07,1.867221e-07,1.867225e-07,1.867228e-07,1.867232e-07,1.867236e-07,1.867239e-07,1.867243e-07,1.867246e-07,1.867250e-07,1.867254e-07,1.867257e-07,1.867261e-07,1.867265e-07,1.867268e-07,1.867272e-07,1.867275e-07,1.867279e-07,1.867283e-07,1.867286e-07,1.867290e-07,1.867294e-07,1.867297e-07,1.867301e-07,1.867305e-07,1.867308e-07,1.867312e-07,1.867315e-07,1.867319e-07,1.867323e-07,1.867326e-07,1.867330e-07,1.867334e-07,1.867337e-07,1.867341e-07,1.867344e-07,1.867348e-07,1.867352e-07,1.867355e-07,1.867359e-07,1.867363e-07,1.867366e-07,1.867370e-07,1.867374e-07,1.867377e-07,1.867381e-07,1.867384e-07,1.867388e-07,1.867392e-07,1.867395e-07,1.867399e-07,1.867403e-07,1.867406e-07,1.867410e-07,1.867413e-07,1.867417e-07,1.867421e-07,1.867424e-07,1.867428e-07,1.867432e-07,1.867435e-07,1.867439e-07,1.867442e-07,1.867446e-07,1.867450e-07,1.867453e-07,1.867457e-07,1.867461e-07,1.867464e-07,1.867468e-07,1.867471e-07,1.867475e-07,1.867479e-07,1.867482e-07,1.867486e-07,1.867490e-07,1.867493e-07,1.867497e-07,1.867500e-07,1.867504e-07,1.867508e-07,1.867511e-07,1.867515e-07,1.867519e-07,1.867522e-07,1.867526e-07,1.867529e-07,1.867533e-07,1.867537e-07,1.867540e-07,1.867544e-07,1.867548e-07,1.867551e-07,1.867555e-07,1.867558e-07,1.867562e-07,1.867566e-07,1.867569e-07,1.867573e-07,1.867577e-07,1.867580e-07,1.867584e-07,1.867587e-07,1.867591e-07,1.867595e-07,1.867598e-07,1.867602e-07,1.867606e-07,1.867609e-07,1.867613e-07,1.867616e-07,1.867620e-07,1.867624e-07,1.867627e-07,1.867631e-07,1.867635e-07,1.867638e-07,1.867642e-07,1.867645e-07,1.867649e-07,1.867653e-07,1.867656e-07,1.867660e-07,1.867663e-07,1.867667e-07,1.867671e-07,1.867674e-07,1.867678e-07,1.867682e-07,1.867685e-07,1.867689e-07,1.867692e-07,1.867696e-07,1.867700e-07,1.867703e-07,1.867707e-07,1.867711e-07,1.867714e-07,1.867718e-07,1.867721e-07,1.867725e-07,1.867729e-07,1.867732e-07,1.867736e-07,1.867739e-07,1.867743e-07,1.867747e-07,1.867750e-07,1.867754e-07,1.867758e-07,1.867761e-07,1.867765e-07,1.867768e-07,1.867772e-07,1.867776e-07,1.867779e-07,1.867783e-07,1.867786e-07,1.867790e-07,1.867794e-07,1.867797e-07,1.867801e-07,1.867805e-07,1.867808e-07,1.867812e-07,1.867815e-07,1.867819e-07,1.867823e-07,1.867826e-07,1.867830e-07,1.867833e-07,1.867837e-07,1.867841e-07,1.867844e-07,1.867848e-07,1.867852e-07,1.867855e-07,1.867859e-07,1.867862e-07,1.867866e-07,1.867870e-07,1.867873e-07,1.867877e-07,1.867880e-07,1.867884e-07,1.867888e-07,1.867891e-07,1.867895e-07,1.867899e-07,1.867902e-07,1.867906e-07,1.867909e-07,1.867913e-07,1.867917e-07,1.867920e-07,1.867924e-07,1.867927e-07,1.867931e-07,1.867935e-07,1.867938e-07,1.867942e-07,1.867945e-07,1.867949e-07,1.867953e-07,1.867956e-07,1.867960e-07,1.867964e-07,1.867967e-07,1.867971e-07,1.867974e-07,1.867978e-07,1.867982e-07,1.867985e-07,1.867989e-07,1.867992e-07,1.867996e-07,1.868000e-07,1.868003e-07,1.868007e-07,1.868010e-07,1.868014e-07,1.868018e-07,1.868021e-07,1.868025e-07,1.868029e-07,1.868032e-07,1.868036e-07,1.868039e-07,1.868043e-07,1.868047e-07,1.868050e-07,1.868054e-07,1.868057e-07,1.868061e-07,1.868065e-07,1.868068e-07,1.868072e-07,1.868075e-07,1.868079e-07,1.868083e-07,1.868086e-07,1.868090e-07,1.868093e-07,1.868097e-07,1.868101e-07,1.868104e-07,1.868108e-07,1.868111e-07,1.868115e-07,1.868119e-07,1.868122e-07,1.868126e-07,1.868129e-07,1.868133e-07,1.868137e-07,1.868140e-07,1.868144e-07,1.868148e-07,1.868151e-07,1.868155e-07,1.868158e-07,1.868162e-07,1.868166e-07,1.868169e-07,1.868173e-07,1.868176e-07,1.868180e-07,1.868184e-07,1.868187e-07,1.868191e-07,1.868194e-07,1.868198e-07,1.868202e-07,1.868205e-07,1.868209e-07,1.868212e-07,1.868216e-07,1.868220e-07,1.868223e-07,1.868227e-07,1.868230e-07,1.868234e-07,1.868238e-07,1.868241e-07,1.868245e-07,1.868248e-07,1.868252e-07,1.868256e-07,1.868259e-07,1.868263e-07,1.868266e-07,1.868270e-07,1.868274e-07,1.868277e-07,1.868281e-07,1.868284e-07,1.868288e-07,1.868292e-07,1.868295e-07,1.868299e-07,1.868302e-07,1.868306e-07,1.868310e-07,1.868313e-07,1.868317e-07,1.868320e-07,1.868324e-07,1.868328e-07,1.868331e-07,1.868335e-07,1.868338e-07,1.868342e-07,1.868346e-07,1.868349e-07,1.868353e-07,1.868356e-07,1.868360e-07,1.868364e-07,1.868367e-07,1.868371e-07,1.868374e-07,1.868378e-07,1.868382e-07,1.868385e-07,1.868389e-07,1.868392e-07,1.868396e-07,1.868400e-07,1.868403e-07,1.868407e-07,1.868410e-07,1.868414e-07,1.868418e-07,1.868421e-07,1.868425e-07,1.868428e-07,1.868432e-07,1.868436e-07,1.868439e-07,1.868443e-07,1.868446e-07,1.868450e-07,1.868454e-07,1.868457e-07,1.868461e-07,1.868464e-07,1.868468e-07,1.868472e-07,1.868475e-07,1.868479e-07,1.868482e-07,1.868486e-07,1.868489e-07,1.868493e-07,1.868497e-07,1.868500e-07,1.868504e-07,1.868507e-07,1.868511e-07,1.868515e-07,1.868518e-07,1.868522e-07,1.868525e-07,1.868529e-07,1.868533e-07,1.868536e-07,1.868540e-07,1.868543e-07,1.868547e-07,1.868551e-07,1.868554e-07,1.868558e-07,1.868561e-07,1.868565e-07,1.868569e-07,1.868572e-07,1.868576e-07,1.868579e-07,1.868583e-07,1.868586e-07,1.868590e-07,1.868594e-07,1.868597e-07,1.868601e-07,1.868604e-07,1.868608e-07,1.868612e-07,1.868615e-07,1.868619e-07,1.868622e-07,1.868626e-07,1.868630e-07,1.868633e-07,1.868637e-07,1.868640e-07,1.868644e-07,1.868648e-07,1.868651e-07,1.868655e-07,1.868658e-07,1.868662e-07,1.868665e-07,1.868669e-07,1.868673e-07,1.868676e-07,1.868680e-07,1.868683e-07,1.868687e-07,1.868691e-07,1.868694e-07,1.868698e-07,1.868701e-07,1.868705e-07,1.868709e-07,1.868712e-07,1.868716e-07,1.868719e-07,1.868723e-07,1.868726e-07,1.868730e-07,1.868734e-07,1.868737e-07,1.868741e-07,1.868744e-07,1.868748e-07,1.868752e-07,1.868755e-07,1.868759e-07,1.868762e-07,1.868766e-07,1.868770e-07,1.868773e-07,1.868777e-07,1.868780e-07,1.868784e-07,1.868787e-07,1.868791e-07,1.868795e-07,1.868798e-07,1.868802e-07,1.868805e-07,1.868809e-07,1.868813e-07,1.868816e-07,1.868820e-07,1.868823e-07,1.868827e-07,1.868830e-07,1.868834e-07,1.868838e-07,1.868841e-07,1.868845e-07,1.868848e-07,1.868852e-07,1.868856e-07,1.868859e-07,1.868863e-07,1.868866e-07,1.868870e-07,1.868873e-07,1.868877e-07,1.868881e-07,1.868884e-07,1.868888e-07,1.868891e-07,1.868895e-07,1.868899e-07,1.868902e-07,1.868906e-07,1.868909e-07,1.868913e-07,1.868916e-07,1.868920e-07,1.868924e-07,1.868927e-07,1.868931e-07,1.868934e-07,1.868938e-07,1.868942e-07,1.868945e-07,1.868949e-07,1.868952e-07,1.868956e-07,1.868959e-07,1.868963e-07,1.868967e-07,1.868970e-07,1.868974e-07,1.868977e-07,1.868981e-07,1.868984e-07,1.868988e-07,1.868992e-07,1.868995e-07,1.868999e-07,1.869002e-07,1.869006e-07,1.869010e-07,1.869013e-07,1.869017e-07,1.869020e-07,1.869024e-07,1.869027e-07,1.869031e-07,1.869035e-07,1.869038e-07,1.869042e-07,1.869045e-07,1.869049e-07,1.869052e-07,1.869056e-07,1.869060e-07,1.869063e-07,1.869067e-07,1.869070e-07,1.869074e-07,1.869077e-07,1.869081e-07,1.869085e-07,1.869088e-07,1.869092e-07,1.869095e-07,1.869099e-07,1.869103e-07,1.869106e-07,1.869110e-07,1.869113e-07,1.869117e-07,1.869120e-07,1.869124e-07,1.869128e-07,1.869131e-07,1.869135e-07,1.869138e-07,1.869142e-07,1.869145e-07,1.869149e-07,1.869153e-07,1.869156e-07,1.869160e-07,1.869163e-07,1.869167e-07,1.869170e-07,1.869174e-07,1.869178e-07,1.869181e-07,1.869185e-07,1.869188e-07,1.869192e-07,1.869195e-07,1.869199e-07,1.869203e-07,1.869206e-07,1.869210e-07,1.869213e-07,1.869217e-07,1.869220e-07,1.869224e-07,1.869228e-07,1.869231e-07,1.869235e-07,1.869238e-07,1.869242e-07,1.869245e-07,1.869249e-07,1.869253e-07,1.869256e-07,1.869260e-07,1.869263e-07,1.869267e-07,1.869270e-07,1.869274e-07,1.869278e-07,1.869281e-07,1.869285e-07,1.869288e-07,1.869292e-07,1.869295e-07,1.869299e-07,1.869303e-07,1.869306e-07,1.869310e-07,1.869313e-07,1.869317e-07,1.869320e-07,1.869324e-07,1.869328e-07,1.869331e-07,1.869335e-07,1.869338e-07,1.869342e-07,1.869345e-07,1.869349e-07,1.869353e-07,1.869356e-07,1.869360e-07,1.869363e-07,1.869367e-07,1.869370e-07,1.869374e-07,1.869378e-07,1.869381e-07,1.869385e-07,1.869388e-07,1.869392e-07,1.869395e-07,1.869399e-07,1.869402e-07,1.869406e-07,1.869410e-07,1.869413e-07,1.869417e-07,1.869420e-07,1.869424e-07,1.869427e-07,1.869431e-07,1.869435e-07,1.869438e-07,1.869442e-07,1.869445e-07,1.869449e-07,1.869452e-07,1.869456e-07,1.869460e-07,1.869463e-07,1.869467e-07,1.869470e-07,1.869474e-07,1.869477e-07,1.869481e-07,1.869484e-07,1.869488e-07,1.869492e-07,1.869495e-07,1.869499e-07,1.869502e-07,1.869506e-07,1.869509e-07,1.869513e-07,1.869517e-07,1.869520e-07,1.869524e-07,1.869527e-07,1.869531e-07,1.869534e-07,1.869538e-07,1.869541e-07,1.869545e-07,1.869549e-07,1.869552e-07,1.869556e-07,1.869559e-07,1.869563e-07,1.869566e-07,1.869570e-07,1.869574e-07,1.869577e-07,1.869581e-07,1.869584e-07,1.869588e-07,1.869591e-07,1.869595e-07,1.869598e-07,1.869602e-07,1.869606e-07,1.869609e-07,1.869613e-07,1.869616e-07,1.869620e-07,1.869623e-07,1.869627e-07,1.869631e-07,1.869634e-07,1.869638e-07,1.869641e-07,1.869645e-07,1.869648e-07,1.869652e-07,1.869655e-07,1.869659e-07,1.869663e-07,1.869666e-07,1.869670e-07,1.869673e-07,1.869677e-07,1.869680e-07,1.869684e-07,1.869687e-07,1.869691e-07,1.869695e-07,1.869698e-07,1.869702e-07,1.869705e-07,1.869709e-07,1.869712e-07,1.869716e-07,1.869719e-07,1.869723e-07,1.869727e-07,1.869730e-07,1.869734e-07,1.869737e-07,1.869741e-07,1.869744e-07,1.869748e-07,1.869751e-07,1.869755e-07,1.869759e-07,1.869762e-07,1.869766e-07,1.869769e-07,1.869773e-07,1.869776e-07,1.869780e-07,1.869783e-07,1.869787e-07,1.869791e-07,1.869794e-07,1.869798e-07,1.869801e-07,1.869805e-07,1.869808e-07,1.869812e-07,1.869815e-07,1.869819e-07,1.869823e-07,1.869826e-07,1.869830e-07,1.869833e-07,1.869837e-07,1.869840e-07,1.869844e-07,1.869847e-07,1.869851e-07,1.869855e-07,1.869858e-07,1.869862e-07,1.869865e-07,1.869869e-07,1.869872e-07,1.869876e-07,1.869879e-07,1.869883e-07,1.869887e-07,1.869890e-07,1.869894e-07,1.869897e-07,1.869901e-07,1.869904e-07,1.869908e-07,1.869911e-07,1.869915e-07,1.869918e-07,1.869922e-07,1.869926e-07,1.869929e-07,1.869933e-07,1.869936e-07,1.869940e-07,1.869943e-07,1.869947e-07,1.869950e-07,1.869954e-07,1.869958e-07,1.869961e-07,1.869965e-07,1.869968e-07,1.869972e-07,1.869975e-07,1.869979e-07,1.869982e-07,1.869986e-07,1.869989e-07,1.869993e-07,1.869997e-07,1.870000e-07,1.870004e-07,1.870007e-07,1.870011e-07,1.870014e-07,1.870018e-07,1.870021e-07,1.870025e-07,1.870028e-07,1.870032e-07,1.870036e-07,1.870039e-07,1.870043e-07,1.870046e-07,1.870050e-07,1.870053e-07,1.870057e-07,1.870060e-07,1.870064e-07,1.870067e-07,1.870071e-07,1.870075e-07,1.870078e-07,1.870082e-07,1.870085e-07,1.870089e-07,1.870092e-07,1.870096e-07,1.870099e-07,1.870103e-07,1.870106e-07,1.870110e-07,1.870114e-07,1.870117e-07,1.870121e-07,1.870124e-07,1.870128e-07,1.870131e-07,1.870135e-07,1.870138e-07,1.870142e-07,1.870145e-07,1.870149e-07,1.870153e-07,1.870156e-07,1.870160e-07,1.870163e-07,1.870167e-07,1.870170e-07,1.870174e-07,1.870177e-07,1.870181e-07,1.870184e-07,1.870188e-07,1.870192e-07,1.870195e-07,1.870199e-07,1.870202e-07,1.870206e-07,1.870209e-07,1.870213e-07,1.870216e-07,1.870220e-07,1.870223e-07,1.870227e-07,1.870231e-07,1.870234e-07,1.870238e-07,1.870241e-07,1.870245e-07,1.870248e-07,1.870252e-07,1.870255e-07,1.870259e-07,1.870262e-07,1.870266e-07,1.870269e-07,1.870273e-07,1.870277e-07,1.870280e-07,1.870284e-07,1.870287e-07,1.870291e-07,1.870294e-07,1.870298e-07,1.870301e-07,1.870305e-07,1.870308e-07,1.870312e-07,1.870315e-07,1.870319e-07,1.870323e-07,1.870326e-07,1.870330e-07,1.870333e-07,1.870337e-07,1.870340e-07,1.870344e-07,1.870347e-07,1.870351e-07,1.870354e-07,1.870358e-07,1.870361e-07,1.870365e-07,1.870369e-07,1.870372e-07,1.870376e-07,1.870379e-07,1.870383e-07,1.870386e-07,1.870390e-07,1.870393e-07,1.870397e-07,1.870400e-07,1.870404e-07,1.870407e-07,1.870411e-07,1.870415e-07,1.870418e-07,1.870422e-07,1.870425e-07,1.870429e-07,1.870432e-07,1.870436e-07,1.870439e-07,1.870443e-07,1.870446e-07,1.870450e-07,1.870453e-07,1.870457e-07,1.870460e-07,1.870464e-07,1.870468e-07,1.870471e-07,1.870475e-07,1.870478e-07,1.870482e-07,1.870485e-07,1.870489e-07,1.870492e-07,1.870496e-07,1.870499e-07,1.870503e-07,1.870506e-07,1.870510e-07,1.870513e-07,1.870517e-07,1.870521e-07,1.870524e-07,1.870528e-07,1.870531e-07,1.870535e-07,1.870538e-07,1.870542e-07,1.870545e-07,1.870549e-07,1.870552e-07,1.870556e-07,1.870559e-07,1.870563e-07,1.870566e-07,1.870570e-07,1.870573e-07,1.870577e-07,1.870581e-07,1.870584e-07,1.870588e-07,1.870591e-07,1.870595e-07,1.870598e-07,1.870602e-07,1.870605e-07,1.870609e-07,1.870612e-07,1.870616e-07,1.870619e-07,1.870623e-07,1.870626e-07,1.870630e-07,1.870634e-07,1.870637e-07,1.870641e-07,1.870644e-07,1.870648e-07,1.870651e-07,1.870655e-07,1.870658e-07,1.870662e-07,1.870665e-07,1.870669e-07,1.870672e-07,1.870676e-07,1.870679e-07,1.870683e-07,1.870686e-07,1.870690e-07,1.870693e-07,1.870697e-07,1.870701e-07,1.870704e-07,1.870708e-07,1.870711e-07,1.870715e-07,1.870718e-07,1.870722e-07,1.870725e-07,1.870729e-07,1.870732e-07,1.870736e-07,1.870739e-07,1.870743e-07,1.870746e-07,1.870750e-07,1.870753e-07,1.870757e-07,1.870760e-07,1.870764e-07,1.870768e-07,1.870771e-07,1.870775e-07,1.870778e-07,1.870782e-07,1.870785e-07,1.870789e-07,1.870792e-07,1.870796e-07,1.870799e-07,1.870803e-07,1.870806e-07,1.870810e-07,1.870813e-07,1.870817e-07,1.870820e-07,1.870824e-07,1.870827e-07,1.870831e-07,1.870834e-07,1.870838e-07,1.870842e-07,1.870845e-07,1.870849e-07,1.870852e-07,1.870856e-07,1.870859e-07,1.870863e-07,1.870866e-07,1.870870e-07,1.870873e-07,1.870877e-07,1.870880e-07,1.870884e-07,1.870887e-07,1.870891e-07,1.870894e-07,1.870898e-07,1.870901e-07,1.870905e-07,1.870908e-07,1.870912e-07,1.870915e-07,1.870919e-07,1.870923e-07,1.870926e-07,1.870930e-07,1.870933e-07,1.870937e-07,1.870940e-07,1.870944e-07,1.870947e-07,1.870951e-07,1.870954e-07,1.870958e-07,1.870961e-07,1.870965e-07,1.870968e-07,1.870972e-07,1.870975e-07,1.870979e-07,1.870982e-07,1.870986e-07,1.870989e-07,1.870993e-07,1.870996e-07,1.871000e-07,1.871003e-07,1.871007e-07,1.871010e-07,1.871014e-07,1.871018e-07,1.871021e-07,1.871025e-07,1.871028e-07,1.871032e-07,1.871035e-07,1.871039e-07,1.871042e-07,1.871046e-07,1.871049e-07,1.871053e-07,1.871056e-07,1.871060e-07,1.871063e-07,1.871067e-07,1.871070e-07,1.871074e-07,1.871077e-07,1.871081e-07,1.871084e-07,1.871088e-07,1.871091e-07,1.871095e-07,1.871098e-07,1.871102e-07,1.871105e-07,1.871109e-07,1.871112e-07,1.871116e-07,1.871119e-07,1.871123e-07,1.871127e-07,1.871130e-07,1.871134e-07,1.871137e-07,1.871141e-07,1.871144e-07,1.871148e-07,1.871151e-07,1.871155e-07,1.871158e-07,1.871162e-07,1.871165e-07,1.871169e-07,1.871172e-07,1.871176e-07,1.871179e-07,1.871183e-07,1.871186e-07,1.871190e-07,1.871193e-07,1.871197e-07,1.871200e-07,1.871204e-07,1.871207e-07,1.871211e-07,1.871214e-07,1.871218e-07,1.871221e-07,1.871225e-07,1.871228e-07,1.871232e-07,1.871235e-07,1.871239e-07,1.871242e-07,1.871246e-07,1.871249e-07,1.871253e-07,1.871256e-07,1.871260e-07,1.871263e-07,1.871267e-07,1.871271e-07,1.871274e-07,1.871278e-07,1.871281e-07,1.871285e-07,1.871288e-07,1.871292e-07,1.871295e-07,1.871299e-07,1.871302e-07,1.871306e-07,1.871309e-07,1.871313e-07,1.871316e-07,1.871320e-07,1.871323e-07,1.871327e-07,1.871330e-07,1.871334e-07,1.871337e-07,1.871341e-07,1.871344e-07,1.871348e-07,1.871351e-07,1.871355e-07,1.871358e-07,1.871362e-07,1.871365e-07,1.871369e-07,1.871372e-07,1.871376e-07,1.871379e-07,1.871383e-07,1.871386e-07,1.871390e-07,1.871393e-07,1.871397e-07,1.871400e-07,1.871404e-07,1.871407e-07,1.871411e-07,1.871414e-07,1.871418e-07,1.871421e-07,1.871425e-07,1.871428e-07,1.871432e-07,1.871435e-07,1.871439e-07,1.871442e-07,1.871446e-07,1.871449e-07,1.871453e-07,1.871456e-07,1.871460e-07,1.871463e-07,1.871467e-07,1.871470e-07,1.871474e-07,1.871477e-07,1.871481e-07,1.871484e-07,1.871488e-07,1.871491e-07,1.871495e-07,1.871498e-07,1.871502e-07,1.871505e-07,1.871509e-07,1.871512e-07,1.871516e-07,1.871519e-07,1.871523e-07,1.871526e-07,1.871530e-07,1.871533e-07,1.871537e-07,1.871540e-07,1.871544e-07,1.871547e-07,1.871551e-07,1.871554e-07,1.871558e-07,1.871561e-07,1.871565e-07,1.871568e-07,1.871572e-07,1.871575e-07,1.871579e-07,1.871582e-07,1.871586e-07,1.871589e-07,1.871593e-07,1.871596e-07,1.871600e-07,1.871603e-07,1.871607e-07,1.871610e-07,1.871614e-07,1.871617e-07,1.871621e-07,1.871624e-07,1.871628e-07,1.871631e-07,1.871635e-07,1.871638e-07,1.871642e-07,1.871645e-07,1.871649e-07,1.871652e-07,1.871656e-07,1.871659e-07,1.871663e-07,1.871666e-07,1.871670e-07,1.871673e-07,1.871677e-07,1.871680e-07,1.871684e-07,1.871687e-07,1.871691e-07,1.871694e-07,1.871698e-07,1.871701e-07,1.871705e-07,1.871708e-07,1.871712e-07,1.871715e-07,1.871719e-07,1.871722e-07,1.871726e-07,1.871729e-07,1.871733e-07,1.871736e-07,1.871740e-07,1.871743e-07,1.871747e-07,1.871750e-07,1.871754e-07,1.871757e-07,1.871761e-07,1.871764e-07,1.871768e-07,1.871771e-07,1.871775e-07,1.871778e-07,1.871782e-07,1.871785e-07,1.871789e-07,1.871792e-07,1.871796e-07,1.871799e-07,1.871803e-07,1.871806e-07,1.871810e-07,1.871813e-07,1.871817e-07,1.871820e-07,1.871824e-07,1.871827e-07,1.871831e-07,1.871834e-07,1.871838e-07,1.871841e-07,1.871845e-07,1.871848e-07,1.871852e-07,1.871855e-07,1.871859e-07,1.871862e-07,1.871866e-07,1.871869e-07,1.871873e-07,1.871876e-07,1.871880e-07,1.871883e-07,1.871887e-07,1.871890e-07,1.871894e-07,1.871897e-07,1.871901e-07,1.871904e-07,1.871908e-07,1.871911e-07,1.871915e-07,1.871918e-07,1.871922e-07,1.871925e-07,1.871929e-07,1.871932e-07,1.871935e-07,1.871939e-07,1.871942e-07,1.871946e-07,1.871949e-07,1.871953e-07,1.871956e-07,1.871960e-07,1.871963e-07,1.871967e-07,1.871970e-07,1.871974e-07,1.871977e-07,1.871981e-07,1.871984e-07,1.871988e-07,1.871991e-07,1.871995e-07,1.871998e-07,1.872002e-07,1.872005e-07,1.872009e-07,1.872012e-07,1.872016e-07,1.872019e-07,1.872023e-07,1.872026e-07,1.872030e-07,1.872033e-07,1.872037e-07,1.872040e-07,1.872044e-07,1.872047e-07,1.872051e-07,1.872054e-07,1.872058e-07,1.872061e-07,1.872065e-07,1.872068e-07,1.872072e-07,1.872075e-07,1.872078e-07,1.872082e-07,1.872085e-07,1.872089e-07,1.872092e-07,1.872096e-07,1.872099e-07,1.872103e-07,1.872106e-07,1.872110e-07,1.872113e-07,1.872117e-07,1.872120e-07,1.872124e-07,1.872127e-07,1.872131e-07,1.872134e-07,1.872138e-07,1.872141e-07,1.872145e-07,1.872148e-07,1.872152e-07,1.872155e-07,1.872159e-07,1.872162e-07,1.872166e-07,1.872169e-07,1.872173e-07,1.872176e-07,1.872180e-07,1.872183e-07,1.872186e-07,1.872190e-07,1.872193e-07,1.872197e-07,1.872200e-07,1.872204e-07,1.872207e-07,1.872211e-07,1.872214e-07,1.872218e-07,1.872221e-07,1.872225e-07,1.872228e-07,1.872232e-07,1.872235e-07,1.872239e-07,1.872242e-07,1.872246e-07,1.872249e-07,1.872253e-07,1.872256e-07,1.872260e-07,1.872263e-07,1.872267e-07,1.872270e-07,1.872274e-07,1.872277e-07,1.872280e-07,1.872284e-07,1.872287e-07,1.872291e-07,1.872294e-07,1.872298e-07,1.872301e-07,1.872305e-07,1.872308e-07,1.872312e-07,1.872315e-07,1.872319e-07,1.872322e-07,1.872326e-07,1.872329e-07,1.872333e-07,1.872336e-07,1.872340e-07,1.872343e-07,1.872347e-07,1.872350e-07,1.872354e-07,1.872357e-07,1.872360e-07,1.872364e-07,1.872367e-07,1.872371e-07,1.872374e-07,1.872378e-07,1.872381e-07,1.872385e-07,1.872388e-07,1.872392e-07,1.872395e-07,1.872399e-07,1.872402e-07,1.872406e-07,1.872409e-07,1.872413e-07,1.872416e-07,1.872420e-07,1.872423e-07,1.872427e-07,1.872430e-07,1.872433e-07,1.872437e-07,1.872440e-07,1.872444e-07,1.872447e-07,1.872451e-07,1.872454e-07,1.872458e-07,1.872461e-07,1.872465e-07,1.872468e-07,1.872472e-07,1.872475e-07,1.872479e-07,1.872482e-07,1.872486e-07,1.872489e-07,1.872493e-07,1.872496e-07,1.872499e-07,1.872503e-07,1.872506e-07,1.872510e-07,1.872513e-07,1.872517e-07,1.872520e-07,1.872524e-07,1.872527e-07,1.872531e-07,1.872534e-07,1.872538e-07,1.872541e-07,1.872545e-07,1.872548e-07,1.872552e-07,1.872555e-07,1.872559e-07,1.872562e-07,1.872565e-07,1.872569e-07,1.872572e-07,1.872576e-07,1.872579e-07,1.872583e-07,1.872586e-07,1.872590e-07,1.872593e-07,1.872597e-07,1.872600e-07,1.872604e-07,1.872607e-07,1.872611e-07,1.872614e-07,1.872618e-07,1.872621e-07,1.872624e-07,1.872628e-07,1.872631e-07,1.872635e-07,1.872638e-07,1.872642e-07,1.872645e-07,1.872649e-07,1.872652e-07,1.872656e-07,1.872659e-07,1.872663e-07,1.872666e-07,1.872670e-07,1.872673e-07,1.872676e-07,1.872680e-07,1.872683e-07,1.872687e-07,1.872690e-07,1.872694e-07,1.872697e-07,1.872701e-07,1.872704e-07,1.872708e-07,1.872711e-07,1.872715e-07,1.872718e-07,1.872722e-07,1.872725e-07,1.872728e-07,1.872732e-07,1.872735e-07,1.872739e-07,1.872742e-07,1.872746e-07,1.872749e-07,1.872753e-07,1.872756e-07,1.872760e-07,1.872763e-07,1.872767e-07,1.872770e-07,1.872774e-07,1.872777e-07,1.872780e-07,1.872784e-07,1.872787e-07,1.872791e-07,1.872794e-07,1.872798e-07,1.872801e-07,1.872805e-07,1.872808e-07,1.872812e-07,1.872815e-07,1.872819e-07,1.872822e-07,1.872825e-07,1.872829e-07,1.872832e-07,1.872836e-07,1.872839e-07,1.872843e-07,1.872846e-07,1.872850e-07,1.872853e-07,1.872857e-07,1.872860e-07,1.872864e-07,1.872867e-07,1.872871e-07,1.872874e-07,1.872877e-07,1.872881e-07,1.872884e-07,1.872888e-07,1.872891e-07,1.872895e-07,1.872898e-07,1.872902e-07,1.872905e-07,1.872909e-07,1.872912e-07,1.872916e-07,1.872919e-07,1.872922e-07,1.872926e-07,1.872929e-07,1.872933e-07,1.872936e-07,1.872940e-07,1.872943e-07,1.872947e-07,1.872950e-07,1.872954e-07,1.872957e-07,1.872960e-07,1.872964e-07,1.872967e-07,1.872971e-07,1.872974e-07,1.872978e-07,1.872981e-07,1.872985e-07,1.872988e-07,1.872992e-07,1.872995e-07,1.872999e-07,1.873002e-07,1.873005e-07,1.873009e-07,1.873012e-07,1.873016e-07,1.873019e-07,1.873023e-07,1.873026e-07,1.873030e-07,1.873033e-07,1.873037e-07,1.873040e-07,1.873043e-07,1.873047e-07,1.873050e-07,1.873054e-07,1.873057e-07,1.873061e-07,1.873064e-07,1.873068e-07,1.873071e-07,1.873075e-07,1.873078e-07,1.873082e-07,1.873085e-07,1.873088e-07,1.873092e-07,1.873095e-07,1.873099e-07,1.873102e-07,1.873106e-07,1.873109e-07,1.873113e-07,1.873116e-07,1.873120e-07,1.873123e-07,1.873126e-07,1.873130e-07,1.873133e-07,1.873137e-07,1.873140e-07,1.873144e-07,1.873147e-07,1.873151e-07,1.873154e-07,1.873158e-07,1.873161e-07,1.873164e-07,1.873168e-07,1.873171e-07,1.873175e-07,1.873178e-07,1.873182e-07,1.873185e-07,1.873189e-07,1.873192e-07,1.873195e-07,1.873199e-07,1.873202e-07,1.873206e-07,1.873209e-07,1.873213e-07,1.873216e-07,1.873220e-07,1.873223e-07,1.873227e-07,1.873230e-07,1.873233e-07,1.873237e-07,1.873240e-07,1.873244e-07,1.873247e-07,1.873251e-07,1.873254e-07,1.873258e-07,1.873261e-07,1.873265e-07,1.873268e-07,1.873271e-07,1.873275e-07,1.873278e-07,1.873282e-07,1.873285e-07,1.873289e-07,1.873292e-07,1.873296e-07,1.873299e-07,1.873302e-07,1.873306e-07,1.873309e-07,1.873313e-07,1.873316e-07,1.873320e-07,1.873323e-07,1.873327e-07,1.873330e-07,1.873334e-07,1.873337e-07,1.873340e-07,1.873344e-07,1.873347e-07,1.873351e-07,1.873354e-07,1.873358e-07,1.873361e-07,1.873365e-07,1.873368e-07,1.873371e-07,1.873375e-07,1.873378e-07,1.873382e-07,1.873385e-07,1.873389e-07,1.873392e-07,1.873396e-07,1.873399e-07,1.873402e-07,1.873406e-07,1.873409e-07,1.873413e-07,1.873416e-07,1.873420e-07,1.873423e-07,1.873427e-07,1.873430e-07,1.873433e-07,1.873437e-07,1.873440e-07,1.873444e-07,1.873447e-07,1.873451e-07,1.873454e-07,1.873458e-07,1.873461e-07,1.873464e-07,1.873468e-07,1.873471e-07,1.873475e-07,1.873478e-07,1.873482e-07,1.873485e-07,1.873489e-07,1.873492e-07,1.873495e-07,1.873499e-07,1.873502e-07,1.873506e-07,1.873509e-07,1.873513e-07,1.873516e-07,1.873520e-07,1.873523e-07,1.873526e-07,1.873530e-07,1.873533e-07,1.873537e-07,1.873540e-07,1.873544e-07,1.873547e-07,1.873551e-07,1.873554e-07,1.873557e-07,1.873561e-07,1.873564e-07,1.873568e-07,1.873571e-07,1.873575e-07,1.873578e-07,1.873582e-07,1.873585e-07,1.873588e-07,1.873592e-07,1.873595e-07,1.873599e-07,1.873602e-07,1.873606e-07,1.873609e-07,1.873612e-07,1.873616e-07,1.873619e-07,1.873623e-07,1.873626e-07,1.873630e-07,1.873633e-07,1.873637e-07,1.873640e-07,1.873643e-07,1.873647e-07,1.873650e-07,1.873654e-07,1.873657e-07,1.873661e-07,1.873664e-07,1.873668e-07,1.873671e-07,1.873674e-07,1.873678e-07,1.873681e-07,1.873685e-07,1.873688e-07,1.873692e-07,1.873695e-07,1.873698e-07,1.873702e-07,1.873705e-07,1.873709e-07,1.873712e-07,1.873716e-07,1.873719e-07,1.873723e-07,1.873726e-07,1.873729e-07,1.873733e-07,1.873736e-07,1.873740e-07,1.873743e-07,1.873747e-07,1.873750e-07,1.873753e-07,1.873757e-07,1.873760e-07,1.873764e-07,1.873767e-07,1.873771e-07,1.873774e-07,1.873778e-07,1.873781e-07,1.873784e-07,1.873788e-07,1.873791e-07,1.873795e-07,1.873798e-07,1.873802e-07,1.873805e-07,1.873808e-07,1.873812e-07,1.873815e-07,1.873819e-07,1.873822e-07,1.873826e-07,1.873829e-07,1.873832e-07,1.873836e-07,1.873839e-07,1.873843e-07,1.873846e-07,1.873850e-07,1.873853e-07,1.873856e-07,1.873860e-07,1.873863e-07,1.873867e-07,1.873870e-07,1.873874e-07,1.873877e-07,1.873881e-07,1.873884e-07,1.873887e-07,1.873891e-07,1.873894e-07,1.873898e-07,1.873901e-07,1.873905e-07,1.873908e-07,1.873911e-07,1.873915e-07,1.873918e-07,1.873922e-07,1.873925e-07,1.873929e-07,1.873932e-07,1.873935e-07,1.873939e-07,1.873942e-07,1.873946e-07,1.873949e-07,1.873953e-07,1.873956e-07,1.873959e-07,1.873963e-07,1.873966e-07,1.873970e-07,1.873973e-07,1.873977e-07,1.873980e-07,1.873983e-07,1.873987e-07,1.873990e-07,1.873994e-07,1.873997e-07,1.874001e-07,1.874004e-07,1.874007e-07,1.874011e-07,1.874014e-07,1.874018e-07,1.874021e-07,1.874025e-07,1.874028e-07,1.874031e-07,1.874035e-07,1.874038e-07,1.874042e-07,1.874045e-07,1.874049e-07,1.874052e-07,1.874055e-07,1.874059e-07,1.874062e-07,1.874066e-07,1.874069e-07,1.874073e-07,1.874076e-07,1.874079e-07,1.874083e-07,1.874086e-07,1.874090e-07,1.874093e-07,1.874097e-07,1.874100e-07,1.874103e-07,1.874107e-07,1.874110e-07,1.874114e-07,1.874117e-07,1.874121e-07,1.874124e-07,1.874127e-07,1.874131e-07,1.874134e-07,1.874138e-07,1.874141e-07,1.874145e-07,1.874148e-07,1.874151e-07,1.874155e-07,1.874158e-07,1.874162e-07,1.874165e-07,1.874168e-07,1.874172e-07,1.874175e-07,1.874179e-07,1.874182e-07,1.874186e-07,1.874189e-07,1.874192e-07,1.874196e-07,1.874199e-07,1.874203e-07,1.874206e-07,1.874210e-07,1.874213e-07,1.874216e-07,1.874220e-07,1.874223e-07,1.874227e-07,1.874230e-07,1.874234e-07,1.874237e-07,1.874240e-07,1.874244e-07,1.874247e-07,1.874251e-07,1.874254e-07,1.874257e-07,1.874261e-07,1.874264e-07,1.874268e-07,1.874271e-07,1.874275e-07,1.874278e-07,1.874281e-07,1.874285e-07,1.874288e-07,1.874292e-07,1.874295e-07,1.874299e-07,1.874302e-07,1.874305e-07,1.874309e-07,1.874312e-07,1.874316e-07,1.874319e-07,1.874322e-07,1.874326e-07,1.874329e-07,1.874333e-07,1.874336e-07,1.874340e-07,1.874343e-07,1.874346e-07,1.874350e-07,1.874353e-07,1.874357e-07,1.874360e-07,1.874363e-07,1.874367e-07,1.874370e-07,1.874374e-07,1.874377e-07,1.874381e-07,1.874384e-07,1.874387e-07,1.874391e-07,1.874394e-07,1.874398e-07,1.874401e-07,1.874404e-07,1.874408e-07,1.874411e-07,1.874415e-07,1.874418e-07,1.874422e-07,1.874425e-07,1.874428e-07,1.874432e-07,1.874435e-07,1.874439e-07,1.874442e-07,1.874445e-07,1.874449e-07,1.874452e-07,1.874456e-07,1.874459e-07,1.874463e-07,1.874466e-07,1.874469e-07,1.874473e-07,1.874476e-07,1.874480e-07,1.874483e-07,1.874486e-07,1.874490e-07,1.874493e-07,1.874497e-07,1.874500e-07,1.874504e-07,1.874507e-07,1.874510e-07,1.874514e-07,1.874517e-07,1.874521e-07,1.874524e-07,1.874527e-07,1.874531e-07,1.874534e-07,1.874538e-07,1.874541e-07,1.874544e-07,1.874548e-07,1.874551e-07,1.874555e-07,1.874558e-07,1.874562e-07,1.874565e-07,1.874568e-07,1.874572e-07,1.874575e-07,1.874579e-07,1.874582e-07,1.874585e-07,1.874589e-07,1.874592e-07,1.874596e-07,1.874599e-07,1.874602e-07,1.874606e-07,1.874609e-07,1.874613e-07,1.874616e-07,1.874620e-07,1.874623e-07,1.874626e-07,1.874630e-07,1.874633e-07,1.874637e-07,1.874640e-07,1.874643e-07,1.874647e-07,1.874650e-07,1.874654e-07,1.874657e-07,1.874660e-07,1.874664e-07,1.874667e-07,1.874671e-07,1.874674e-07,1.874678e-07,1.874681e-07,1.874684e-07,1.874688e-07,1.874691e-07,1.874695e-07,1.874698e-07,1.874701e-07,1.874705e-07,1.874708e-07,1.874712e-07,1.874715e-07,1.874718e-07,1.874722e-07,1.874725e-07,1.874729e-07,1.874732e-07,1.874735e-07,1.874739e-07,1.874742e-07,1.874746e-07,1.874749e-07,1.874752e-07,1.874756e-07,1.874759e-07,1.874763e-07,1.874766e-07,1.874770e-07,1.874773e-07,1.874776e-07,1.874780e-07,1.874783e-07,1.874787e-07,1.874790e-07,1.874793e-07,1.874797e-07,1.874800e-07,1.874804e-07,1.874807e-07,1.874810e-07,1.874814e-07,1.874817e-07,1.874821e-07,1.874824e-07,1.874827e-07,1.874831e-07,1.874834e-07,1.874838e-07,1.874841e-07,1.874844e-07,1.874848e-07,1.874851e-07,1.874855e-07,1.874858e-07,1.874861e-07,1.874865e-07,1.874868e-07,1.874872e-07,1.874875e-07,1.874878e-07,1.874882e-07,1.874885e-07,1.874889e-07,1.874892e-07,1.874895e-07,1.874899e-07,1.874902e-07,1.874906e-07,1.874909e-07,1.874912e-07,1.874916e-07,1.874919e-07,1.874923e-07,1.874926e-07,1.874929e-07,1.874933e-07,1.874936e-07,1.874940e-07,1.874943e-07,1.874947e-07,1.874950e-07,1.874953e-07,1.874957e-07,1.874960e-07,1.874964e-07,1.874967e-07,1.874970e-07,1.874974e-07,1.874977e-07,1.874981e-07,1.874984e-07,1.874987e-07,1.874991e-07,1.874994e-07,1.874998e-07,1.875001e-07,1.875004e-07,1.875008e-07,1.875011e-07,1.875015e-07,1.875018e-07,1.875021e-07,1.875025e-07,1.875028e-07,1.875032e-07,1.875035e-07,1.875038e-07,1.875042e-07,1.875045e-07,1.875048e-07,1.875052e-07,1.875055e-07,1.875059e-07,1.875062e-07,1.875065e-07,1.875069e-07,1.875072e-07,1.875076e-07,1.875079e-07,1.875082e-07,1.875086e-07,1.875089e-07,1.875093e-07,1.875096e-07,1.875099e-07,1.875103e-07,1.875106e-07,1.875110e-07,1.875113e-07,1.875116e-07,1.875120e-07,1.875123e-07,1.875127e-07,1.875130e-07,1.875133e-07,1.875137e-07,1.875140e-07,1.875144e-07,1.875147e-07,1.875150e-07,1.875154e-07,1.875157e-07,1.875161e-07,1.875164e-07,1.875167e-07,1.875171e-07,1.875174e-07,1.875178e-07,1.875181e-07,1.875184e-07,1.875188e-07,1.875191e-07,1.875195e-07,1.875198e-07,1.875201e-07,1.875205e-07,1.875208e-07,1.875211e-07,1.875215e-07,1.875218e-07,1.875222e-07,1.875225e-07,1.875228e-07,1.875232e-07,1.875235e-07,1.875239e-07,1.875242e-07,1.875245e-07,1.875249e-07,1.875252e-07,1.875256e-07,1.875259e-07,1.875262e-07,1.875266e-07,1.875269e-07,1.875273e-07,1.875276e-07,1.875279e-07,1.875283e-07,1.875286e-07,1.875290e-07,1.875293e-07,1.875296e-07,1.875300e-07,1.875303e-07,1.875306e-07,1.875310e-07,1.875313e-07,1.875317e-07,1.875320e-07,1.875323e-07,1.875327e-07,1.875330e-07,1.875334e-07,1.875337e-07,1.875340e-07,1.875344e-07,1.875347e-07,1.875351e-07,1.875354e-07,1.875357e-07,1.875361e-07,1.875364e-07,1.875367e-07,1.875371e-07,1.875374e-07,1.875378e-07,1.875381e-07,1.875384e-07,1.875388e-07,1.875391e-07,1.875395e-07,1.875398e-07,1.875401e-07,1.875405e-07,1.875408e-07,1.875412e-07,1.875415e-07,1.875418e-07,1.875422e-07,1.875425e-07,1.875428e-07,1.875432e-07,1.875435e-07,1.875439e-07,1.875442e-07,1.875445e-07,1.875449e-07,1.875452e-07,1.875456e-07,1.875459e-07,1.875462e-07,1.875466e-07,1.875469e-07,1.875472e-07,1.875476e-07,1.875479e-07,1.875483e-07,1.875486e-07,1.875489e-07,1.875493e-07,1.875496e-07,1.875500e-07,1.875503e-07,1.875506e-07,1.875510e-07,1.875513e-07,1.875516e-07,1.875520e-07,1.875523e-07,1.875527e-07,1.875530e-07,1.875533e-07,1.875537e-07,1.875540e-07,1.875544e-07,1.875547e-07,1.875550e-07,1.875554e-07,1.875557e-07,1.875560e-07,1.875564e-07,1.875567e-07,1.875571e-07,1.875574e-07,1.875577e-07,1.875581e-07,1.875584e-07,1.875588e-07,1.875591e-07,1.875594e-07,1.875598e-07,1.875601e-07,1.875604e-07,1.875608e-07,1.875611e-07,1.875615e-07,1.875618e-07,1.875621e-07,1.875625e-07,1.875628e-07,1.875632e-07,1.875635e-07,1.875638e-07,1.875642e-07,1.875645e-07,1.875648e-07,1.875652e-07,1.875655e-07,1.875659e-07,1.875662e-07,1.875665e-07,1.875669e-07,1.875672e-07,1.875675e-07,1.875679e-07,1.875682e-07,1.875686e-07,1.875689e-07,1.875692e-07,1.875696e-07,1.875699e-07,1.875702e-07,1.875706e-07,1.875709e-07,1.875713e-07,1.875716e-07,1.875719e-07,1.875723e-07,1.875726e-07,1.875730e-07,1.875733e-07,1.875736e-07,1.875740e-07,1.875743e-07,1.875746e-07,1.875750e-07,1.875753e-07,1.875757e-07,1.875760e-07,1.875763e-07,1.875767e-07,1.875770e-07,1.875773e-07,1.875777e-07,1.875780e-07,1.875784e-07,1.875787e-07,1.875790e-07,1.875794e-07,1.875797e-07,1.875800e-07,1.875804e-07,1.875807e-07,1.875811e-07,1.875814e-07,1.875817e-07,1.875821e-07,1.875824e-07,1.875827e-07,1.875831e-07,1.875834e-07,1.875838e-07,1.875841e-07,1.875844e-07,1.875848e-07,1.875851e-07,1.875854e-07,1.875858e-07,1.875861e-07,1.875865e-07,1.875868e-07,1.875871e-07,1.875875e-07,1.875878e-07,1.875881e-07,1.875885e-07,1.875888e-07,1.875892e-07,1.875895e-07,1.875898e-07,1.875902e-07,1.875905e-07,1.875908e-07,1.875912e-07,1.875915e-07,1.875919e-07,1.875922e-07,1.875925e-07,1.875929e-07,1.875932e-07,1.875935e-07,1.875939e-07,1.875942e-07,1.875946e-07,1.875949e-07,1.875952e-07,1.875956e-07,1.875959e-07,1.875962e-07,1.875966e-07,1.875969e-07,1.875973e-07,1.875976e-07,1.875979e-07,1.875983e-07,1.875986e-07,1.875989e-07,1.875993e-07,1.875996e-07,1.875999e-07,1.876003e-07,1.876006e-07,1.876010e-07,1.876013e-07,1.876016e-07,1.876020e-07,1.876023e-07,1.876026e-07,1.876030e-07,1.876033e-07,1.876037e-07,1.876040e-07,1.876043e-07,1.876047e-07,1.876050e-07,1.876053e-07,1.876057e-07,1.876060e-07,1.876064e-07,1.876067e-07,1.876070e-07,1.876074e-07,1.876077e-07,1.876080e-07,1.876084e-07,1.876087e-07,1.876090e-07,1.876094e-07,1.876097e-07,1.876101e-07,1.876104e-07,1.876107e-07,1.876111e-07,1.876114e-07,1.876117e-07,1.876121e-07,1.876124e-07,1.876127e-07,1.876131e-07,1.876134e-07,1.876138e-07,1.876141e-07,1.876144e-07,1.876148e-07,1.876151e-07,1.876154e-07,1.876158e-07,1.876161e-07,1.876165e-07,1.876168e-07,1.876171e-07,1.876175e-07,1.876178e-07,1.876181e-07,1.876185e-07,1.876188e-07,1.876191e-07,1.876195e-07,1.876198e-07,1.876202e-07,1.876205e-07,1.876208e-07,1.876212e-07,1.876215e-07,1.876218e-07,1.876222e-07,1.876225e-07,1.876228e-07,1.876232e-07,1.876235e-07,1.876239e-07,1.876242e-07,1.876245e-07,1.876249e-07,1.876252e-07,1.876255e-07,1.876259e-07,1.876262e-07,1.876265e-07,1.876269e-07,1.876272e-07,1.876276e-07,1.876279e-07,1.876282e-07,1.876286e-07,1.876289e-07,1.876292e-07,1.876296e-07,1.876299e-07,1.876302e-07,1.876306e-07,1.876309e-07,1.876313e-07,1.876316e-07,1.876319e-07,1.876323e-07,1.876326e-07,1.876329e-07,1.876333e-07,1.876336e-07,1.876339e-07,1.876343e-07,1.876346e-07,1.876350e-07,1.876353e-07,1.876356e-07,1.876360e-07,1.876363e-07,1.876366e-07,1.876370e-07,1.876373e-07,1.876376e-07,1.876380e-07,1.876383e-07,1.876386e-07,1.876390e-07,1.876393e-07,1.876397e-07,1.876400e-07,1.876403e-07,1.876407e-07,1.876410e-07,1.876413e-07,1.876417e-07,1.876420e-07,1.876423e-07,1.876427e-07,1.876430e-07,1.876433e-07,1.876437e-07,1.876440e-07,1.876444e-07,1.876447e-07,1.876450e-07,1.876454e-07,1.876457e-07,1.876460e-07,1.876464e-07,1.876467e-07,1.876470e-07,1.876474e-07,1.876477e-07,1.876480e-07,1.876484e-07,1.876487e-07,1.876491e-07,1.876494e-07,1.876497e-07,1.876501e-07,1.876504e-07,1.876507e-07,1.876511e-07,1.876514e-07,1.876517e-07,1.876521e-07,1.876524e-07,1.876527e-07,1.876531e-07,1.876534e-07,1.876538e-07,1.876541e-07,1.876544e-07,1.876548e-07,1.876551e-07,1.876554e-07,1.876558e-07,1.876561e-07,1.876564e-07,1.876568e-07,1.876571e-07,1.876574e-07,1.876578e-07,1.876581e-07,1.876584e-07,1.876588e-07,1.876591e-07,1.876595e-07,1.876598e-07,1.876601e-07,1.876605e-07,1.876608e-07,1.876611e-07,1.876615e-07,1.876618e-07,1.876621e-07,1.876625e-07,1.876628e-07,1.876631e-07,1.876635e-07,1.876638e-07,1.876641e-07,1.876645e-07,1.876648e-07,1.876652e-07,1.876655e-07,1.876658e-07,1.876662e-07,1.876665e-07,1.876668e-07,1.876672e-07,1.876675e-07,1.876678e-07,1.876682e-07,1.876685e-07,1.876688e-07,1.876692e-07,1.876695e-07,1.876698e-07,1.876702e-07,1.876705e-07,1.876709e-07,1.876712e-07,1.876715e-07,1.876719e-07,1.876722e-07,1.876725e-07,1.876729e-07,1.876732e-07,1.876735e-07,1.876739e-07,1.876742e-07,1.876745e-07,1.876749e-07,1.876752e-07,1.876755e-07,1.876759e-07,1.876762e-07,1.876765e-07,1.876769e-07,1.876772e-07,1.876776e-07,1.876779e-07,1.876782e-07,1.876786e-07,1.876789e-07,1.876792e-07,1.876796e-07,1.876799e-07,1.876802e-07,1.876806e-07,1.876809e-07,1.876812e-07,1.876816e-07,1.876819e-07,1.876822e-07,1.876826e-07,1.876829e-07,1.876832e-07,1.876836e-07,1.876839e-07,1.876842e-07,1.876846e-07,1.876849e-07,1.876852e-07,1.876856e-07,1.876859e-07,1.876863e-07,1.876866e-07,1.876869e-07,1.876873e-07,1.876876e-07,1.876879e-07,1.876883e-07,1.876886e-07,1.876889e-07,1.876893e-07,1.876896e-07,1.876899e-07,1.876903e-07,1.876906e-07,1.876909e-07,1.876913e-07,1.876916e-07,1.876919e-07,1.876923e-07,1.876926e-07,1.876929e-07,1.876933e-07,1.876936e-07,1.876939e-07,1.876943e-07,1.876946e-07,1.876949e-07,1.876953e-07,1.876956e-07,1.876960e-07,1.876963e-07,1.876966e-07,1.876970e-07,1.876973e-07,1.876976e-07,1.876980e-07,1.876983e-07,1.876986e-07,1.876990e-07,1.876993e-07,1.876996e-07,1.877000e-07,1.877003e-07,1.877006e-07,1.877010e-07,1.877013e-07,1.877016e-07,1.877020e-07,1.877023e-07,1.877026e-07,1.877030e-07,1.877033e-07,1.877036e-07,1.877040e-07,1.877043e-07,1.877046e-07,1.877050e-07,1.877053e-07,1.877056e-07,1.877060e-07,1.877063e-07,1.877066e-07,1.877070e-07,1.877073e-07,1.877076e-07,1.877080e-07,1.877083e-07,1.877086e-07,1.877090e-07,1.877093e-07,1.877096e-07,1.877100e-07,1.877103e-07,1.877107e-07,1.877110e-07,1.877113e-07,1.877117e-07,1.877120e-07,1.877123e-07,1.877127e-07,1.877130e-07,1.877133e-07,1.877137e-07,1.877140e-07,1.877143e-07,1.877147e-07,1.877150e-07,1.877153e-07,1.877157e-07,1.877160e-07,1.877163e-07,1.877167e-07,1.877170e-07,1.877173e-07,1.877177e-07,1.877180e-07,1.877183e-07,1.877187e-07,1.877190e-07,1.877193e-07,1.877197e-07,1.877200e-07,1.877203e-07,1.877207e-07,1.877210e-07,1.877213e-07,1.877217e-07,1.877220e-07,1.877223e-07,1.877227e-07,1.877230e-07,1.877233e-07,1.877237e-07,1.877240e-07,1.877243e-07,1.877247e-07,1.877250e-07,1.877253e-07,1.877257e-07,1.877260e-07,1.877263e-07,1.877267e-07,1.877270e-07,1.877273e-07,1.877277e-07,1.877280e-07,1.877283e-07,1.877287e-07,1.877290e-07,1.877293e-07,1.877297e-07,1.877300e-07,1.877303e-07,1.877307e-07,1.877310e-07,1.877313e-07,1.877317e-07,1.877320e-07,1.877323e-07,1.877327e-07,1.877330e-07,1.877333e-07,1.877337e-07,1.877340e-07,1.877343e-07,1.877347e-07,1.877350e-07,1.877353e-07,1.877357e-07,1.877360e-07,1.877363e-07,1.877367e-07,1.877370e-07,1.877373e-07,1.877377e-07,1.877380e-07,1.877383e-07,1.877387e-07,1.877390e-07,1.877393e-07,1.877397e-07,1.877400e-07,1.877403e-07,1.877407e-07,1.877410e-07,1.877413e-07,1.877417e-07,1.877420e-07,1.877423e-07,1.877427e-07,1.877430e-07,1.877433e-07,1.877437e-07,1.877440e-07,1.877443e-07,1.877447e-07,1.877450e-07,1.877453e-07,1.877457e-07,1.877460e-07,1.877463e-07,1.877467e-07,1.877470e-07,1.877473e-07,1.877477e-07,1.877480e-07,1.877483e-07,1.877487e-07,1.877490e-07,1.877493e-07,1.877497e-07,1.877500e-07,1.877503e-07,1.877506e-07,1.877510e-07,1.877513e-07,1.877516e-07,1.877520e-07,1.877523e-07,1.877526e-07,1.877530e-07,1.877533e-07,1.877536e-07,1.877540e-07,1.877543e-07,1.877546e-07,1.877550e-07,1.877553e-07,1.877556e-07,1.877560e-07,1.877563e-07,1.877566e-07,1.877570e-07,1.877573e-07,1.877576e-07,1.877580e-07,1.877583e-07,1.877586e-07,1.877590e-07,1.877593e-07,1.877596e-07,1.877600e-07,1.877603e-07,1.877606e-07,1.877610e-07,1.877613e-07,1.877616e-07,1.877620e-07,1.877623e-07,1.877626e-07,1.877630e-07,1.877633e-07,1.877636e-07,1.877640e-07,1.877643e-07,1.877646e-07,1.877649e-07,1.877653e-07,1.877656e-07,1.877659e-07,1.877663e-07,1.877666e-07,1.877669e-07,1.877673e-07,1.877676e-07,1.877679e-07,1.877683e-07,1.877686e-07,1.877689e-07,1.877693e-07,1.877696e-07,1.877699e-07,1.877703e-07,1.877706e-07,1.877709e-07,1.877713e-07,1.877716e-07,1.877719e-07,1.877723e-07,1.877726e-07,1.877729e-07,1.877733e-07,1.877736e-07,1.877739e-07,1.877742e-07,1.877746e-07,1.877749e-07,1.877752e-07,1.877756e-07,1.877759e-07,1.877762e-07,1.877766e-07,1.877769e-07,1.877772e-07,1.877776e-07,1.877779e-07,1.877782e-07,1.877786e-07,1.877789e-07,1.877792e-07,1.877796e-07,1.877799e-07,1.877802e-07,1.877806e-07,1.877809e-07,1.877812e-07,1.877816e-07,1.877819e-07,1.877822e-07,1.877825e-07,1.877829e-07,1.877832e-07,1.877835e-07,1.877839e-07,1.877842e-07,1.877845e-07,1.877849e-07,1.877852e-07,1.877855e-07,1.877859e-07,1.877862e-07,1.877865e-07,1.877869e-07,1.877872e-07,1.877875e-07,1.877879e-07,1.877882e-07,1.877885e-07,1.877889e-07,1.877892e-07,1.877895e-07,1.877898e-07,1.877902e-07,1.877905e-07,1.877908e-07,1.877912e-07,1.877915e-07,1.877918e-07,1.877922e-07,1.877925e-07,1.877928e-07,1.877932e-07,1.877935e-07,1.877938e-07,1.877942e-07,1.877945e-07,1.877948e-07,1.877952e-07,1.877955e-07,1.877958e-07,1.877961e-07,1.877965e-07,1.877968e-07,1.877971e-07,1.877975e-07,1.877978e-07,1.877981e-07,1.877985e-07,1.877988e-07,1.877991e-07,1.877995e-07,1.877998e-07,1.878001e-07,1.878005e-07,1.878008e-07,1.878011e-07,1.878014e-07,1.878018e-07,1.878021e-07,1.878024e-07,1.878028e-07,1.878031e-07,1.878034e-07,1.878038e-07,1.878041e-07,1.878044e-07,1.878048e-07,1.878051e-07,1.878054e-07,1.878058e-07,1.878061e-07,1.878064e-07,1.878067e-07,1.878071e-07,1.878074e-07,1.878077e-07,1.878081e-07,1.878084e-07,1.878087e-07,1.878091e-07,1.878094e-07,1.878097e-07,1.878101e-07,1.878104e-07,1.878107e-07,1.878111e-07,1.878114e-07,1.878117e-07,1.878120e-07,1.878124e-07,1.878127e-07,1.878130e-07,1.878134e-07,1.878137e-07,1.878140e-07,1.878144e-07,1.878147e-07,1.878150e-07,1.878154e-07,1.878157e-07,1.878160e-07,1.878163e-07,1.878167e-07,1.878170e-07,1.878173e-07,1.878177e-07,1.878180e-07,1.878183e-07,1.878187e-07,1.878190e-07,1.878193e-07,1.878197e-07,1.878200e-07,1.878203e-07,1.878206e-07,1.878210e-07,1.878213e-07,1.878216e-07,1.878220e-07,1.878223e-07,1.878226e-07,1.878230e-07,1.878233e-07,1.878236e-07,1.878240e-07,1.878243e-07,1.878246e-07,1.878249e-07,1.878253e-07,1.878256e-07,1.878259e-07,1.878263e-07,1.878266e-07,1.878269e-07,1.878273e-07,1.878276e-07,1.878279e-07,1.878283e-07,1.878286e-07,1.878289e-07,1.878292e-07,1.878296e-07,1.878299e-07,1.878302e-07,1.878306e-07,1.878309e-07,1.878312e-07,1.878316e-07,1.878319e-07,1.878322e-07,1.878325e-07,1.878329e-07,1.878332e-07,1.878335e-07,1.878339e-07,1.878342e-07,1.878345e-07,1.878349e-07,1.878352e-07,1.878355e-07,1.878359e-07,1.878362e-07,1.878365e-07,1.878368e-07,1.878372e-07,1.878375e-07,1.878378e-07,1.878382e-07,1.878385e-07,1.878388e-07,1.878392e-07,1.878395e-07,1.878398e-07,1.878401e-07,1.878405e-07,1.878408e-07,1.878411e-07,1.878415e-07,1.878418e-07,1.878421e-07,1.878425e-07,1.878428e-07,1.878431e-07,1.878434e-07,1.878438e-07,1.878441e-07,1.878444e-07,1.878448e-07,1.878451e-07,1.878454e-07,1.878458e-07,1.878461e-07,1.878464e-07,1.878467e-07,1.878471e-07,1.878474e-07,1.878477e-07,1.878481e-07,1.878484e-07,1.878487e-07,1.878491e-07,1.878494e-07,1.878497e-07,1.878500e-07,1.878504e-07,1.878507e-07,1.878510e-07,1.878514e-07,1.878517e-07,1.878520e-07,1.878524e-07,1.878527e-07,1.878530e-07,1.878533e-07,1.878537e-07,1.878540e-07,1.878543e-07,1.878547e-07,1.878550e-07,1.878553e-07,1.878557e-07,1.878560e-07,1.878563e-07,1.878566e-07,1.878570e-07,1.878573e-07,1.878576e-07,1.878580e-07,1.878583e-07,1.878586e-07,1.878590e-07,1.878593e-07,1.878596e-07,1.878599e-07,1.878603e-07,1.878606e-07,1.878609e-07,1.878613e-07,1.878616e-07,1.878619e-07,1.878622e-07,1.878626e-07,1.878629e-07,1.878632e-07,1.878636e-07,1.878639e-07,1.878642e-07,1.878646e-07,1.878649e-07,1.878652e-07,1.878655e-07,1.878659e-07,1.878662e-07,1.878665e-07,1.878669e-07,1.878672e-07,1.878675e-07,1.878678e-07,1.878682e-07,1.878685e-07,1.878688e-07,1.878692e-07,1.878695e-07,1.878698e-07,1.878702e-07,1.878705e-07,1.878708e-07,1.878711e-07,1.878715e-07,1.878718e-07,1.878721e-07,1.878725e-07,1.878728e-07,1.878731e-07,1.878734e-07,1.878738e-07,1.878741e-07,1.878744e-07,1.878748e-07,1.878751e-07,1.878754e-07,1.878758e-07,1.878761e-07,1.878764e-07,1.878767e-07,1.878771e-07,1.878774e-07,1.878777e-07,1.878781e-07,1.878784e-07,1.878787e-07,1.878790e-07,1.878794e-07,1.878797e-07,1.878800e-07,1.878804e-07,1.878807e-07,1.878810e-07,1.878813e-07,1.878817e-07,1.878820e-07,1.878823e-07,1.878827e-07,1.878830e-07,1.878833e-07,1.878836e-07,1.878840e-07,1.878843e-07,1.878846e-07,1.878850e-07,1.878853e-07,1.878856e-07,1.878860e-07,1.878863e-07,1.878866e-07,1.878869e-07,1.878873e-07,1.878876e-07,1.878879e-07,1.878883e-07,1.878886e-07,1.878889e-07,1.878892e-07,1.878896e-07,1.878899e-07,1.878902e-07,1.878906e-07,1.878909e-07,1.878912e-07,1.878915e-07,1.878919e-07,1.878922e-07,1.878925e-07,1.878929e-07,1.878932e-07,1.878935e-07,1.878938e-07,1.878942e-07,1.878945e-07,1.878948e-07,1.878952e-07,1.878955e-07,1.878958e-07,1.878961e-07,1.878965e-07,1.878968e-07,1.878971e-07,1.878975e-07,1.878978e-07,1.878981e-07,1.878984e-07,1.878988e-07,1.878991e-07,1.878994e-07,1.878998e-07,1.879001e-07,1.879004e-07,1.879007e-07,1.879011e-07,1.879014e-07,1.879017e-07,1.879021e-07,1.879024e-07,1.879027e-07,1.879030e-07,1.879034e-07,1.879037e-07,1.879040e-07,1.879044e-07,1.879047e-07,1.879050e-07,1.879053e-07,1.879057e-07,1.879060e-07,1.879063e-07,1.879067e-07,1.879070e-07,1.879073e-07,1.879076e-07,1.879080e-07,1.879083e-07,1.879086e-07,1.879090e-07,1.879093e-07,1.879096e-07,1.879099e-07,1.879103e-07,1.879106e-07,1.879109e-07,1.879113e-07,1.879116e-07,1.879119e-07,1.879122e-07,1.879126e-07,1.879129e-07,1.879132e-07,1.879135e-07,1.879139e-07,1.879142e-07,1.879145e-07,1.879149e-07,1.879152e-07,1.879155e-07,1.879158e-07,1.879162e-07,1.879165e-07,1.879168e-07,1.879172e-07,1.879175e-07,1.879178e-07,1.879181e-07,1.879185e-07,1.879188e-07,1.879191e-07,1.879195e-07,1.879198e-07,1.879201e-07,1.879204e-07,1.879208e-07,1.879211e-07,1.879214e-07,1.879217e-07,1.879221e-07,1.879224e-07,1.879227e-07,1.879231e-07,1.879234e-07,1.879237e-07,1.879240e-07,1.879244e-07,1.879247e-07,1.879250e-07,1.879254e-07,1.879257e-07,1.879260e-07,1.879263e-07,1.879267e-07,1.879270e-07,1.879273e-07,1.879276e-07,1.879280e-07,1.879283e-07,1.879286e-07,1.879290e-07,1.879293e-07,1.879296e-07,1.879299e-07,1.879303e-07,1.879306e-07,1.879309e-07,1.879313e-07,1.879316e-07,1.879319e-07,1.879322e-07,1.879326e-07,1.879329e-07,1.879332e-07,1.879335e-07,1.879339e-07,1.879342e-07,1.879345e-07,1.879349e-07,1.879352e-07,1.879355e-07,1.879358e-07,1.879362e-07,1.879365e-07,1.879368e-07,1.879371e-07,1.879375e-07,1.879378e-07,1.879381e-07,1.879385e-07,1.879388e-07,1.879391e-07,1.879394e-07,1.879398e-07,1.879401e-07,1.879404e-07,1.879408e-07,1.879411e-07,1.879414e-07,1.879417e-07,1.879421e-07,1.879424e-07,1.879427e-07,1.879430e-07,1.879434e-07,1.879437e-07,1.879440e-07,1.879444e-07,1.879447e-07,1.879450e-07,1.879453e-07,1.879457e-07,1.879460e-07,1.879463e-07,1.879466e-07,1.879470e-07,1.879473e-07,1.879476e-07,1.879480e-07,1.879483e-07,1.879486e-07,1.879489e-07,1.879493e-07,1.879496e-07,1.879499e-07,1.879502e-07,1.879506e-07,1.879509e-07,1.879512e-07,1.879515e-07,1.879519e-07,1.879522e-07,1.879525e-07,1.879529e-07,1.879532e-07,1.879535e-07,1.879538e-07,1.879542e-07,1.879545e-07,1.879548e-07,1.879551e-07,1.879555e-07,1.879558e-07,1.879561e-07,1.879565e-07,1.879568e-07,1.879571e-07,1.879574e-07,1.879578e-07,1.879581e-07,1.879584e-07,1.879587e-07,1.879591e-07,1.879594e-07,1.879597e-07,1.879600e-07,1.879604e-07,1.879607e-07,1.879610e-07,1.879614e-07,1.879617e-07,1.879620e-07,1.879623e-07,1.879627e-07,1.879630e-07,1.879633e-07,1.879636e-07,1.879640e-07,1.879643e-07,1.879646e-07,1.879650e-07,1.879653e-07,1.879656e-07,1.879659e-07,1.879663e-07,1.879666e-07,1.879669e-07,1.879672e-07,1.879676e-07,1.879679e-07,1.879682e-07,1.879685e-07,1.879689e-07,1.879692e-07,1.879695e-07,1.879699e-07,1.879702e-07,1.879705e-07,1.879708e-07,1.879712e-07,1.879715e-07,1.879718e-07,1.879721e-07,1.879725e-07,1.879728e-07,1.879731e-07,1.879734e-07,1.879738e-07,1.879741e-07,1.879744e-07,1.879747e-07,1.879751e-07,1.879754e-07,1.879757e-07,1.879761e-07,1.879764e-07,1.879767e-07,1.879770e-07,1.879774e-07,1.879777e-07,1.879780e-07,1.879783e-07,1.879787e-07,1.879790e-07,1.879793e-07,1.879796e-07,1.879800e-07,1.879803e-07,1.879806e-07,1.879809e-07,1.879813e-07,1.879816e-07,1.879819e-07,1.879823e-07,1.879826e-07,1.879829e-07,1.879832e-07,1.879836e-07,1.879839e-07,1.879842e-07,1.879845e-07,1.879849e-07,1.879852e-07,1.879855e-07,1.879858e-07,1.879862e-07,1.879865e-07,1.879868e-07,1.879871e-07,1.879875e-07,1.879878e-07,1.879881e-07,1.879884e-07,1.879888e-07,1.879891e-07,1.879894e-07,1.879898e-07,1.879901e-07,1.879904e-07,1.879907e-07,1.879911e-07,1.879914e-07,1.879917e-07,1.879920e-07,1.879924e-07,1.879927e-07,1.879930e-07,1.879933e-07,1.879937e-07,1.879940e-07,1.879943e-07,1.879946e-07,1.879950e-07,1.879953e-07,1.879956e-07,1.879959e-07,1.879963e-07,1.879966e-07,1.879969e-07,1.879972e-07,1.879976e-07,1.879979e-07,1.879982e-07,1.879986e-07,1.879989e-07,1.879992e-07,1.879995e-07,1.879999e-07,1.880002e-07,1.880005e-07,1.880008e-07,1.880012e-07,1.880015e-07,1.880018e-07,1.880021e-07,1.880025e-07,1.880028e-07,1.880031e-07,1.880034e-07,1.880038e-07,1.880041e-07,1.880044e-07,1.880047e-07,1.880051e-07,1.880054e-07,1.880057e-07,1.880060e-07,1.880064e-07,1.880067e-07,1.880070e-07,1.880073e-07,1.880077e-07,1.880080e-07,1.880083e-07,1.880086e-07,1.880090e-07,1.880093e-07,1.880096e-07,1.880099e-07,1.880103e-07,1.880106e-07,1.880109e-07,1.880112e-07,1.880116e-07,1.880119e-07,1.880122e-07,1.880126e-07,1.880129e-07,1.880132e-07,1.880135e-07,1.880139e-07,1.880142e-07,1.880145e-07,1.880148e-07,1.880152e-07,1.880155e-07,1.880158e-07,1.880161e-07,1.880165e-07,1.880168e-07,1.880171e-07,1.880174e-07,1.880178e-07,1.880181e-07,1.880184e-07,1.880187e-07,1.880191e-07,1.880194e-07,1.880197e-07,1.880200e-07,1.880204e-07,1.880207e-07,1.880210e-07,1.880213e-07,1.880217e-07,1.880220e-07,1.880223e-07,1.880226e-07,1.880230e-07,1.880233e-07,1.880236e-07,1.880239e-07,1.880243e-07,1.880246e-07,1.880249e-07,1.880252e-07,1.880256e-07,1.880259e-07,1.880262e-07,1.880265e-07,1.880269e-07,1.880272e-07,1.880275e-07,1.880278e-07,1.880282e-07,1.880285e-07,1.880288e-07,1.880291e-07,1.880295e-07,1.880298e-07,1.880301e-07,1.880304e-07,1.880308e-07,1.880311e-07,1.880314e-07,1.880317e-07,1.880321e-07,1.880324e-07,1.880327e-07,1.880330e-07,1.880334e-07,1.880337e-07,1.880340e-07,1.880343e-07,1.880347e-07,1.880350e-07,1.880353e-07,1.880356e-07,1.880360e-07,1.880363e-07,1.880366e-07,1.880369e-07,1.880373e-07,1.880376e-07,1.880379e-07,1.880382e-07,1.880386e-07,1.880389e-07,1.880392e-07,1.880395e-07,1.880398e-07,1.880402e-07,1.880405e-07,1.880408e-07,1.880411e-07,1.880415e-07,1.880418e-07,1.880421e-07,1.880424e-07,1.880428e-07,1.880431e-07,1.880434e-07,1.880437e-07,1.880441e-07,1.880444e-07,1.880447e-07,1.880450e-07,1.880454e-07,1.880457e-07,1.880460e-07,1.880463e-07,1.880467e-07,1.880470e-07,1.880473e-07,1.880476e-07,1.880480e-07,1.880483e-07,1.880486e-07,1.880489e-07,1.880493e-07,1.880496e-07,1.880499e-07,1.880502e-07,1.880506e-07,1.880509e-07,1.880512e-07,1.880515e-07,1.880519e-07,1.880522e-07,1.880525e-07,1.880528e-07,1.880532e-07,1.880535e-07,1.880538e-07,1.880541e-07,1.880544e-07,1.880548e-07,1.880551e-07,1.880554e-07,1.880557e-07,1.880561e-07,1.880564e-07,1.880567e-07,1.880570e-07,1.880574e-07,1.880577e-07,1.880580e-07,1.880583e-07,1.880587e-07,1.880590e-07,1.880593e-07,1.880596e-07,1.880600e-07,1.880603e-07,1.880606e-07,1.880609e-07,1.880613e-07,1.880616e-07,1.880619e-07,1.880622e-07,1.880625e-07,1.880629e-07,1.880632e-07,1.880635e-07,1.880638e-07,1.880642e-07,1.880645e-07,1.880648e-07,1.880651e-07,1.880655e-07,1.880658e-07,1.880661e-07,1.880664e-07,1.880668e-07,1.880671e-07,1.880674e-07,1.880677e-07,1.880681e-07,1.880684e-07,1.880687e-07,1.880690e-07,1.880694e-07,1.880697e-07,1.880700e-07,1.880703e-07,1.880706e-07,1.880710e-07,1.880713e-07,1.880716e-07,1.880719e-07,1.880723e-07,1.880726e-07,1.880729e-07,1.880732e-07,1.880736e-07,1.880739e-07,1.880742e-07,1.880745e-07,1.880749e-07,1.880752e-07,1.880755e-07,1.880758e-07,1.880761e-07,1.880765e-07,1.880768e-07,1.880771e-07,1.880774e-07,1.880778e-07,1.880781e-07,1.880784e-07,1.880787e-07,1.880791e-07,1.880794e-07,1.880797e-07,1.880800e-07,1.880804e-07,1.880807e-07,1.880810e-07,1.880813e-07,1.880816e-07,1.880820e-07,1.880823e-07,1.880826e-07,1.880829e-07,1.880833e-07,1.880836e-07,1.880839e-07,1.880842e-07,1.880846e-07,1.880849e-07,1.880852e-07,1.880855e-07,1.880859e-07,1.880862e-07,1.880865e-07,1.880868e-07,1.880871e-07,1.880875e-07,1.880878e-07,1.880881e-07,1.880884e-07,1.880888e-07,1.880891e-07,1.880894e-07,1.880897e-07,1.880901e-07,1.880904e-07,1.880907e-07,1.880910e-07,1.880913e-07,1.880917e-07,1.880920e-07,1.880923e-07,1.880926e-07,1.880930e-07,1.880933e-07,1.880936e-07,1.880939e-07,1.880943e-07,1.880946e-07,1.880949e-07,1.880952e-07,1.880955e-07,1.880959e-07,1.880962e-07,1.880965e-07,1.880968e-07,1.880972e-07,1.880975e-07,1.880978e-07,1.880981e-07,1.880985e-07,1.880988e-07,1.880991e-07,1.880994e-07,1.880997e-07,1.881001e-07,1.881004e-07,1.881007e-07,1.881010e-07,1.881014e-07,1.881017e-07,1.881020e-07,1.881023e-07,1.881027e-07,1.881030e-07,1.881033e-07,1.881036e-07,1.881039e-07,1.881043e-07,1.881046e-07,1.881049e-07,1.881052e-07,1.881056e-07,1.881059e-07,1.881062e-07,1.881065e-07,1.881068e-07,1.881072e-07,1.881075e-07,1.881078e-07,1.881081e-07,1.881085e-07,1.881088e-07,1.881091e-07,1.881094e-07,1.881098e-07,1.881101e-07,1.881104e-07,1.881107e-07,1.881110e-07,1.881114e-07,1.881117e-07,1.881120e-07,1.881123e-07,1.881127e-07,1.881130e-07,1.881133e-07,1.881136e-07,1.881139e-07,1.881143e-07,1.881146e-07,1.881149e-07,1.881152e-07,1.881156e-07,1.881159e-07,1.881162e-07,1.881165e-07,1.881169e-07,1.881172e-07,1.881175e-07,1.881178e-07,1.881181e-07,1.881185e-07,1.881188e-07,1.881191e-07,1.881194e-07,1.881198e-07,1.881201e-07,1.881204e-07,1.881207e-07,1.881210e-07,1.881214e-07,1.881217e-07,1.881220e-07,1.881223e-07,1.881227e-07,1.881230e-07,1.881233e-07,1.881236e-07,1.881239e-07,1.881243e-07,1.881246e-07,1.881249e-07,1.881252e-07,1.881256e-07,1.881259e-07,1.881262e-07,1.881265e-07,1.881268e-07,1.881272e-07,1.881275e-07,1.881278e-07,1.881281e-07,1.881285e-07,1.881288e-07,1.881291e-07,1.881294e-07,1.881297e-07,1.881301e-07,1.881304e-07,1.881307e-07,1.881310e-07,1.881314e-07,1.881317e-07,1.881320e-07,1.881323e-07,1.881326e-07,1.881330e-07,1.881333e-07,1.881336e-07,1.881339e-07,1.881343e-07,1.881346e-07,1.881349e-07,1.881352e-07,1.881355e-07,1.881359e-07,1.881362e-07,1.881365e-07,1.881368e-07,1.881371e-07,1.881375e-07,1.881378e-07,1.881381e-07,1.881384e-07,1.881388e-07,1.881391e-07,1.881394e-07,1.881397e-07,1.881400e-07,1.881404e-07,1.881407e-07,1.881410e-07,1.881413e-07,1.881417e-07,1.881420e-07,1.881423e-07,1.881426e-07,1.881429e-07,1.881433e-07,1.881436e-07,1.881439e-07,1.881442e-07,1.881446e-07,1.881449e-07,1.881452e-07,1.881455e-07,1.881458e-07,1.881462e-07,1.881465e-07,1.881468e-07,1.881471e-07,1.881474e-07,1.881478e-07,1.881481e-07,1.881484e-07,1.881487e-07,1.881491e-07,1.881494e-07,1.881497e-07,1.881500e-07,1.881503e-07,1.881507e-07,1.881510e-07,1.881513e-07,1.881516e-07,1.881519e-07,1.881523e-07,1.881526e-07,1.881529e-07,1.881532e-07,1.881536e-07,1.881539e-07,1.881542e-07,1.881545e-07,1.881548e-07,1.881552e-07,1.881555e-07,1.881558e-07,1.881561e-07,1.881564e-07,1.881568e-07,1.881571e-07,1.881574e-07,1.881577e-07,1.881581e-07,1.881584e-07,1.881587e-07,1.881590e-07,1.881593e-07,1.881597e-07,1.881600e-07,1.881603e-07,1.881606e-07,1.881609e-07,1.881613e-07,1.881616e-07,1.881619e-07,1.881622e-07,1.881626e-07,1.881629e-07,1.881632e-07,1.881635e-07,1.881638e-07,1.881642e-07,1.881645e-07,1.881648e-07,1.881651e-07,1.881654e-07,1.881658e-07,1.881661e-07,1.881664e-07,1.881667e-07,1.881670e-07,1.881674e-07,1.881677e-07,1.881680e-07,1.881683e-07,1.881687e-07,1.881690e-07,1.881693e-07,1.881696e-07,1.881699e-07,1.881703e-07,1.881706e-07,1.881709e-07,1.881712e-07,1.881715e-07,1.881719e-07,1.881722e-07,1.881725e-07,1.881728e-07,1.881731e-07,1.881735e-07,1.881738e-07,1.881741e-07,1.881744e-07,1.881748e-07,1.881751e-07,1.881754e-07,1.881757e-07,1.881760e-07,1.881764e-07,1.881767e-07,1.881770e-07,1.881773e-07,1.881776e-07,1.881780e-07,1.881783e-07,1.881786e-07,1.881789e-07,1.881792e-07,1.881796e-07,1.881799e-07,1.881802e-07,1.881805e-07,1.881808e-07,1.881812e-07,1.881815e-07,1.881818e-07,1.881821e-07,1.881825e-07,1.881828e-07,1.881831e-07,1.881834e-07,1.881837e-07,1.881841e-07,1.881844e-07,1.881847e-07,1.881850e-07,1.881853e-07,1.881857e-07,1.881860e-07,1.881863e-07,1.881866e-07,1.881869e-07,1.881873e-07,1.881876e-07,1.881879e-07,1.881882e-07,1.881885e-07,1.881889e-07,1.881892e-07,1.881895e-07,1.881898e-07,1.881901e-07,1.881905e-07,1.881908e-07,1.881911e-07,1.881914e-07,1.881917e-07,1.881921e-07,1.881924e-07,1.881927e-07,1.881930e-07,1.881933e-07,1.881937e-07,1.881940e-07,1.881943e-07,1.881946e-07,1.881949e-07,1.881953e-07,1.881956e-07,1.881959e-07,1.881962e-07,1.881966e-07,1.881969e-07,1.881972e-07,1.881975e-07,1.881978e-07,1.881982e-07,1.881985e-07,1.881988e-07,1.881991e-07,1.881994e-07,1.881998e-07,1.882001e-07,1.882004e-07,1.882007e-07,1.882010e-07,1.882014e-07,1.882017e-07,1.882020e-07,1.882023e-07,1.882026e-07,1.882030e-07,1.882033e-07,1.882036e-07,1.882039e-07,1.882042e-07,1.882046e-07,1.882049e-07,1.882052e-07,1.882055e-07,1.882058e-07,1.882062e-07,1.882065e-07,1.882068e-07,1.882071e-07,1.882074e-07,1.882078e-07,1.882081e-07,1.882084e-07,1.882087e-07,1.882090e-07,1.882094e-07,1.882097e-07,1.882100e-07,1.882103e-07,1.882106e-07,1.882110e-07,1.882113e-07,1.882116e-07,1.882119e-07,1.882122e-07,1.882126e-07,1.882129e-07,1.882132e-07,1.882135e-07,1.882138e-07,1.882142e-07,1.882145e-07,1.882148e-07,1.882151e-07,1.882154e-07,1.882158e-07,1.882161e-07,1.882164e-07,1.882167e-07,1.882170e-07,1.882174e-07,1.882177e-07,1.882180e-07,1.882183e-07,1.882186e-07,1.882189e-07,1.882193e-07,1.882196e-07,1.882199e-07,1.882202e-07,1.882205e-07,1.882209e-07,1.882212e-07,1.882215e-07,1.882218e-07,1.882221e-07,1.882225e-07,1.882228e-07,1.882231e-07,1.882234e-07,1.882237e-07,1.882241e-07,1.882244e-07,1.882247e-07,1.882250e-07,1.882253e-07,1.882257e-07,1.882260e-07,1.882263e-07,1.882266e-07,1.882269e-07,1.882273e-07,1.882276e-07,1.882279e-07,1.882282e-07,1.882285e-07,1.882289e-07,1.882292e-07,1.882295e-07,1.882298e-07,1.882301e-07,1.882305e-07,1.882308e-07,1.882311e-07,1.882314e-07,1.882317e-07,1.882320e-07,1.882324e-07,1.882327e-07,1.882330e-07,1.882333e-07,1.882336e-07,1.882340e-07,1.882343e-07,1.882346e-07,1.882349e-07,1.882352e-07,1.882356e-07,1.882359e-07,1.882362e-07,1.882365e-07,1.882368e-07,1.882372e-07,1.882375e-07,1.882378e-07,1.882381e-07,1.882384e-07,1.882388e-07,1.882391e-07,1.882394e-07,1.882397e-07,1.882400e-07,1.882403e-07,1.882407e-07,1.882410e-07,1.882413e-07,1.882416e-07,1.882419e-07,1.882423e-07,1.882426e-07,1.882429e-07,1.882432e-07,1.882435e-07,1.882439e-07,1.882442e-07,1.882445e-07,1.882448e-07,1.882451e-07,1.882455e-07,1.882458e-07,1.882461e-07,1.882464e-07,1.882467e-07,1.882470e-07,1.882474e-07,1.882477e-07,1.882480e-07,1.882483e-07,1.882486e-07,1.882490e-07,1.882493e-07,1.882496e-07,1.882499e-07,1.882502e-07,1.882506e-07,1.882509e-07,1.882512e-07,1.882515e-07,1.882518e-07,1.882521e-07,1.882525e-07,1.882528e-07,1.882531e-07,1.882534e-07,1.882537e-07,1.882541e-07,1.882544e-07,1.882547e-07,1.882550e-07,1.882553e-07,1.882557e-07,1.882560e-07,1.882563e-07,1.882566e-07,1.882569e-07,1.882572e-07,1.882576e-07,1.882579e-07,1.882582e-07,1.882585e-07,1.882588e-07,1.882592e-07,1.882595e-07,1.882598e-07,1.882601e-07,1.882604e-07,1.882608e-07,1.882611e-07,1.882614e-07,1.882617e-07,1.882620e-07,1.882623e-07,1.882627e-07,1.882630e-07,1.882633e-07,1.882636e-07,1.882639e-07,1.882643e-07,1.882646e-07,1.882649e-07,1.882652e-07,1.882655e-07,1.882658e-07,1.882662e-07,1.882665e-07,1.882668e-07,1.882671e-07,1.882674e-07,1.882678e-07,1.882681e-07,1.882684e-07,1.882687e-07,1.882690e-07,1.882693e-07,1.882697e-07,1.882700e-07,1.882703e-07,1.882706e-07,1.882709e-07,1.882713e-07,1.882716e-07,1.882719e-07,1.882722e-07,1.882725e-07,1.882728e-07,1.882732e-07,1.882735e-07,1.882738e-07,1.882741e-07,1.882744e-07,1.882748e-07,1.882751e-07,1.882754e-07,1.882757e-07,1.882760e-07,1.882763e-07,1.882767e-07,1.882770e-07,1.882773e-07,1.882776e-07,1.882779e-07,1.882783e-07,1.882786e-07,1.882789e-07,1.882792e-07,1.882795e-07,1.882798e-07,1.882802e-07,1.882805e-07,1.882808e-07,1.882811e-07,1.882814e-07,1.882818e-07,1.882821e-07,1.882824e-07,1.882827e-07,1.882830e-07,1.882833e-07,1.882837e-07,1.882840e-07,1.882843e-07,1.882846e-07,1.882849e-07,1.882853e-07,1.882856e-07,1.882859e-07,1.882862e-07,1.882865e-07,1.882868e-07,1.882872e-07,1.882875e-07,1.882878e-07,1.882881e-07,1.882884e-07,1.882887e-07,1.882891e-07,1.882894e-07,1.882897e-07,1.882900e-07,1.882903e-07,1.882907e-07,1.882910e-07,1.882913e-07,1.882916e-07,1.882919e-07,1.882922e-07,1.882926e-07,1.882929e-07,1.882932e-07,1.882935e-07,1.882938e-07,1.882941e-07,1.882945e-07,1.882948e-07,1.882951e-07,1.882954e-07,1.882957e-07,1.882961e-07,1.882964e-07,1.882967e-07,1.882970e-07,1.882973e-07,1.882976e-07,1.882980e-07,1.882983e-07,1.882986e-07,1.882989e-07,1.882992e-07,1.882995e-07,1.882999e-07,1.883002e-07,1.883005e-07,1.883008e-07,1.883011e-07,1.883015e-07,1.883018e-07,1.883021e-07,1.883024e-07,1.883027e-07,1.883030e-07,1.883034e-07,1.883037e-07,1.883040e-07,1.883043e-07,1.883046e-07,1.883049e-07,1.883053e-07,1.883056e-07,1.883059e-07,1.883062e-07,1.883065e-07,1.883068e-07,1.883072e-07,1.883075e-07,1.883078e-07,1.883081e-07,1.883084e-07,1.883087e-07,1.883091e-07,1.883094e-07,1.883097e-07,1.883100e-07,1.883103e-07,1.883107e-07,1.883110e-07,1.883113e-07,1.883116e-07,1.883119e-07,1.883122e-07,1.883126e-07,1.883129e-07,1.883132e-07,1.883135e-07,1.883138e-07,1.883141e-07,1.883145e-07,1.883148e-07,1.883151e-07,1.883154e-07,1.883157e-07,1.883160e-07,1.883164e-07,1.883167e-07,1.883170e-07,1.883173e-07,1.883176e-07,1.883179e-07,1.883183e-07,1.883186e-07,1.883189e-07,1.883192e-07,1.883195e-07,1.883198e-07,1.883202e-07,1.883205e-07,1.883208e-07,1.883211e-07,1.883214e-07,1.883217e-07,1.883221e-07,1.883224e-07,1.883227e-07,1.883230e-07,1.883233e-07,1.883236e-07,1.883240e-07,1.883243e-07,1.883246e-07,1.883249e-07,1.883252e-07,1.883256e-07,1.883259e-07,1.883262e-07,1.883265e-07,1.883268e-07,1.883271e-07,1.883275e-07,1.883278e-07,1.883281e-07,1.883284e-07,1.883287e-07,1.883290e-07,1.883294e-07,1.883297e-07,1.883300e-07,1.883303e-07,1.883306e-07,1.883309e-07,1.883313e-07,1.883316e-07,1.883319e-07,1.883322e-07,1.883325e-07,1.883328e-07,1.883331e-07,1.883335e-07,1.883338e-07,1.883341e-07,1.883344e-07,1.883347e-07,1.883350e-07,1.883354e-07,1.883357e-07,1.883360e-07,1.883363e-07,1.883366e-07,1.883369e-07,1.883373e-07,1.883376e-07,1.883379e-07,1.883382e-07,1.883385e-07,1.883388e-07,1.883392e-07,1.883395e-07,1.883398e-07,1.883401e-07,1.883404e-07,1.883407e-07,1.883411e-07,1.883414e-07,1.883417e-07,1.883420e-07,1.883423e-07,1.883426e-07,1.883430e-07,1.883433e-07,1.883436e-07,1.883439e-07,1.883442e-07,1.883445e-07,1.883449e-07,1.883452e-07,1.883455e-07,1.883458e-07,1.883461e-07,1.883464e-07,1.883468e-07,1.883471e-07,1.883474e-07,1.883477e-07,1.883480e-07,1.883483e-07,1.883487e-07,1.883490e-07,1.883493e-07,1.883496e-07,1.883499e-07,1.883502e-07,1.883505e-07,1.883509e-07,1.883512e-07,1.883515e-07,1.883518e-07,1.883521e-07,1.883524e-07,1.883528e-07,1.883531e-07,1.883534e-07,1.883537e-07,1.883540e-07,1.883543e-07,1.883547e-07,1.883550e-07,1.883553e-07,1.883556e-07,1.883559e-07,1.883562e-07,1.883566e-07,1.883569e-07,1.883572e-07,1.883575e-07,1.883578e-07,1.883581e-07,1.883584e-07,1.883588e-07,1.883591e-07,1.883594e-07,1.883597e-07,1.883600e-07,1.883603e-07,1.883607e-07,1.883610e-07,1.883613e-07,1.883616e-07,1.883619e-07,1.883622e-07,1.883626e-07,1.883629e-07,1.883632e-07,1.883635e-07,1.883638e-07,1.883641e-07,1.883644e-07,1.883648e-07,1.883651e-07,1.883654e-07,1.883657e-07,1.883660e-07,1.883663e-07,1.883667e-07,1.883670e-07,1.883673e-07,1.883676e-07,1.883679e-07,1.883682e-07,1.883686e-07,1.883689e-07,1.883692e-07,1.883695e-07,1.883698e-07,1.883701e-07,1.883704e-07,1.883708e-07,1.883711e-07,1.883714e-07,1.883717e-07,1.883720e-07,1.883723e-07,1.883727e-07,1.883730e-07,1.883733e-07,1.883736e-07,1.883739e-07,1.883742e-07,1.883745e-07,1.883749e-07,1.883752e-07,1.883755e-07,1.883758e-07,1.883761e-07,1.883764e-07,1.883768e-07,1.883771e-07,1.883774e-07,1.883777e-07,1.883780e-07,1.883783e-07,1.883786e-07,1.883790e-07,1.883793e-07,1.883796e-07,1.883799e-07,1.883802e-07,1.883805e-07,1.883809e-07,1.883812e-07,1.883815e-07,1.883818e-07,1.883821e-07,1.883824e-07,1.883827e-07,1.883831e-07,1.883834e-07,1.883837e-07,1.883840e-07,1.883843e-07,1.883846e-07,1.883850e-07,1.883853e-07,1.883856e-07,1.883859e-07,1.883862e-07,1.883865e-07,1.883868e-07,1.883872e-07,1.883875e-07,1.883878e-07,1.883881e-07,1.883884e-07,1.883887e-07,1.883890e-07,1.883894e-07,1.883897e-07,1.883900e-07,1.883903e-07,1.883906e-07,1.883909e-07,1.883913e-07,1.883916e-07,1.883919e-07,1.883922e-07,1.883925e-07,1.883928e-07,1.883931e-07,1.883935e-07,1.883938e-07,1.883941e-07,1.883944e-07,1.883947e-07,1.883950e-07,1.883953e-07,1.883957e-07,1.883960e-07,1.883963e-07,1.883966e-07,1.883969e-07,1.883972e-07,1.883976e-07,1.883979e-07,1.883982e-07,1.883985e-07,1.883988e-07,1.883991e-07,1.883994e-07,1.883998e-07,1.884001e-07,1.884004e-07,1.884007e-07,1.884010e-07,1.884013e-07,1.884016e-07,1.884020e-07,1.884023e-07,1.884026e-07,1.884029e-07,1.884032e-07,1.884035e-07,1.884038e-07,1.884042e-07,1.884045e-07,1.884048e-07,1.884051e-07,1.884054e-07,1.884057e-07,1.884060e-07,1.884064e-07,1.884067e-07,1.884070e-07,1.884073e-07,1.884076e-07,1.884079e-07,1.884082e-07,1.884086e-07,1.884089e-07,1.884092e-07,1.884095e-07,1.884098e-07,1.884101e-07,1.884105e-07,1.884108e-07,1.884111e-07,1.884114e-07,1.884117e-07,1.884120e-07,1.884123e-07,1.884127e-07,1.884130e-07,1.884133e-07,1.884136e-07,1.884139e-07,1.884142e-07,1.884145e-07,1.884149e-07,1.884152e-07,1.884155e-07,1.884158e-07,1.884161e-07,1.884164e-07,1.884167e-07,1.884171e-07,1.884174e-07,1.884177e-07,1.884180e-07,1.884183e-07,1.884186e-07,1.884189e-07,1.884193e-07,1.884196e-07,1.884199e-07,1.884202e-07,1.884205e-07,1.884208e-07,1.884211e-07,1.884215e-07,1.884218e-07,1.884221e-07,1.884224e-07,1.884227e-07,1.884230e-07,1.884233e-07,1.884237e-07,1.884240e-07,1.884243e-07,1.884246e-07,1.884249e-07,1.884252e-07,1.884255e-07,1.884258e-07,1.884262e-07,1.884265e-07,1.884268e-07,1.884271e-07,1.884274e-07,1.884277e-07,1.884280e-07,1.884284e-07,1.884287e-07,1.884290e-07,1.884293e-07,1.884296e-07,1.884299e-07,1.884302e-07,1.884306e-07,1.884309e-07,1.884312e-07,1.884315e-07,1.884318e-07,1.884321e-07,1.884324e-07,1.884328e-07,1.884331e-07,1.884334e-07,1.884337e-07,1.884340e-07,1.884343e-07,1.884346e-07,1.884350e-07,1.884353e-07,1.884356e-07,1.884359e-07,1.884362e-07,1.884365e-07,1.884368e-07,1.884371e-07,1.884375e-07,1.884378e-07,1.884381e-07,1.884384e-07,1.884387e-07,1.884390e-07,1.884393e-07,1.884397e-07,1.884400e-07,1.884403e-07,1.884406e-07,1.884409e-07,1.884412e-07,1.884415e-07,1.884419e-07,1.884422e-07,1.884425e-07,1.884428e-07,1.884431e-07,1.884434e-07,1.884437e-07,1.884441e-07,1.884444e-07,1.884447e-07,1.884450e-07,1.884453e-07,1.884456e-07,1.884459e-07,1.884462e-07,1.884466e-07,1.884469e-07,1.884472e-07,1.884475e-07,1.884478e-07,1.884481e-07,1.884484e-07,1.884488e-07,1.884491e-07,1.884494e-07,1.884497e-07,1.884500e-07,1.884503e-07,1.884506e-07,1.884509e-07,1.884513e-07,1.884516e-07,1.884519e-07,1.884522e-07,1.884525e-07,1.884528e-07,1.884531e-07,1.884535e-07,1.884538e-07,1.884541e-07,1.884544e-07,1.884547e-07,1.884550e-07,1.884553e-07,1.884556e-07,1.884560e-07,1.884563e-07,1.884566e-07,1.884569e-07,1.884572e-07,1.884575e-07,1.884578e-07,1.884582e-07,1.884585e-07,1.884588e-07,1.884591e-07,1.884594e-07,1.884597e-07,1.884600e-07,1.884603e-07,1.884607e-07,1.884610e-07,1.884613e-07,1.884616e-07,1.884619e-07,1.884622e-07,1.884625e-07,1.884628e-07,1.884632e-07,1.884635e-07,1.884638e-07,1.884641e-07,1.884644e-07,1.884647e-07,1.884650e-07,1.884654e-07,1.884657e-07,1.884660e-07,1.884663e-07,1.884666e-07,1.884669e-07,1.884672e-07,1.884675e-07,1.884679e-07,1.884682e-07,1.884685e-07,1.884688e-07,1.884691e-07,1.884694e-07,1.884697e-07,1.884700e-07,1.884704e-07,1.884707e-07,1.884710e-07,1.884713e-07,1.884716e-07,1.884719e-07,1.884722e-07,1.884726e-07,1.884729e-07,1.884732e-07,1.884735e-07,1.884738e-07,1.884741e-07,1.884744e-07,1.884747e-07,1.884751e-07,1.884754e-07,1.884757e-07,1.884760e-07,1.884763e-07,1.884766e-07,1.884769e-07,1.884772e-07,1.884776e-07,1.884779e-07,1.884782e-07,1.884785e-07,1.884788e-07,1.884791e-07,1.884794e-07,1.884797e-07,1.884801e-07,1.884804e-07,1.884807e-07,1.884810e-07,1.884813e-07,1.884816e-07,1.884819e-07,1.884822e-07,1.884826e-07,1.884829e-07,1.884832e-07,1.884835e-07,1.884838e-07,1.884841e-07,1.884844e-07,1.884847e-07,1.884851e-07,1.884854e-07,1.884857e-07,1.884860e-07,1.884863e-07,1.884866e-07,1.884869e-07,1.884872e-07,1.884876e-07,1.884879e-07,1.884882e-07,1.884885e-07,1.884888e-07,1.884891e-07,1.884894e-07,1.884897e-07,1.884901e-07,1.884904e-07,1.884907e-07,1.884910e-07,1.884913e-07,1.884916e-07,1.884919e-07,1.884922e-07,1.884926e-07,1.884929e-07,1.884932e-07,1.884935e-07,1.884938e-07,1.884941e-07,1.884944e-07,1.884947e-07,1.884951e-07,1.884954e-07,1.884957e-07,1.884960e-07,1.884963e-07,1.884966e-07,1.884969e-07,1.884972e-07,1.884975e-07,1.884979e-07,1.884982e-07,1.884985e-07,1.884988e-07,1.884991e-07,1.884994e-07,1.884997e-07,1.885000e-07,1.885004e-07,1.885007e-07,1.885010e-07,1.885013e-07,1.885016e-07,1.885019e-07,1.885022e-07,1.885025e-07,1.885029e-07,1.885032e-07,1.885035e-07,1.885038e-07,1.885041e-07,1.885044e-07,1.885047e-07,1.885050e-07,1.885053e-07,1.885057e-07,1.885060e-07,1.885063e-07,1.885066e-07,1.885069e-07,1.885072e-07,1.885075e-07,1.885078e-07,1.885082e-07,1.885085e-07,1.885088e-07,1.885091e-07,1.885094e-07,1.885097e-07,1.885100e-07,1.885103e-07,1.885107e-07,1.885110e-07,1.885113e-07,1.885116e-07,1.885119e-07,1.885122e-07,1.885125e-07,1.885128e-07,1.885131e-07,1.885135e-07,1.885138e-07,1.885141e-07,1.885144e-07,1.885147e-07,1.885150e-07,1.885153e-07,1.885156e-07,1.885159e-07,1.885163e-07,1.885166e-07,1.885169e-07,1.885172e-07,1.885175e-07,1.885178e-07,1.885181e-07,1.885184e-07,1.885188e-07,1.885191e-07,1.885194e-07,1.885197e-07,1.885200e-07,1.885203e-07,1.885206e-07,1.885209e-07,1.885212e-07,1.885216e-07,1.885219e-07,1.885222e-07,1.885225e-07,1.885228e-07,1.885231e-07,1.885234e-07,1.885237e-07,1.885240e-07,1.885244e-07,1.885247e-07,1.885250e-07,1.885253e-07,1.885256e-07,1.885259e-07,1.885262e-07,1.885265e-07,1.885269e-07,1.885272e-07,1.885275e-07,1.885278e-07,1.885281e-07,1.885284e-07,1.885287e-07,1.885290e-07,1.885293e-07,1.885297e-07,1.885300e-07,1.885303e-07,1.885306e-07,1.885309e-07,1.885312e-07,1.885315e-07,1.885318e-07,1.885321e-07,1.885325e-07,1.885328e-07,1.885331e-07,1.885334e-07,1.885337e-07,1.885340e-07,1.885343e-07,1.885346e-07,1.885349e-07,1.885353e-07,1.885356e-07,1.885359e-07,1.885362e-07,1.885365e-07,1.885368e-07,1.885371e-07,1.885374e-07,1.885377e-07,1.885381e-07,1.885384e-07,1.885387e-07,1.885390e-07,1.885393e-07,1.885396e-07,1.885399e-07,1.885402e-07,1.885405e-07,1.885409e-07,1.885412e-07,1.885415e-07,1.885418e-07,1.885421e-07,1.885424e-07,1.885427e-07,1.885430e-07,1.885433e-07,1.885437e-07,1.885440e-07,1.885443e-07,1.885446e-07,1.885449e-07,1.885452e-07,1.885455e-07,1.885458e-07,1.885461e-07,1.885465e-07,1.885468e-07,1.885471e-07,1.885474e-07,1.885477e-07,1.885480e-07,1.885483e-07,1.885486e-07,1.885489e-07,1.885492e-07,1.885496e-07,1.885499e-07,1.885502e-07,1.885505e-07,1.885508e-07,1.885511e-07,1.885514e-07,1.885517e-07,1.885520e-07,1.885524e-07,1.885527e-07,1.885530e-07,1.885533e-07,1.885536e-07,1.885539e-07,1.885542e-07,1.885545e-07,1.885548e-07,1.885552e-07,1.885555e-07,1.885558e-07,1.885561e-07,1.885564e-07,1.885567e-07,1.885570e-07,1.885573e-07,1.885576e-07,1.885579e-07,1.885583e-07,1.885586e-07,1.885589e-07,1.885592e-07,1.885595e-07,1.885598e-07,1.885601e-07,1.885604e-07,1.885607e-07,1.885611e-07,1.885614e-07,1.885617e-07,1.885620e-07,1.885623e-07,1.885626e-07,1.885629e-07,1.885632e-07,1.885635e-07,1.885638e-07,1.885642e-07,1.885645e-07,1.885648e-07,1.885651e-07,1.885654e-07,1.885657e-07,1.885660e-07,1.885663e-07,1.885666e-07,1.885669e-07,1.885673e-07,1.885676e-07,1.885679e-07,1.885682e-07,1.885685e-07,1.885688e-07,1.885691e-07,1.885694e-07,1.885697e-07,1.885701e-07,1.885704e-07,1.885707e-07,1.885710e-07,1.885713e-07,1.885716e-07,1.885719e-07,1.885722e-07,1.885725e-07,1.885728e-07,1.885732e-07,1.885735e-07,1.885738e-07,1.885741e-07,1.885744e-07,1.885747e-07,1.885750e-07,1.885753e-07,1.885756e-07,1.885759e-07,1.885763e-07,1.885766e-07,1.885769e-07,1.885772e-07,1.885775e-07,1.885778e-07,1.885781e-07,1.885784e-07,1.885787e-07,1.885790e-07,1.885794e-07,1.885797e-07,1.885800e-07,1.885803e-07,1.885806e-07,1.885809e-07,1.885812e-07,1.885815e-07,1.885818e-07,1.885821e-07,1.885825e-07,1.885828e-07,1.885831e-07,1.885834e-07,1.885837e-07,1.885840e-07,1.885843e-07,1.885846e-07,1.885849e-07,1.885852e-07,1.885856e-07,1.885859e-07,1.885862e-07,1.885865e-07,1.885868e-07,1.885871e-07,1.885874e-07,1.885877e-07,1.885880e-07,1.885883e-07,1.885886e-07,1.885890e-07,1.885893e-07,1.885896e-07,1.885899e-07,1.885902e-07,1.885905e-07,1.885908e-07,1.885911e-07,1.885914e-07,1.885917e-07,1.885921e-07,1.885924e-07,1.885927e-07,1.885930e-07,1.885933e-07,1.885936e-07,1.885939e-07,1.885942e-07,1.885945e-07,1.885948e-07,1.885951e-07,1.885955e-07,1.885958e-07,1.885961e-07,1.885964e-07,1.885967e-07,1.885970e-07,1.885973e-07,1.885976e-07,1.885979e-07,1.885982e-07,1.885986e-07,1.885989e-07,1.885992e-07,1.885995e-07,1.885998e-07,1.886001e-07,1.886004e-07,1.886007e-07,1.886010e-07,1.886013e-07,1.886016e-07,1.886020e-07,1.886023e-07,1.886026e-07,1.886029e-07,1.886032e-07,1.886035e-07,1.886038e-07,1.886041e-07,1.886044e-07,1.886047e-07,1.886051e-07,1.886054e-07,1.886057e-07,1.886060e-07,1.886063e-07,1.886066e-07,1.886069e-07,1.886072e-07,1.886075e-07,1.886078e-07,1.886081e-07,1.886085e-07,1.886088e-07,1.886091e-07,1.886094e-07,1.886097e-07,1.886100e-07,1.886103e-07,1.886106e-07,1.886109e-07,1.886112e-07,1.886115e-07,1.886119e-07,1.886122e-07,1.886125e-07,1.886128e-07,1.886131e-07,1.886134e-07,1.886137e-07,1.886140e-07,1.886143e-07,1.886146e-07,1.886149e-07,1.886153e-07,1.886156e-07,1.886159e-07,1.886162e-07,1.886165e-07,1.886168e-07,1.886171e-07,1.886174e-07,1.886177e-07,1.886180e-07,1.886183e-07,1.886187e-07,1.886190e-07,1.886193e-07,1.886196e-07,1.886199e-07,1.886202e-07,1.886205e-07,1.886208e-07,1.886211e-07,1.886214e-07,1.886217e-07,1.886220e-07,1.886224e-07,1.886227e-07,1.886230e-07,1.886233e-07,1.886236e-07,1.886239e-07,1.886242e-07,1.886245e-07,1.886248e-07,1.886251e-07,1.886254e-07,1.886258e-07,1.886261e-07,1.886264e-07,1.886267e-07,1.886270e-07,1.886273e-07,1.886276e-07,1.886279e-07,1.886282e-07,1.886285e-07,1.886288e-07,1.886291e-07,1.886295e-07,1.886298e-07,1.886301e-07,1.886304e-07,1.886307e-07,1.886310e-07,1.886313e-07,1.886316e-07,1.886319e-07,1.886322e-07,1.886325e-07,1.886329e-07,1.886332e-07,1.886335e-07,1.886338e-07,1.886341e-07,1.886344e-07,1.886347e-07,1.886350e-07,1.886353e-07,1.886356e-07,1.886359e-07,1.886362e-07,1.886366e-07,1.886369e-07,1.886372e-07,1.886375e-07,1.886378e-07,1.886381e-07,1.886384e-07,1.886387e-07,1.886390e-07,1.886393e-07,1.886396e-07,1.886399e-07,1.886403e-07,1.886406e-07,1.886409e-07,1.886412e-07,1.886415e-07,1.886418e-07,1.886421e-07,1.886424e-07,1.886427e-07,1.886430e-07,1.886433e-07,1.886436e-07,1.886440e-07,1.886443e-07,1.886446e-07,1.886449e-07,1.886452e-07,1.886455e-07,1.886458e-07,1.886461e-07,1.886464e-07,1.886467e-07,1.886470e-07,1.886473e-07,1.886477e-07,1.886480e-07,1.886483e-07,1.886486e-07,1.886489e-07,1.886492e-07,1.886495e-07,1.886498e-07,1.886501e-07,1.886504e-07,1.886507e-07,1.886510e-07,1.886514e-07,1.886517e-07,1.886520e-07,1.886523e-07,1.886526e-07,1.886529e-07,1.886532e-07,1.886535e-07,1.886538e-07,1.886541e-07,1.886544e-07,1.886547e-07,1.886550e-07,1.886554e-07,1.886557e-07,1.886560e-07,1.886563e-07,1.886566e-07,1.886569e-07,1.886572e-07,1.886575e-07,1.886578e-07,1.886581e-07,1.886584e-07,1.886587e-07,1.886590e-07,1.886594e-07,1.886597e-07,1.886600e-07,1.886603e-07,1.886606e-07,1.886609e-07,1.886612e-07,1.886615e-07,1.886618e-07,1.886621e-07,1.886624e-07,1.886627e-07,1.886631e-07,1.886634e-07,1.886637e-07,1.886640e-07,1.886643e-07,1.886646e-07,1.886649e-07,1.886652e-07,1.886655e-07,1.886658e-07,1.886661e-07,1.886664e-07,1.886667e-07,1.886671e-07,1.886674e-07,1.886677e-07,1.886680e-07,1.886683e-07,1.886686e-07,1.886689e-07,1.886692e-07,1.886695e-07,1.886698e-07,1.886701e-07,1.886704e-07,1.886707e-07,1.886710e-07,1.886714e-07,1.886717e-07,1.886720e-07,1.886723e-07,1.886726e-07,1.886729e-07,1.886732e-07,1.886735e-07,1.886738e-07,1.886741e-07,1.886744e-07,1.886747e-07,1.886750e-07,1.886754e-07,1.886757e-07,1.886760e-07,1.886763e-07,1.886766e-07,1.886769e-07,1.886772e-07,1.886775e-07,1.886778e-07,1.886781e-07,1.886784e-07,1.886787e-07,1.886790e-07,1.886794e-07,1.886797e-07,1.886800e-07,1.886803e-07,1.886806e-07,1.886809e-07,1.886812e-07,1.886815e-07,1.886818e-07,1.886821e-07,1.886824e-07,1.886827e-07,1.886830e-07,1.886833e-07,1.886837e-07,1.886840e-07,1.886843e-07,1.886846e-07,1.886849e-07,1.886852e-07,1.886855e-07,1.886858e-07,1.886861e-07,1.886864e-07,1.886867e-07,1.886870e-07,1.886873e-07,1.886876e-07,1.886880e-07,1.886883e-07,1.886886e-07,1.886889e-07,1.886892e-07,1.886895e-07,1.886898e-07,1.886901e-07,1.886904e-07,1.886907e-07,1.886910e-07,1.886913e-07,1.886916e-07,1.886919e-07,1.886923e-07,1.886926e-07,1.886929e-07,1.886932e-07,1.886935e-07,1.886938e-07,1.886941e-07,1.886944e-07,1.886947e-07,1.886950e-07,1.886953e-07,1.886956e-07,1.886959e-07,1.886962e-07,1.886965e-07,1.886969e-07,1.886972e-07,1.886975e-07,1.886978e-07,1.886981e-07,1.886984e-07,1.886987e-07,1.886990e-07,1.886993e-07,1.886996e-07,1.886999e-07,1.887002e-07,1.887005e-07,1.887008e-07,1.887011e-07,1.887015e-07,1.887018e-07,1.887021e-07,1.887024e-07,1.887027e-07,1.887030e-07,1.887033e-07,1.887036e-07,1.887039e-07,1.887042e-07,1.887045e-07,1.887048e-07,1.887051e-07,1.887054e-07,1.887057e-07,1.887061e-07,1.887064e-07,1.887067e-07,1.887070e-07,1.887073e-07,1.887076e-07,1.887079e-07,1.887082e-07,1.887085e-07,1.887088e-07,1.887091e-07,1.887094e-07,1.887097e-07,1.887100e-07,1.887103e-07,1.887107e-07,1.887110e-07,1.887113e-07,1.887116e-07,1.887119e-07,1.887122e-07,1.887125e-07,1.887128e-07,1.887131e-07,1.887134e-07,1.887137e-07,1.887140e-07,1.887143e-07,1.887146e-07,1.887149e-07,1.887153e-07,1.887156e-07,1.887159e-07,1.887162e-07,1.887165e-07,1.887168e-07,1.887171e-07,1.887174e-07,1.887177e-07,1.887180e-07,1.887183e-07,1.887186e-07,1.887189e-07,1.887192e-07,1.887195e-07,1.887198e-07,1.887202e-07,1.887205e-07,1.887208e-07,1.887211e-07,1.887214e-07,1.887217e-07,1.887220e-07,1.887223e-07,1.887226e-07,1.887229e-07,1.887232e-07,1.887235e-07,1.887238e-07,1.887241e-07,1.887244e-07,1.887247e-07,1.887251e-07,1.887254e-07,1.887257e-07,1.887260e-07,1.887263e-07,1.887266e-07,1.887269e-07,1.887272e-07,1.887275e-07,1.887278e-07,1.887281e-07,1.887284e-07,1.887287e-07,1.887290e-07,1.887293e-07,1.887296e-07,1.887299e-07,1.887303e-07,1.887306e-07,1.887309e-07,1.887312e-07,1.887315e-07,1.887318e-07,1.887321e-07,1.887324e-07,1.887327e-07,1.887330e-07,1.887333e-07,1.887336e-07,1.887339e-07,1.887342e-07,1.887345e-07,1.887348e-07,1.887351e-07,1.887355e-07,1.887358e-07,1.887361e-07,1.887364e-07,1.887367e-07,1.887370e-07,1.887373e-07,1.887376e-07,1.887379e-07,1.887382e-07,1.887385e-07,1.887388e-07,1.887391e-07,1.887394e-07,1.887397e-07,1.887400e-07,1.887403e-07,1.887407e-07,1.887410e-07,1.887413e-07,1.887416e-07,1.887419e-07,1.887422e-07,1.887425e-07,1.887428e-07,1.887431e-07,1.887434e-07,1.887437e-07,1.887440e-07,1.887443e-07,1.887446e-07,1.887449e-07,1.887452e-07,1.887455e-07,1.887458e-07,1.887462e-07,1.887465e-07,1.887468e-07,1.887471e-07,1.887474e-07,1.887477e-07,1.887480e-07,1.887483e-07,1.887486e-07,1.887489e-07,1.887492e-07,1.887495e-07,1.887498e-07,1.887501e-07,1.887504e-07,1.887507e-07,1.887510e-07,1.887513e-07,1.887517e-07,1.887520e-07,1.887523e-07,1.887526e-07,1.887529e-07,1.887532e-07,1.887535e-07,1.887538e-07,1.887541e-07,1.887544e-07,1.887547e-07,1.887550e-07,1.887553e-07,1.887556e-07,1.887559e-07,1.887562e-07,1.887565e-07,1.887568e-07,1.887571e-07,1.887575e-07,1.887578e-07,1.887581e-07,1.887584e-07,1.887587e-07,1.887590e-07,1.887593e-07,1.887596e-07,1.887599e-07,1.887602e-07,1.887605e-07,1.887608e-07,1.887611e-07,1.887614e-07,1.887617e-07,1.887620e-07,1.887623e-07,1.887626e-07,1.887629e-07,1.887633e-07,1.887636e-07,1.887639e-07,1.887642e-07,1.887645e-07,1.887648e-07,1.887651e-07,1.887654e-07,1.887657e-07,1.887660e-07,1.887663e-07,1.887666e-07,1.887669e-07,1.887672e-07,1.887675e-07,1.887678e-07,1.887681e-07,1.887684e-07,1.887687e-07,1.887690e-07,1.887694e-07,1.887697e-07,1.887700e-07,1.887703e-07,1.887706e-07,1.887709e-07,1.887712e-07,1.887715e-07,1.887718e-07,1.887721e-07,1.887724e-07,1.887727e-07,1.887730e-07,1.887733e-07,1.887736e-07,1.887739e-07,1.887742e-07,1.887745e-07,1.887748e-07,1.887751e-07,1.887755e-07,1.887758e-07,1.887761e-07,1.887764e-07,1.887767e-07,1.887770e-07,1.887773e-07,1.887776e-07,1.887779e-07,1.887782e-07,1.887785e-07,1.887788e-07,1.887791e-07,1.887794e-07,1.887797e-07,1.887800e-07,1.887803e-07,1.887806e-07,1.887809e-07,1.887812e-07,1.887815e-07,1.887819e-07,1.887822e-07,1.887825e-07,1.887828e-07,1.887831e-07,1.887834e-07,1.887837e-07,1.887840e-07,1.887843e-07,1.887846e-07,1.887849e-07,1.887852e-07,1.887855e-07,1.887858e-07,1.887861e-07,1.887864e-07,1.887867e-07,1.887870e-07,1.887873e-07,1.887876e-07,1.887879e-07,1.887882e-07,1.887886e-07,1.887889e-07,1.887892e-07,1.887895e-07,1.887898e-07,1.887901e-07,1.887904e-07,1.887907e-07,1.887910e-07,1.887913e-07,1.887916e-07,1.887919e-07,1.887922e-07,1.887925e-07,1.887928e-07,1.887931e-07,1.887934e-07,1.887937e-07,1.887940e-07,1.887943e-07,1.887946e-07,1.887949e-07,1.887952e-07,1.887956e-07,1.887959e-07,1.887962e-07,1.887965e-07,1.887968e-07,1.887971e-07,1.887974e-07,1.887977e-07,1.887980e-07,1.887983e-07,1.887986e-07,1.887989e-07,1.887992e-07,1.887995e-07,1.887998e-07,1.888001e-07,1.888004e-07,1.888007e-07,1.888010e-07,1.888013e-07,1.888016e-07,1.888019e-07,1.888022e-07,1.888025e-07,1.888029e-07,1.888032e-07,1.888035e-07,1.888038e-07,1.888041e-07,1.888044e-07,1.888047e-07,1.888050e-07,1.888053e-07,1.888056e-07,1.888059e-07,1.888062e-07,1.888065e-07,1.888068e-07,1.888071e-07,1.888074e-07,1.888077e-07,1.888080e-07,1.888083e-07,1.888086e-07,1.888089e-07,1.888092e-07,1.888095e-07,1.888098e-07,1.888101e-07,1.888105e-07,1.888108e-07,1.888111e-07,1.888114e-07,1.888117e-07,1.888120e-07,1.888123e-07,1.888126e-07,1.888129e-07,1.888132e-07,1.888135e-07,1.888138e-07,1.888141e-07,1.888144e-07,1.888147e-07,1.888150e-07,1.888153e-07,1.888156e-07,1.888159e-07,1.888162e-07,1.888165e-07,1.888168e-07,1.888171e-07,1.888174e-07,1.888177e-07,1.888180e-07,1.888183e-07,1.888187e-07,1.888190e-07,1.888193e-07,1.888196e-07,1.888199e-07,1.888202e-07,1.888205e-07,1.888208e-07,1.888211e-07,1.888214e-07,1.888217e-07,1.888220e-07,1.888223e-07,1.888226e-07,1.888229e-07,1.888232e-07,1.888235e-07,1.888238e-07,1.888241e-07,1.888244e-07,1.888247e-07,1.888250e-07,1.888253e-07,1.888256e-07,1.888259e-07,1.888262e-07,1.888265e-07,1.888269e-07,1.888272e-07,1.888275e-07,1.888278e-07,1.888281e-07,1.888284e-07,1.888287e-07,1.888290e-07,1.888293e-07,1.888296e-07,1.888299e-07,1.888302e-07,1.888305e-07,1.888308e-07,1.888311e-07,1.888314e-07,1.888317e-07,1.888320e-07,1.888323e-07,1.888326e-07,1.888329e-07,1.888332e-07,1.888335e-07,1.888338e-07,1.888341e-07,1.888344e-07,1.888347e-07,1.888350e-07,1.888353e-07,1.888356e-07,1.888360e-07,1.888363e-07,1.888366e-07,1.888369e-07,1.888372e-07,1.888375e-07,1.888378e-07,1.888381e-07,1.888384e-07,1.888387e-07,1.888390e-07,1.888393e-07,1.888396e-07,1.888399e-07,1.888402e-07,1.888405e-07,1.888408e-07,1.888411e-07,1.888414e-07,1.888417e-07,1.888420e-07,1.888423e-07,1.888426e-07,1.888429e-07,1.888432e-07,1.888435e-07,1.888438e-07,1.888441e-07,1.888444e-07,1.888447e-07,1.888450e-07,1.888453e-07,1.888456e-07,1.888460e-07,1.888463e-07,1.888466e-07,1.888469e-07,1.888472e-07,1.888475e-07,1.888478e-07,1.888481e-07,1.888484e-07,1.888487e-07,1.888490e-07,1.888493e-07,1.888496e-07,1.888499e-07,1.888502e-07,1.888505e-07,1.888508e-07,1.888511e-07,1.888514e-07,1.888517e-07,1.888520e-07,1.888523e-07,1.888526e-07,1.888529e-07,1.888532e-07,1.888535e-07,1.888538e-07,1.888541e-07,1.888544e-07,1.888547e-07,1.888550e-07,1.888553e-07,1.888556e-07,1.888559e-07,1.888562e-07,1.888566e-07,1.888569e-07,1.888572e-07,1.888575e-07,1.888578e-07,1.888581e-07,1.888584e-07,1.888587e-07,1.888590e-07,1.888593e-07,1.888596e-07,1.888599e-07,1.888602e-07,1.888605e-07,1.888608e-07,1.888611e-07,1.888614e-07,1.888617e-07,1.888620e-07,1.888623e-07,1.888626e-07,1.888629e-07,1.888632e-07,1.888635e-07,1.888638e-07,1.888641e-07,1.888644e-07,1.888647e-07,1.888650e-07,1.888653e-07,1.888656e-07,1.888659e-07,1.888662e-07,1.888665e-07,1.888668e-07,1.888671e-07,1.888674e-07,1.888677e-07,1.888680e-07,1.888684e-07,1.888687e-07,1.888690e-07,1.888693e-07,1.888696e-07,1.888699e-07,1.888702e-07,1.888705e-07,1.888708e-07,1.888711e-07,1.888714e-07,1.888717e-07,1.888720e-07,1.888723e-07,1.888726e-07,1.888729e-07,1.888732e-07,1.888735e-07,1.888738e-07,1.888741e-07,1.888744e-07,1.888747e-07,1.888750e-07,1.888753e-07,1.888756e-07,1.888759e-07,1.888762e-07,1.888765e-07,1.888768e-07,1.888771e-07,1.888774e-07,1.888777e-07,1.888780e-07,1.888783e-07,1.888786e-07,1.888789e-07,1.888792e-07,1.888795e-07,1.888798e-07,1.888801e-07,1.888804e-07,1.888807e-07,1.888810e-07,1.888813e-07,1.888816e-07,1.888820e-07,1.888823e-07,1.888826e-07,1.888829e-07,1.888832e-07,1.888835e-07,1.888838e-07,1.888841e-07,1.888844e-07,1.888847e-07,1.888850e-07,1.888853e-07,1.888856e-07,1.888859e-07,1.888862e-07,1.888865e-07,1.888868e-07,1.888871e-07,1.888874e-07,1.888877e-07,1.888880e-07,1.888883e-07,1.888886e-07,1.888889e-07,1.888892e-07,1.888895e-07,1.888898e-07,1.888901e-07,1.888904e-07,1.888907e-07,1.888910e-07,1.888913e-07,1.888916e-07,1.888919e-07,1.888922e-07,1.888925e-07,1.888928e-07,1.888931e-07,1.888934e-07,1.888937e-07,1.888940e-07,1.888943e-07,1.888946e-07,1.888949e-07,1.888952e-07,1.888955e-07,1.888958e-07,1.888961e-07,1.888964e-07,1.888967e-07,1.888970e-07,1.888973e-07,1.888976e-07,1.888979e-07,1.888982e-07,1.888986e-07,1.888989e-07,1.888992e-07,1.888995e-07,1.888998e-07,1.889001e-07,1.889004e-07,1.889007e-07,1.889010e-07,1.889013e-07,1.889016e-07,1.889019e-07,1.889022e-07,1.889025e-07,1.889028e-07,1.889031e-07,1.889034e-07,1.889037e-07,1.889040e-07,1.889043e-07,1.889046e-07,1.889049e-07,1.889052e-07,1.889055e-07,1.889058e-07,1.889061e-07,1.889064e-07,1.889067e-07,1.889070e-07,1.889073e-07,1.889076e-07,1.889079e-07,1.889082e-07,1.889085e-07,1.889088e-07,1.889091e-07,1.889094e-07,1.889097e-07,1.889100e-07,1.889103e-07,1.889106e-07,1.889109e-07,1.889112e-07,1.889115e-07,1.889118e-07,1.889121e-07,1.889124e-07,1.889127e-07,1.889130e-07,1.889133e-07,1.889136e-07,1.889139e-07,1.889142e-07,1.889145e-07,1.889148e-07,1.889151e-07,1.889154e-07,1.889157e-07,1.889160e-07,1.889163e-07,1.889166e-07,1.889169e-07,1.889172e-07,1.889175e-07,1.889178e-07,1.889181e-07,1.889184e-07,1.889187e-07,1.889190e-07,1.889193e-07,1.889196e-07,1.889199e-07,1.889202e-07,1.889205e-07,1.889208e-07,1.889211e-07,1.889215e-07,1.889218e-07,1.889221e-07,1.889224e-07,1.889227e-07,1.889230e-07,1.889233e-07,1.889236e-07,1.889239e-07,1.889242e-07,1.889245e-07,1.889248e-07,1.889251e-07,1.889254e-07,1.889257e-07,1.889260e-07,1.889263e-07,1.889266e-07,1.889269e-07,1.889272e-07,1.889275e-07,1.889278e-07,1.889281e-07,1.889284e-07,1.889287e-07,1.889290e-07,1.889293e-07,1.889296e-07,1.889299e-07,1.889302e-07,1.889305e-07,1.889308e-07,1.889311e-07,1.889314e-07,1.889317e-07,1.889320e-07,1.889323e-07,1.889326e-07,1.889329e-07,1.889332e-07,1.889335e-07,1.889338e-07,1.889341e-07,1.889344e-07,1.889347e-07,1.889350e-07,1.889353e-07,1.889356e-07,1.889359e-07,1.889362e-07,1.889365e-07,1.889368e-07,1.889371e-07,1.889374e-07,1.889377e-07,1.889380e-07,1.889383e-07,1.889386e-07,1.889389e-07,1.889392e-07,1.889395e-07,1.889398e-07,1.889401e-07,1.889404e-07,1.889407e-07,1.889410e-07,1.889413e-07,1.889416e-07,1.889419e-07,1.889422e-07,1.889425e-07,1.889428e-07,1.889431e-07,1.889434e-07,1.889437e-07,1.889440e-07,1.889443e-07,1.889446e-07,1.889449e-07,1.889452e-07,1.889455e-07,1.889458e-07,1.889461e-07,1.889464e-07,1.889467e-07,1.889470e-07,1.889473e-07,1.889476e-07,1.889479e-07,1.889482e-07,1.889485e-07,1.889488e-07,1.889491e-07,1.889494e-07,1.889497e-07,1.889500e-07,1.889503e-07,1.889506e-07,1.889509e-07,1.889512e-07,1.889515e-07,1.889518e-07,1.889521e-07,1.889524e-07,1.889527e-07,1.889530e-07,1.889533e-07,1.889536e-07,1.889539e-07,1.889542e-07,1.889545e-07,1.889548e-07,1.889551e-07,1.889554e-07,1.889557e-07,1.889560e-07,1.889563e-07,1.889566e-07,1.889569e-07,1.889572e-07,1.889575e-07,1.889578e-07,1.889581e-07,1.889584e-07,1.889587e-07,1.889590e-07,1.889593e-07,1.889596e-07,1.889599e-07,1.889602e-07,1.889605e-07,1.889608e-07,1.889611e-07,1.889614e-07,1.889617e-07,1.889620e-07,1.889623e-07,1.889626e-07,1.889629e-07,1.889632e-07,1.889635e-07,1.889638e-07,1.889641e-07,1.889644e-07,1.889647e-07,1.889650e-07,1.889653e-07,1.889656e-07,1.889659e-07,1.889662e-07,1.889665e-07,1.889668e-07,1.889671e-07,1.889674e-07,1.889677e-07,1.889680e-07,1.889683e-07,1.889686e-07,1.889689e-07,1.889692e-07,1.889695e-07,1.889698e-07,1.889701e-07,1.889704e-07,1.889707e-07,1.889710e-07,1.889713e-07,1.889716e-07,1.889719e-07,1.889722e-07,1.889725e-07,1.889728e-07,1.889731e-07,1.889734e-07,1.889737e-07,1.889740e-07,1.889743e-07,1.889746e-07,1.889749e-07,1.889752e-07,1.889755e-07,1.889758e-07,1.889761e-07,1.889764e-07,1.889767e-07,1.889770e-07,1.889773e-07,1.889776e-07,1.889779e-07,1.889782e-07,1.889785e-07,1.889788e-07,1.889791e-07,1.889794e-07,1.889797e-07,1.889800e-07,1.889803e-07,1.889806e-07,1.889809e-07,1.889812e-07,1.889815e-07,1.889818e-07,1.889821e-07,1.889824e-07,1.889827e-07,1.889830e-07,1.889833e-07,1.889836e-07,1.889839e-07,1.889842e-07,1.889845e-07,1.889848e-07,1.889851e-07,1.889854e-07,1.889857e-07,1.889860e-07,1.889863e-07,1.889866e-07,1.889869e-07,1.889872e-07,1.889875e-07,1.889878e-07,1.889881e-07,1.889884e-07,1.889887e-07,1.889890e-07,1.889893e-07,1.889896e-07,1.889899e-07,1.889902e-07,1.889905e-07,1.889908e-07,1.889911e-07,1.889914e-07,1.889917e-07,1.889920e-07,1.889923e-07,1.889926e-07,1.889929e-07,1.889932e-07,1.889935e-07,1.889938e-07,1.889941e-07,1.889944e-07,1.889947e-07,1.889950e-07,1.889953e-07,1.889956e-07,1.889959e-07,1.889962e-07,1.889965e-07,1.889968e-07,1.889971e-07,1.889974e-07,1.889977e-07,1.889980e-07,1.889983e-07,1.889986e-07,1.889989e-07,1.889992e-07,1.889995e-07,1.889998e-07,1.890001e-07,1.890004e-07,1.890006e-07,1.890009e-07,1.890012e-07,1.890015e-07,1.890018e-07,1.890021e-07,1.890024e-07,1.890027e-07,1.890030e-07,1.890033e-07,1.890036e-07,1.890039e-07,1.890042e-07,1.890045e-07,1.890048e-07,1.890051e-07,1.890054e-07,1.890057e-07,1.890060e-07,1.890063e-07,1.890066e-07,1.890069e-07,1.890072e-07,1.890075e-07,1.890078e-07,1.890081e-07,1.890084e-07,1.890087e-07,1.890090e-07,1.890093e-07,1.890096e-07,1.890099e-07,1.890102e-07,1.890105e-07,1.890108e-07,1.890111e-07,1.890114e-07,1.890117e-07,1.890120e-07,1.890123e-07,1.890126e-07,1.890129e-07,1.890132e-07,1.890135e-07,1.890138e-07,1.890141e-07,1.890144e-07,1.890147e-07,1.890150e-07,1.890153e-07,1.890156e-07,1.890159e-07,1.890162e-07,1.890165e-07,1.890168e-07,1.890171e-07,1.890174e-07,1.890177e-07,1.890180e-07,1.890183e-07,1.890186e-07,1.890189e-07,1.890192e-07,1.890195e-07,1.890198e-07,1.890201e-07,1.890204e-07,1.890207e-07,1.890210e-07,1.890213e-07,1.890216e-07,1.890219e-07,1.890222e-07,1.890225e-07,1.890228e-07,1.890231e-07,1.890234e-07,1.890236e-07,1.890239e-07,1.890242e-07,1.890245e-07,1.890248e-07,1.890251e-07,1.890254e-07,1.890257e-07,1.890260e-07,1.890263e-07,1.890266e-07,1.890269e-07,1.890272e-07,1.890275e-07,1.890278e-07,1.890281e-07,1.890284e-07,1.890287e-07,1.890290e-07,1.890293e-07,1.890296e-07,1.890299e-07,1.890302e-07,1.890305e-07,1.890308e-07,1.890311e-07,1.890314e-07,1.890317e-07,1.890320e-07,1.890323e-07,1.890326e-07,1.890329e-07,1.890332e-07,1.890335e-07,1.890338e-07,1.890341e-07,1.890344e-07,1.890347e-07,1.890350e-07,1.890353e-07,1.890356e-07,1.890359e-07,1.890362e-07,1.890365e-07,1.890368e-07,1.890371e-07,1.890374e-07,1.890377e-07,1.890380e-07,1.890383e-07,1.890386e-07,1.890389e-07,1.890392e-07,1.890395e-07,1.890398e-07,1.890400e-07,1.890403e-07,1.890406e-07,1.890409e-07,1.890412e-07,1.890415e-07,1.890418e-07,1.890421e-07,1.890424e-07,1.890427e-07,1.890430e-07,1.890433e-07,1.890436e-07,1.890439e-07,1.890442e-07,1.890445e-07,1.890448e-07,1.890451e-07,1.890454e-07,1.890457e-07,1.890460e-07,1.890463e-07,1.890466e-07,1.890469e-07,1.890472e-07,1.890475e-07,1.890478e-07,1.890481e-07,1.890484e-07,1.890487e-07,1.890490e-07,1.890493e-07,1.890496e-07,1.890499e-07,1.890502e-07,1.890505e-07,1.890508e-07,1.890511e-07,1.890514e-07,1.890517e-07,1.890520e-07,1.890523e-07,1.890526e-07,1.890529e-07,1.890532e-07,1.890535e-07,1.890537e-07,1.890540e-07,1.890543e-07,1.890546e-07,1.890549e-07,1.890552e-07,1.890555e-07,1.890558e-07,1.890561e-07,1.890564e-07,1.890567e-07,1.890570e-07,1.890573e-07,1.890576e-07,1.890579e-07,1.890582e-07,1.890585e-07,1.890588e-07,1.890591e-07,1.890594e-07,1.890597e-07,1.890600e-07,1.890603e-07,1.890606e-07,1.890609e-07,1.890612e-07,1.890615e-07,1.890618e-07,1.890621e-07,1.890624e-07,1.890627e-07,1.890630e-07,1.890633e-07,1.890636e-07,1.890639e-07,1.890642e-07,1.890645e-07,1.890648e-07,1.890651e-07,1.890654e-07,1.890656e-07,1.890659e-07,1.890662e-07,1.890665e-07,1.890668e-07,1.890671e-07,1.890674e-07,1.890677e-07,1.890680e-07,1.890683e-07,1.890686e-07,1.890689e-07,1.890692e-07,1.890695e-07,1.890698e-07,1.890701e-07,1.890704e-07,1.890707e-07,1.890710e-07,1.890713e-07,1.890716e-07,1.890719e-07,1.890722e-07,1.890725e-07,1.890728e-07,1.890731e-07,1.890734e-07,1.890737e-07,1.890740e-07,1.890743e-07,1.890746e-07,1.890749e-07,1.890752e-07,1.890755e-07,1.890758e-07,1.890760e-07,1.890763e-07,1.890766e-07,1.890769e-07,1.890772e-07,1.890775e-07,1.890778e-07,1.890781e-07,1.890784e-07,1.890787e-07,1.890790e-07,1.890793e-07,1.890796e-07,1.890799e-07,1.890802e-07,1.890805e-07,1.890808e-07,1.890811e-07,1.890814e-07,1.890817e-07,1.890820e-07,1.890823e-07,1.890826e-07,1.890829e-07,1.890832e-07,1.890835e-07,1.890838e-07,1.890841e-07,1.890844e-07,1.890847e-07,1.890850e-07,1.890853e-07,1.890856e-07,1.890858e-07,1.890861e-07,1.890864e-07,1.890867e-07,1.890870e-07,1.890873e-07,1.890876e-07,1.890879e-07,1.890882e-07,1.890885e-07,1.890888e-07,1.890891e-07,1.890894e-07,1.890897e-07,1.890900e-07,1.890903e-07,1.890906e-07,1.890909e-07,1.890912e-07,1.890915e-07,1.890918e-07,1.890921e-07,1.890924e-07,1.890927e-07,1.890930e-07,1.890933e-07,1.890936e-07,1.890939e-07,1.890942e-07,1.890945e-07,1.890947e-07,1.890950e-07,1.890953e-07,1.890956e-07,1.890959e-07,1.890962e-07,1.890965e-07,1.890968e-07,1.890971e-07,1.890974e-07,1.890977e-07,1.890980e-07,1.890983e-07,1.890986e-07,1.890989e-07,1.890992e-07,1.890995e-07,1.890998e-07,1.891001e-07,1.891004e-07,1.891007e-07,1.891010e-07,1.891013e-07,1.891016e-07,1.891019e-07,1.891022e-07,1.891025e-07,1.891028e-07,1.891031e-07,1.891033e-07,1.891036e-07,1.891039e-07,1.891042e-07,1.891045e-07,1.891048e-07,1.891051e-07,1.891054e-07,1.891057e-07,1.891060e-07,1.891063e-07,1.891066e-07,1.891069e-07,1.891072e-07,1.891075e-07,1.891078e-07,1.891081e-07,1.891084e-07,1.891087e-07,1.891090e-07,1.891093e-07,1.891096e-07,1.891099e-07,1.891102e-07,1.891105e-07,1.891108e-07,1.891111e-07,1.891113e-07,1.891116e-07,1.891119e-07,1.891122e-07,1.891125e-07,1.891128e-07,1.891131e-07,1.891134e-07,1.891137e-07,1.891140e-07,1.891143e-07,1.891146e-07,1.891149e-07,1.891152e-07,1.891155e-07,1.891158e-07,1.891161e-07,1.891164e-07,1.891167e-07,1.891170e-07,1.891173e-07,1.891176e-07,1.891179e-07,1.891182e-07,1.891185e-07,1.891187e-07,1.891190e-07,1.891193e-07,1.891196e-07,1.891199e-07,1.891202e-07,1.891205e-07,1.891208e-07,1.891211e-07,1.891214e-07,1.891217e-07,1.891220e-07,1.891223e-07,1.891226e-07,1.891229e-07,1.891232e-07,1.891235e-07,1.891238e-07,1.891241e-07,1.891244e-07,1.891247e-07,1.891250e-07,1.891253e-07,1.891256e-07,1.891258e-07,1.891261e-07,1.891264e-07,1.891267e-07,1.891270e-07,1.891273e-07,1.891276e-07,1.891279e-07,1.891282e-07,1.891285e-07,1.891288e-07,1.891291e-07,1.891294e-07,1.891297e-07,1.891300e-07,1.891303e-07,1.891306e-07,1.891309e-07,1.891312e-07,1.891315e-07,1.891318e-07,1.891321e-07,1.891324e-07,1.891327e-07,1.891329e-07,1.891332e-07,1.891335e-07,1.891338e-07,1.891341e-07,1.891344e-07,1.891347e-07,1.891350e-07,1.891353e-07,1.891356e-07,1.891359e-07,1.891362e-07,1.891365e-07,1.891368e-07,1.891371e-07,1.891374e-07,1.891377e-07,1.891380e-07,1.891383e-07,1.891386e-07,1.891389e-07,1.891392e-07,1.891394e-07,1.891397e-07,1.891400e-07,1.891403e-07,1.891406e-07,1.891409e-07,1.891412e-07,1.891415e-07,1.891418e-07,1.891421e-07,1.891424e-07,1.891427e-07,1.891430e-07,1.891433e-07,1.891436e-07,1.891439e-07,1.891442e-07,1.891445e-07,1.891448e-07,1.891451e-07,1.891454e-07,1.891457e-07,1.891459e-07,1.891462e-07,1.891465e-07,1.891468e-07,1.891471e-07,1.891474e-07,1.891477e-07,1.891480e-07,1.891483e-07,1.891486e-07,1.891489e-07,1.891492e-07,1.891495e-07,1.891498e-07,1.891501e-07,1.891504e-07,1.891507e-07,1.891510e-07,1.891513e-07,1.891516e-07,1.891519e-07,1.891521e-07,1.891524e-07,1.891527e-07,1.891530e-07,1.891533e-07,1.891536e-07,1.891539e-07,1.891542e-07,1.891545e-07,1.891548e-07,1.891551e-07,1.891554e-07,1.891557e-07,1.891560e-07,1.891563e-07,1.891566e-07,1.891569e-07,1.891572e-07,1.891575e-07,1.891578e-07,1.891580e-07,1.891583e-07,1.891586e-07,1.891589e-07,1.891592e-07,1.891595e-07,1.891598e-07,1.891601e-07,1.891604e-07,1.891607e-07,1.891610e-07,1.891613e-07,1.891616e-07,1.891619e-07,1.891622e-07,1.891625e-07,1.891628e-07,1.891631e-07,1.891634e-07,1.891637e-07,1.891639e-07,1.891642e-07,1.891645e-07,1.891648e-07,1.891651e-07,1.891654e-07,1.891657e-07,1.891660e-07,1.891663e-07,1.891666e-07,1.891669e-07,1.891672e-07,1.891675e-07,1.891678e-07,1.891681e-07,1.891684e-07,1.891687e-07,1.891690e-07,1.891693e-07,1.891695e-07,1.891698e-07,1.891701e-07,1.891704e-07,1.891707e-07,1.891710e-07,1.891713e-07,1.891716e-07,1.891719e-07,1.891722e-07,1.891725e-07,1.891728e-07,1.891731e-07,1.891734e-07,1.891737e-07,1.891740e-07,1.891743e-07,1.891746e-07,1.891748e-07,1.891751e-07,1.891754e-07,1.891757e-07,1.891760e-07,1.891763e-07,1.891766e-07,1.891769e-07,1.891772e-07,1.891775e-07,1.891778e-07,1.891781e-07,1.891784e-07,1.891787e-07,1.891790e-07,1.891793e-07,1.891796e-07,1.891799e-07,1.891802e-07,1.891804e-07,1.891807e-07,1.891810e-07,1.891813e-07,1.891816e-07,1.891819e-07,1.891822e-07,1.891825e-07,1.891828e-07,1.891831e-07,1.891834e-07,1.891837e-07,1.891840e-07,1.891843e-07,1.891846e-07,1.891849e-07,1.891852e-07,1.891854e-07,1.891857e-07,1.891860e-07,1.891863e-07,1.891866e-07,1.891869e-07,1.891872e-07,1.891875e-07,1.891878e-07,1.891881e-07,1.891884e-07,1.891887e-07,1.891890e-07,1.891893e-07,1.891896e-07,1.891899e-07,1.891902e-07,1.891905e-07,1.891907e-07,1.891910e-07,1.891913e-07,1.891916e-07,1.891919e-07,1.891922e-07,1.891925e-07,1.891928e-07,1.891931e-07,1.891934e-07,1.891937e-07,1.891940e-07,1.891943e-07,1.891946e-07,1.891949e-07,1.891952e-07,1.891955e-07,1.891957e-07,1.891960e-07,1.891963e-07,1.891966e-07,1.891969e-07,1.891972e-07,1.891975e-07,1.891978e-07,1.891981e-07,1.891984e-07,1.891987e-07,1.891990e-07,1.891993e-07,1.891996e-07,1.891999e-07,1.892002e-07,1.892004e-07,1.892007e-07,1.892010e-07,1.892013e-07,1.892016e-07,1.892019e-07,1.892022e-07,1.892025e-07,1.892028e-07,1.892031e-07,1.892034e-07,1.892037e-07,1.892040e-07,1.892043e-07,1.892046e-07,1.892049e-07,1.892051e-07,1.892054e-07,1.892057e-07,1.892060e-07,1.892063e-07,1.892066e-07,1.892069e-07,1.892072e-07,1.892075e-07,1.892078e-07,1.892081e-07,1.892084e-07,1.892087e-07,1.892090e-07,1.892093e-07,1.892096e-07,1.892098e-07,1.892101e-07,1.892104e-07,1.892107e-07,1.892110e-07,1.892113e-07,1.892116e-07,1.892119e-07,1.892122e-07,1.892125e-07,1.892128e-07,1.892131e-07,1.892134e-07,1.892137e-07,1.892140e-07,1.892143e-07,1.892145e-07,1.892148e-07,1.892151e-07,1.892154e-07,1.892157e-07,1.892160e-07,1.892163e-07,1.892166e-07,1.892169e-07,1.892172e-07,1.892175e-07,1.892178e-07,1.892181e-07,1.892184e-07,1.892187e-07,1.892190e-07,1.892192e-07,1.892195e-07,1.892198e-07,1.892201e-07,1.892204e-07,1.892207e-07,1.892210e-07,1.892213e-07,1.892216e-07,1.892219e-07,1.892222e-07,1.892225e-07,1.892228e-07,1.892231e-07,1.892234e-07,1.892236e-07,1.892239e-07,1.892242e-07,1.892245e-07,1.892248e-07,1.892251e-07,1.892254e-07,1.892257e-07,1.892260e-07,1.892263e-07,1.892266e-07,1.892269e-07,1.892272e-07,1.892275e-07,1.892278e-07,1.892280e-07,1.892283e-07,1.892286e-07,1.892289e-07,1.892292e-07,1.892295e-07,1.892298e-07,1.892301e-07,1.892304e-07,1.892307e-07,1.892310e-07,1.892313e-07,1.892316e-07,1.892319e-07,1.892321e-07,1.892324e-07,1.892327e-07,1.892330e-07,1.892333e-07,1.892336e-07,1.892339e-07,1.892342e-07,1.892345e-07,1.892348e-07,1.892351e-07,1.892354e-07,1.892357e-07,1.892360e-07,1.892363e-07,1.892365e-07,1.892368e-07,1.892371e-07,1.892374e-07,1.892377e-07,1.892380e-07,1.892383e-07,1.892386e-07,1.892389e-07,1.892392e-07,1.892395e-07,1.892398e-07,1.892401e-07,1.892404e-07,1.892406e-07,1.892409e-07,1.892412e-07,1.892415e-07,1.892418e-07,1.892421e-07,1.892424e-07,1.892427e-07,1.892430e-07,1.892433e-07,1.892436e-07,1.892439e-07,1.892442e-07,1.892445e-07,1.892447e-07,1.892450e-07,1.892453e-07,1.892456e-07,1.892459e-07,1.892462e-07,1.892465e-07,1.892468e-07,1.892471e-07,1.892474e-07,1.892477e-07,1.892480e-07,1.892483e-07,1.892486e-07,1.892488e-07,1.892491e-07,1.892494e-07,1.892497e-07,1.892500e-07,1.892503e-07,1.892506e-07,1.892509e-07,1.892512e-07,1.892515e-07,1.892518e-07,1.892521e-07,1.892524e-07,1.892526e-07,1.892529e-07,1.892532e-07,1.892535e-07,1.892538e-07,1.892541e-07,1.892544e-07,1.892547e-07,1.892550e-07,1.892553e-07,1.892556e-07,1.892559e-07,1.892562e-07,1.892565e-07,1.892567e-07,1.892570e-07,1.892573e-07,1.892576e-07,1.892579e-07,1.892582e-07,1.892585e-07,1.892588e-07,1.892591e-07,1.892594e-07,1.892597e-07,1.892600e-07,1.892603e-07,1.892605e-07,1.892608e-07,1.892611e-07,1.892614e-07,1.892617e-07,1.892620e-07,1.892623e-07,1.892626e-07,1.892629e-07,1.892632e-07,1.892635e-07,1.892638e-07,1.892641e-07,1.892643e-07,1.892646e-07,1.892649e-07,1.892652e-07,1.892655e-07,1.892658e-07,1.892661e-07,1.892664e-07,1.892667e-07,1.892670e-07,1.892673e-07,1.892676e-07,1.892679e-07,1.892681e-07,1.892684e-07,1.892687e-07,1.892690e-07,1.892693e-07,1.892696e-07,1.892699e-07,1.892702e-07,1.892705e-07,1.892708e-07,1.892711e-07,1.892714e-07,1.892717e-07,1.892719e-07,1.892722e-07,1.892725e-07,1.892728e-07,1.892731e-07,1.892734e-07,1.892737e-07,1.892740e-07,1.892743e-07,1.892746e-07,1.892749e-07,1.892752e-07,1.892754e-07,1.892757e-07,1.892760e-07,1.892763e-07,1.892766e-07,1.892769e-07,1.892772e-07,1.892775e-07,1.892778e-07,1.892781e-07,1.892784e-07,1.892787e-07,1.892790e-07,1.892792e-07,1.892795e-07,1.892798e-07,1.892801e-07,1.892804e-07,1.892807e-07,1.892810e-07,1.892813e-07,1.892816e-07,1.892819e-07,1.892822e-07,1.892825e-07,1.892827e-07,1.892830e-07,1.892833e-07,1.892836e-07,1.892839e-07,1.892842e-07,1.892845e-07,1.892848e-07,1.892851e-07,1.892854e-07,1.892857e-07,1.892860e-07,1.892863e-07,1.892865e-07,1.892868e-07,1.892871e-07,1.892874e-07,1.892877e-07,1.892880e-07,1.892883e-07,1.892886e-07,1.892889e-07,1.892892e-07,1.892895e-07,1.892898e-07,1.892900e-07,1.892903e-07,1.892906e-07,1.892909e-07,1.892912e-07,1.892915e-07,1.892918e-07,1.892921e-07,1.892924e-07,1.892927e-07,1.892930e-07,1.892933e-07,1.892935e-07,1.892938e-07,1.892941e-07,1.892944e-07,1.892947e-07,1.892950e-07,1.892953e-07,1.892956e-07,1.892959e-07,1.892962e-07,1.892965e-07,1.892967e-07,1.892970e-07,1.892973e-07,1.892976e-07,1.892979e-07,1.892982e-07,1.892985e-07,1.892988e-07,1.892991e-07,1.892994e-07,1.892997e-07,1.893000e-07,1.893002e-07,1.893005e-07,1.893008e-07,1.893011e-07,1.893014e-07,1.893017e-07,1.893020e-07,1.893023e-07,1.893026e-07,1.893029e-07,1.893032e-07,1.893035e-07,1.893037e-07,1.893040e-07,1.893043e-07,1.893046e-07,1.893049e-07,1.893052e-07,1.893055e-07,1.893058e-07,1.893061e-07,1.893064e-07,1.893067e-07,1.893069e-07,1.893072e-07,1.893075e-07,1.893078e-07,1.893081e-07,1.893084e-07,1.893087e-07,1.893090e-07,1.893093e-07,1.893096e-07,1.893099e-07,1.893102e-07,1.893104e-07,1.893107e-07,1.893110e-07,1.893113e-07,1.893116e-07,1.893119e-07,1.893122e-07,1.893125e-07,1.893128e-07,1.893131e-07,1.893134e-07,1.893136e-07,1.893139e-07,1.893142e-07,1.893145e-07,1.893148e-07,1.893151e-07,1.893154e-07,1.893157e-07,1.893160e-07,1.893163e-07,1.893166e-07,1.893168e-07,1.893171e-07,1.893174e-07,1.893177e-07,1.893180e-07,1.893183e-07,1.893186e-07,1.893189e-07,1.893192e-07,1.893195e-07,1.893198e-07,1.893200e-07,1.893203e-07,1.893206e-07,1.893209e-07,1.893212e-07,1.893215e-07,1.893218e-07,1.893221e-07,1.893224e-07,1.893227e-07,1.893230e-07,1.893232e-07,1.893235e-07,1.893238e-07,1.893241e-07,1.893244e-07,1.893247e-07,1.893250e-07,1.893253e-07,1.893256e-07,1.893259e-07,1.893262e-07,1.893264e-07,1.893267e-07,1.893270e-07,1.893273e-07,1.893276e-07,1.893279e-07,1.893282e-07,1.893285e-07,1.893288e-07,1.893291e-07,1.893294e-07,1.893296e-07,1.893299e-07,1.893302e-07,1.893305e-07,1.893308e-07,1.893311e-07,1.893314e-07,1.893317e-07,1.893320e-07,1.893323e-07,1.893325e-07,1.893328e-07,1.893331e-07,1.893334e-07,1.893337e-07,1.893340e-07,1.893343e-07,1.893346e-07,1.893349e-07,1.893352e-07,1.893355e-07,1.893357e-07,1.893360e-07,1.893363e-07,1.893366e-07,1.893369e-07,1.893372e-07,1.893375e-07,1.893378e-07,1.893381e-07,1.893384e-07,1.893387e-07,1.893389e-07,1.893392e-07,1.893395e-07,1.893398e-07,1.893401e-07,1.893404e-07,1.893407e-07,1.893410e-07,1.893413e-07,1.893416e-07,1.893418e-07,1.893421e-07,1.893424e-07,1.893427e-07,1.893430e-07,1.893433e-07,1.893436e-07,1.893439e-07,1.893442e-07,1.893445e-07,1.893447e-07,1.893450e-07,1.893453e-07,1.893456e-07,1.893459e-07,1.893462e-07,1.893465e-07,1.893468e-07,1.893471e-07,1.893474e-07,1.893477e-07,1.893479e-07,1.893482e-07,1.893485e-07,1.893488e-07,1.893491e-07,1.893494e-07,1.893497e-07,1.893500e-07,1.893503e-07,1.893506e-07,1.893508e-07,1.893511e-07,1.893514e-07,1.893517e-07,1.893520e-07,1.893523e-07,1.893526e-07,1.893529e-07,1.893532e-07,1.893535e-07,1.893537e-07,1.893540e-07,1.893543e-07,1.893546e-07,1.893549e-07,1.893552e-07,1.893555e-07,1.893558e-07,1.893561e-07,1.893564e-07,1.893566e-07,1.893569e-07,1.893572e-07,1.893575e-07,1.893578e-07,1.893581e-07,1.893584e-07,1.893587e-07,1.893590e-07,1.893593e-07,1.893595e-07,1.893598e-07,1.893601e-07,1.893604e-07,1.893607e-07,1.893610e-07,1.893613e-07,1.893616e-07,1.893619e-07,1.893622e-07,1.893624e-07,1.893627e-07,1.893630e-07,1.893633e-07,1.893636e-07,1.893639e-07,1.893642e-07,1.893645e-07,1.893648e-07,1.893651e-07,1.893653e-07,1.893656e-07,1.893659e-07,1.893662e-07,1.893665e-07,1.893668e-07,1.893671e-07,1.893674e-07,1.893677e-07,1.893680e-07,1.893682e-07,1.893685e-07,1.893688e-07,1.893691e-07,1.893694e-07,1.893697e-07,1.893700e-07,1.893703e-07,1.893706e-07,1.893708e-07,1.893711e-07,1.893714e-07,1.893717e-07,1.893720e-07,1.893723e-07,1.893726e-07,1.893729e-07,1.893732e-07,1.893735e-07,1.893737e-07,1.893740e-07,1.893743e-07,1.893746e-07,1.893749e-07,1.893752e-07,1.893755e-07,1.893758e-07,1.893761e-07,1.893764e-07,1.893766e-07,1.893769e-07,1.893772e-07,1.893775e-07,1.893778e-07,1.893781e-07,1.893784e-07,1.893787e-07,1.893790e-07,1.893792e-07,1.893795e-07,1.893798e-07,1.893801e-07,1.893804e-07,1.893807e-07,1.893810e-07,1.893813e-07,1.893816e-07,1.893818e-07,1.893821e-07,1.893824e-07,1.893827e-07,1.893830e-07,1.893833e-07,1.893836e-07,1.893839e-07,1.893842e-07,1.893845e-07,1.893847e-07,1.893850e-07,1.893853e-07,1.893856e-07,1.893859e-07,1.893862e-07,1.893865e-07,1.893868e-07,1.893871e-07,1.893873e-07,1.893876e-07,1.893879e-07,1.893882e-07,1.893885e-07,1.893888e-07,1.893891e-07,1.893894e-07,1.893897e-07,1.893900e-07,1.893902e-07,1.893905e-07,1.893908e-07,1.893911e-07,1.893914e-07,1.893917e-07,1.893920e-07,1.893923e-07,1.893926e-07,1.893928e-07,1.893931e-07,1.893934e-07,1.893937e-07,1.893940e-07,1.893943e-07,1.893946e-07,1.893949e-07,1.893952e-07,1.893954e-07,1.893957e-07,1.893960e-07,1.893963e-07,1.893966e-07,1.893969e-07,1.893972e-07,1.893975e-07,1.893978e-07,1.893980e-07,1.893983e-07,1.893986e-07,1.893989e-07,1.893992e-07,1.893995e-07,1.893998e-07,1.894001e-07,1.894004e-07,1.894006e-07,1.894009e-07,1.894012e-07,1.894015e-07,1.894018e-07,1.894021e-07,1.894024e-07,1.894027e-07,1.894030e-07,1.894032e-07,1.894035e-07,1.894038e-07,1.894041e-07,1.894044e-07,1.894047e-07,1.894050e-07,1.894053e-07,1.894056e-07,1.894058e-07,1.894061e-07,1.894064e-07,1.894067e-07,1.894070e-07,1.894073e-07,1.894076e-07,1.894079e-07,1.894082e-07,1.894084e-07,1.894087e-07,1.894090e-07,1.894093e-07,1.894096e-07,1.894099e-07,1.894102e-07,1.894105e-07,1.894108e-07,1.894110e-07,1.894113e-07,1.894116e-07,1.894119e-07,1.894122e-07,1.894125e-07,1.894128e-07,1.894131e-07,1.894134e-07,1.894136e-07,1.894139e-07,1.894142e-07,1.894145e-07,1.894148e-07,1.894151e-07,1.894154e-07,1.894157e-07,1.894159e-07,1.894162e-07,1.894165e-07,1.894168e-07,1.894171e-07,1.894174e-07,1.894177e-07,1.894180e-07,1.894183e-07,1.894185e-07,1.894188e-07,1.894191e-07,1.894194e-07,1.894197e-07,1.894200e-07,1.894203e-07,1.894206e-07,1.894209e-07,1.894211e-07,1.894214e-07,1.894217e-07,1.894220e-07,1.894223e-07,1.894226e-07,1.894229e-07,1.894232e-07,1.894234e-07,1.894237e-07,1.894240e-07,1.894243e-07,1.894246e-07,1.894249e-07,1.894252e-07,1.894255e-07,1.894258e-07,1.894260e-07,1.894263e-07,1.894266e-07,1.894269e-07,1.894272e-07,1.894275e-07,1.894278e-07,1.894281e-07,1.894283e-07,1.894286e-07,1.894289e-07,1.894292e-07,1.894295e-07,1.894298e-07,1.894301e-07,1.894304e-07,1.894307e-07,1.894309e-07,1.894312e-07,1.894315e-07,1.894318e-07,1.894321e-07,1.894324e-07,1.894327e-07,1.894330e-07,1.894332e-07,1.894335e-07,1.894338e-07,1.894341e-07,1.894344e-07,1.894347e-07,1.894350e-07,1.894353e-07,1.894356e-07,1.894358e-07,1.894361e-07,1.894364e-07,1.894367e-07,1.894370e-07,1.894373e-07,1.894376e-07,1.894379e-07,1.894381e-07,1.894384e-07,1.894387e-07,1.894390e-07,1.894393e-07,1.894396e-07,1.894399e-07,1.894402e-07,1.894404e-07,1.894407e-07,1.894410e-07,1.894413e-07,1.894416e-07,1.894419e-07,1.894422e-07,1.894425e-07,1.894428e-07,1.894430e-07,1.894433e-07,1.894436e-07,1.894439e-07,1.894442e-07,1.894445e-07,1.894448e-07,1.894451e-07,1.894453e-07,1.894456e-07,1.894459e-07,1.894462e-07,1.894465e-07,1.894468e-07,1.894471e-07,1.894474e-07,1.894476e-07,1.894479e-07,1.894482e-07,1.894485e-07,1.894488e-07,1.894491e-07,1.894494e-07,1.894497e-07,1.894499e-07,1.894502e-07,1.894505e-07,1.894508e-07,1.894511e-07,1.894514e-07,1.894517e-07,1.894520e-07,1.894522e-07,1.894525e-07,1.894528e-07,1.894531e-07,1.894534e-07,1.894537e-07,1.894540e-07,1.894543e-07,1.894546e-07,1.894548e-07,1.894551e-07,1.894554e-07,1.894557e-07,1.894560e-07,1.894563e-07,1.894566e-07,1.894569e-07,1.894571e-07,1.894574e-07,1.894577e-07,1.894580e-07,1.894583e-07,1.894586e-07,1.894589e-07,1.894592e-07,1.894594e-07,1.894597e-07,1.894600e-07,1.894603e-07,1.894606e-07,1.894609e-07,1.894612e-07,1.894615e-07,1.894617e-07,1.894620e-07,1.894623e-07,1.894626e-07,1.894629e-07,1.894632e-07,1.894635e-07,1.894637e-07,1.894640e-07,1.894643e-07,1.894646e-07,1.894649e-07,1.894652e-07,1.894655e-07,1.894658e-07,1.894660e-07,1.894663e-07,1.894666e-07,1.894669e-07,1.894672e-07,1.894675e-07,1.894678e-07,1.894681e-07,1.894683e-07,1.894686e-07,1.894689e-07,1.894692e-07,1.894695e-07,1.894698e-07,1.894701e-07,1.894704e-07,1.894706e-07,1.894709e-07,1.894712e-07,1.894715e-07,1.894718e-07,1.894721e-07,1.894724e-07,1.894727e-07,1.894729e-07,1.894732e-07,1.894735e-07,1.894738e-07,1.894741e-07,1.894744e-07,1.894747e-07,1.894750e-07,1.894752e-07,1.894755e-07,1.894758e-07,1.894761e-07,1.894764e-07,1.894767e-07,1.894770e-07,1.894772e-07,1.894775e-07,1.894778e-07,1.894781e-07,1.894784e-07,1.894787e-07,1.894790e-07,1.894793e-07,1.894795e-07,1.894798e-07,1.894801e-07,1.894804e-07,1.894807e-07,1.894810e-07,1.894813e-07,1.894816e-07,1.894818e-07,1.894821e-07,1.894824e-07,1.894827e-07,1.894830e-07,1.894833e-07,1.894836e-07,1.894838e-07,1.894841e-07,1.894844e-07,1.894847e-07,1.894850e-07,1.894853e-07,1.894856e-07,1.894859e-07,1.894861e-07,1.894864e-07,1.894867e-07,1.894870e-07,1.894873e-07,1.894876e-07,1.894879e-07,1.894882e-07,1.894884e-07,1.894887e-07,1.894890e-07,1.894893e-07,1.894896e-07,1.894899e-07,1.894902e-07,1.894904e-07,1.894907e-07,1.894910e-07,1.894913e-07,1.894916e-07,1.894919e-07,1.894922e-07,1.894925e-07,1.894927e-07,1.894930e-07,1.894933e-07,1.894936e-07,1.894939e-07,1.894942e-07,1.894945e-07,1.894947e-07,1.894950e-07,1.894953e-07,1.894956e-07,1.894959e-07,1.894962e-07,1.894965e-07,1.894968e-07,1.894970e-07,1.894973e-07,1.894976e-07,1.894979e-07,1.894982e-07,1.894985e-07,1.894988e-07,1.894990e-07,1.894993e-07,1.894996e-07,1.894999e-07,1.895002e-07,1.895005e-07,1.895008e-07,1.895010e-07,1.895013e-07,1.895016e-07,1.895019e-07,1.895022e-07,1.895025e-07,1.895028e-07,1.895031e-07,1.895033e-07,1.895036e-07,1.895039e-07,1.895042e-07,1.895045e-07,1.895048e-07,1.895051e-07,1.895053e-07,1.895056e-07,1.895059e-07,1.895062e-07,1.895065e-07,1.895068e-07,1.895071e-07,1.895073e-07,1.895076e-07,1.895079e-07,1.895082e-07,1.895085e-07,1.895088e-07,1.895091e-07,1.895094e-07,1.895096e-07,1.895099e-07,1.895102e-07,1.895105e-07,1.895108e-07,1.895111e-07,1.895114e-07,1.895116e-07,1.895119e-07,1.895122e-07,1.895125e-07,1.895128e-07,1.895131e-07,1.895134e-07,1.895136e-07,1.895139e-07,1.895142e-07,1.895145e-07,1.895148e-07,1.895151e-07,1.895154e-07,1.895156e-07,1.895159e-07,1.895162e-07,1.895165e-07,1.895168e-07,1.895171e-07,1.895174e-07,1.895177e-07,1.895179e-07,1.895182e-07,1.895185e-07,1.895188e-07,1.895191e-07,1.895194e-07,1.895197e-07,1.895199e-07,1.895202e-07,1.895205e-07,1.895208e-07,1.895211e-07,1.895214e-07,1.895217e-07,1.895219e-07,1.895222e-07,1.895225e-07,1.895228e-07,1.895231e-07,1.895234e-07,1.895237e-07,1.895239e-07,1.895242e-07,1.895245e-07,1.895248e-07,1.895251e-07,1.895254e-07,1.895257e-07,1.895259e-07,1.895262e-07,1.895265e-07,1.895268e-07,1.895271e-07,1.895274e-07,1.895277e-07,1.895279e-07,1.895282e-07,1.895285e-07,1.895288e-07,1.895291e-07,1.895294e-07,1.895297e-07,1.895299e-07,1.895302e-07,1.895305e-07,1.895308e-07,1.895311e-07,1.895314e-07,1.895317e-07,1.895319e-07,1.895322e-07,1.895325e-07,1.895328e-07,1.895331e-07,1.895334e-07,1.895337e-07,1.895339e-07,1.895342e-07,1.895345e-07,1.895348e-07,1.895351e-07,1.895354e-07,1.895357e-07,1.895359e-07,1.895362e-07,1.895365e-07,1.895368e-07,1.895371e-07,1.895374e-07,1.895377e-07,1.895379e-07,1.895382e-07,1.895385e-07,1.895388e-07,1.895391e-07,1.895394e-07,1.895397e-07,1.895399e-07,1.895402e-07,1.895405e-07,1.895408e-07,1.895411e-07,1.895414e-07,1.895417e-07,1.895419e-07,1.895422e-07,1.895425e-07,1.895428e-07,1.895431e-07,1.895434e-07,1.895437e-07,1.895439e-07,1.895442e-07,1.895445e-07,1.895448e-07,1.895451e-07,1.895454e-07,1.895457e-07,1.895459e-07,1.895462e-07,1.895465e-07,1.895468e-07,1.895471e-07,1.895474e-07,1.895476e-07,1.895479e-07,1.895482e-07,1.895485e-07,1.895488e-07,1.895491e-07,1.895494e-07,1.895496e-07,1.895499e-07,1.895502e-07,1.895505e-07,1.895508e-07,1.895511e-07,1.895514e-07,1.895516e-07,1.895519e-07,1.895522e-07,1.895525e-07,1.895528e-07,1.895531e-07,1.895534e-07,1.895536e-07,1.895539e-07,1.895542e-07,1.895545e-07,1.895548e-07,1.895551e-07,1.895553e-07,1.895556e-07,1.895559e-07,1.895562e-07,1.895565e-07,1.895568e-07,1.895571e-07,1.895573e-07,1.895576e-07,1.895579e-07,1.895582e-07,1.895585e-07,1.895588e-07,1.895591e-07,1.895593e-07,1.895596e-07,1.895599e-07,1.895602e-07,1.895605e-07,1.895608e-07,1.895610e-07,1.895613e-07,1.895616e-07,1.895619e-07,1.895622e-07,1.895625e-07,1.895628e-07,1.895630e-07,1.895633e-07,1.895636e-07,1.895639e-07,1.895642e-07,1.895645e-07,1.895648e-07,1.895650e-07,1.895653e-07,1.895656e-07,1.895659e-07,1.895662e-07,1.895665e-07,1.895667e-07,1.895670e-07,1.895673e-07,1.895676e-07,1.895679e-07,1.895682e-07,1.895685e-07,1.895687e-07,1.895690e-07,1.895693e-07,1.895696e-07,1.895699e-07,1.895702e-07,1.895705e-07,1.895707e-07,1.895710e-07,1.895713e-07,1.895716e-07,1.895719e-07,1.895722e-07,1.895724e-07,1.895727e-07,1.895730e-07,1.895733e-07,1.895736e-07,1.895739e-07,1.895742e-07,1.895744e-07,1.895747e-07,1.895750e-07,1.895753e-07,1.895756e-07,1.895759e-07,1.895761e-07,1.895764e-07,1.895767e-07,1.895770e-07,1.895773e-07,1.895776e-07,1.895779e-07,1.895781e-07,1.895784e-07,1.895787e-07,1.895790e-07,1.895793e-07,1.895796e-07,1.895798e-07,1.895801e-07,1.895804e-07,1.895807e-07,1.895810e-07,1.895813e-07,1.895816e-07,1.895818e-07,1.895821e-07,1.895824e-07,1.895827e-07,1.895830e-07,1.895833e-07,1.895835e-07,1.895838e-07,1.895841e-07,1.895844e-07,1.895847e-07,1.895850e-07,1.895852e-07,1.895855e-07,1.895858e-07,1.895861e-07,1.895864e-07,1.895867e-07,1.895870e-07,1.895872e-07,1.895875e-07,1.895878e-07,1.895881e-07,1.895884e-07,1.895887e-07,1.895889e-07,1.895892e-07,1.895895e-07,1.895898e-07,1.895901e-07,1.895904e-07,1.895907e-07,1.895909e-07,1.895912e-07,1.895915e-07,1.895918e-07,1.895921e-07,1.895924e-07,1.895926e-07,1.895929e-07,1.895932e-07,1.895935e-07,1.895938e-07,1.895941e-07,1.895943e-07,1.895946e-07,1.895949e-07,1.895952e-07,1.895955e-07,1.895958e-07,1.895961e-07,1.895963e-07,1.895966e-07,1.895969e-07,1.895972e-07,1.895975e-07,1.895978e-07,1.895980e-07,1.895983e-07,1.895986e-07,1.895989e-07,1.895992e-07,1.895995e-07,1.895997e-07,1.896000e-07,1.896003e-07,1.896006e-07,1.896009e-07,1.896012e-07,1.896014e-07,1.896017e-07,1.896020e-07,1.896023e-07,1.896026e-07,1.896029e-07,1.896032e-07,1.896034e-07,1.896037e-07,1.896040e-07,1.896043e-07,1.896046e-07,1.896049e-07,1.896051e-07,1.896054e-07,1.896057e-07,1.896060e-07,1.896063e-07,1.896066e-07,1.896068e-07,1.896071e-07,1.896074e-07,1.896077e-07,1.896080e-07,1.896083e-07,1.896085e-07,1.896088e-07,1.896091e-07,1.896094e-07,1.896097e-07,1.896100e-07,1.896102e-07,1.896105e-07,1.896108e-07,1.896111e-07,1.896114e-07,1.896117e-07,1.896120e-07,1.896122e-07,1.896125e-07,1.896128e-07,1.896131e-07,1.896134e-07,1.896137e-07,1.896139e-07,1.896142e-07,1.896145e-07,1.896148e-07,1.896151e-07,1.896154e-07,1.896156e-07,1.896159e-07,1.896162e-07,1.896165e-07,1.896168e-07,1.896171e-07,1.896173e-07,1.896176e-07,1.896179e-07,1.896182e-07,1.896185e-07,1.896188e-07,1.896190e-07,1.896193e-07,1.896196e-07,1.896199e-07,1.896202e-07,1.896205e-07,1.896207e-07,1.896210e-07,1.896213e-07,1.896216e-07,1.896219e-07,1.896222e-07,1.896224e-07,1.896227e-07,1.896230e-07,1.896233e-07,1.896236e-07,1.896239e-07,1.896241e-07,1.896244e-07,1.896247e-07,1.896250e-07,1.896253e-07,1.896256e-07,1.896258e-07,1.896261e-07,1.896264e-07,1.896267e-07,1.896270e-07,1.896273e-07,1.896275e-07,1.896278e-07,1.896281e-07,1.896284e-07,1.896287e-07,1.896290e-07,1.896292e-07,1.896295e-07,1.896298e-07,1.896301e-07,1.896304e-07,1.896307e-07,1.896309e-07,1.896312e-07,1.896315e-07,1.896318e-07,1.896321e-07,1.896324e-07,1.896326e-07,1.896329e-07,1.896332e-07,1.896335e-07,1.896338e-07,1.896341e-07,1.896343e-07,1.896346e-07,1.896349e-07,1.896352e-07,1.896355e-07,1.896358e-07,1.896360e-07,1.896363e-07,1.896366e-07,1.896369e-07,1.896372e-07,1.896375e-07,1.896377e-07,1.896380e-07,1.896383e-07,1.896386e-07,1.896389e-07,1.896392e-07,1.896394e-07,1.896397e-07,1.896400e-07,1.896403e-07,1.896406e-07,1.896409e-07,1.896411e-07,1.896414e-07,1.896417e-07,1.896420e-07,1.896423e-07,1.896426e-07,1.896428e-07,1.896431e-07,1.896434e-07,1.896437e-07,1.896440e-07,1.896443e-07,1.896445e-07,1.896448e-07,1.896451e-07,1.896454e-07,1.896457e-07,1.896460e-07,1.896462e-07,1.896465e-07,1.896468e-07,1.896471e-07,1.896474e-07,1.896476e-07,1.896479e-07,1.896482e-07,1.896485e-07,1.896488e-07,1.896491e-07,1.896493e-07,1.896496e-07,1.896499e-07,1.896502e-07,1.896505e-07,1.896508e-07,1.896510e-07,1.896513e-07,1.896516e-07,1.896519e-07,1.896522e-07,1.896525e-07,1.896527e-07,1.896530e-07,1.896533e-07,1.896536e-07,1.896539e-07,1.896542e-07,1.896544e-07,1.896547e-07,1.896550e-07,1.896553e-07,1.896556e-07,1.896559e-07,1.896561e-07,1.896564e-07,1.896567e-07,1.896570e-07,1.896573e-07,1.896575e-07,1.896578e-07,1.896581e-07,1.896584e-07,1.896587e-07,1.896590e-07,1.896592e-07,1.896595e-07,1.896598e-07,1.896601e-07,1.896604e-07,1.896607e-07,1.896609e-07,1.896612e-07,1.896615e-07,1.896618e-07,1.896621e-07,1.896624e-07,1.896626e-07,1.896629e-07,1.896632e-07,1.896635e-07,1.896638e-07,1.896640e-07,1.896643e-07,1.896646e-07,1.896649e-07,1.896652e-07,1.896655e-07,1.896657e-07,1.896660e-07,1.896663e-07,1.896666e-07,1.896669e-07,1.896672e-07,1.896674e-07,1.896677e-07,1.896680e-07,1.896683e-07,1.896686e-07,1.896688e-07,1.896691e-07,1.896694e-07,1.896697e-07,1.896700e-07,1.896703e-07,1.896705e-07,1.896708e-07,1.896711e-07,1.896714e-07,1.896717e-07,1.896720e-07,1.896722e-07,1.896725e-07,1.896728e-07,1.896731e-07,1.896734e-07,1.896736e-07,1.896739e-07,1.896742e-07,1.896745e-07,1.896748e-07,1.896751e-07,1.896753e-07,1.896756e-07,1.896759e-07,1.896762e-07,1.896765e-07,1.896768e-07,1.896770e-07,1.896773e-07,1.896776e-07,1.896779e-07,1.896782e-07,1.896784e-07,1.896787e-07,1.896790e-07,1.896793e-07,1.896796e-07,1.896799e-07,1.896801e-07,1.896804e-07,1.896807e-07,1.896810e-07,1.896813e-07,1.896815e-07,1.896818e-07,1.896821e-07,1.896824e-07,1.896827e-07,1.896830e-07,1.896832e-07,1.896835e-07,1.896838e-07,1.896841e-07,1.896844e-07,1.896846e-07,1.896849e-07,1.896852e-07,1.896855e-07,1.896858e-07,1.896861e-07,1.896863e-07,1.896866e-07,1.896869e-07,1.896872e-07,1.896875e-07,1.896878e-07,1.896880e-07,1.896883e-07,1.896886e-07,1.896889e-07,1.896892e-07,1.896894e-07,1.896897e-07,1.896900e-07,1.896903e-07,1.896906e-07,1.896909e-07,1.896911e-07,1.896914e-07,1.896917e-07,1.896920e-07,1.896923e-07,1.896925e-07,1.896928e-07,1.896931e-07,1.896934e-07,1.896937e-07,1.896940e-07,1.896942e-07,1.896945e-07,1.896948e-07,1.896951e-07,1.896954e-07,1.896956e-07,1.896959e-07,1.896962e-07,1.896965e-07,1.896968e-07,1.896971e-07,1.896973e-07,1.896976e-07,1.896979e-07,1.896982e-07,1.896985e-07,1.896987e-07,1.896990e-07,1.896993e-07,1.896996e-07,1.896999e-07,1.897001e-07,1.897004e-07,1.897007e-07,1.897010e-07,1.897013e-07,1.897016e-07,1.897018e-07,1.897021e-07,1.897024e-07,1.897027e-07,1.897030e-07,1.897032e-07,1.897035e-07,1.897038e-07,1.897041e-07,1.897044e-07,1.897047e-07,1.897049e-07,1.897052e-07,1.897055e-07,1.897058e-07,1.897061e-07,1.897063e-07,1.897066e-07,1.897069e-07,1.897072e-07,1.897075e-07,1.897077e-07,1.897080e-07,1.897083e-07,1.897086e-07,1.897089e-07,1.897092e-07,1.897094e-07,1.897097e-07,1.897100e-07,1.897103e-07,1.897106e-07,1.897108e-07,1.897111e-07,1.897114e-07,1.897117e-07,1.897120e-07,1.897123e-07,1.897125e-07,1.897128e-07,1.897131e-07,1.897134e-07,1.897137e-07,1.897139e-07,1.897142e-07,1.897145e-07,1.897148e-07,1.897151e-07,1.897153e-07,1.897156e-07,1.897159e-07,1.897162e-07,1.897165e-07,1.897168e-07,1.897170e-07,1.897173e-07,1.897176e-07,1.897179e-07,1.897182e-07,1.897184e-07,1.897187e-07,1.897190e-07,1.897193e-07,1.897196e-07,1.897198e-07,1.897201e-07,1.897204e-07,1.897207e-07,1.897210e-07,1.897213e-07,1.897215e-07,1.897218e-07,1.897221e-07,1.897224e-07,1.897227e-07,1.897229e-07,1.897232e-07,1.897235e-07,1.897238e-07,1.897241e-07,1.897243e-07,1.897246e-07,1.897249e-07,1.897252e-07,1.897255e-07,1.897257e-07,1.897260e-07,1.897263e-07,1.897266e-07,1.897269e-07,1.897272e-07,1.897274e-07,1.897277e-07,1.897280e-07,1.897283e-07,1.897286e-07,1.897288e-07,1.897291e-07,1.897294e-07,1.897297e-07,1.897300e-07,1.897302e-07,1.897305e-07,1.897308e-07,1.897311e-07,1.897314e-07,1.897316e-07,1.897319e-07,1.897322e-07,1.897325e-07,1.897328e-07,1.897331e-07,1.897333e-07,1.897336e-07,1.897339e-07,1.897342e-07,1.897345e-07,1.897347e-07,1.897350e-07,1.897353e-07,1.897356e-07,1.897359e-07,1.897361e-07,1.897364e-07,1.897367e-07,1.897370e-07,1.897373e-07,1.897375e-07,1.897378e-07,1.897381e-07,1.897384e-07,1.897387e-07,1.897389e-07,1.897392e-07,1.897395e-07,1.897398e-07,1.897401e-07,1.897404e-07,1.897406e-07,1.897409e-07,1.897412e-07,1.897415e-07,1.897418e-07,1.897420e-07,1.897423e-07,1.897426e-07,1.897429e-07,1.897432e-07,1.897434e-07,1.897437e-07,1.897440e-07,1.897443e-07,1.897446e-07,1.897448e-07,1.897451e-07,1.897454e-07,1.897457e-07,1.897460e-07,1.897462e-07,1.897465e-07,1.897468e-07,1.897471e-07,1.897474e-07,1.897476e-07,1.897479e-07,1.897482e-07,1.897485e-07,1.897488e-07,1.897490e-07,1.897493e-07,1.897496e-07,1.897499e-07,1.897502e-07,1.897504e-07,1.897507e-07,1.897510e-07,1.897513e-07,1.897516e-07,1.897519e-07,1.897521e-07,1.897524e-07,1.897527e-07,1.897530e-07,1.897533e-07,1.897535e-07,1.897538e-07,1.897541e-07,1.897544e-07,1.897547e-07,1.897549e-07,1.897552e-07,1.897555e-07,1.897558e-07,1.897561e-07,1.897563e-07,1.897566e-07,1.897569e-07,1.897572e-07,1.897575e-07,1.897577e-07,1.897580e-07,1.897583e-07,1.897586e-07,1.897589e-07,1.897591e-07,1.897594e-07,1.897597e-07,1.897600e-07,1.897603e-07,1.897605e-07,1.897608e-07,1.897611e-07,1.897614e-07,1.897617e-07,1.897619e-07,1.897622e-07,1.897625e-07,1.897628e-07,1.897631e-07,1.897633e-07,1.897636e-07,1.897639e-07,1.897642e-07,1.897645e-07,1.897647e-07,1.897650e-07,1.897653e-07,1.897656e-07,1.897659e-07,1.897661e-07,1.897664e-07,1.897667e-07,1.897670e-07,1.897673e-07,1.897675e-07,1.897678e-07,1.897681e-07,1.897684e-07,1.897687e-07,1.897689e-07,1.897692e-07,1.897695e-07,1.897698e-07,1.897701e-07,1.897703e-07,1.897706e-07,1.897709e-07,1.897712e-07,1.897715e-07,1.897717e-07,1.897720e-07,1.897723e-07,1.897726e-07,1.897729e-07,1.897731e-07,1.897734e-07,1.897737e-07,1.897740e-07,1.897743e-07,1.897745e-07,1.897748e-07,1.897751e-07,1.897754e-07,1.897757e-07,1.897759e-07,1.897762e-07,1.897765e-07,1.897768e-07,1.897771e-07,1.897773e-07,1.897776e-07,1.897779e-07,1.897782e-07,1.897785e-07,1.897787e-07,1.897790e-07,1.897793e-07,1.897796e-07,1.897799e-07,1.897801e-07,1.897804e-07,1.897807e-07,1.897810e-07,1.897813e-07,1.897815e-07,1.897818e-07,1.897821e-07,1.897824e-07,1.897827e-07,1.897829e-07,1.897832e-07,1.897835e-07,1.897838e-07,1.897841e-07,1.897843e-07,1.897846e-07,1.897849e-07,1.897852e-07,1.897854e-07,1.897857e-07,1.897860e-07,1.897863e-07,1.897866e-07,1.897868e-07,1.897871e-07,1.897874e-07,1.897877e-07,1.897880e-07,1.897882e-07,1.897885e-07,1.897888e-07,1.897891e-07,1.897894e-07,1.897896e-07,1.897899e-07,1.897902e-07,1.897905e-07,1.897908e-07,1.897910e-07,1.897913e-07,1.897916e-07,1.897919e-07,1.897922e-07,1.897924e-07,1.897927e-07,1.897930e-07,1.897933e-07,1.897936e-07,1.897938e-07,1.897941e-07,1.897944e-07,1.897947e-07,1.897949e-07,1.897952e-07,1.897955e-07,1.897958e-07,1.897961e-07,1.897963e-07,1.897966e-07,1.897969e-07,1.897972e-07,1.897975e-07,1.897977e-07,1.897980e-07,1.897983e-07,1.897986e-07,1.897989e-07,1.897991e-07,1.897994e-07,1.897997e-07,1.898000e-07,1.898003e-07,1.898005e-07,1.898008e-07,1.898011e-07,1.898014e-07,1.898017e-07,1.898019e-07,1.898022e-07,1.898025e-07,1.898028e-07,1.898030e-07,1.898033e-07,1.898036e-07,1.898039e-07,1.898042e-07,1.898044e-07,1.898047e-07,1.898050e-07,1.898053e-07,1.898056e-07,1.898058e-07,1.898061e-07,1.898064e-07,1.898067e-07,1.898070e-07,1.898072e-07,1.898075e-07,1.898078e-07,1.898081e-07,1.898084e-07,1.898086e-07,1.898089e-07,1.898092e-07,1.898095e-07,1.898097e-07,1.898100e-07,1.898103e-07,1.898106e-07,1.898109e-07,1.898111e-07,1.898114e-07,1.898117e-07,1.898120e-07,1.898123e-07,1.898125e-07,1.898128e-07,1.898131e-07,1.898134e-07,1.898137e-07,1.898139e-07,1.898142e-07,1.898145e-07,1.898148e-07,1.898150e-07,1.898153e-07,1.898156e-07,1.898159e-07,1.898162e-07,1.898164e-07,1.898167e-07,1.898170e-07,1.898173e-07,1.898176e-07,1.898178e-07,1.898181e-07,1.898184e-07,1.898187e-07,1.898189e-07,1.898192e-07,1.898195e-07,1.898198e-07,1.898201e-07,1.898203e-07,1.898206e-07,1.898209e-07,1.898212e-07,1.898215e-07,1.898217e-07,1.898220e-07,1.898223e-07,1.898226e-07,1.898229e-07,1.898231e-07,1.898234e-07,1.898237e-07,1.898240e-07,1.898242e-07,1.898245e-07,1.898248e-07,1.898251e-07,1.898254e-07,1.898256e-07,1.898259e-07,1.898262e-07,1.898265e-07,1.898268e-07,1.898270e-07,1.898273e-07,1.898276e-07,1.898279e-07,1.898281e-07,1.898284e-07,1.898287e-07,1.898290e-07,1.898293e-07,1.898295e-07,1.898298e-07,1.898301e-07,1.898304e-07,1.898307e-07,1.898309e-07,1.898312e-07,1.898315e-07,1.898318e-07,1.898320e-07,1.898323e-07,1.898326e-07,1.898329e-07,1.898332e-07,1.898334e-07,1.898337e-07,1.898340e-07,1.898343e-07,1.898345e-07,1.898348e-07,1.898351e-07,1.898354e-07,1.898357e-07,1.898359e-07,1.898362e-07,1.898365e-07,1.898368e-07,1.898371e-07,1.898373e-07,1.898376e-07,1.898379e-07,1.898382e-07,1.898384e-07,1.898387e-07,1.898390e-07,1.898393e-07,1.898396e-07,1.898398e-07,1.898401e-07,1.898404e-07,1.898407e-07,1.898410e-07,1.898412e-07,1.898415e-07,1.898418e-07,1.898421e-07,1.898423e-07,1.898426e-07,1.898429e-07,1.898432e-07,1.898435e-07,1.898437e-07,1.898440e-07,1.898443e-07,1.898446e-07,1.898448e-07,1.898451e-07,1.898454e-07,1.898457e-07,1.898460e-07,1.898462e-07,1.898465e-07,1.898468e-07,1.898471e-07,1.898473e-07,1.898476e-07,1.898479e-07,1.898482e-07,1.898485e-07,1.898487e-07,1.898490e-07,1.898493e-07,1.898496e-07,1.898499e-07,1.898501e-07,1.898504e-07,1.898507e-07,1.898510e-07,1.898512e-07,1.898515e-07,1.898518e-07,1.898521e-07,1.898524e-07,1.898526e-07,1.898529e-07,1.898532e-07,1.898535e-07,1.898537e-07,1.898540e-07,1.898543e-07,1.898546e-07,1.898549e-07,1.898551e-07,1.898554e-07,1.898557e-07,1.898560e-07,1.898562e-07,1.898565e-07,1.898568e-07,1.898571e-07,1.898574e-07,1.898576e-07,1.898579e-07,1.898582e-07,1.898585e-07,1.898587e-07,1.898590e-07,1.898593e-07,1.898596e-07,1.898599e-07,1.898601e-07,1.898604e-07,1.898607e-07,1.898610e-07,1.898612e-07,1.898615e-07,1.898618e-07,1.898621e-07,1.898624e-07,1.898626e-07,1.898629e-07,1.898632e-07,1.898635e-07,1.898637e-07,1.898640e-07,1.898643e-07,1.898646e-07,1.898649e-07,1.898651e-07,1.898654e-07,1.898657e-07,1.898660e-07,1.898662e-07,1.898665e-07,1.898668e-07,1.898671e-07,1.898674e-07,1.898676e-07,1.898679e-07,1.898682e-07,1.898685e-07,1.898687e-07,1.898690e-07,1.898693e-07,1.898696e-07,1.898699e-07,1.898701e-07,1.898704e-07,1.898707e-07,1.898710e-07,1.898712e-07,1.898715e-07,1.898718e-07,1.898721e-07,1.898724e-07,1.898726e-07,1.898729e-07,1.898732e-07,1.898735e-07,1.898737e-07,1.898740e-07,1.898743e-07,1.898746e-07,1.898748e-07,1.898751e-07,1.898754e-07,1.898757e-07,1.898760e-07,1.898762e-07,1.898765e-07,1.898768e-07,1.898771e-07,1.898773e-07,1.898776e-07,1.898779e-07,1.898782e-07,1.898785e-07,1.898787e-07,1.898790e-07,1.898793e-07,1.898796e-07,1.898798e-07,1.898801e-07,1.898804e-07,1.898807e-07,1.898810e-07,1.898812e-07,1.898815e-07,1.898818e-07,1.898821e-07,1.898823e-07,1.898826e-07,1.898829e-07,1.898832e-07,1.898834e-07,1.898837e-07,1.898840e-07,1.898843e-07,1.898846e-07,1.898848e-07,1.898851e-07,1.898854e-07,1.898857e-07,1.898859e-07,1.898862e-07,1.898865e-07,1.898868e-07,1.898870e-07,1.898873e-07,1.898876e-07,1.898879e-07,1.898882e-07,1.898884e-07,1.898887e-07,1.898890e-07,1.898893e-07,1.898895e-07,1.898898e-07,1.898901e-07,1.898904e-07,1.898907e-07,1.898909e-07,1.898912e-07,1.898915e-07,1.898918e-07,1.898920e-07,1.898923e-07,1.898926e-07,1.898929e-07,1.898931e-07,1.898934e-07,1.898937e-07,1.898940e-07,1.898943e-07,1.898945e-07,1.898948e-07,1.898951e-07,1.898954e-07,1.898956e-07,1.898959e-07,1.898962e-07,1.898965e-07,1.898967e-07,1.898970e-07,1.898973e-07,1.898976e-07,1.898979e-07,1.898981e-07,1.898984e-07,1.898987e-07,1.898990e-07,1.898992e-07,1.898995e-07,1.898998e-07,1.899001e-07,1.899003e-07,1.899006e-07,1.899009e-07,1.899012e-07,1.899015e-07,1.899017e-07,1.899020e-07,1.899023e-07,1.899026e-07,1.899028e-07,1.899031e-07,1.899034e-07,1.899037e-07,1.899039e-07,1.899042e-07,1.899045e-07,1.899048e-07,1.899051e-07,1.899053e-07,1.899056e-07,1.899059e-07,1.899062e-07,1.899064e-07,1.899067e-07,1.899070e-07,1.899073e-07,1.899075e-07,1.899078e-07,1.899081e-07,1.899084e-07,1.899086e-07,1.899089e-07,1.899092e-07,1.899095e-07,1.899098e-07,1.899100e-07,1.899103e-07,1.899106e-07,1.899109e-07,1.899111e-07,1.899114e-07,1.899117e-07,1.899120e-07,1.899122e-07,1.899125e-07,1.899128e-07,1.899131e-07,1.899133e-07,1.899136e-07,1.899139e-07,1.899142e-07,1.899145e-07,1.899147e-07,1.899150e-07,1.899153e-07,1.899156e-07,1.899158e-07,1.899161e-07,1.899164e-07,1.899167e-07,1.899169e-07,1.899172e-07,1.899175e-07,1.899178e-07,1.899180e-07,1.899183e-07,1.899186e-07,1.899189e-07,1.899192e-07,1.899194e-07,1.899197e-07,1.899200e-07,1.899203e-07,1.899205e-07,1.899208e-07,1.899211e-07,1.899214e-07,1.899216e-07,1.899219e-07,1.899222e-07,1.899225e-07,1.899227e-07,1.899230e-07,1.899233e-07,1.899236e-07,1.899239e-07,1.899241e-07,1.899244e-07,1.899247e-07,1.899250e-07,1.899252e-07,1.899255e-07,1.899258e-07,1.899261e-07,1.899263e-07,1.899266e-07,1.899269e-07,1.899272e-07,1.899274e-07,1.899277e-07,1.899280e-07,1.899283e-07,1.899285e-07,1.899288e-07,1.899291e-07,1.899294e-07,1.899297e-07,1.899299e-07,1.899302e-07,1.899305e-07,1.899308e-07,1.899310e-07,1.899313e-07,1.899316e-07,1.899319e-07,1.899321e-07,1.899324e-07,1.899327e-07,1.899330e-07,1.899332e-07,1.899335e-07,1.899338e-07,1.899341e-07,1.899343e-07,1.899346e-07,1.899349e-07,1.899352e-07,1.899355e-07,1.899357e-07,1.899360e-07,1.899363e-07,1.899366e-07,1.899368e-07,1.899371e-07,1.899374e-07,1.899377e-07,1.899379e-07,1.899382e-07,1.899385e-07,1.899388e-07,1.899390e-07,1.899393e-07,1.899396e-07,1.899399e-07,1.899401e-07,1.899404e-07,1.899407e-07,1.899410e-07,1.899412e-07,1.899415e-07,1.899418e-07,1.899421e-07,1.899423e-07,1.899426e-07,1.899429e-07,1.899432e-07,1.899435e-07,1.899437e-07,1.899440e-07,1.899443e-07,1.899446e-07,1.899448e-07,1.899451e-07,1.899454e-07,1.899457e-07,1.899459e-07,1.899462e-07,1.899465e-07,1.899468e-07,1.899470e-07,1.899473e-07,1.899476e-07,1.899479e-07,1.899481e-07,1.899484e-07,1.899487e-07,1.899490e-07,1.899492e-07,1.899495e-07,1.899498e-07,1.899501e-07,1.899503e-07,1.899506e-07,1.899509e-07,1.899512e-07,1.899514e-07,1.899517e-07,1.899520e-07,1.899523e-07,1.899526e-07,1.899528e-07,1.899531e-07,1.899534e-07,1.899537e-07,1.899539e-07,1.899542e-07,1.899545e-07,1.899548e-07,1.899550e-07,1.899553e-07,1.899556e-07,1.899559e-07,1.899561e-07,1.899564e-07,1.899567e-07,1.899570e-07,1.899572e-07,1.899575e-07,1.899578e-07,1.899581e-07,1.899583e-07,1.899586e-07,1.899589e-07,1.899592e-07,1.899594e-07,1.899597e-07,1.899600e-07,1.899603e-07,1.899605e-07,1.899608e-07,1.899611e-07,1.899614e-07,1.899616e-07,1.899619e-07,1.899622e-07,1.899625e-07,1.899627e-07,1.899630e-07,1.899633e-07,1.899636e-07,1.899638e-07,1.899641e-07,1.899644e-07,1.899647e-07,1.899649e-07,1.899652e-07,1.899655e-07,1.899658e-07,1.899660e-07,1.899663e-07,1.899666e-07,1.899669e-07,1.899671e-07,1.899674e-07,1.899677e-07,1.899680e-07,1.899682e-07,1.899685e-07,1.899688e-07,1.899691e-07,1.899693e-07,1.899696e-07,1.899699e-07,1.899702e-07,1.899705e-07,1.899707e-07,1.899710e-07,1.899713e-07,1.899716e-07,1.899718e-07,1.899721e-07,1.899724e-07,1.899727e-07,1.899729e-07,1.899732e-07,1.899735e-07,1.899738e-07,1.899740e-07,1.899743e-07,1.899746e-07,1.899749e-07,1.899751e-07,1.899754e-07,1.899757e-07,1.899760e-07,1.899762e-07,1.899765e-07,1.899768e-07,1.899771e-07,1.899773e-07,1.899776e-07,1.899779e-07,1.899782e-07,1.899784e-07,1.899787e-07,1.899790e-07,1.899793e-07,1.899795e-07,1.899798e-07,1.899801e-07,1.899804e-07,1.899806e-07,1.899809e-07,1.899812e-07,1.899815e-07,1.899817e-07,1.899820e-07,1.899823e-07,1.899826e-07,1.899828e-07,1.899831e-07,1.899834e-07,1.899837e-07,1.899839e-07,1.899842e-07,1.899845e-07,1.899848e-07,1.899850e-07,1.899853e-07,1.899856e-07,1.899859e-07,1.899861e-07,1.899864e-07,1.899867e-07,1.899869e-07,1.899872e-07,1.899875e-07,1.899878e-07,1.899880e-07,1.899883e-07,1.899886e-07,1.899889e-07,1.899891e-07,1.899894e-07,1.899897e-07,1.899900e-07,1.899902e-07,1.899905e-07,1.899908e-07,1.899911e-07,1.899913e-07,1.899916e-07,1.899919e-07,1.899922e-07,1.899924e-07,1.899927e-07,1.899930e-07,1.899933e-07,1.899935e-07,1.899938e-07,1.899941e-07,1.899944e-07,1.899946e-07,1.899949e-07,1.899952e-07,1.899955e-07,1.899957e-07,1.899960e-07,1.899963e-07,1.899966e-07,1.899968e-07,1.899971e-07,1.899974e-07,1.899977e-07,1.899979e-07,1.899982e-07,1.899985e-07,1.899988e-07,1.899990e-07,1.899993e-07,1.899996e-07,1.899999e-07,1.900001e-07,1.900004e-07,1.900007e-07,1.900010e-07,1.900012e-07,1.900015e-07,1.900018e-07,1.900021e-07,1.900023e-07,1.900026e-07,1.900029e-07,1.900032e-07,1.900034e-07,1.900037e-07,1.900040e-07,1.900042e-07,1.900045e-07,1.900048e-07,1.900051e-07,1.900053e-07,1.900056e-07,1.900059e-07,1.900062e-07,1.900064e-07,1.900067e-07,1.900070e-07,1.900073e-07,1.900075e-07,1.900078e-07,1.900081e-07,1.900084e-07,1.900086e-07,1.900089e-07,1.900092e-07,1.900095e-07,1.900097e-07,1.900100e-07,1.900103e-07,1.900106e-07,1.900108e-07,1.900111e-07,1.900114e-07,1.900117e-07,1.900119e-07,1.900122e-07,1.900125e-07,1.900128e-07,1.900130e-07,1.900133e-07,1.900136e-07,1.900138e-07,1.900141e-07,1.900144e-07,1.900147e-07,1.900149e-07,1.900152e-07,1.900155e-07,1.900158e-07,1.900160e-07,1.900163e-07,1.900166e-07,1.900169e-07,1.900171e-07,1.900174e-07,1.900177e-07,1.900180e-07,1.900182e-07,1.900185e-07,1.900188e-07,1.900191e-07,1.900193e-07,1.900196e-07,1.900199e-07,1.900202e-07,1.900204e-07,1.900207e-07,1.900210e-07,1.900212e-07,1.900215e-07,1.900218e-07,1.900221e-07,1.900223e-07,1.900226e-07,1.900229e-07,1.900232e-07,1.900234e-07,1.900237e-07,1.900240e-07,1.900243e-07,1.900245e-07,1.900248e-07,1.900251e-07,1.900254e-07,1.900256e-07,1.900259e-07,1.900262e-07,1.900265e-07,1.900267e-07,1.900270e-07,1.900273e-07,1.900275e-07,1.900278e-07,1.900281e-07,1.900284e-07,1.900286e-07,1.900289e-07,1.900292e-07,1.900295e-07,1.900297e-07,1.900300e-07,1.900303e-07,1.900306e-07,1.900308e-07,1.900311e-07,1.900314e-07,1.900317e-07,1.900319e-07,1.900322e-07,1.900325e-07,1.900328e-07,1.900330e-07,1.900333e-07,1.900336e-07,1.900338e-07,1.900341e-07,1.900344e-07,1.900347e-07,1.900349e-07,1.900352e-07,1.900355e-07,1.900358e-07,1.900360e-07,1.900363e-07,1.900366e-07,1.900369e-07,1.900371e-07,1.900374e-07,1.900377e-07,1.900380e-07,1.900382e-07,1.900385e-07,1.900388e-07,1.900390e-07,1.900393e-07,1.900396e-07,1.900399e-07,1.900401e-07,1.900404e-07,1.900407e-07,1.900410e-07,1.900412e-07,1.900415e-07,1.900418e-07,1.900421e-07,1.900423e-07,1.900426e-07,1.900429e-07,1.900431e-07,1.900434e-07,1.900437e-07,1.900440e-07,1.900442e-07,1.900445e-07,1.900448e-07,1.900451e-07,1.900453e-07,1.900456e-07,1.900459e-07,1.900462e-07,1.900464e-07,1.900467e-07,1.900470e-07,1.900472e-07,1.900475e-07,1.900478e-07,1.900481e-07,1.900483e-07,1.900486e-07,1.900489e-07,1.900492e-07,1.900494e-07,1.900497e-07,1.900500e-07,1.900503e-07,1.900505e-07,1.900508e-07,1.900511e-07,1.900513e-07,1.900516e-07,1.900519e-07,1.900522e-07,1.900524e-07,1.900527e-07,1.900530e-07,1.900533e-07,1.900535e-07,1.900538e-07,1.900541e-07,1.900544e-07,1.900546e-07,1.900549e-07,1.900552e-07,1.900554e-07,1.900557e-07,1.900560e-07,1.900563e-07,1.900565e-07,1.900568e-07,1.900571e-07,1.900574e-07,1.900576e-07,1.900579e-07,1.900582e-07,1.900585e-07,1.900587e-07,1.900590e-07,1.900593e-07,1.900595e-07,1.900598e-07,1.900601e-07,1.900604e-07,1.900606e-07,1.900609e-07,1.900612e-07,1.900615e-07,1.900617e-07,1.900620e-07,1.900623e-07,1.900625e-07,1.900628e-07,1.900631e-07,1.900634e-07,1.900636e-07,1.900639e-07,1.900642e-07,1.900645e-07,1.900647e-07,1.900650e-07,1.900653e-07,1.900656e-07,1.900658e-07,1.900661e-07,1.900664e-07,1.900666e-07,1.900669e-07,1.900672e-07,1.900675e-07,1.900677e-07,1.900680e-07,1.900683e-07,1.900686e-07,1.900688e-07,1.900691e-07,1.900694e-07,1.900696e-07,1.900699e-07,1.900702e-07,1.900705e-07,1.900707e-07,1.900710e-07,1.900713e-07,1.900716e-07,1.900718e-07,1.900721e-07,1.900724e-07,1.900726e-07,1.900729e-07,1.900732e-07,1.900735e-07,1.900737e-07,1.900740e-07,1.900743e-07,1.900746e-07,1.900748e-07,1.900751e-07,1.900754e-07,1.900756e-07,1.900759e-07,1.900762e-07,1.900765e-07,1.900767e-07,1.900770e-07,1.900773e-07,1.900776e-07,1.900778e-07,1.900781e-07,1.900784e-07,1.900786e-07,1.900789e-07,1.900792e-07,1.900795e-07,1.900797e-07,1.900800e-07,1.900803e-07,1.900806e-07,1.900808e-07,1.900811e-07,1.900814e-07,1.900816e-07,1.900819e-07,1.900822e-07,1.900825e-07,1.900827e-07,1.900830e-07,1.900833e-07,1.900836e-07,1.900838e-07,1.900841e-07,1.900844e-07,1.900846e-07,1.900849e-07,1.900852e-07,1.900855e-07,1.900857e-07,1.900860e-07,1.900863e-07,1.900865e-07,1.900868e-07,1.900871e-07,1.900874e-07,1.900876e-07,1.900879e-07,1.900882e-07,1.900885e-07,1.900887e-07,1.900890e-07,1.900893e-07,1.900895e-07,1.900898e-07,1.900901e-07,1.900904e-07,1.900906e-07,1.900909e-07,1.900912e-07,1.900915e-07,1.900917e-07,1.900920e-07,1.900923e-07,1.900925e-07,1.900928e-07,1.900931e-07,1.900934e-07,1.900936e-07,1.900939e-07,1.900942e-07,1.900944e-07,1.900947e-07,1.900950e-07,1.900953e-07,1.900955e-07,1.900958e-07,1.900961e-07,1.900964e-07,1.900966e-07,1.900969e-07,1.900972e-07,1.900974e-07,1.900977e-07,1.900980e-07,1.900983e-07,1.900985e-07,1.900988e-07,1.900991e-07,1.900993e-07,1.900996e-07,1.900999e-07,1.901002e-07,1.901004e-07,1.901007e-07,1.901010e-07,1.901013e-07,1.901015e-07,1.901018e-07,1.901021e-07,1.901023e-07,1.901026e-07,1.901029e-07,1.901032e-07,1.901034e-07,1.901037e-07,1.901040e-07,1.901042e-07,1.901045e-07,1.901048e-07,1.901051e-07,1.901053e-07,1.901056e-07,1.901059e-07,1.901062e-07,1.901064e-07,1.901067e-07,1.901070e-07,1.901072e-07,1.901075e-07,1.901078e-07,1.901081e-07,1.901083e-07,1.901086e-07,1.901089e-07,1.901091e-07,1.901094e-07,1.901097e-07,1.901100e-07,1.901102e-07,1.901105e-07,1.901108e-07,1.901110e-07,1.901113e-07,1.901116e-07,1.901119e-07,1.901121e-07,1.901124e-07,1.901127e-07,1.901129e-07,1.901132e-07,1.901135e-07,1.901138e-07,1.901140e-07,1.901143e-07,1.901146e-07,1.901149e-07,1.901151e-07,1.901154e-07,1.901157e-07,1.901159e-07,1.901162e-07,1.901165e-07,1.901168e-07,1.901170e-07,1.901173e-07,1.901176e-07,1.901178e-07,1.901181e-07,1.901184e-07,1.901187e-07,1.901189e-07,1.901192e-07,1.901195e-07,1.901197e-07,1.901200e-07,1.901203e-07,1.901206e-07,1.901208e-07,1.901211e-07,1.901214e-07,1.901216e-07,1.901219e-07,1.901222e-07,1.901225e-07,1.901227e-07,1.901230e-07,1.901233e-07,1.901235e-07,1.901238e-07,1.901241e-07,1.901244e-07,1.901246e-07,1.901249e-07,1.901252e-07,1.901254e-07,1.901257e-07,1.901260e-07,1.901263e-07,1.901265e-07,1.901268e-07,1.901271e-07,1.901273e-07,1.901276e-07,1.901279e-07,1.901282e-07,1.901284e-07,1.901287e-07,1.901290e-07,1.901292e-07,1.901295e-07,1.901298e-07,1.901301e-07,1.901303e-07,1.901306e-07,1.901309e-07,1.901311e-07,1.901314e-07,1.901317e-07,1.901320e-07,1.901322e-07,1.901325e-07,1.901328e-07,1.901330e-07,1.901333e-07,1.901336e-07,1.901339e-07,1.901341e-07,1.901344e-07,1.901347e-07,1.901349e-07,1.901352e-07,1.901355e-07,1.901358e-07,1.901360e-07,1.901363e-07,1.901366e-07,1.901368e-07,1.901371e-07,1.901374e-07,1.901377e-07,1.901379e-07,1.901382e-07,1.901385e-07,1.901387e-07,1.901390e-07,1.901393e-07,1.901396e-07,1.901398e-07,1.901401e-07,1.901404e-07,1.901406e-07,1.901409e-07,1.901412e-07,1.901415e-07,1.901417e-07,1.901420e-07,1.901423e-07,1.901425e-07,1.901428e-07,1.901431e-07,1.901434e-07,1.901436e-07,1.901439e-07,1.901442e-07,1.901444e-07,1.901447e-07,1.901450e-07,1.901453e-07,1.901455e-07,1.901458e-07,1.901461e-07,1.901463e-07,1.901466e-07,1.901469e-07,1.901472e-07,1.901474e-07,1.901477e-07,1.901480e-07,1.901482e-07,1.901485e-07,1.901488e-07,1.901490e-07,1.901493e-07,1.901496e-07,1.901499e-07,1.901501e-07,1.901504e-07,1.901507e-07,1.901509e-07,1.901512e-07,1.901515e-07,1.901518e-07,1.901520e-07,1.901523e-07,1.901526e-07,1.901528e-07,1.901531e-07,1.901534e-07,1.901537e-07,1.901539e-07,1.901542e-07,1.901545e-07,1.901547e-07,1.901550e-07,1.901553e-07,1.901556e-07,1.901558e-07,1.901561e-07,1.901564e-07,1.901566e-07,1.901569e-07,1.901572e-07,1.901574e-07,1.901577e-07,1.901580e-07,1.901583e-07,1.901585e-07,1.901588e-07,1.901591e-07,1.901593e-07,1.901596e-07,1.901599e-07,1.901602e-07,1.901604e-07,1.901607e-07,1.901610e-07,1.901612e-07,1.901615e-07,1.901618e-07,1.901620e-07,1.901623e-07,1.901626e-07,1.901629e-07,1.901631e-07,1.901634e-07,1.901637e-07,1.901639e-07,1.901642e-07,1.901645e-07,1.901648e-07,1.901650e-07,1.901653e-07,1.901656e-07,1.901658e-07,1.901661e-07,1.901664e-07,1.901667e-07,1.901669e-07,1.901672e-07,1.901675e-07,1.901677e-07,1.901680e-07,1.901683e-07,1.901685e-07,1.901688e-07,1.901691e-07,1.901694e-07,1.901696e-07,1.901699e-07,1.901702e-07,1.901704e-07,1.901707e-07,1.901710e-07,1.901713e-07,1.901715e-07,1.901718e-07,1.901721e-07,1.901723e-07,1.901726e-07,1.901729e-07,1.901731e-07,1.901734e-07,1.901737e-07,1.901740e-07,1.901742e-07,1.901745e-07,1.901748e-07,1.901750e-07,1.901753e-07,1.901756e-07,1.901758e-07,1.901761e-07,1.901764e-07,1.901767e-07,1.901769e-07,1.901772e-07,1.901775e-07,1.901777e-07,1.901780e-07,1.901783e-07,1.901786e-07,1.901788e-07,1.901791e-07,1.901794e-07,1.901796e-07,1.901799e-07,1.901802e-07,1.901804e-07,1.901807e-07,1.901810e-07,1.901813e-07,1.901815e-07,1.901818e-07,1.901821e-07,1.901823e-07,1.901826e-07,1.901829e-07,1.901831e-07,1.901834e-07,1.901837e-07,1.901840e-07,1.901842e-07,1.901845e-07,1.901848e-07,1.901850e-07,1.901853e-07,1.901856e-07,1.901858e-07,1.901861e-07,1.901864e-07,1.901867e-07,1.901869e-07,1.901872e-07,1.901875e-07,1.901877e-07,1.901880e-07,1.901883e-07,1.901885e-07,1.901888e-07,1.901891e-07,1.901894e-07,1.901896e-07,1.901899e-07,1.901902e-07,1.901904e-07,1.901907e-07,1.901910e-07,1.901912e-07,1.901915e-07,1.901918e-07,1.901921e-07,1.901923e-07,1.901926e-07,1.901929e-07,1.901931e-07,1.901934e-07,1.901937e-07,1.901939e-07,1.901942e-07,1.901945e-07,1.901948e-07,1.901950e-07,1.901953e-07,1.901956e-07,1.901958e-07,1.901961e-07,1.901964e-07,1.901966e-07,1.901969e-07,1.901972e-07,1.901975e-07,1.901977e-07,1.901980e-07,1.901983e-07,1.901985e-07,1.901988e-07,1.901991e-07,1.901993e-07,1.901996e-07,1.901999e-07,1.902002e-07,1.902004e-07,1.902007e-07,1.902010e-07,1.902012e-07,1.902015e-07,1.902018e-07,1.902020e-07,1.902023e-07,1.902026e-07,1.902029e-07,1.902031e-07,1.902034e-07,1.902037e-07,1.902039e-07,1.902042e-07,1.902045e-07,1.902047e-07,1.902050e-07,1.902053e-07,1.902056e-07,1.902058e-07,1.902061e-07,1.902064e-07,1.902066e-07,1.902069e-07,1.902072e-07,1.902074e-07,1.902077e-07,1.902080e-07,1.902082e-07,1.902085e-07,1.902088e-07,1.902091e-07,1.902093e-07,1.902096e-07,1.902099e-07,1.902101e-07,1.902104e-07,1.902107e-07,1.902109e-07,1.902112e-07,1.902115e-07,1.902118e-07,1.902120e-07,1.902123e-07,1.902126e-07,1.902128e-07,1.902131e-07,1.902134e-07,1.902136e-07,1.902139e-07,1.902142e-07,1.902144e-07,1.902147e-07,1.902150e-07,1.902153e-07,1.902155e-07,1.902158e-07,1.902161e-07,1.902163e-07,1.902166e-07,1.902169e-07,1.902171e-07,1.902174e-07,1.902177e-07,1.902180e-07,1.902182e-07,1.902185e-07,1.902188e-07,1.902190e-07,1.902193e-07,1.902196e-07,1.902198e-07,1.902201e-07,1.902204e-07,1.902206e-07,1.902209e-07,1.902212e-07,1.902215e-07,1.902217e-07,1.902220e-07,1.902223e-07,1.902225e-07,1.902228e-07,1.902231e-07,1.902233e-07,1.902236e-07,1.902239e-07,1.902241e-07,1.902244e-07,1.902247e-07,1.902250e-07,1.902252e-07,1.902255e-07,1.902258e-07,1.902260e-07,1.902263e-07,1.902266e-07,1.902268e-07,1.902271e-07,1.902274e-07,1.902276e-07,1.902279e-07,1.902282e-07,1.902285e-07,1.902287e-07,1.902290e-07,1.902293e-07,1.902295e-07,1.902298e-07,1.902301e-07,1.902303e-07,1.902306e-07,1.902309e-07,1.902311e-07,1.902314e-07,1.902317e-07,1.902320e-07,1.902322e-07,1.902325e-07,1.902328e-07,1.902330e-07,1.902333e-07,1.902336e-07,1.902338e-07,1.902341e-07,1.902344e-07,1.902346e-07,1.902349e-07,1.902352e-07,1.902355e-07,1.902357e-07,1.902360e-07,1.902363e-07,1.902365e-07,1.902368e-07,1.902371e-07,1.902373e-07,1.902376e-07,1.902379e-07,1.902381e-07,1.902384e-07,1.902387e-07,1.902389e-07,1.902392e-07,1.902395e-07,1.902398e-07,1.902400e-07,1.902403e-07,1.902406e-07,1.902408e-07,1.902411e-07,1.902414e-07,1.902416e-07,1.902419e-07,1.902422e-07,1.902424e-07,1.902427e-07,1.902430e-07,1.902433e-07,1.902435e-07,1.902438e-07,1.902441e-07,1.902443e-07,1.902446e-07,1.902449e-07,1.902451e-07,1.902454e-07,1.902457e-07,1.902459e-07,1.902462e-07,1.902465e-07,1.902467e-07,1.902470e-07,1.902473e-07,1.902476e-07,1.902478e-07,1.902481e-07,1.902484e-07,1.902486e-07,1.902489e-07,1.902492e-07,1.902494e-07,1.902497e-07,1.902500e-07,1.902502e-07,1.902505e-07,1.902508e-07,1.902510e-07,1.902513e-07,1.902516e-07,1.902519e-07,1.902521e-07,1.902524e-07,1.902527e-07,1.902529e-07,1.902532e-07,1.902535e-07,1.902537e-07,1.902540e-07,1.902543e-07,1.902545e-07,1.902548e-07,1.902551e-07,1.902553e-07,1.902556e-07,1.902559e-07,1.902561e-07,1.902564e-07,1.902567e-07,1.902570e-07,1.902572e-07,1.902575e-07,1.902578e-07,1.902580e-07,1.902583e-07,1.902586e-07,1.902588e-07,1.902591e-07,1.902594e-07,1.902596e-07,1.902599e-07,1.902602e-07,1.902604e-07,1.902607e-07,1.902610e-07,1.902612e-07,1.902615e-07,1.902618e-07,1.902621e-07,1.902623e-07,1.902626e-07,1.902629e-07,1.902631e-07,1.902634e-07,1.902637e-07,1.902639e-07,1.902642e-07,1.902645e-07,1.902647e-07,1.902650e-07,1.902653e-07,1.902655e-07,1.902658e-07,1.902661e-07,1.902663e-07,1.902666e-07,1.902669e-07,1.902672e-07,1.902674e-07,1.902677e-07,1.902680e-07,1.902682e-07,1.902685e-07,1.902688e-07,1.902690e-07,1.902693e-07,1.902696e-07,1.902698e-07,1.902701e-07,1.902704e-07,1.902706e-07,1.902709e-07,1.902712e-07,1.902714e-07,1.902717e-07,1.902720e-07,1.902722e-07,1.902725e-07,1.902728e-07,1.902731e-07,1.902733e-07,1.902736e-07,1.902739e-07,1.902741e-07,1.902744e-07,1.902747e-07,1.902749e-07,1.902752e-07,1.902755e-07,1.902757e-07,1.902760e-07,1.902763e-07,1.902765e-07,1.902768e-07,1.902771e-07,1.902773e-07,1.902776e-07,1.902779e-07,1.902781e-07,1.902784e-07,1.902787e-07,1.902790e-07,1.902792e-07,1.902795e-07,1.902798e-07,1.902800e-07,1.902803e-07,1.902806e-07,1.902808e-07,1.902811e-07,1.902814e-07,1.902816e-07,1.902819e-07,1.902822e-07,1.902824e-07,1.902827e-07,1.902830e-07,1.902832e-07,1.902835e-07,1.902838e-07,1.902840e-07,1.902843e-07,1.902846e-07,1.902848e-07,1.902851e-07,1.902854e-07,1.902856e-07,1.902859e-07,1.902862e-07,1.902865e-07,1.902867e-07,1.902870e-07,1.902873e-07,1.902875e-07,1.902878e-07,1.902881e-07,1.902883e-07,1.902886e-07,1.902889e-07,1.902891e-07,1.902894e-07,1.902897e-07,1.902899e-07,1.902902e-07,1.902905e-07,1.902907e-07,1.902910e-07,1.902913e-07,1.902915e-07,1.902918e-07,1.902921e-07,1.902923e-07,1.902926e-07,1.902929e-07,1.902931e-07,1.902934e-07,1.902937e-07,1.902940e-07,1.902942e-07,1.902945e-07,1.902948e-07,1.902950e-07,1.902953e-07,1.902956e-07,1.902958e-07,1.902961e-07,1.902964e-07,1.902966e-07,1.902969e-07,1.902972e-07,1.902974e-07,1.902977e-07,1.902980e-07,1.902982e-07,1.902985e-07,1.902988e-07,1.902990e-07,1.902993e-07,1.902996e-07,1.902998e-07,1.903001e-07,1.903004e-07,1.903006e-07,1.903009e-07,1.903012e-07,1.903014e-07,1.903017e-07,1.903020e-07,1.903022e-07,1.903025e-07,1.903028e-07,1.903030e-07,1.903033e-07,1.903036e-07,1.903039e-07,1.903041e-07,1.903044e-07,1.903047e-07,1.903049e-07,1.903052e-07,1.903055e-07,1.903057e-07,1.903060e-07,1.903063e-07,1.903065e-07,1.903068e-07,1.903071e-07,1.903073e-07,1.903076e-07,1.903079e-07,1.903081e-07,1.903084e-07,1.903087e-07,1.903089e-07,1.903092e-07,1.903095e-07,1.903097e-07,1.903100e-07,1.903103e-07,1.903105e-07,1.903108e-07,1.903111e-07,1.903113e-07,1.903116e-07,1.903119e-07,1.903121e-07,1.903124e-07,1.903127e-07,1.903129e-07,1.903132e-07,1.903135e-07,1.903137e-07,1.903140e-07,1.903143e-07,1.903145e-07,1.903148e-07,1.903151e-07,1.903153e-07,1.903156e-07,1.903159e-07,1.903161e-07,1.903164e-07,1.903167e-07,1.903169e-07,1.903172e-07,1.903175e-07,1.903177e-07,1.903180e-07,1.903183e-07,1.903186e-07,1.903188e-07,1.903191e-07,1.903194e-07,1.903196e-07,1.903199e-07,1.903202e-07,1.903204e-07,1.903207e-07,1.903210e-07,1.903212e-07,1.903215e-07,1.903218e-07,1.903220e-07,1.903223e-07,1.903226e-07,1.903228e-07,1.903231e-07,1.903234e-07,1.903236e-07,1.903239e-07,1.903242e-07,1.903244e-07,1.903247e-07,1.903250e-07,1.903252e-07,1.903255e-07,1.903258e-07,1.903260e-07,1.903263e-07,1.903266e-07,1.903268e-07,1.903271e-07,1.903274e-07,1.903276e-07,1.903279e-07,1.903282e-07,1.903284e-07,1.903287e-07,1.903290e-07,1.903292e-07,1.903295e-07,1.903298e-07,1.903300e-07,1.903303e-07,1.903306e-07,1.903308e-07,1.903311e-07,1.903314e-07,1.903316e-07,1.903319e-07,1.903322e-07,1.903324e-07,1.903327e-07,1.903330e-07,1.903332e-07,1.903335e-07,1.903338e-07,1.903340e-07,1.903343e-07,1.903346e-07,1.903348e-07,1.903351e-07,1.903354e-07,1.903356e-07,1.903359e-07,1.903362e-07,1.903364e-07,1.903367e-07,1.903370e-07,1.903372e-07,1.903375e-07,1.903378e-07,1.903380e-07,1.903383e-07,1.903386e-07,1.903388e-07,1.903391e-07,1.903394e-07,1.903396e-07,1.903399e-07,1.903402e-07,1.903404e-07,1.903407e-07,1.903410e-07,1.903412e-07,1.903415e-07,1.903418e-07,1.903420e-07,1.903423e-07,1.903426e-07,1.903428e-07,1.903431e-07,1.903434e-07,1.903436e-07,1.903439e-07,1.903442e-07,1.903444e-07,1.903447e-07,1.903450e-07,1.903452e-07,1.903455e-07,1.903458e-07,1.903460e-07,1.903463e-07,1.903466e-07,1.903468e-07,1.903471e-07,1.903474e-07,1.903476e-07,1.903479e-07,1.903482e-07,1.903484e-07,1.903487e-07,1.903490e-07,1.903492e-07,1.903495e-07,1.903498e-07,1.903500e-07,1.903503e-07,1.903506e-07,1.903508e-07,1.903511e-07,1.903514e-07,1.903516e-07,1.903519e-07,1.903522e-07,1.903524e-07,1.903527e-07,1.903530e-07,1.903532e-07,1.903535e-07,1.903538e-07,1.903540e-07,1.903543e-07,1.903546e-07,1.903548e-07,1.903551e-07,1.903554e-07,1.903556e-07,1.903559e-07,1.903562e-07,1.903564e-07,1.903567e-07,1.903570e-07,1.903572e-07,1.903575e-07,1.903577e-07,1.903580e-07,1.903583e-07,1.903585e-07,1.903588e-07,1.903591e-07,1.903593e-07,1.903596e-07,1.903599e-07,1.903601e-07,1.903604e-07,1.903607e-07,1.903609e-07,1.903612e-07,1.903615e-07,1.903617e-07,1.903620e-07,1.903623e-07,1.903625e-07,1.903628e-07,1.903631e-07,1.903633e-07,1.903636e-07,1.903639e-07,1.903641e-07,1.903644e-07,1.903647e-07,1.903649e-07,1.903652e-07,1.903655e-07,1.903657e-07,1.903660e-07,1.903663e-07,1.903665e-07,1.903668e-07,1.903671e-07,1.903673e-07,1.903676e-07,1.903679e-07,1.903681e-07,1.903684e-07,1.903687e-07,1.903689e-07,1.903692e-07,1.903695e-07,1.903697e-07,1.903700e-07,1.903703e-07,1.903705e-07,1.903708e-07,1.903711e-07,1.903713e-07,1.903716e-07,1.903719e-07,1.903721e-07,1.903724e-07,1.903726e-07,1.903729e-07,1.903732e-07,1.903734e-07,1.903737e-07,1.903740e-07,1.903742e-07,1.903745e-07,1.903748e-07,1.903750e-07,1.903753e-07,1.903756e-07,1.903758e-07,1.903761e-07,1.903764e-07,1.903766e-07,1.903769e-07,1.903772e-07,1.903774e-07,1.903777e-07,1.903780e-07,1.903782e-07,1.903785e-07,1.903788e-07,1.903790e-07,1.903793e-07,1.903796e-07,1.903798e-07,1.903801e-07,1.903804e-07,1.903806e-07,1.903809e-07,1.903812e-07,1.903814e-07,1.903817e-07,1.903820e-07,1.903822e-07,1.903825e-07,1.903827e-07,1.903830e-07,1.903833e-07,1.903835e-07,1.903838e-07,1.903841e-07,1.903843e-07,1.903846e-07,1.903849e-07,1.903851e-07,1.903854e-07,1.903857e-07,1.903859e-07,1.903862e-07,1.903865e-07,1.903867e-07,1.903870e-07,1.903873e-07,1.903875e-07,1.903878e-07,1.903881e-07,1.903883e-07,1.903886e-07,1.903889e-07,1.903891e-07,1.903894e-07,1.903897e-07,1.903899e-07,1.903902e-07,1.903904e-07,1.903907e-07,1.903910e-07,1.903912e-07,1.903915e-07,1.903918e-07,1.903920e-07,1.903923e-07,1.903926e-07,1.903928e-07,1.903931e-07,1.903934e-07,1.903936e-07,1.903939e-07,1.903942e-07,1.903944e-07,1.903947e-07,1.903950e-07,1.903952e-07,1.903955e-07,1.903958e-07,1.903960e-07,1.903963e-07,1.903966e-07,1.903968e-07,1.903971e-07,1.903973e-07,1.903976e-07,1.903979e-07,1.903981e-07,1.903984e-07,1.903987e-07,1.903989e-07,1.903992e-07,1.903995e-07,1.903997e-07,1.904000e-07,1.904003e-07,1.904005e-07,1.904008e-07,1.904011e-07,1.904013e-07,1.904016e-07,1.904019e-07,1.904021e-07,1.904024e-07,1.904027e-07,1.904029e-07,1.904032e-07,1.904034e-07,1.904037e-07,1.904040e-07,1.904042e-07,1.904045e-07,1.904048e-07,1.904050e-07,1.904053e-07,1.904056e-07,1.904058e-07,1.904061e-07,1.904064e-07,1.904066e-07,1.904069e-07,1.904072e-07,1.904074e-07,1.904077e-07,1.904080e-07,1.904082e-07,1.904085e-07,1.904088e-07,1.904090e-07,1.904093e-07,1.904095e-07,1.904098e-07,1.904101e-07,1.904103e-07,1.904106e-07,1.904109e-07,1.904111e-07,1.904114e-07,1.904117e-07,1.904119e-07,1.904122e-07,1.904125e-07,1.904127e-07,1.904130e-07,1.904133e-07,1.904135e-07,1.904138e-07,1.904141e-07,1.904143e-07,1.904146e-07,1.904148e-07,1.904151e-07,1.904154e-07,1.904156e-07,1.904159e-07,1.904162e-07,1.904164e-07,1.904167e-07,1.904170e-07,1.904172e-07,1.904175e-07,1.904178e-07,1.904180e-07,1.904183e-07,1.904186e-07,1.904188e-07,1.904191e-07,1.904193e-07,1.904196e-07,1.904199e-07,1.904201e-07,1.904204e-07,1.904207e-07,1.904209e-07,1.904212e-07,1.904215e-07,1.904217e-07,1.904220e-07,1.904223e-07,1.904225e-07,1.904228e-07,1.904231e-07,1.904233e-07,1.904236e-07,1.904239e-07,1.904241e-07,1.904244e-07,1.904246e-07,1.904249e-07,1.904252e-07,1.904254e-07,1.904257e-07,1.904260e-07,1.904262e-07,1.904265e-07,1.904268e-07,1.904270e-07,1.904273e-07,1.904276e-07,1.904278e-07,1.904281e-07,1.904283e-07,1.904286e-07,1.904289e-07,1.904291e-07,1.904294e-07,1.904297e-07,1.904299e-07,1.904302e-07,1.904305e-07,1.904307e-07,1.904310e-07,1.904313e-07,1.904315e-07,1.904318e-07,1.904321e-07,1.904323e-07,1.904326e-07,1.904328e-07,1.904331e-07,1.904334e-07,1.904336e-07,1.904339e-07,1.904342e-07,1.904344e-07,1.904347e-07,1.904350e-07,1.904352e-07,1.904355e-07,1.904358e-07,1.904360e-07,1.904363e-07,1.904365e-07,1.904368e-07,1.904371e-07,1.904373e-07,1.904376e-07,1.904379e-07,1.904381e-07,1.904384e-07,1.904387e-07,1.904389e-07,1.904392e-07,1.904395e-07,1.904397e-07,1.904400e-07,1.904403e-07,1.904405e-07,1.904408e-07,1.904410e-07,1.904413e-07,1.904416e-07,1.904418e-07,1.904421e-07,1.904424e-07,1.904426e-07,1.904429e-07,1.904432e-07,1.904434e-07,1.904437e-07,1.904440e-07,1.904442e-07,1.904445e-07,1.904447e-07,1.904450e-07,1.904453e-07,1.904455e-07,1.904458e-07,1.904461e-07,1.904463e-07,1.904466e-07,1.904469e-07,1.904471e-07,1.904474e-07,1.904477e-07,1.904479e-07,1.904482e-07,1.904484e-07,1.904487e-07,1.904490e-07,1.904492e-07,1.904495e-07,1.904498e-07,1.904500e-07,1.904503e-07,1.904506e-07,1.904508e-07,1.904511e-07,1.904513e-07,1.904516e-07,1.904519e-07,1.904521e-07,1.904524e-07,1.904527e-07,1.904529e-07,1.904532e-07,1.904535e-07,1.904537e-07,1.904540e-07,1.904543e-07,1.904545e-07,1.904548e-07,1.904550e-07,1.904553e-07,1.904556e-07,1.904558e-07,1.904561e-07,1.904564e-07,1.904566e-07,1.904569e-07,1.904572e-07,1.904574e-07,1.904577e-07,1.904579e-07,1.904582e-07,1.904585e-07,1.904587e-07,1.904590e-07,1.904593e-07,1.904595e-07,1.904598e-07,1.904601e-07,1.904603e-07,1.904606e-07,1.904609e-07,1.904611e-07,1.904614e-07,1.904616e-07,1.904619e-07,1.904622e-07,1.904624e-07,1.904627e-07,1.904630e-07,1.904632e-07,1.904635e-07,1.904638e-07,1.904640e-07,1.904643e-07,1.904645e-07,1.904648e-07,1.904651e-07,1.904653e-07,1.904656e-07,1.904659e-07,1.904661e-07,1.904664e-07,1.904667e-07,1.904669e-07,1.904672e-07,1.904674e-07,1.904677e-07,1.904680e-07,1.904682e-07,1.904685e-07,1.904688e-07,1.904690e-07,1.904693e-07,1.904696e-07,1.904698e-07,1.904701e-07,1.904703e-07,1.904706e-07,1.904709e-07,1.904711e-07,1.904714e-07,1.904717e-07,1.904719e-07,1.904722e-07,1.904725e-07,1.904727e-07,1.904730e-07,1.904732e-07,1.904735e-07,1.904738e-07,1.904740e-07,1.904743e-07,1.904746e-07,1.904748e-07,1.904751e-07,1.904754e-07,1.904756e-07,1.904759e-07,1.904761e-07,1.904764e-07,1.904767e-07,1.904769e-07,1.904772e-07,1.904775e-07,1.904777e-07,1.904780e-07,1.904783e-07,1.904785e-07,1.904788e-07,1.904790e-07,1.904793e-07,1.904796e-07,1.904798e-07,1.904801e-07,1.904804e-07,1.904806e-07,1.904809e-07,1.904812e-07,1.904814e-07,1.904817e-07,1.904819e-07,1.904822e-07,1.904825e-07,1.904827e-07,1.904830e-07,1.904833e-07,1.904835e-07,1.904838e-07,1.904841e-07,1.904843e-07,1.904846e-07,1.904848e-07,1.904851e-07,1.904854e-07,1.904856e-07,1.904859e-07,1.904862e-07,1.904864e-07,1.904867e-07,1.904869e-07,1.904872e-07,1.904875e-07,1.904877e-07,1.904880e-07,1.904883e-07,1.904885e-07,1.904888e-07,1.904891e-07,1.904893e-07,1.904896e-07,1.904898e-07,1.904901e-07,1.904904e-07,1.904906e-07,1.904909e-07,1.904912e-07,1.904914e-07,1.904917e-07,1.904919e-07,1.904922e-07,1.904925e-07,1.904927e-07,1.904930e-07,1.904933e-07,1.904935e-07,1.904938e-07,1.904941e-07,1.904943e-07,1.904946e-07,1.904948e-07,1.904951e-07,1.904954e-07,1.904956e-07,1.904959e-07,1.904962e-07,1.904964e-07,1.904967e-07,1.904969e-07,1.904972e-07,1.904975e-07,1.904977e-07,1.904980e-07,1.904983e-07,1.904985e-07,1.904988e-07,1.904991e-07,1.904993e-07,1.904996e-07,1.904998e-07,1.905001e-07,1.905004e-07,1.905006e-07,1.905009e-07,1.905012e-07,1.905014e-07,1.905017e-07,1.905019e-07,1.905022e-07,1.905025e-07,1.905027e-07,1.905030e-07,1.905033e-07,1.905035e-07,1.905038e-07,1.905040e-07,1.905043e-07,1.905046e-07,1.905048e-07,1.905051e-07,1.905054e-07,1.905056e-07,1.905059e-07,1.905062e-07,1.905064e-07,1.905067e-07,1.905069e-07,1.905072e-07,1.905075e-07,1.905077e-07,1.905080e-07,1.905083e-07,1.905085e-07,1.905088e-07,1.905090e-07,1.905093e-07,1.905096e-07,1.905098e-07,1.905101e-07,1.905104e-07,1.905106e-07,1.905109e-07,1.905111e-07,1.905114e-07,1.905117e-07,1.905119e-07,1.905122e-07,1.905125e-07,1.905127e-07,1.905130e-07,1.905132e-07,1.905135e-07,1.905138e-07,1.905140e-07,1.905143e-07,1.905146e-07,1.905148e-07,1.905151e-07,1.905153e-07,1.905156e-07,1.905159e-07,1.905161e-07,1.905164e-07,1.905167e-07,1.905169e-07,1.905172e-07,1.905174e-07,1.905177e-07,1.905180e-07,1.905182e-07,1.905185e-07,1.905188e-07,1.905190e-07,1.905193e-07,1.905195e-07,1.905198e-07,1.905201e-07,1.905203e-07,1.905206e-07,1.905209e-07,1.905211e-07,1.905214e-07,1.905216e-07,1.905219e-07,1.905222e-07,1.905224e-07,1.905227e-07,1.905230e-07,1.905232e-07,1.905235e-07,1.905237e-07,1.905240e-07,1.905243e-07,1.905245e-07,1.905248e-07,1.905251e-07,1.905253e-07,1.905256e-07,1.905258e-07,1.905261e-07,1.905264e-07,1.905266e-07,1.905269e-07,1.905272e-07,1.905274e-07,1.905277e-07,1.905279e-07,1.905282e-07,1.905285e-07,1.905287e-07,1.905290e-07,1.905293e-07,1.905295e-07,1.905298e-07,1.905300e-07,1.905303e-07,1.905306e-07,1.905308e-07,1.905311e-07,1.905314e-07,1.905316e-07,1.905319e-07,1.905321e-07,1.905324e-07,1.905327e-07,1.905329e-07,1.905332e-07,1.905335e-07,1.905337e-07,1.905340e-07,1.905342e-07,1.905345e-07,1.905348e-07,1.905350e-07,1.905353e-07,1.905356e-07,1.905358e-07,1.905361e-07,1.905363e-07,1.905366e-07,1.905369e-07,1.905371e-07,1.905374e-07,1.905377e-07,1.905379e-07,1.905382e-07,1.905384e-07,1.905387e-07,1.905390e-07,1.905392e-07,1.905395e-07,1.905397e-07,1.905400e-07,1.905403e-07,1.905405e-07,1.905408e-07,1.905411e-07,1.905413e-07,1.905416e-07,1.905418e-07,1.905421e-07,1.905424e-07,1.905426e-07,1.905429e-07,1.905432e-07,1.905434e-07,1.905437e-07,1.905439e-07,1.905442e-07,1.905445e-07,1.905447e-07,1.905450e-07,1.905453e-07,1.905455e-07,1.905458e-07,1.905460e-07,1.905463e-07,1.905466e-07,1.905468e-07,1.905471e-07,1.905473e-07,1.905476e-07,1.905479e-07,1.905481e-07,1.905484e-07,1.905487e-07,1.905489e-07,1.905492e-07,1.905494e-07,1.905497e-07,1.905500e-07,1.905502e-07,1.905505e-07,1.905508e-07,1.905510e-07,1.905513e-07,1.905515e-07,1.905518e-07,1.905521e-07,1.905523e-07,1.905526e-07,1.905528e-07,1.905531e-07,1.905534e-07,1.905536e-07,1.905539e-07,1.905542e-07,1.905544e-07,1.905547e-07,1.905549e-07,1.905552e-07,1.905555e-07,1.905557e-07,1.905560e-07,1.905562e-07,1.905565e-07,1.905568e-07,1.905570e-07,1.905573e-07,1.905576e-07,1.905578e-07,1.905581e-07,1.905583e-07,1.905586e-07,1.905589e-07,1.905591e-07,1.905594e-07,1.905597e-07,1.905599e-07,1.905602e-07,1.905604e-07,1.905607e-07,1.905610e-07,1.905612e-07,1.905615e-07,1.905617e-07,1.905620e-07,1.905623e-07,1.905625e-07,1.905628e-07,1.905631e-07,1.905633e-07,1.905636e-07,1.905638e-07,1.905641e-07,1.905644e-07,1.905646e-07,1.905649e-07,1.905651e-07,1.905654e-07,1.905657e-07,1.905659e-07,1.905662e-07,1.905665e-07,1.905667e-07,1.905670e-07,1.905672e-07,1.905675e-07,1.905678e-07,1.905680e-07,1.905683e-07,1.905685e-07,1.905688e-07,1.905691e-07,1.905693e-07,1.905696e-07,1.905699e-07,1.905701e-07,1.905704e-07,1.905706e-07,1.905709e-07,1.905712e-07,1.905714e-07,1.905717e-07,1.905719e-07,1.905722e-07,1.905725e-07,1.905727e-07,1.905730e-07,1.905733e-07,1.905735e-07,1.905738e-07,1.905740e-07,1.905743e-07,1.905746e-07,1.905748e-07,1.905751e-07,1.905753e-07,1.905756e-07,1.905759e-07,1.905761e-07,1.905764e-07,1.905766e-07,1.905769e-07,1.905772e-07,1.905774e-07,1.905777e-07,1.905780e-07,1.905782e-07,1.905785e-07,1.905787e-07,1.905790e-07,1.905793e-07,1.905795e-07,1.905798e-07,1.905800e-07,1.905803e-07,1.905806e-07,1.905808e-07,1.905811e-07,1.905813e-07,1.905816e-07,1.905819e-07,1.905821e-07,1.905824e-07,1.905827e-07,1.905829e-07,1.905832e-07,1.905834e-07,1.905837e-07,1.905840e-07,1.905842e-07,1.905845e-07,1.905847e-07,1.905850e-07,1.905853e-07,1.905855e-07,1.905858e-07,1.905860e-07,1.905863e-07,1.905866e-07,1.905868e-07,1.905871e-07,1.905874e-07,1.905876e-07,1.905879e-07,1.905881e-07,1.905884e-07,1.905887e-07,1.905889e-07,1.905892e-07,1.905894e-07,1.905897e-07,1.905900e-07,1.905902e-07,1.905905e-07,1.905907e-07,1.905910e-07,1.905913e-07,1.905915e-07,1.905918e-07,1.905921e-07,1.905923e-07,1.905926e-07,1.905928e-07,1.905931e-07,1.905934e-07,1.905936e-07,1.905939e-07,1.905941e-07,1.905944e-07,1.905947e-07,1.905949e-07,1.905952e-07,1.905954e-07,1.905957e-07,1.905960e-07,1.905962e-07,1.905965e-07,1.905967e-07,1.905970e-07,1.905973e-07,1.905975e-07,1.905978e-07,1.905981e-07,1.905983e-07,1.905986e-07,1.905988e-07,1.905991e-07,1.905994e-07,1.905996e-07,1.905999e-07,1.906001e-07,1.906004e-07,1.906007e-07,1.906009e-07,1.906012e-07,1.906014e-07,1.906017e-07,1.906020e-07,1.906022e-07,1.906025e-07,1.906027e-07,1.906030e-07,1.906033e-07,1.906035e-07,1.906038e-07,1.906040e-07,1.906043e-07,1.906046e-07,1.906048e-07,1.906051e-07,1.906054e-07,1.906056e-07,1.906059e-07,1.906061e-07,1.906064e-07,1.906067e-07,1.906069e-07,1.906072e-07,1.906074e-07,1.906077e-07,1.906080e-07,1.906082e-07,1.906085e-07,1.906087e-07,1.906090e-07,1.906093e-07,1.906095e-07,1.906098e-07,1.906100e-07,1.906103e-07,1.906106e-07,1.906108e-07,1.906111e-07,1.906113e-07,1.906116e-07,1.906119e-07,1.906121e-07,1.906124e-07,1.906126e-07,1.906129e-07,1.906132e-07,1.906134e-07,1.906137e-07,1.906140e-07,1.906142e-07,1.906145e-07,1.906147e-07,1.906150e-07,1.906153e-07,1.906155e-07,1.906158e-07,1.906160e-07,1.906163e-07,1.906166e-07,1.906168e-07,1.906171e-07,1.906173e-07,1.906176e-07,1.906179e-07,1.906181e-07,1.906184e-07,1.906186e-07,1.906189e-07,1.906192e-07,1.906194e-07,1.906197e-07,1.906199e-07,1.906202e-07,1.906205e-07,1.906207e-07,1.906210e-07,1.906212e-07,1.906215e-07,1.906218e-07,1.906220e-07,1.906223e-07,1.906225e-07,1.906228e-07,1.906231e-07,1.906233e-07,1.906236e-07,1.906238e-07,1.906241e-07,1.906244e-07,1.906246e-07,1.906249e-07,1.906251e-07,1.906254e-07,1.906257e-07,1.906259e-07,1.906262e-07,1.906264e-07,1.906267e-07,1.906270e-07,1.906272e-07,1.906275e-07,1.906277e-07,1.906280e-07,1.906283e-07,1.906285e-07,1.906288e-07,1.906290e-07,1.906293e-07,1.906296e-07,1.906298e-07,1.906301e-07,1.906303e-07,1.906306e-07,1.906309e-07,1.906311e-07,1.906314e-07,1.906316e-07,1.906319e-07,1.906322e-07,1.906324e-07,1.906327e-07,1.906329e-07,1.906332e-07,1.906335e-07,1.906337e-07,1.906340e-07,1.906342e-07,1.906345e-07,1.906348e-07,1.906350e-07,1.906353e-07,1.906355e-07,1.906358e-07,1.906361e-07,1.906363e-07,1.906366e-07,1.906368e-07,1.906371e-07,1.906374e-07,1.906376e-07,1.906379e-07,1.906381e-07,1.906384e-07,1.906387e-07,1.906389e-07,1.906392e-07,1.906394e-07,1.906397e-07,1.906400e-07,1.906402e-07,1.906405e-07,1.906407e-07,1.906410e-07,1.906413e-07,1.906415e-07,1.906418e-07,1.906420e-07,1.906423e-07,1.906426e-07,1.906428e-07,1.906431e-07,1.906433e-07,1.906436e-07,1.906439e-07,1.906441e-07,1.906444e-07,1.906446e-07,1.906449e-07,1.906452e-07,1.906454e-07,1.906457e-07,1.906459e-07,1.906462e-07,1.906465e-07,1.906467e-07,1.906470e-07,1.906472e-07,1.906475e-07,1.906478e-07,1.906480e-07,1.906483e-07,1.906485e-07,1.906488e-07,1.906491e-07,1.906493e-07,1.906496e-07,1.906498e-07,1.906501e-07,1.906504e-07,1.906506e-07,1.906509e-07,1.906511e-07,1.906514e-07,1.906517e-07,1.906519e-07,1.906522e-07,1.906524e-07,1.906527e-07,1.906530e-07,1.906532e-07,1.906535e-07,1.906537e-07,1.906540e-07,1.906543e-07,1.906545e-07,1.906548e-07,1.906550e-07,1.906553e-07,1.906555e-07,1.906558e-07,1.906561e-07,1.906563e-07,1.906566e-07,1.906568e-07,1.906571e-07,1.906574e-07,1.906576e-07,1.906579e-07,1.906581e-07,1.906584e-07,1.906587e-07,1.906589e-07,1.906592e-07,1.906594e-07,1.906597e-07,1.906600e-07,1.906602e-07,1.906605e-07,1.906607e-07,1.906610e-07,1.906613e-07,1.906615e-07,1.906618e-07,1.906620e-07,1.906623e-07,1.906626e-07,1.906628e-07,1.906631e-07,1.906633e-07,1.906636e-07,1.906638e-07,1.906641e-07,1.906644e-07,1.906646e-07,1.906649e-07,1.906651e-07,1.906654e-07,1.906657e-07,1.906659e-07,1.906662e-07,1.906664e-07,1.906667e-07,1.906670e-07,1.906672e-07,1.906675e-07,1.906677e-07,1.906680e-07,1.906683e-07,1.906685e-07,1.906688e-07,1.906690e-07,1.906693e-07,1.906696e-07,1.906698e-07,1.906701e-07,1.906703e-07,1.906706e-07,1.906708e-07,1.906711e-07,1.906714e-07,1.906716e-07,1.906719e-07,1.906721e-07,1.906724e-07,1.906727e-07,1.906729e-07,1.906732e-07,1.906734e-07,1.906737e-07,1.906740e-07,1.906742e-07,1.906745e-07,1.906747e-07,1.906750e-07,1.906753e-07,1.906755e-07,1.906758e-07,1.906760e-07,1.906763e-07,1.906766e-07,1.906768e-07,1.906771e-07,1.906773e-07,1.906776e-07,1.906778e-07,1.906781e-07,1.906784e-07,1.906786e-07,1.906789e-07,1.906791e-07,1.906794e-07,1.906797e-07,1.906799e-07,1.906802e-07,1.906804e-07,1.906807e-07,1.906810e-07,1.906812e-07,1.906815e-07,1.906817e-07,1.906820e-07,1.906822e-07,1.906825e-07,1.906828e-07,1.906830e-07,1.906833e-07,1.906835e-07,1.906838e-07,1.906841e-07,1.906843e-07,1.906846e-07,1.906848e-07,1.906851e-07,1.906854e-07,1.906856e-07,1.906859e-07,1.906861e-07,1.906864e-07,1.906866e-07,1.906869e-07,1.906872e-07,1.906874e-07,1.906877e-07,1.906879e-07,1.906882e-07,1.906885e-07,1.906887e-07,1.906890e-07,1.906892e-07,1.906895e-07,1.906898e-07,1.906900e-07,1.906903e-07,1.906905e-07,1.906908e-07,1.906910e-07,1.906913e-07,1.906916e-07,1.906918e-07,1.906921e-07,1.906923e-07,1.906926e-07,1.906929e-07,1.906931e-07,1.906934e-07,1.906936e-07,1.906939e-07,1.906942e-07,1.906944e-07,1.906947e-07,1.906949e-07,1.906952e-07,1.906954e-07,1.906957e-07,1.906960e-07,1.906962e-07,1.906965e-07,1.906967e-07,1.906970e-07,1.906973e-07,1.906975e-07,1.906978e-07,1.906980e-07,1.906983e-07,1.906985e-07,1.906988e-07,1.906991e-07,1.906993e-07,1.906996e-07,1.906998e-07,1.907001e-07,1.907004e-07,1.907006e-07,1.907009e-07,1.907011e-07,1.907014e-07,1.907017e-07,1.907019e-07,1.907022e-07,1.907024e-07,1.907027e-07,1.907029e-07,1.907032e-07,1.907035e-07,1.907037e-07,1.907040e-07,1.907042e-07,1.907045e-07,1.907048e-07,1.907050e-07,1.907053e-07,1.907055e-07,1.907058e-07,1.907060e-07,1.907063e-07,1.907066e-07,1.907068e-07,1.907071e-07,1.907073e-07,1.907076e-07,1.907079e-07,1.907081e-07,1.907084e-07,1.907086e-07,1.907089e-07,1.907091e-07,1.907094e-07,1.907097e-07,1.907099e-07,1.907102e-07,1.907104e-07,1.907107e-07,1.907110e-07,1.907112e-07,1.907115e-07,1.907117e-07,1.907120e-07,1.907122e-07,1.907125e-07,1.907128e-07,1.907130e-07,1.907133e-07,1.907135e-07,1.907138e-07,1.907141e-07,1.907143e-07,1.907146e-07,1.907148e-07,1.907151e-07,1.907153e-07,1.907156e-07,1.907159e-07,1.907161e-07,1.907164e-07,1.907166e-07,1.907169e-07,1.907172e-07,1.907174e-07,1.907177e-07,1.907179e-07,1.907182e-07,1.907184e-07,1.907187e-07,1.907190e-07,1.907192e-07,1.907195e-07,1.907197e-07,1.907200e-07,1.907202e-07,1.907205e-07,1.907208e-07,1.907210e-07,1.907213e-07,1.907215e-07,1.907218e-07,1.907221e-07,1.907223e-07,1.907226e-07,1.907228e-07,1.907231e-07,1.907233e-07,1.907236e-07,1.907239e-07,1.907241e-07,1.907244e-07,1.907246e-07,1.907249e-07,1.907252e-07,1.907254e-07,1.907257e-07,1.907259e-07,1.907262e-07,1.907264e-07,1.907267e-07,1.907270e-07,1.907272e-07,1.907275e-07,1.907277e-07,1.907280e-07,1.907282e-07,1.907285e-07,1.907288e-07,1.907290e-07,1.907293e-07,1.907295e-07,1.907298e-07,1.907301e-07,1.907303e-07,1.907306e-07,1.907308e-07,1.907311e-07,1.907313e-07,1.907316e-07,1.907319e-07,1.907321e-07,1.907324e-07,1.907326e-07,1.907329e-07,1.907331e-07,1.907334e-07,1.907337e-07,1.907339e-07,1.907342e-07,1.907344e-07,1.907347e-07,1.907350e-07,1.907352e-07,1.907355e-07,1.907357e-07,1.907360e-07,1.907362e-07,1.907365e-07,1.907368e-07,1.907370e-07,1.907373e-07,1.907375e-07,1.907378e-07,1.907380e-07,1.907383e-07,1.907386e-07,1.907388e-07,1.907391e-07,1.907393e-07,1.907396e-07,1.907398e-07,1.907401e-07,1.907404e-07,1.907406e-07,1.907409e-07,1.907411e-07,1.907414e-07,1.907417e-07,1.907419e-07,1.907422e-07,1.907424e-07,1.907427e-07,1.907429e-07,1.907432e-07,1.907435e-07,1.907437e-07,1.907440e-07,1.907442e-07,1.907445e-07,1.907447e-07,1.907450e-07,1.907453e-07,1.907455e-07,1.907458e-07,1.907460e-07,1.907463e-07,1.907465e-07,1.907468e-07,1.907471e-07,1.907473e-07,1.907476e-07,1.907478e-07,1.907481e-07,1.907483e-07,1.907486e-07,1.907489e-07,1.907491e-07,1.907494e-07,1.907496e-07,1.907499e-07,1.907501e-07,1.907504e-07,1.907507e-07,1.907509e-07,1.907512e-07,1.907514e-07,1.907517e-07,1.907520e-07,1.907522e-07,1.907525e-07,1.907527e-07,1.907530e-07,1.907532e-07,1.907535e-07,1.907538e-07,1.907540e-07,1.907543e-07,1.907545e-07,1.907548e-07,1.907550e-07,1.907553e-07,1.907556e-07,1.907558e-07,1.907561e-07,1.907563e-07,1.907566e-07,1.907568e-07,1.907571e-07,1.907574e-07,1.907576e-07,1.907579e-07,1.907581e-07,1.907584e-07,1.907586e-07,1.907589e-07,1.907592e-07,1.907594e-07,1.907597e-07,1.907599e-07,1.907602e-07,1.907604e-07,1.907607e-07,1.907610e-07,1.907612e-07,1.907615e-07,1.907617e-07,1.907620e-07,1.907622e-07,1.907625e-07,1.907628e-07,1.907630e-07,1.907633e-07,1.907635e-07,1.907638e-07,1.907640e-07,1.907643e-07,1.907646e-07,1.907648e-07,1.907651e-07,1.907653e-07,1.907656e-07,1.907658e-07,1.907661e-07,1.907664e-07,1.907666e-07,1.907669e-07,1.907671e-07,1.907674e-07,1.907676e-07,1.907679e-07,1.907682e-07,1.907684e-07,1.907687e-07,1.907689e-07,1.907692e-07,1.907694e-07,1.907697e-07,1.907700e-07,1.907702e-07,1.907705e-07,1.907707e-07,1.907710e-07,1.907712e-07,1.907715e-07,1.907718e-07,1.907720e-07,1.907723e-07,1.907725e-07,1.907728e-07,1.907730e-07,1.907733e-07,1.907736e-07,1.907738e-07,1.907741e-07,1.907743e-07,1.907746e-07,1.907748e-07,1.907751e-07,1.907754e-07,1.907756e-07,1.907759e-07,1.907761e-07,1.907764e-07,1.907766e-07,1.907769e-07,1.907771e-07,1.907774e-07,1.907777e-07,1.907779e-07,1.907782e-07,1.907784e-07,1.907787e-07,1.907789e-07,1.907792e-07,1.907795e-07,1.907797e-07,1.907800e-07,1.907802e-07,1.907805e-07,1.907807e-07,1.907810e-07,1.907813e-07,1.907815e-07,1.907818e-07,1.907820e-07,1.907823e-07,1.907825e-07,1.907828e-07,1.907831e-07,1.907833e-07,1.907836e-07,1.907838e-07,1.907841e-07,1.907843e-07,1.907846e-07,1.907849e-07,1.907851e-07,1.907854e-07,1.907856e-07,1.907859e-07,1.907861e-07,1.907864e-07,1.907866e-07,1.907869e-07,1.907872e-07,1.907874e-07,1.907877e-07,1.907879e-07,1.907882e-07,1.907884e-07,1.907887e-07,1.907890e-07,1.907892e-07,1.907895e-07,1.907897e-07,1.907900e-07,1.907902e-07,1.907905e-07,1.907908e-07,1.907910e-07,1.907913e-07,1.907915e-07,1.907918e-07,1.907920e-07,1.907923e-07,1.907925e-07,1.907928e-07,1.907931e-07,1.907933e-07,1.907936e-07,1.907938e-07,1.907941e-07,1.907943e-07,1.907946e-07,1.907949e-07,1.907951e-07,1.907954e-07,1.907956e-07,1.907959e-07,1.907961e-07,1.907964e-07,1.907967e-07,1.907969e-07,1.907972e-07,1.907974e-07,1.907977e-07,1.907979e-07,1.907982e-07,1.907984e-07,1.907987e-07,1.907990e-07,1.907992e-07,1.907995e-07,1.907997e-07,1.908000e-07,1.908002e-07,1.908005e-07,1.908008e-07,1.908010e-07,1.908013e-07,1.908015e-07,1.908018e-07,1.908020e-07,1.908023e-07,1.908025e-07,1.908028e-07,1.908031e-07,1.908033e-07,1.908036e-07,1.908038e-07,1.908041e-07,1.908043e-07,1.908046e-07,1.908049e-07,1.908051e-07,1.908054e-07,1.908056e-07,1.908059e-07,1.908061e-07,1.908064e-07,1.908066e-07,1.908069e-07,1.908072e-07,1.908074e-07,1.908077e-07,1.908079e-07,1.908082e-07,1.908084e-07,1.908087e-07,1.908090e-07,1.908092e-07,1.908095e-07,1.908097e-07,1.908100e-07,1.908102e-07,1.908105e-07,1.908107e-07,1.908110e-07,1.908113e-07,1.908115e-07,1.908118e-07,1.908120e-07,1.908123e-07,1.908125e-07,1.908128e-07,1.908131e-07,1.908133e-07,1.908136e-07,1.908138e-07,1.908141e-07,1.908143e-07,1.908146e-07,1.908148e-07,1.908151e-07,1.908154e-07,1.908156e-07,1.908159e-07,1.908161e-07,1.908164e-07,1.908166e-07,1.908169e-07,1.908171e-07,1.908174e-07,1.908177e-07,1.908179e-07,1.908182e-07,1.908184e-07,1.908187e-07,1.908189e-07,1.908192e-07,1.908194e-07,1.908197e-07,1.908200e-07,1.908202e-07,1.908205e-07,1.908207e-07,1.908210e-07,1.908212e-07,1.908215e-07,1.908218e-07,1.908220e-07,1.908223e-07,1.908225e-07,1.908228e-07,1.908230e-07,1.908233e-07,1.908235e-07,1.908238e-07,1.908241e-07,1.908243e-07,1.908246e-07,1.908248e-07,1.908251e-07,1.908253e-07,1.908256e-07,1.908258e-07,1.908261e-07,1.908264e-07,1.908266e-07,1.908269e-07,1.908271e-07,1.908274e-07,1.908276e-07,1.908279e-07,1.908281e-07,1.908284e-07,1.908287e-07,1.908289e-07,1.908292e-07,1.908294e-07,1.908297e-07,1.908299e-07,1.908302e-07,1.908304e-07,1.908307e-07,1.908310e-07,1.908312e-07,1.908315e-07,1.908317e-07,1.908320e-07,1.908322e-07,1.908325e-07,1.908327e-07,1.908330e-07,1.908333e-07,1.908335e-07,1.908338e-07,1.908340e-07,1.908343e-07,1.908345e-07,1.908348e-07,1.908350e-07,1.908353e-07,1.908356e-07,1.908358e-07,1.908361e-07,1.908363e-07,1.908366e-07,1.908368e-07,1.908371e-07,1.908373e-07,1.908376e-07,1.908379e-07,1.908381e-07,1.908384e-07,1.908386e-07,1.908389e-07,1.908391e-07,1.908394e-07,1.908396e-07,1.908399e-07,1.908402e-07,1.908404e-07,1.908407e-07,1.908409e-07,1.908412e-07,1.908414e-07,1.908417e-07,1.908419e-07,1.908422e-07,1.908425e-07,1.908427e-07,1.908430e-07,1.908432e-07,1.908435e-07,1.908437e-07,1.908440e-07,1.908442e-07,1.908445e-07,1.908448e-07,1.908450e-07,1.908453e-07,1.908455e-07,1.908458e-07,1.908460e-07,1.908463e-07,1.908465e-07,1.908468e-07,1.908471e-07,1.908473e-07,1.908476e-07,1.908478e-07,1.908481e-07,1.908483e-07,1.908486e-07,1.908488e-07,1.908491e-07,1.908494e-07,1.908496e-07,1.908499e-07,1.908501e-07,1.908504e-07,1.908506e-07,1.908509e-07,1.908511e-07,1.908514e-07,1.908516e-07,1.908519e-07,1.908522e-07,1.908524e-07,1.908527e-07,1.908529e-07,1.908532e-07,1.908534e-07,1.908537e-07,1.908539e-07,1.908542e-07,1.908545e-07,1.908547e-07,1.908550e-07,1.908552e-07,1.908555e-07,1.908557e-07,1.908560e-07,1.908562e-07,1.908565e-07,1.908568e-07,1.908570e-07,1.908573e-07,1.908575e-07,1.908578e-07,1.908580e-07,1.908583e-07,1.908585e-07,1.908588e-07,1.908590e-07,1.908593e-07,1.908596e-07,1.908598e-07,1.908601e-07,1.908603e-07,1.908606e-07,1.908608e-07,1.908611e-07,1.908613e-07,1.908616e-07,1.908619e-07,1.908621e-07,1.908624e-07,1.908626e-07,1.908629e-07,1.908631e-07,1.908634e-07,1.908636e-07,1.908639e-07,1.908641e-07,1.908644e-07,1.908647e-07,1.908649e-07,1.908652e-07,1.908654e-07,1.908657e-07,1.908659e-07,1.908662e-07,1.908664e-07,1.908667e-07,1.908670e-07,1.908672e-07,1.908675e-07,1.908677e-07,1.908680e-07,1.908682e-07,1.908685e-07,1.908687e-07,1.908690e-07,1.908692e-07,1.908695e-07,1.908698e-07,1.908700e-07,1.908703e-07,1.908705e-07,1.908708e-07,1.908710e-07,1.908713e-07,1.908715e-07,1.908718e-07,1.908720e-07,1.908723e-07,1.908726e-07,1.908728e-07,1.908731e-07,1.908733e-07,1.908736e-07,1.908738e-07,1.908741e-07,1.908743e-07,1.908746e-07,1.908749e-07,1.908751e-07,1.908754e-07,1.908756e-07,1.908759e-07,1.908761e-07,1.908764e-07,1.908766e-07,1.908769e-07,1.908771e-07,1.908774e-07,1.908777e-07,1.908779e-07,1.908782e-07,1.908784e-07,1.908787e-07,1.908789e-07,1.908792e-07,1.908794e-07,1.908797e-07,1.908799e-07,1.908802e-07,1.908805e-07,1.908807e-07,1.908810e-07,1.908812e-07,1.908815e-07,1.908817e-07,1.908820e-07,1.908822e-07,1.908825e-07,1.908827e-07,1.908830e-07,1.908833e-07,1.908835e-07,1.908838e-07,1.908840e-07,1.908843e-07,1.908845e-07,1.908848e-07,1.908850e-07,1.908853e-07,1.908855e-07,1.908858e-07,1.908861e-07,1.908863e-07,1.908866e-07,1.908868e-07,1.908871e-07,1.908873e-07,1.908876e-07,1.908878e-07,1.908881e-07,1.908883e-07,1.908886e-07,1.908889e-07,1.908891e-07,1.908894e-07,1.908896e-07,1.908899e-07,1.908901e-07,1.908904e-07,1.908906e-07,1.908909e-07,1.908911e-07,1.908914e-07,1.908916e-07,1.908919e-07,1.908922e-07,1.908924e-07,1.908927e-07,1.908929e-07,1.908932e-07,1.908934e-07,1.908937e-07,1.908939e-07,1.908942e-07,1.908944e-07,1.908947e-07,1.908950e-07,1.908952e-07,1.908955e-07,1.908957e-07,1.908960e-07,1.908962e-07,1.908965e-07,1.908967e-07,1.908970e-07,1.908972e-07,1.908975e-07,1.908978e-07,1.908980e-07,1.908983e-07,1.908985e-07,1.908988e-07,1.908990e-07,1.908993e-07,1.908995e-07,1.908998e-07,1.909000e-07,1.909003e-07,1.909005e-07,1.909008e-07,1.909011e-07,1.909013e-07,1.909016e-07,1.909018e-07,1.909021e-07,1.909023e-07,1.909026e-07,1.909028e-07,1.909031e-07,1.909033e-07,1.909036e-07,1.909039e-07,1.909041e-07,1.909044e-07,1.909046e-07,1.909049e-07,1.909051e-07,1.909054e-07,1.909056e-07,1.909059e-07,1.909061e-07,1.909064e-07,1.909066e-07,1.909069e-07,1.909072e-07,1.909074e-07,1.909077e-07,1.909079e-07,1.909082e-07,1.909084e-07,1.909087e-07,1.909089e-07,1.909092e-07,1.909094e-07,1.909097e-07,1.909099e-07,1.909102e-07,1.909105e-07,1.909107e-07,1.909110e-07,1.909112e-07,1.909115e-07,1.909117e-07,1.909120e-07,1.909122e-07,1.909125e-07,1.909127e-07,1.909130e-07,1.909132e-07,1.909135e-07,1.909138e-07,1.909140e-07,1.909143e-07,1.909145e-07,1.909148e-07,1.909150e-07,1.909153e-07,1.909155e-07,1.909158e-07,1.909160e-07,1.909163e-07,1.909165e-07,1.909168e-07,1.909171e-07,1.909173e-07,1.909176e-07,1.909178e-07,1.909181e-07,1.909183e-07,1.909186e-07,1.909188e-07,1.909191e-07,1.909193e-07,1.909196e-07,1.909198e-07,1.909201e-07,1.909204e-07,1.909206e-07,1.909209e-07,1.909211e-07,1.909214e-07,1.909216e-07,1.909219e-07,1.909221e-07,1.909224e-07,1.909226e-07,1.909229e-07,1.909231e-07,1.909234e-07,1.909237e-07,1.909239e-07,1.909242e-07,1.909244e-07,1.909247e-07,1.909249e-07,1.909252e-07,1.909254e-07,1.909257e-07,1.909259e-07,1.909262e-07,1.909264e-07,1.909267e-07,1.909269e-07,1.909272e-07,1.909275e-07,1.909277e-07,1.909280e-07,1.909282e-07,1.909285e-07,1.909287e-07,1.909290e-07,1.909292e-07,1.909295e-07,1.909297e-07,1.909300e-07,1.909302e-07,1.909305e-07,1.909308e-07,1.909310e-07,1.909313e-07,1.909315e-07,1.909318e-07,1.909320e-07,1.909323e-07,1.909325e-07,1.909328e-07,1.909330e-07,1.909333e-07,1.909335e-07,1.909338e-07,1.909340e-07,1.909343e-07,1.909346e-07,1.909348e-07,1.909351e-07,1.909353e-07,1.909356e-07,1.909358e-07,1.909361e-07,1.909363e-07,1.909366e-07,1.909368e-07,1.909371e-07,1.909373e-07,1.909376e-07,1.909378e-07,1.909381e-07,1.909384e-07,1.909386e-07,1.909389e-07,1.909391e-07,1.909394e-07,1.909396e-07,1.909399e-07,1.909401e-07,1.909404e-07,1.909406e-07,1.909409e-07,1.909411e-07,1.909414e-07,1.909416e-07,1.909419e-07,1.909422e-07,1.909424e-07,1.909427e-07,1.909429e-07,1.909432e-07,1.909434e-07,1.909437e-07,1.909439e-07,1.909442e-07,1.909444e-07,1.909447e-07,1.909449e-07,1.909452e-07,1.909454e-07,1.909457e-07,1.909459e-07,1.909462e-07,1.909465e-07,1.909467e-07,1.909470e-07,1.909472e-07,1.909475e-07,1.909477e-07,1.909480e-07,1.909482e-07,1.909485e-07,1.909487e-07,1.909490e-07,1.909492e-07,1.909495e-07,1.909497e-07,1.909500e-07,1.909503e-07,1.909505e-07,1.909508e-07,1.909510e-07,1.909513e-07,1.909515e-07,1.909518e-07,1.909520e-07,1.909523e-07,1.909525e-07,1.909528e-07,1.909530e-07,1.909533e-07,1.909535e-07,1.909538e-07,1.909540e-07,1.909543e-07,1.909546e-07,1.909548e-07,1.909551e-07,1.909553e-07,1.909556e-07,1.909558e-07,1.909561e-07,1.909563e-07,1.909566e-07,1.909568e-07,1.909571e-07,1.909573e-07,1.909576e-07,1.909578e-07,1.909581e-07,1.909583e-07,1.909586e-07,1.909589e-07,1.909591e-07,1.909594e-07,1.909596e-07,1.909599e-07,1.909601e-07,1.909604e-07,1.909606e-07,1.909609e-07,1.909611e-07,1.909614e-07,1.909616e-07,1.909619e-07,1.909621e-07,1.909624e-07,1.909626e-07,1.909629e-07,1.909632e-07,1.909634e-07,1.909637e-07,1.909639e-07,1.909642e-07,1.909644e-07,1.909647e-07,1.909649e-07,1.909652e-07,1.909654e-07,1.909657e-07,1.909659e-07,1.909662e-07,1.909664e-07,1.909667e-07,1.909669e-07,1.909672e-07,1.909674e-07,1.909677e-07,1.909680e-07,1.909682e-07,1.909685e-07,1.909687e-07,1.909690e-07,1.909692e-07,1.909695e-07,1.909697e-07,1.909700e-07,1.909702e-07,1.909705e-07,1.909707e-07,1.909710e-07,1.909712e-07,1.909715e-07,1.909717e-07,1.909720e-07,1.909722e-07,1.909725e-07,1.909728e-07,1.909730e-07,1.909733e-07,1.909735e-07,1.909738e-07,1.909740e-07,1.909743e-07,1.909745e-07,1.909748e-07,1.909750e-07,1.909753e-07,1.909755e-07,1.909758e-07,1.909760e-07,1.909763e-07,1.909765e-07,1.909768e-07,1.909770e-07,1.909773e-07,1.909776e-07,1.909778e-07,1.909781e-07,1.909783e-07,1.909786e-07,1.909788e-07,1.909791e-07,1.909793e-07,1.909796e-07,1.909798e-07,1.909801e-07,1.909803e-07,1.909806e-07,1.909808e-07,1.909811e-07,1.909813e-07,1.909816e-07,1.909818e-07,1.909821e-07,1.909823e-07,1.909826e-07,1.909829e-07,1.909831e-07,1.909834e-07,1.909836e-07,1.909839e-07,1.909841e-07,1.909844e-07,1.909846e-07,1.909849e-07,1.909851e-07,1.909854e-07,1.909856e-07,1.909859e-07,1.909861e-07,1.909864e-07,1.909866e-07,1.909869e-07,1.909871e-07,1.909874e-07,1.909876e-07,1.909879e-07,1.909882e-07,1.909884e-07,1.909887e-07,1.909889e-07,1.909892e-07,1.909894e-07,1.909897e-07,1.909899e-07,1.909902e-07,1.909904e-07,1.909907e-07,1.909909e-07,1.909912e-07,1.909914e-07,1.909917e-07,1.909919e-07,1.909922e-07,1.909924e-07,1.909927e-07,1.909929e-07,1.909932e-07,1.909934e-07,1.909937e-07,1.909940e-07,1.909942e-07,1.909945e-07,1.909947e-07,1.909950e-07,1.909952e-07,1.909955e-07,1.909957e-07,1.909960e-07,1.909962e-07,1.909965e-07,1.909967e-07,1.909970e-07,1.909972e-07,1.909975e-07,1.909977e-07,1.909980e-07,1.909982e-07,1.909985e-07,1.909987e-07,1.909990e-07,1.909992e-07,1.909995e-07,1.909997e-07,1.910000e-07,1.910003e-07,1.910005e-07,1.910008e-07,1.910010e-07,1.910013e-07,1.910015e-07,1.910018e-07,1.910020e-07,1.910023e-07,1.910025e-07,1.910028e-07,1.910030e-07,1.910033e-07,1.910035e-07,1.910038e-07,1.910040e-07,1.910043e-07,1.910045e-07,1.910048e-07,1.910050e-07,1.910053e-07,1.910055e-07,1.910058e-07,1.910060e-07,1.910063e-07,1.910066e-07,1.910068e-07,1.910071e-07,1.910073e-07,1.910076e-07,1.910078e-07,1.910081e-07,1.910083e-07,1.910086e-07,1.910088e-07,1.910091e-07,1.910093e-07,1.910096e-07,1.910098e-07,1.910101e-07,1.910103e-07,1.910106e-07,1.910108e-07,1.910111e-07,1.910113e-07,1.910116e-07,1.910118e-07,1.910121e-07,1.910123e-07,1.910126e-07,1.910128e-07,1.910131e-07,1.910133e-07,1.910136e-07,1.910139e-07,1.910141e-07,1.910144e-07,1.910146e-07,1.910149e-07,1.910151e-07,1.910154e-07,1.910156e-07,1.910159e-07,1.910161e-07,1.910164e-07,1.910166e-07,1.910169e-07,1.910171e-07,1.910174e-07,1.910176e-07,1.910179e-07,1.910181e-07,1.910184e-07,1.910186e-07,1.910189e-07,1.910191e-07,1.910194e-07,1.910196e-07,1.910199e-07,1.910201e-07,1.910204e-07,1.910206e-07,1.910209e-07,1.910211e-07,1.910214e-07,1.910217e-07,1.910219e-07,1.910222e-07,1.910224e-07,1.910227e-07,1.910229e-07,1.910232e-07,1.910234e-07,1.910237e-07,1.910239e-07,1.910242e-07,1.910244e-07,1.910247e-07,1.910249e-07,1.910252e-07,1.910254e-07,1.910257e-07,1.910259e-07,1.910262e-07,1.910264e-07,1.910267e-07,1.910269e-07,1.910272e-07,1.910274e-07,1.910277e-07,1.910279e-07,1.910282e-07,1.910284e-07,1.910287e-07,1.910289e-07,1.910292e-07,1.910294e-07,1.910297e-07,1.910299e-07,1.910302e-07,1.910305e-07,1.910307e-07,1.910310e-07,1.910312e-07,1.910315e-07,1.910317e-07,1.910320e-07,1.910322e-07,1.910325e-07,1.910327e-07,1.910330e-07,1.910332e-07,1.910335e-07,1.910337e-07,1.910340e-07,1.910342e-07,1.910345e-07,1.910347e-07,1.910350e-07,1.910352e-07,1.910355e-07,1.910357e-07,1.910360e-07,1.910362e-07,1.910365e-07,1.910367e-07,1.910370e-07,1.910372e-07,1.910375e-07,1.910377e-07,1.910380e-07,1.910382e-07,1.910385e-07,1.910387e-07,1.910390e-07,1.910392e-07,1.910395e-07,1.910397e-07,1.910400e-07,1.910402e-07,1.910405e-07,1.910408e-07,1.910410e-07,1.910413e-07,1.910415e-07,1.910418e-07,1.910420e-07,1.910423e-07,1.910425e-07,1.910428e-07,1.910430e-07,1.910433e-07,1.910435e-07,1.910438e-07,1.910440e-07,1.910443e-07,1.910445e-07,1.910448e-07,1.910450e-07,1.910453e-07,1.910455e-07,1.910458e-07,1.910460e-07,1.910463e-07,1.910465e-07,1.910468e-07,1.910470e-07,1.910473e-07,1.910475e-07,1.910478e-07,1.910480e-07,1.910483e-07,1.910485e-07,1.910488e-07,1.910490e-07,1.910493e-07,1.910495e-07,1.910498e-07,1.910500e-07,1.910503e-07,1.910505e-07,1.910508e-07,1.910510e-07,1.910513e-07,1.910515e-07,1.910518e-07,1.910520e-07,1.910523e-07,1.910525e-07,1.910528e-07,1.910530e-07,1.910533e-07,1.910536e-07,1.910538e-07,1.910541e-07,1.910543e-07,1.910546e-07,1.910548e-07,1.910551e-07,1.910553e-07,1.910556e-07,1.910558e-07,1.910561e-07,1.910563e-07,1.910566e-07,1.910568e-07,1.910571e-07,1.910573e-07,1.910576e-07,1.910578e-07,1.910581e-07,1.910583e-07,1.910586e-07,1.910588e-07,1.910591e-07,1.910593e-07,1.910596e-07,1.910598e-07,1.910601e-07,1.910603e-07,1.910606e-07,1.910608e-07,1.910611e-07,1.910613e-07,1.910616e-07,1.910618e-07,1.910621e-07,1.910623e-07,1.910626e-07,1.910628e-07,1.910631e-07,1.910633e-07,1.910636e-07,1.910638e-07,1.910641e-07,1.910643e-07,1.910646e-07,1.910648e-07,1.910651e-07,1.910653e-07,1.910656e-07,1.910658e-07,1.910661e-07,1.910663e-07,1.910666e-07,1.910668e-07,1.910671e-07,1.910673e-07,1.910676e-07,1.910678e-07,1.910681e-07,1.910683e-07,1.910686e-07,1.910688e-07,1.910691e-07,1.910693e-07,1.910696e-07,1.910698e-07,1.910701e-07,1.910703e-07,1.910706e-07,1.910708e-07,1.910711e-07,1.910713e-07,1.910716e-07,1.910718e-07,1.910721e-07,1.910723e-07,1.910726e-07,1.910728e-07,1.910731e-07,1.910734e-07,1.910736e-07,1.910739e-07,1.910741e-07,1.910744e-07,1.910746e-07,1.910749e-07,1.910751e-07,1.910754e-07,1.910756e-07,1.910759e-07,1.910761e-07,1.910764e-07,1.910766e-07,1.910769e-07,1.910771e-07,1.910774e-07,1.910776e-07,1.910779e-07,1.910781e-07,1.910784e-07,1.910786e-07,1.910789e-07,1.910791e-07,1.910794e-07,1.910796e-07,1.910799e-07,1.910801e-07,1.910804e-07,1.910806e-07,1.910809e-07,1.910811e-07,1.910814e-07,1.910816e-07,1.910819e-07,1.910821e-07,1.910824e-07,1.910826e-07,1.910829e-07,1.910831e-07,1.910834e-07,1.910836e-07,1.910839e-07,1.910841e-07,1.910844e-07,1.910846e-07,1.910849e-07,1.910851e-07,1.910854e-07,1.910856e-07,1.910859e-07,1.910861e-07,1.910864e-07,1.910866e-07,1.910869e-07,1.910871e-07,1.910874e-07,1.910876e-07,1.910879e-07,1.910881e-07,1.910884e-07,1.910886e-07,1.910889e-07,1.910891e-07,1.910894e-07,1.910896e-07,1.910899e-07,1.910901e-07,1.910904e-07,1.910906e-07,1.910909e-07,1.910911e-07,1.910914e-07,1.910916e-07,1.910919e-07,1.910921e-07,1.910924e-07,1.910926e-07,1.910929e-07,1.910931e-07,1.910934e-07,1.910936e-07,1.910939e-07,1.910941e-07,1.910944e-07,1.910946e-07,1.910949e-07,1.910951e-07,1.910954e-07,1.910956e-07,1.910959e-07,1.910961e-07,1.910964e-07,1.910966e-07,1.910969e-07,1.910971e-07,1.910974e-07,1.910976e-07,1.910979e-07,1.910981e-07,1.910984e-07,1.910986e-07,1.910989e-07,1.910991e-07,1.910994e-07,1.910996e-07,1.910999e-07,1.911001e-07,1.911004e-07,1.911006e-07,1.911009e-07,1.911011e-07,1.911014e-07,1.911016e-07,1.911019e-07,1.911021e-07,1.911024e-07,1.911026e-07,1.911029e-07,1.911031e-07,1.911034e-07,1.911036e-07,1.911039e-07,1.911041e-07,1.911044e-07,1.911046e-07,1.911049e-07,1.911051e-07,1.911054e-07,1.911056e-07,1.911059e-07,1.911061e-07,1.911064e-07,1.911066e-07,1.911069e-07,1.911071e-07,1.911074e-07,1.911076e-07,1.911079e-07,1.911081e-07,1.911084e-07,1.911086e-07,1.911089e-07,1.911091e-07,1.911094e-07,1.911096e-07,1.911099e-07,1.911101e-07,1.911104e-07,1.911106e-07,1.911109e-07,1.911111e-07,1.911114e-07,1.911116e-07,1.911119e-07,1.911121e-07,1.911124e-07,1.911126e-07,1.911128e-07,1.911131e-07,1.911133e-07,1.911136e-07,1.911138e-07,1.911141e-07,1.911143e-07,1.911146e-07,1.911148e-07,1.911151e-07,1.911153e-07,1.911156e-07,1.911158e-07,1.911161e-07,1.911163e-07,1.911166e-07,1.911168e-07,1.911171e-07,1.911173e-07,1.911176e-07,1.911178e-07,1.911181e-07,1.911183e-07,1.911186e-07,1.911188e-07,1.911191e-07,1.911193e-07,1.911196e-07,1.911198e-07,1.911201e-07,1.911203e-07,1.911206e-07,1.911208e-07,1.911211e-07,1.911213e-07,1.911216e-07,1.911218e-07,1.911221e-07,1.911223e-07,1.911226e-07,1.911228e-07,1.911231e-07,1.911233e-07,1.911236e-07,1.911238e-07,1.911241e-07,1.911243e-07,1.911246e-07,1.911248e-07,1.911251e-07,1.911253e-07,1.911256e-07,1.911258e-07,1.911261e-07,1.911263e-07,1.911266e-07,1.911268e-07,1.911271e-07,1.911273e-07,1.911276e-07,1.911278e-07,1.911281e-07,1.911283e-07,1.911286e-07,1.911288e-07,1.911291e-07,1.911293e-07,1.911296e-07,1.911298e-07,1.911301e-07,1.911303e-07,1.911306e-07,1.911308e-07,1.911311e-07,1.911313e-07,1.911316e-07,1.911318e-07,1.911321e-07,1.911323e-07,1.911325e-07,1.911328e-07,1.911330e-07,1.911333e-07,1.911335e-07,1.911338e-07,1.911340e-07,1.911343e-07,1.911345e-07,1.911348e-07,1.911350e-07,1.911353e-07,1.911355e-07,1.911358e-07,1.911360e-07,1.911363e-07,1.911365e-07,1.911368e-07,1.911370e-07,1.911373e-07,1.911375e-07,1.911378e-07,1.911380e-07,1.911383e-07,1.911385e-07,1.911388e-07,1.911390e-07,1.911393e-07,1.911395e-07,1.911398e-07,1.911400e-07,1.911403e-07,1.911405e-07,1.911408e-07,1.911410e-07,1.911413e-07,1.911415e-07,1.911418e-07,1.911420e-07,1.911423e-07,1.911425e-07,1.911428e-07,1.911430e-07,1.911433e-07,1.911435e-07,1.911438e-07,1.911440e-07,1.911443e-07,1.911445e-07,1.911448e-07,1.911450e-07,1.911452e-07,1.911455e-07,1.911457e-07,1.911460e-07,1.911462e-07,1.911465e-07,1.911467e-07,1.911470e-07,1.911472e-07,1.911475e-07,1.911477e-07,1.911480e-07,1.911482e-07,1.911485e-07,1.911487e-07,1.911490e-07,1.911492e-07,1.911495e-07,1.911497e-07,1.911500e-07,1.911502e-07,1.911505e-07,1.911507e-07,1.911510e-07,1.911512e-07,1.911515e-07,1.911517e-07,1.911520e-07,1.911522e-07,1.911525e-07,1.911527e-07,1.911530e-07,1.911532e-07,1.911535e-07,1.911537e-07,1.911540e-07,1.911542e-07,1.911545e-07,1.911547e-07,1.911550e-07,1.911552e-07,1.911554e-07,1.911557e-07,1.911559e-07,1.911562e-07,1.911564e-07,1.911567e-07,1.911569e-07,1.911572e-07,1.911574e-07,1.911577e-07,1.911579e-07,1.911582e-07,1.911584e-07,1.911587e-07,1.911589e-07,1.911592e-07,1.911594e-07,1.911597e-07,1.911599e-07,1.911602e-07,1.911604e-07,1.911607e-07,1.911609e-07,1.911612e-07,1.911614e-07,1.911617e-07,1.911619e-07,1.911622e-07,1.911624e-07,1.911627e-07,1.911629e-07,1.911632e-07,1.911634e-07,1.911637e-07,1.911639e-07,1.911641e-07,1.911644e-07,1.911646e-07,1.911649e-07,1.911651e-07,1.911654e-07,1.911656e-07,1.911659e-07,1.911661e-07,1.911664e-07,1.911666e-07,1.911669e-07,1.911671e-07,1.911674e-07,1.911676e-07,1.911679e-07,1.911681e-07,1.911684e-07,1.911686e-07,1.911689e-07,1.911691e-07,1.911694e-07,1.911696e-07,1.911699e-07,1.911701e-07,1.911704e-07,1.911706e-07,1.911709e-07,1.911711e-07,1.911714e-07,1.911716e-07,1.911718e-07,1.911721e-07,1.911723e-07,1.911726e-07,1.911728e-07,1.911731e-07,1.911733e-07,1.911736e-07,1.911738e-07,1.911741e-07,1.911743e-07,1.911746e-07,1.911748e-07,1.911751e-07,1.911753e-07,1.911756e-07,1.911758e-07,1.911761e-07,1.911763e-07,1.911766e-07,1.911768e-07,1.911771e-07,1.911773e-07,1.911776e-07,1.911778e-07,1.911781e-07,1.911783e-07,1.911786e-07,1.911788e-07,1.911790e-07,1.911793e-07,1.911795e-07,1.911798e-07,1.911800e-07,1.911803e-07,1.911805e-07,1.911808e-07,1.911810e-07,1.911813e-07,1.911815e-07,1.911818e-07,1.911820e-07,1.911823e-07,1.911825e-07,1.911828e-07,1.911830e-07,1.911833e-07,1.911835e-07,1.911838e-07,1.911840e-07,1.911843e-07,1.911845e-07,1.911848e-07,1.911850e-07,1.911852e-07,1.911855e-07,1.911857e-07,1.911860e-07,1.911862e-07,1.911865e-07,1.911867e-07,1.911870e-07,1.911872e-07,1.911875e-07,1.911877e-07,1.911880e-07,1.911882e-07,1.911885e-07,1.911887e-07,1.911890e-07,1.911892e-07,1.911895e-07,1.911897e-07,1.911900e-07,1.911902e-07,1.911905e-07,1.911907e-07,1.911910e-07,1.911912e-07,1.911914e-07,1.911917e-07,1.911919e-07,1.911922e-07,1.911924e-07,1.911927e-07,1.911929e-07,1.911932e-07,1.911934e-07,1.911937e-07,1.911939e-07,1.911942e-07,1.911944e-07,1.911947e-07,1.911949e-07,1.911952e-07,1.911954e-07,1.911957e-07,1.911959e-07,1.911962e-07,1.911964e-07,1.911967e-07,1.911969e-07,1.911971e-07,1.911974e-07,1.911976e-07,1.911979e-07,1.911981e-07,1.911984e-07,1.911986e-07,1.911989e-07,1.911991e-07,1.911994e-07,1.911996e-07,1.911999e-07,1.912001e-07,1.912004e-07,1.912006e-07,1.912009e-07,1.912011e-07,1.912014e-07,1.912016e-07,1.912019e-07,1.912021e-07,1.912024e-07,1.912026e-07,1.912028e-07,1.912031e-07,1.912033e-07,1.912036e-07,1.912038e-07,1.912041e-07,1.912043e-07,1.912046e-07,1.912048e-07,1.912051e-07,1.912053e-07,1.912056e-07,1.912058e-07,1.912061e-07,1.912063e-07,1.912066e-07,1.912068e-07,1.912071e-07,1.912073e-07,1.912076e-07,1.912078e-07,1.912080e-07,1.912083e-07,1.912085e-07,1.912088e-07,1.912090e-07,1.912093e-07,1.912095e-07,1.912098e-07,1.912100e-07,1.912103e-07,1.912105e-07,1.912108e-07,1.912110e-07,1.912113e-07,1.912115e-07,1.912118e-07,1.912120e-07,1.912123e-07,1.912125e-07,1.912127e-07,1.912130e-07,1.912132e-07,1.912135e-07,1.912137e-07,1.912140e-07,1.912142e-07,1.912145e-07,1.912147e-07,1.912150e-07,1.912152e-07,1.912155e-07,1.912157e-07,1.912160e-07,1.912162e-07,1.912165e-07,1.912167e-07,1.912170e-07,1.912172e-07,1.912174e-07,1.912177e-07,1.912179e-07,1.912182e-07,1.912184e-07,1.912187e-07,1.912189e-07,1.912192e-07,1.912194e-07,1.912197e-07,1.912199e-07,1.912202e-07,1.912204e-07,1.912207e-07,1.912209e-07,1.912212e-07,1.912214e-07,1.912217e-07,1.912219e-07,1.912221e-07,1.912224e-07,1.912226e-07,1.912229e-07,1.912231e-07,1.912234e-07,1.912236e-07,1.912239e-07,1.912241e-07,1.912244e-07,1.912246e-07,1.912249e-07,1.912251e-07,1.912254e-07,1.912256e-07,1.912259e-07,1.912261e-07,1.912263e-07,1.912266e-07,1.912268e-07,1.912271e-07,1.912273e-07,1.912276e-07,1.912278e-07,1.912281e-07,1.912283e-07,1.912286e-07,1.912288e-07,1.912291e-07,1.912293e-07,1.912296e-07,1.912298e-07,1.912301e-07,1.912303e-07,1.912306e-07,1.912308e-07,1.912310e-07,1.912313e-07,1.912315e-07,1.912318e-07,1.912320e-07,1.912323e-07,1.912325e-07,1.912328e-07,1.912330e-07,1.912333e-07,1.912335e-07,1.912338e-07,1.912340e-07,1.912343e-07,1.912345e-07,1.912348e-07,1.912350e-07,1.912352e-07,1.912355e-07,1.912357e-07,1.912360e-07,1.912362e-07,1.912365e-07,1.912367e-07,1.912370e-07,1.912372e-07,1.912375e-07,1.912377e-07,1.912380e-07,1.912382e-07,1.912385e-07,1.912387e-07,1.912389e-07,1.912392e-07,1.912394e-07,1.912397e-07,1.912399e-07,1.912402e-07,1.912404e-07,1.912407e-07,1.912409e-07,1.912412e-07,1.912414e-07,1.912417e-07,1.912419e-07,1.912422e-07,1.912424e-07,1.912427e-07,1.912429e-07,1.912431e-07,1.912434e-07,1.912436e-07,1.912439e-07,1.912441e-07,1.912444e-07,1.912446e-07,1.912449e-07,1.912451e-07,1.912454e-07,1.912456e-07,1.912459e-07,1.912461e-07,1.912464e-07,1.912466e-07,1.912468e-07,1.912471e-07,1.912473e-07,1.912476e-07,1.912478e-07,1.912481e-07,1.912483e-07,1.912486e-07,1.912488e-07,1.912491e-07,1.912493e-07,1.912496e-07,1.912498e-07,1.912501e-07,1.912503e-07,1.912505e-07,1.912508e-07,1.912510e-07,1.912513e-07,1.912515e-07,1.912518e-07,1.912520e-07,1.912523e-07,1.912525e-07,1.912528e-07,1.912530e-07,1.912533e-07,1.912535e-07,1.912538e-07,1.912540e-07,1.912542e-07,1.912545e-07,1.912547e-07,1.912550e-07,1.912552e-07,1.912555e-07,1.912557e-07,1.912560e-07,1.912562e-07,1.912565e-07,1.912567e-07,1.912570e-07,1.912572e-07,1.912575e-07,1.912577e-07,1.912579e-07,1.912582e-07,1.912584e-07,1.912587e-07,1.912589e-07,1.912592e-07,1.912594e-07,1.912597e-07,1.912599e-07,1.912602e-07,1.912604e-07,1.912607e-07,1.912609e-07,1.912611e-07,1.912614e-07,1.912616e-07,1.912619e-07,1.912621e-07,1.912624e-07,1.912626e-07,1.912629e-07,1.912631e-07,1.912634e-07,1.912636e-07,1.912639e-07,1.912641e-07,1.912644e-07,1.912646e-07,1.912648e-07,1.912651e-07,1.912653e-07,1.912656e-07,1.912658e-07,1.912661e-07,1.912663e-07,1.912666e-07,1.912668e-07,1.912671e-07,1.912673e-07,1.912676e-07,1.912678e-07,1.912680e-07,1.912683e-07,1.912685e-07,1.912688e-07,1.912690e-07,1.912693e-07,1.912695e-07,1.912698e-07,1.912700e-07,1.912703e-07,1.912705e-07,1.912708e-07,1.912710e-07,1.912712e-07,1.912715e-07,1.912717e-07,1.912720e-07,1.912722e-07,1.912725e-07,1.912727e-07,1.912730e-07,1.912732e-07,1.912735e-07,1.912737e-07,1.912740e-07,1.912742e-07,1.912744e-07,1.912747e-07,1.912749e-07,1.912752e-07,1.912754e-07,1.912757e-07,1.912759e-07,1.912762e-07,1.912764e-07,1.912767e-07,1.912769e-07,1.912772e-07,1.912774e-07,1.912776e-07,1.912779e-07,1.912781e-07,1.912784e-07,1.912786e-07,1.912789e-07,1.912791e-07,1.912794e-07,1.912796e-07,1.912799e-07,1.912801e-07,1.912804e-07,1.912806e-07,1.912808e-07,1.912811e-07,1.912813e-07,1.912816e-07,1.912818e-07,1.912821e-07,1.912823e-07,1.912826e-07,1.912828e-07,1.912831e-07,1.912833e-07,1.912836e-07,1.912838e-07,1.912840e-07,1.912843e-07,1.912845e-07,1.912848e-07,1.912850e-07,1.912853e-07,1.912855e-07,1.912858e-07,1.912860e-07,1.912863e-07,1.912865e-07,1.912867e-07,1.912870e-07,1.912872e-07,1.912875e-07,1.912877e-07,1.912880e-07,1.912882e-07,1.912885e-07,1.912887e-07,1.912890e-07,1.912892e-07,1.912895e-07,1.912897e-07,1.912899e-07,1.912902e-07,1.912904e-07,1.912907e-07,1.912909e-07,1.912912e-07,1.912914e-07,1.912917e-07,1.912919e-07,1.912922e-07,1.912924e-07,1.912926e-07,1.912929e-07,1.912931e-07,1.912934e-07,1.912936e-07,1.912939e-07,1.912941e-07,1.912944e-07,1.912946e-07,1.912949e-07,1.912951e-07,1.912954e-07,1.912956e-07,1.912958e-07,1.912961e-07,1.912963e-07,1.912966e-07,1.912968e-07,1.912971e-07,1.912973e-07,1.912976e-07,1.912978e-07,1.912981e-07,1.912983e-07,1.912985e-07,1.912988e-07,1.912990e-07,1.912993e-07,1.912995e-07,1.912998e-07,1.913000e-07,1.913003e-07,1.913005e-07,1.913008e-07,1.913010e-07,1.913012e-07,1.913015e-07,1.913017e-07,1.913020e-07,1.913022e-07,1.913025e-07,1.913027e-07,1.913030e-07,1.913032e-07,1.913035e-07,1.913037e-07,1.913039e-07,1.913042e-07,1.913044e-07,1.913047e-07,1.913049e-07,1.913052e-07,1.913054e-07,1.913057e-07,1.913059e-07,1.913062e-07,1.913064e-07,1.913066e-07,1.913069e-07,1.913071e-07,1.913074e-07,1.913076e-07,1.913079e-07,1.913081e-07,1.913084e-07,1.913086e-07,1.913089e-07,1.913091e-07,1.913093e-07,1.913096e-07,1.913098e-07,1.913101e-07,1.913103e-07,1.913106e-07,1.913108e-07,1.913111e-07,1.913113e-07,1.913116e-07,1.913118e-07,1.913120e-07,1.913123e-07,1.913125e-07,1.913128e-07,1.913130e-07,1.913133e-07,1.913135e-07,1.913138e-07,1.913140e-07,1.913143e-07,1.913145e-07,1.913147e-07,1.913150e-07,1.913152e-07,1.913155e-07,1.913157e-07,1.913160e-07,1.913162e-07,1.913165e-07,1.913167e-07,1.913170e-07,1.913172e-07,1.913174e-07,1.913177e-07,1.913179e-07,1.913182e-07,1.913184e-07,1.913187e-07,1.913189e-07,1.913192e-07,1.913194e-07,1.913196e-07,1.913199e-07,1.913201e-07,1.913204e-07,1.913206e-07,1.913209e-07,1.913211e-07,1.913214e-07,1.913216e-07,1.913219e-07,1.913221e-07,1.913223e-07,1.913226e-07,1.913228e-07,1.913231e-07,1.913233e-07,1.913236e-07,1.913238e-07,1.913241e-07,1.913243e-07,1.913246e-07,1.913248e-07,1.913250e-07,1.913253e-07,1.913255e-07,1.913258e-07,1.913260e-07,1.913263e-07,1.913265e-07,1.913268e-07,1.913270e-07,1.913272e-07,1.913275e-07,1.913277e-07,1.913280e-07,1.913282e-07,1.913285e-07,1.913287e-07,1.913290e-07,1.913292e-07,1.913295e-07,1.913297e-07,1.913299e-07,1.913302e-07,1.913304e-07,1.913307e-07,1.913309e-07,1.913312e-07,1.913314e-07,1.913317e-07,1.913319e-07,1.913321e-07,1.913324e-07,1.913326e-07,1.913329e-07,1.913331e-07,1.913334e-07,1.913336e-07,1.913339e-07,1.913341e-07,1.913344e-07,1.913346e-07,1.913348e-07,1.913351e-07,1.913353e-07,1.913356e-07,1.913358e-07,1.913361e-07,1.913363e-07,1.913366e-07,1.913368e-07,1.913370e-07,1.913373e-07,1.913375e-07,1.913378e-07,1.913380e-07,1.913383e-07,1.913385e-07,1.913388e-07,1.913390e-07,1.913392e-07,1.913395e-07,1.913397e-07,1.913400e-07,1.913402e-07,1.913405e-07,1.913407e-07,1.913410e-07,1.913412e-07,1.913415e-07,1.913417e-07,1.913419e-07,1.913422e-07,1.913424e-07,1.913427e-07,1.913429e-07,1.913432e-07,1.913434e-07,1.913437e-07,1.913439e-07,1.913441e-07,1.913444e-07,1.913446e-07,1.913449e-07,1.913451e-07,1.913454e-07,1.913456e-07,1.913459e-07,1.913461e-07,1.913463e-07,1.913466e-07,1.913468e-07,1.913471e-07,1.913473e-07,1.913476e-07,1.913478e-07,1.913481e-07,1.913483e-07,1.913485e-07,1.913488e-07,1.913490e-07,1.913493e-07,1.913495e-07,1.913498e-07,1.913500e-07,1.913503e-07,1.913505e-07,1.913507e-07,1.913510e-07,1.913512e-07,1.913515e-07,1.913517e-07,1.913520e-07,1.913522e-07,1.913525e-07,1.913527e-07,1.913529e-07,1.913532e-07,1.913534e-07,1.913537e-07,1.913539e-07,1.913542e-07,1.913544e-07,1.913547e-07,1.913549e-07,1.913551e-07,1.913554e-07,1.913556e-07,1.913559e-07,1.913561e-07,1.913564e-07,1.913566e-07,1.913569e-07,1.913571e-07,1.913573e-07,1.913576e-07,1.913578e-07,1.913581e-07,1.913583e-07,1.913586e-07,1.913588e-07,1.913591e-07,1.913593e-07,1.913595e-07,1.913598e-07,1.913600e-07,1.913603e-07,1.913605e-07,1.913608e-07,1.913610e-07,1.913613e-07,1.913615e-07,1.913617e-07,1.913620e-07,1.913622e-07,1.913625e-07,1.913627e-07,1.913630e-07,1.913632e-07,1.913635e-07,1.913637e-07,1.913639e-07,1.913642e-07,1.913644e-07,1.913647e-07,1.913649e-07,1.913652e-07,1.913654e-07,1.913657e-07,1.913659e-07,1.913661e-07,1.913664e-07,1.913666e-07,1.913669e-07,1.913671e-07,1.913674e-07,1.913676e-07,1.913679e-07,1.913681e-07,1.913683e-07,1.913686e-07,1.913688e-07,1.913691e-07,1.913693e-07,1.913696e-07,1.913698e-07,1.913701e-07,1.913703e-07,1.913705e-07,1.913708e-07,1.913710e-07,1.913713e-07,1.913715e-07,1.913718e-07,1.913720e-07,1.913722e-07,1.913725e-07,1.913727e-07,1.913730e-07,1.913732e-07,1.913735e-07,1.913737e-07,1.913740e-07,1.913742e-07,1.913744e-07,1.913747e-07,1.913749e-07,1.913752e-07,1.913754e-07,1.913757e-07,1.913759e-07,1.913762e-07,1.913764e-07,1.913766e-07,1.913769e-07,1.913771e-07,1.913774e-07,1.913776e-07,1.913779e-07,1.913781e-07,1.913783e-07,1.913786e-07,1.913788e-07,1.913791e-07,1.913793e-07,1.913796e-07,1.913798e-07,1.913801e-07,1.913803e-07,1.913805e-07,1.913808e-07,1.913810e-07,1.913813e-07,1.913815e-07,1.913818e-07,1.913820e-07,1.913823e-07,1.913825e-07,1.913827e-07,1.913830e-07,1.913832e-07,1.913835e-07,1.913837e-07,1.913840e-07,1.913842e-07,1.913844e-07,1.913847e-07,1.913849e-07,1.913852e-07,1.913854e-07,1.913857e-07,1.913859e-07,1.913862e-07,1.913864e-07,1.913866e-07,1.913869e-07,1.913871e-07,1.913874e-07,1.913876e-07,1.913879e-07,1.913881e-07,1.913883e-07,1.913886e-07,1.913888e-07,1.913891e-07,1.913893e-07,1.913896e-07,1.913898e-07,1.913901e-07,1.913903e-07,1.913905e-07,1.913908e-07,1.913910e-07,1.913913e-07,1.913915e-07,1.913918e-07,1.913920e-07,1.913922e-07,1.913925e-07,1.913927e-07,1.913930e-07,1.913932e-07,1.913935e-07,1.913937e-07,1.913940e-07,1.913942e-07,1.913944e-07,1.913947e-07,1.913949e-07,1.913952e-07,1.913954e-07,1.913957e-07,1.913959e-07,1.913961e-07,1.913964e-07,1.913966e-07,1.913969e-07,1.913971e-07,1.913974e-07,1.913976e-07,1.913979e-07,1.913981e-07,1.913983e-07,1.913986e-07,1.913988e-07,1.913991e-07,1.913993e-07,1.913996e-07,1.913998e-07,1.914000e-07,1.914003e-07,1.914005e-07,1.914008e-07,1.914010e-07,1.914013e-07,1.914015e-07,1.914017e-07,1.914020e-07,1.914022e-07,1.914025e-07,1.914027e-07,1.914030e-07,1.914032e-07,1.914035e-07,1.914037e-07,1.914039e-07,1.914042e-07,1.914044e-07,1.914047e-07,1.914049e-07,1.914052e-07,1.914054e-07,1.914056e-07,1.914059e-07,1.914061e-07,1.914064e-07,1.914066e-07,1.914069e-07,1.914071e-07,1.914073e-07,1.914076e-07,1.914078e-07,1.914081e-07,1.914083e-07,1.914086e-07,1.914088e-07,1.914090e-07,1.914093e-07,1.914095e-07,1.914098e-07,1.914100e-07,1.914103e-07,1.914105e-07,1.914108e-07,1.914110e-07,1.914112e-07,1.914115e-07,1.914117e-07,1.914120e-07,1.914122e-07,1.914125e-07,1.914127e-07,1.914129e-07,1.914132e-07,1.914134e-07,1.914137e-07,1.914139e-07,1.914142e-07,1.914144e-07,1.914146e-07,1.914149e-07,1.914151e-07,1.914154e-07,1.914156e-07,1.914159e-07,1.914161e-07,1.914163e-07,1.914166e-07,1.914168e-07,1.914171e-07,1.914173e-07,1.914176e-07,1.914178e-07,1.914180e-07,1.914183e-07,1.914185e-07,1.914188e-07,1.914190e-07,1.914193e-07,1.914195e-07,1.914198e-07,1.914200e-07,1.914202e-07,1.914205e-07,1.914207e-07,1.914210e-07,1.914212e-07,1.914215e-07,1.914217e-07,1.914219e-07,1.914222e-07,1.914224e-07,1.914227e-07,1.914229e-07,1.914232e-07,1.914234e-07,1.914236e-07,1.914239e-07,1.914241e-07,1.914244e-07,1.914246e-07,1.914249e-07,1.914251e-07,1.914253e-07,1.914256e-07,1.914258e-07,1.914261e-07,1.914263e-07,1.914266e-07,1.914268e-07,1.914270e-07,1.914273e-07,1.914275e-07,1.914278e-07,1.914280e-07,1.914283e-07,1.914285e-07,1.914287e-07,1.914290e-07,1.914292e-07,1.914295e-07,1.914297e-07,1.914300e-07,1.914302e-07,1.914304e-07,1.914307e-07,1.914309e-07,1.914312e-07,1.914314e-07,1.914317e-07,1.914319e-07,1.914321e-07,1.914324e-07,1.914326e-07,1.914329e-07,1.914331e-07,1.914334e-07,1.914336e-07,1.914338e-07,1.914341e-07,1.914343e-07,1.914346e-07,1.914348e-07,1.914351e-07,1.914353e-07,1.914355e-07,1.914358e-07,1.914360e-07,1.914363e-07,1.914365e-07,1.914368e-07,1.914370e-07,1.914372e-07,1.914375e-07,1.914377e-07,1.914380e-07,1.914382e-07,1.914385e-07,1.914387e-07,1.914389e-07,1.914392e-07,1.914394e-07,1.914397e-07,1.914399e-07,1.914402e-07,1.914404e-07,1.914406e-07,1.914409e-07,1.914411e-07,1.914414e-07,1.914416e-07,1.914419e-07,1.914421e-07,1.914423e-07,1.914426e-07,1.914428e-07,1.914431e-07,1.914433e-07,1.914436e-07,1.914438e-07,1.914440e-07,1.914443e-07,1.914445e-07,1.914448e-07,1.914450e-07,1.914452e-07,1.914455e-07,1.914457e-07,1.914460e-07,1.914462e-07,1.914465e-07,1.914467e-07,1.914469e-07,1.914472e-07,1.914474e-07,1.914477e-07,1.914479e-07,1.914482e-07,1.914484e-07,1.914486e-07,1.914489e-07,1.914491e-07,1.914494e-07,1.914496e-07,1.914499e-07,1.914501e-07,1.914503e-07,1.914506e-07,1.914508e-07,1.914511e-07,1.914513e-07,1.914516e-07,1.914518e-07,1.914520e-07,1.914523e-07,1.914525e-07,1.914528e-07,1.914530e-07,1.914533e-07,1.914535e-07,1.914537e-07,1.914540e-07,1.914542e-07,1.914545e-07,1.914547e-07,1.914549e-07,1.914552e-07,1.914554e-07,1.914557e-07,1.914559e-07,1.914562e-07,1.914564e-07,1.914566e-07,1.914569e-07,1.914571e-07,1.914574e-07,1.914576e-07,1.914579e-07,1.914581e-07,1.914583e-07,1.914586e-07,1.914588e-07,1.914591e-07,1.914593e-07,1.914596e-07,1.914598e-07,1.914600e-07,1.914603e-07,1.914605e-07,1.914608e-07,1.914610e-07,1.914612e-07,1.914615e-07,1.914617e-07,1.914620e-07,1.914622e-07,1.914625e-07,1.914627e-07,1.914629e-07,1.914632e-07,1.914634e-07,1.914637e-07,1.914639e-07,1.914642e-07,1.914644e-07,1.914646e-07,1.914649e-07,1.914651e-07,1.914654e-07,1.914656e-07,1.914658e-07,1.914661e-07,1.914663e-07,1.914666e-07,1.914668e-07,1.914671e-07,1.914673e-07,1.914675e-07,1.914678e-07,1.914680e-07,1.914683e-07,1.914685e-07,1.914688e-07,1.914690e-07,1.914692e-07,1.914695e-07,1.914697e-07,1.914700e-07,1.914702e-07,1.914704e-07,1.914707e-07,1.914709e-07,1.914712e-07,1.914714e-07,1.914717e-07,1.914719e-07,1.914721e-07,1.914724e-07,1.914726e-07,1.914729e-07,1.914731e-07,1.914734e-07,1.914736e-07,1.914738e-07,1.914741e-07,1.914743e-07,1.914746e-07,1.914748e-07,1.914750e-07,1.914753e-07,1.914755e-07,1.914758e-07,1.914760e-07,1.914763e-07,1.914765e-07,1.914767e-07,1.914770e-07,1.914772e-07,1.914775e-07,1.914777e-07,1.914780e-07,1.914782e-07,1.914784e-07,1.914787e-07,1.914789e-07,1.914792e-07,1.914794e-07,1.914796e-07,1.914799e-07,1.914801e-07,1.914804e-07,1.914806e-07,1.914809e-07,1.914811e-07,1.914813e-07,1.914816e-07,1.914818e-07,1.914821e-07,1.914823e-07,1.914825e-07,1.914828e-07,1.914830e-07,1.914833e-07,1.914835e-07,1.914838e-07,1.914840e-07,1.914842e-07,1.914845e-07,1.914847e-07,1.914850e-07,1.914852e-07,1.914854e-07,1.914857e-07,1.914859e-07,1.914862e-07,1.914864e-07,1.914867e-07,1.914869e-07,1.914871e-07,1.914874e-07,1.914876e-07,1.914879e-07,1.914881e-07,1.914883e-07,1.914886e-07,1.914888e-07,1.914891e-07,1.914893e-07,1.914896e-07,1.914898e-07,1.914900e-07,1.914903e-07,1.914905e-07,1.914908e-07,1.914910e-07,1.914912e-07,1.914915e-07,1.914917e-07,1.914920e-07,1.914922e-07,1.914925e-07,1.914927e-07,1.914929e-07,1.914932e-07,1.914934e-07,1.914937e-07,1.914939e-07,1.914941e-07,1.914944e-07,1.914946e-07,1.914949e-07,1.914951e-07,1.914954e-07,1.914956e-07,1.914958e-07,1.914961e-07,1.914963e-07,1.914966e-07,1.914968e-07,1.914970e-07,1.914973e-07,1.914975e-07,1.914978e-07,1.914980e-07,1.914983e-07,1.914985e-07,1.914987e-07,1.914990e-07,1.914992e-07,1.914995e-07,1.914997e-07,1.914999e-07,1.915002e-07,1.915004e-07,1.915007e-07,1.915009e-07,1.915012e-07,1.915014e-07,1.915016e-07,1.915019e-07,1.915021e-07,1.915024e-07,1.915026e-07,1.915028e-07,1.915031e-07,1.915033e-07,1.915036e-07,1.915038e-07,1.915040e-07,1.915043e-07,1.915045e-07,1.915048e-07,1.915050e-07,1.915053e-07,1.915055e-07,1.915057e-07,1.915060e-07,1.915062e-07,1.915065e-07,1.915067e-07,1.915069e-07,1.915072e-07,1.915074e-07,1.915077e-07,1.915079e-07,1.915081e-07,1.915084e-07,1.915086e-07,1.915089e-07,1.915091e-07,1.915094e-07,1.915096e-07,1.915098e-07,1.915101e-07,1.915103e-07,1.915106e-07,1.915108e-07,1.915110e-07,1.915113e-07,1.915115e-07,1.915118e-07,1.915120e-07,1.915123e-07,1.915125e-07,1.915127e-07,1.915130e-07,1.915132e-07,1.915135e-07,1.915137e-07,1.915139e-07,1.915142e-07,1.915144e-07,1.915147e-07,1.915149e-07,1.915151e-07,1.915154e-07,1.915156e-07,1.915159e-07,1.915161e-07,1.915163e-07,1.915166e-07,1.915168e-07,1.915171e-07,1.915173e-07,1.915176e-07,1.915178e-07,1.915180e-07,1.915183e-07,1.915185e-07,1.915188e-07,1.915190e-07,1.915192e-07,1.915195e-07,1.915197e-07,1.915200e-07,1.915202e-07,1.915204e-07,1.915207e-07,1.915209e-07,1.915212e-07,1.915214e-07,1.915217e-07,1.915219e-07,1.915221e-07,1.915224e-07,1.915226e-07,1.915229e-07,1.915231e-07,1.915233e-07,1.915236e-07,1.915238e-07,1.915241e-07,1.915243e-07,1.915245e-07,1.915248e-07,1.915250e-07,1.915253e-07,1.915255e-07,1.915257e-07,1.915260e-07,1.915262e-07,1.915265e-07,1.915267e-07,1.915270e-07,1.915272e-07,1.915274e-07,1.915277e-07,1.915279e-07,1.915282e-07,1.915284e-07,1.915286e-07,1.915289e-07,1.915291e-07,1.915294e-07,1.915296e-07,1.915298e-07,1.915301e-07,1.915303e-07,1.915306e-07,1.915308e-07,1.915310e-07,1.915313e-07,1.915315e-07,1.915318e-07,1.915320e-07,1.915323e-07,1.915325e-07,1.915327e-07,1.915330e-07,1.915332e-07,1.915335e-07,1.915337e-07,1.915339e-07,1.915342e-07,1.915344e-07,1.915347e-07,1.915349e-07,1.915351e-07,1.915354e-07,1.915356e-07,1.915359e-07,1.915361e-07,1.915363e-07,1.915366e-07,1.915368e-07,1.915371e-07,1.915373e-07,1.915375e-07,1.915378e-07,1.915380e-07,1.915383e-07,1.915385e-07,1.915388e-07,1.915390e-07,1.915392e-07,1.915395e-07,1.915397e-07,1.915400e-07,1.915402e-07,1.915404e-07,1.915407e-07,1.915409e-07,1.915412e-07,1.915414e-07,1.915416e-07,1.915419e-07,1.915421e-07,1.915424e-07,1.915426e-07,1.915428e-07,1.915431e-07,1.915433e-07,1.915436e-07,1.915438e-07,1.915440e-07,1.915443e-07,1.915445e-07,1.915448e-07,1.915450e-07,1.915452e-07,1.915455e-07,1.915457e-07,1.915460e-07,1.915462e-07,1.915464e-07,1.915467e-07,1.915469e-07,1.915472e-07,1.915474e-07,1.915477e-07,1.915479e-07,1.915481e-07,1.915484e-07,1.915486e-07,1.915489e-07,1.915491e-07,1.915493e-07,1.915496e-07,1.915498e-07,1.915501e-07,1.915503e-07,1.915505e-07,1.915508e-07,1.915510e-07,1.915513e-07,1.915515e-07,1.915517e-07,1.915520e-07,1.915522e-07,1.915525e-07,1.915527e-07,1.915529e-07,1.915532e-07,1.915534e-07,1.915537e-07,1.915539e-07,1.915541e-07,1.915544e-07,1.915546e-07,1.915549e-07,1.915551e-07,1.915553e-07,1.915556e-07,1.915558e-07,1.915561e-07,1.915563e-07,1.915565e-07,1.915568e-07,1.915570e-07,1.915573e-07,1.915575e-07,1.915577e-07,1.915580e-07,1.915582e-07,1.915585e-07,1.915587e-07,1.915589e-07,1.915592e-07,1.915594e-07,1.915597e-07,1.915599e-07,1.915601e-07,1.915604e-07,1.915606e-07,1.915609e-07,1.915611e-07,1.915613e-07,1.915616e-07,1.915618e-07,1.915621e-07,1.915623e-07,1.915626e-07,1.915628e-07,1.915630e-07,1.915633e-07,1.915635e-07,1.915638e-07,1.915640e-07,1.915642e-07,1.915645e-07,1.915647e-07,1.915650e-07,1.915652e-07,1.915654e-07,1.915657e-07,1.915659e-07,1.915662e-07,1.915664e-07,1.915666e-07,1.915669e-07,1.915671e-07,1.915674e-07,1.915676e-07,1.915678e-07,1.915681e-07,1.915683e-07,1.915686e-07,1.915688e-07,1.915690e-07,1.915693e-07,1.915695e-07,1.915698e-07,1.915700e-07,1.915702e-07,1.915705e-07,1.915707e-07,1.915710e-07,1.915712e-07,1.915714e-07,1.915717e-07,1.915719e-07,1.915722e-07,1.915724e-07,1.915726e-07,1.915729e-07,1.915731e-07,1.915734e-07,1.915736e-07,1.915738e-07,1.915741e-07,1.915743e-07,1.915746e-07,1.915748e-07,1.915750e-07,1.915753e-07,1.915755e-07,1.915758e-07,1.915760e-07,1.915762e-07,1.915765e-07,1.915767e-07,1.915770e-07,1.915772e-07,1.915774e-07,1.915777e-07,1.915779e-07,1.915782e-07,1.915784e-07,1.915786e-07,1.915789e-07,1.915791e-07,1.915793e-07,1.915796e-07,1.915798e-07,1.915801e-07,1.915803e-07,1.915805e-07,1.915808e-07,1.915810e-07,1.915813e-07,1.915815e-07,1.915817e-07,1.915820e-07,1.915822e-07,1.915825e-07,1.915827e-07,1.915829e-07,1.915832e-07,1.915834e-07,1.915837e-07,1.915839e-07,1.915841e-07,1.915844e-07,1.915846e-07,1.915849e-07,1.915851e-07,1.915853e-07,1.915856e-07,1.915858e-07,1.915861e-07,1.915863e-07,1.915865e-07,1.915868e-07,1.915870e-07,1.915873e-07,1.915875e-07,1.915877e-07,1.915880e-07,1.915882e-07,1.915885e-07,1.915887e-07,1.915889e-07,1.915892e-07,1.915894e-07,1.915897e-07,1.915899e-07,1.915901e-07,1.915904e-07,1.915906e-07,1.915909e-07,1.915911e-07,1.915913e-07,1.915916e-07,1.915918e-07,1.915921e-07,1.915923e-07,1.915925e-07,1.915928e-07,1.915930e-07,1.915933e-07,1.915935e-07,1.915937e-07,1.915940e-07,1.915942e-07,1.915944e-07,1.915947e-07,1.915949e-07,1.915952e-07,1.915954e-07,1.915956e-07,1.915959e-07,1.915961e-07,1.915964e-07,1.915966e-07,1.915968e-07,1.915971e-07,1.915973e-07,1.915976e-07,1.915978e-07,1.915980e-07,1.915983e-07,1.915985e-07,1.915988e-07,1.915990e-07,1.915992e-07,1.915995e-07,1.915997e-07,1.916000e-07,1.916002e-07,1.916004e-07,1.916007e-07,1.916009e-07,1.916012e-07,1.916014e-07,1.916016e-07,1.916019e-07,1.916021e-07,1.916023e-07,1.916026e-07,1.916028e-07,1.916031e-07,1.916033e-07,1.916035e-07,1.916038e-07,1.916040e-07,1.916043e-07,1.916045e-07,1.916047e-07,1.916050e-07,1.916052e-07,1.916055e-07,1.916057e-07,1.916059e-07,1.916062e-07,1.916064e-07,1.916067e-07,1.916069e-07,1.916071e-07,1.916074e-07,1.916076e-07,1.916079e-07,1.916081e-07,1.916083e-07,1.916086e-07,1.916088e-07,1.916090e-07,1.916093e-07,1.916095e-07,1.916098e-07,1.916100e-07,1.916102e-07,1.916105e-07,1.916107e-07,1.916110e-07,1.916112e-07,1.916114e-07,1.916117e-07,1.916119e-07,1.916122e-07,1.916124e-07,1.916126e-07,1.916129e-07,1.916131e-07,1.916134e-07,1.916136e-07,1.916138e-07,1.916141e-07,1.916143e-07,1.916145e-07,1.916148e-07,1.916150e-07,1.916153e-07,1.916155e-07,1.916157e-07,1.916160e-07,1.916162e-07,1.916165e-07,1.916167e-07,1.916169e-07,1.916172e-07,1.916174e-07,1.916177e-07,1.916179e-07,1.916181e-07,1.916184e-07,1.916186e-07,1.916189e-07,1.916191e-07,1.916193e-07,1.916196e-07,1.916198e-07,1.916200e-07,1.916203e-07,1.916205e-07,1.916208e-07,1.916210e-07,1.916212e-07,1.916215e-07,1.916217e-07,1.916220e-07,1.916222e-07,1.916224e-07,1.916227e-07,1.916229e-07,1.916232e-07,1.916234e-07,1.916236e-07,1.916239e-07,1.916241e-07,1.916243e-07,1.916246e-07,1.916248e-07,1.916251e-07,1.916253e-07,1.916255e-07,1.916258e-07,1.916260e-07,1.916263e-07,1.916265e-07,1.916267e-07,1.916270e-07,1.916272e-07,1.916275e-07,1.916277e-07,1.916279e-07,1.916282e-07,1.916284e-07,1.916286e-07,1.916289e-07,1.916291e-07,1.916294e-07,1.916296e-07,1.916298e-07,1.916301e-07,1.916303e-07,1.916306e-07,1.916308e-07,1.916310e-07,1.916313e-07,1.916315e-07,1.916318e-07,1.916320e-07,1.916322e-07,1.916325e-07,1.916327e-07,1.916329e-07,1.916332e-07,1.916334e-07,1.916337e-07,1.916339e-07,1.916341e-07,1.916344e-07,1.916346e-07,1.916349e-07,1.916351e-07,1.916353e-07,1.916356e-07,1.916358e-07,1.916360e-07,1.916363e-07,1.916365e-07,1.916368e-07,1.916370e-07,1.916372e-07,1.916375e-07,1.916377e-07,1.916380e-07,1.916382e-07,1.916384e-07,1.916387e-07,1.916389e-07,1.916391e-07,1.916394e-07,1.916396e-07,1.916399e-07,1.916401e-07,1.916403e-07,1.916406e-07,1.916408e-07,1.916411e-07,1.916413e-07,1.916415e-07,1.916418e-07,1.916420e-07,1.916423e-07,1.916425e-07,1.916427e-07,1.916430e-07,1.916432e-07,1.916434e-07,1.916437e-07,1.916439e-07,1.916442e-07,1.916444e-07,1.916446e-07,1.916449e-07,1.916451e-07,1.916454e-07,1.916456e-07,1.916458e-07,1.916461e-07,1.916463e-07,1.916465e-07,1.916468e-07,1.916470e-07,1.916473e-07,1.916475e-07,1.916477e-07,1.916480e-07,1.916482e-07,1.916485e-07,1.916487e-07,1.916489e-07,1.916492e-07,1.916494e-07,1.916496e-07,1.916499e-07,1.916501e-07,1.916504e-07,1.916506e-07,1.916508e-07,1.916511e-07,1.916513e-07,1.916515e-07,1.916518e-07,1.916520e-07,1.916523e-07,1.916525e-07,1.916527e-07,1.916530e-07,1.916532e-07,1.916535e-07,1.916537e-07,1.916539e-07,1.916542e-07,1.916544e-07,1.916546e-07,1.916549e-07,1.916551e-07,1.916554e-07,1.916556e-07,1.916558e-07,1.916561e-07,1.916563e-07,1.916566e-07,1.916568e-07,1.916570e-07,1.916573e-07,1.916575e-07,1.916577e-07,1.916580e-07,1.916582e-07,1.916585e-07,1.916587e-07,1.916589e-07,1.916592e-07,1.916594e-07,1.916596e-07,1.916599e-07,1.916601e-07,1.916604e-07,1.916606e-07,1.916608e-07,1.916611e-07,1.916613e-07,1.916616e-07,1.916618e-07,1.916620e-07,1.916623e-07,1.916625e-07,1.916627e-07,1.916630e-07,1.916632e-07,1.916635e-07,1.916637e-07,1.916639e-07,1.916642e-07,1.916644e-07,1.916647e-07,1.916649e-07,1.916651e-07,1.916654e-07,1.916656e-07,1.916658e-07,1.916661e-07,1.916663e-07,1.916666e-07,1.916668e-07,1.916670e-07,1.916673e-07,1.916675e-07,1.916677e-07,1.916680e-07,1.916682e-07,1.916685e-07,1.916687e-07,1.916689e-07,1.916692e-07,1.916694e-07,1.916696e-07,1.916699e-07,1.916701e-07,1.916704e-07,1.916706e-07,1.916708e-07,1.916711e-07,1.916713e-07,1.916716e-07,1.916718e-07,1.916720e-07,1.916723e-07,1.916725e-07,1.916727e-07,1.916730e-07,1.916732e-07,1.916735e-07,1.916737e-07,1.916739e-07,1.916742e-07,1.916744e-07,1.916746e-07,1.916749e-07,1.916751e-07,1.916754e-07,1.916756e-07,1.916758e-07,1.916761e-07,1.916763e-07,1.916765e-07,1.916768e-07,1.916770e-07,1.916773e-07,1.916775e-07,1.916777e-07,1.916780e-07,1.916782e-07,1.916785e-07,1.916787e-07,1.916789e-07,1.916792e-07,1.916794e-07,1.916796e-07,1.916799e-07,1.916801e-07,1.916804e-07,1.916806e-07,1.916808e-07,1.916811e-07,1.916813e-07,1.916815e-07,1.916818e-07,1.916820e-07,1.916823e-07,1.916825e-07,1.916827e-07,1.916830e-07,1.916832e-07,1.916834e-07,1.916837e-07,1.916839e-07,1.916842e-07,1.916844e-07,1.916846e-07,1.916849e-07,1.916851e-07,1.916853e-07,1.916856e-07,1.916858e-07,1.916861e-07,1.916863e-07,1.916865e-07,1.916868e-07,1.916870e-07,1.916872e-07,1.916875e-07,1.916877e-07,1.916880e-07,1.916882e-07,1.916884e-07,1.916887e-07,1.916889e-07,1.916891e-07,1.916894e-07,1.916896e-07,1.916899e-07,1.916901e-07,1.916903e-07,1.916906e-07,1.916908e-07,1.916910e-07,1.916913e-07,1.916915e-07,1.916918e-07,1.916920e-07,1.916922e-07,1.916925e-07,1.916927e-07,1.916929e-07,1.916932e-07,1.916934e-07,1.916937e-07,1.916939e-07,1.916941e-07,1.916944e-07,1.916946e-07,1.916948e-07,1.916951e-07,1.916953e-07,1.916956e-07,1.916958e-07,1.916960e-07,1.916963e-07,1.916965e-07,1.916967e-07,1.916970e-07,1.916972e-07,1.916975e-07,1.916977e-07,1.916979e-07,1.916982e-07,1.916984e-07,1.916986e-07,1.916989e-07,1.916991e-07,1.916994e-07,1.916996e-07,1.916998e-07,1.917001e-07,1.917003e-07,1.917005e-07,1.917008e-07,1.917010e-07,1.917013e-07,1.917015e-07,1.917017e-07,1.917020e-07,1.917022e-07,1.917024e-07,1.917027e-07,1.917029e-07,1.917032e-07,1.917034e-07,1.917036e-07,1.917039e-07,1.917041e-07,1.917043e-07,1.917046e-07,1.917048e-07,1.917051e-07,1.917053e-07,1.917055e-07,1.917058e-07,1.917060e-07,1.917062e-07,1.917065e-07,1.917067e-07,1.917069e-07,1.917072e-07,1.917074e-07,1.917077e-07,1.917079e-07,1.917081e-07,1.917084e-07,1.917086e-07,1.917088e-07,1.917091e-07,1.917093e-07,1.917096e-07,1.917098e-07,1.917100e-07,1.917103e-07,1.917105e-07,1.917107e-07,1.917110e-07,1.917112e-07,1.917115e-07,1.917117e-07,1.917119e-07,1.917122e-07,1.917124e-07,1.917126e-07,1.917129e-07,1.917131e-07,1.917134e-07,1.917136e-07,1.917138e-07,1.917141e-07,1.917143e-07,1.917145e-07,1.917148e-07,1.917150e-07,1.917152e-07,1.917155e-07,1.917157e-07,1.917160e-07,1.917162e-07,1.917164e-07,1.917167e-07,1.917169e-07,1.917171e-07,1.917174e-07,1.917176e-07,1.917179e-07,1.917181e-07,1.917183e-07,1.917186e-07,1.917188e-07,1.917190e-07,1.917193e-07,1.917195e-07,1.917198e-07,1.917200e-07,1.917202e-07,1.917205e-07,1.917207e-07,1.917209e-07,1.917212e-07,1.917214e-07,1.917216e-07,1.917219e-07,1.917221e-07,1.917224e-07,1.917226e-07,1.917228e-07,1.917231e-07,1.917233e-07,1.917235e-07,1.917238e-07,1.917240e-07,1.917243e-07,1.917245e-07,1.917247e-07,1.917250e-07,1.917252e-07,1.917254e-07,1.917257e-07,1.917259e-07,1.917261e-07,1.917264e-07,1.917266e-07,1.917269e-07,1.917271e-07,1.917273e-07,1.917276e-07,1.917278e-07,1.917280e-07,1.917283e-07,1.917285e-07,1.917288e-07,1.917290e-07,1.917292e-07,1.917295e-07,1.917297e-07,1.917299e-07,1.917302e-07,1.917304e-07,1.917306e-07,1.917309e-07,1.917311e-07,1.917314e-07,1.917316e-07,1.917318e-07,1.917321e-07,1.917323e-07,1.917325e-07,1.917328e-07,1.917330e-07,1.917333e-07,1.917335e-07,1.917337e-07,1.917340e-07,1.917342e-07,1.917344e-07,1.917347e-07,1.917349e-07,1.917351e-07,1.917354e-07,1.917356e-07,1.917359e-07,1.917361e-07,1.917363e-07,1.917366e-07,1.917368e-07,1.917370e-07,1.917373e-07,1.917375e-07,1.917377e-07,1.917380e-07,1.917382e-07,1.917385e-07,1.917387e-07,1.917389e-07,1.917392e-07,1.917394e-07,1.917396e-07,1.917399e-07,1.917401e-07,1.917403e-07,1.917406e-07,1.917408e-07,1.917411e-07,1.917413e-07,1.917415e-07,1.917418e-07,1.917420e-07,1.917422e-07,1.917425e-07,1.917427e-07,1.917430e-07,1.917432e-07,1.917434e-07,1.917437e-07,1.917439e-07,1.917441e-07,1.917444e-07,1.917446e-07,1.917448e-07,1.917451e-07,1.917453e-07,1.917456e-07,1.917458e-07,1.917460e-07,1.917463e-07,1.917465e-07,1.917467e-07,1.917470e-07,1.917472e-07,1.917474e-07,1.917477e-07,1.917479e-07,1.917482e-07,1.917484e-07,1.917486e-07,1.917489e-07,1.917491e-07,1.917493e-07,1.917496e-07,1.917498e-07,1.917500e-07,1.917503e-07,1.917505e-07,1.917508e-07,1.917510e-07,1.917512e-07,1.917515e-07,1.917517e-07,1.917519e-07,1.917522e-07,1.917524e-07,1.917526e-07,1.917529e-07,1.917531e-07,1.917534e-07,1.917536e-07,1.917538e-07,1.917541e-07,1.917543e-07,1.917545e-07,1.917548e-07,1.917550e-07,1.917552e-07,1.917555e-07,1.917557e-07,1.917559e-07,1.917562e-07,1.917564e-07,1.917567e-07,1.917569e-07,1.917571e-07,1.917574e-07,1.917576e-07,1.917578e-07,1.917581e-07,1.917583e-07,1.917585e-07,1.917588e-07,1.917590e-07,1.917593e-07,1.917595e-07,1.917597e-07,1.917600e-07,1.917602e-07,1.917604e-07,1.917607e-07,1.917609e-07,1.917611e-07,1.917614e-07,1.917616e-07,1.917619e-07,1.917621e-07,1.917623e-07,1.917626e-07,1.917628e-07,1.917630e-07,1.917633e-07,1.917635e-07,1.917637e-07,1.917640e-07,1.917642e-07,1.917645e-07,1.917647e-07,1.917649e-07,1.917652e-07,1.917654e-07,1.917656e-07,1.917659e-07,1.917661e-07,1.917663e-07,1.917666e-07,1.917668e-07,1.917670e-07,1.917673e-07,1.917675e-07,1.917678e-07,1.917680e-07,1.917682e-07,1.917685e-07,1.917687e-07,1.917689e-07,1.917692e-07,1.917694e-07,1.917696e-07,1.917699e-07,1.917701e-07,1.917703e-07,1.917706e-07,1.917708e-07,1.917711e-07,1.917713e-07,1.917715e-07,1.917718e-07,1.917720e-07,1.917722e-07,1.917725e-07,1.917727e-07,1.917729e-07,1.917732e-07,1.917734e-07,1.917737e-07,1.917739e-07,1.917741e-07,1.917744e-07,1.917746e-07,1.917748e-07,1.917751e-07,1.917753e-07,1.917755e-07,1.917758e-07,1.917760e-07,1.917762e-07,1.917765e-07,1.917767e-07,1.917770e-07,1.917772e-07,1.917774e-07,1.917777e-07,1.917779e-07,1.917781e-07,1.917784e-07,1.917786e-07,1.917788e-07,1.917791e-07,1.917793e-07,1.917795e-07,1.917798e-07,1.917800e-07,1.917803e-07,1.917805e-07,1.917807e-07,1.917810e-07,1.917812e-07,1.917814e-07,1.917817e-07,1.917819e-07,1.917821e-07,1.917824e-07,1.917826e-07,1.917828e-07,1.917831e-07,1.917833e-07,1.917836e-07,1.917838e-07,1.917840e-07,1.917843e-07,1.917845e-07,1.917847e-07,1.917850e-07,1.917852e-07,1.917854e-07,1.917857e-07,1.917859e-07,1.917861e-07,1.917864e-07,1.917866e-07,1.917869e-07,1.917871e-07,1.917873e-07,1.917876e-07,1.917878e-07,1.917880e-07,1.917883e-07,1.917885e-07,1.917887e-07,1.917890e-07,1.917892e-07,1.917894e-07,1.917897e-07,1.917899e-07,1.917902e-07,1.917904e-07,1.917906e-07,1.917909e-07,1.917911e-07,1.917913e-07,1.917916e-07,1.917918e-07,1.917920e-07,1.917923e-07,1.917925e-07,1.917927e-07,1.917930e-07,1.917932e-07,1.917934e-07,1.917937e-07,1.917939e-07,1.917942e-07,1.917944e-07,1.917946e-07,1.917949e-07,1.917951e-07,1.917953e-07,1.917956e-07,1.917958e-07,1.917960e-07,1.917963e-07,1.917965e-07,1.917967e-07,1.917970e-07,1.917972e-07,1.917975e-07,1.917977e-07,1.917979e-07,1.917982e-07,1.917984e-07,1.917986e-07,1.917989e-07,1.917991e-07,1.917993e-07,1.917996e-07,1.917998e-07,1.918000e-07,1.918003e-07,1.918005e-07,1.918007e-07,1.918010e-07,1.918012e-07,1.918015e-07,1.918017e-07,1.918019e-07,1.918022e-07,1.918024e-07,1.918026e-07,1.918029e-07,1.918031e-07,1.918033e-07,1.918036e-07,1.918038e-07,1.918040e-07,1.918043e-07,1.918045e-07,1.918047e-07,1.918050e-07,1.918052e-07,1.918055e-07,1.918057e-07,1.918059e-07,1.918062e-07,1.918064e-07,1.918066e-07,1.918069e-07,1.918071e-07,1.918073e-07,1.918076e-07,1.918078e-07,1.918080e-07,1.918083e-07,1.918085e-07,1.918087e-07,1.918090e-07,1.918092e-07,1.918094e-07,1.918097e-07,1.918099e-07,1.918102e-07,1.918104e-07,1.918106e-07,1.918109e-07,1.918111e-07,1.918113e-07,1.918116e-07,1.918118e-07,1.918120e-07,1.918123e-07,1.918125e-07,1.918127e-07,1.918130e-07,1.918132e-07,1.918134e-07,1.918137e-07,1.918139e-07,1.918142e-07,1.918144e-07,1.918146e-07,1.918149e-07,1.918151e-07,1.918153e-07,1.918156e-07,1.918158e-07,1.918160e-07,1.918163e-07,1.918165e-07,1.918167e-07,1.918170e-07,1.918172e-07,1.918174e-07,1.918177e-07,1.918179e-07,1.918181e-07,1.918184e-07,1.918186e-07,1.918189e-07,1.918191e-07,1.918193e-07,1.918196e-07,1.918198e-07,1.918200e-07,1.918203e-07,1.918205e-07,1.918207e-07,1.918210e-07,1.918212e-07,1.918214e-07,1.918217e-07,1.918219e-07,1.918221e-07,1.918224e-07,1.918226e-07,1.918228e-07,1.918231e-07,1.918233e-07,1.918235e-07,1.918238e-07,1.918240e-07,1.918243e-07,1.918245e-07,1.918247e-07,1.918250e-07,1.918252e-07,1.918254e-07,1.918257e-07,1.918259e-07,1.918261e-07,1.918264e-07,1.918266e-07,1.918268e-07,1.918271e-07,1.918273e-07,1.918275e-07,1.918278e-07,1.918280e-07,1.918282e-07,1.918285e-07,1.918287e-07,1.918289e-07,1.918292e-07,1.918294e-07,1.918297e-07,1.918299e-07,1.918301e-07,1.918304e-07,1.918306e-07,1.918308e-07,1.918311e-07,1.918313e-07,1.918315e-07,1.918318e-07,1.918320e-07,1.918322e-07,1.918325e-07,1.918327e-07,1.918329e-07,1.918332e-07,1.918334e-07,1.918336e-07,1.918339e-07,1.918341e-07,1.918343e-07,1.918346e-07,1.918348e-07,1.918351e-07,1.918353e-07,1.918355e-07,1.918358e-07,1.918360e-07,1.918362e-07,1.918365e-07,1.918367e-07,1.918369e-07,1.918372e-07,1.918374e-07,1.918376e-07,1.918379e-07,1.918381e-07,1.918383e-07,1.918386e-07,1.918388e-07,1.918390e-07,1.918393e-07,1.918395e-07,1.918397e-07,1.918400e-07,1.918402e-07,1.918404e-07,1.918407e-07,1.918409e-07,1.918411e-07,1.918414e-07,1.918416e-07,1.918419e-07,1.918421e-07,1.918423e-07,1.918426e-07,1.918428e-07,1.918430e-07,1.918433e-07,1.918435e-07,1.918437e-07,1.918440e-07,1.918442e-07,1.918444e-07,1.918447e-07,1.918449e-07,1.918451e-07,1.918454e-07,1.918456e-07,1.918458e-07,1.918461e-07,1.918463e-07,1.918465e-07,1.918468e-07,1.918470e-07,1.918472e-07,1.918475e-07,1.918477e-07,1.918479e-07,1.918482e-07,1.918484e-07,1.918487e-07,1.918489e-07,1.918491e-07,1.918494e-07,1.918496e-07,1.918498e-07,1.918501e-07,1.918503e-07,1.918505e-07,1.918508e-07,1.918510e-07,1.918512e-07,1.918515e-07,1.918517e-07,1.918519e-07,1.918522e-07,1.918524e-07,1.918526e-07,1.918529e-07,1.918531e-07,1.918533e-07,1.918536e-07,1.918538e-07,1.918540e-07,1.918543e-07,1.918545e-07,1.918547e-07,1.918550e-07,1.918552e-07,1.918554e-07,1.918557e-07,1.918559e-07,1.918561e-07,1.918564e-07,1.918566e-07,1.918569e-07,1.918571e-07,1.918573e-07,1.918576e-07,1.918578e-07,1.918580e-07,1.918583e-07,1.918585e-07,1.918587e-07,1.918590e-07,1.918592e-07,1.918594e-07,1.918597e-07,1.918599e-07,1.918601e-07,1.918604e-07,1.918606e-07,1.918608e-07,1.918611e-07,1.918613e-07,1.918615e-07,1.918618e-07,1.918620e-07,1.918622e-07,1.918625e-07,1.918627e-07,1.918629e-07,1.918632e-07,1.918634e-07,1.918636e-07,1.918639e-07,1.918641e-07,1.918643e-07,1.918646e-07,1.918648e-07,1.918650e-07,1.918653e-07,1.918655e-07,1.918657e-07,1.918660e-07,1.918662e-07,1.918664e-07,1.918667e-07,1.918669e-07,1.918672e-07,1.918674e-07,1.918676e-07,1.918679e-07,1.918681e-07,1.918683e-07,1.918686e-07,1.918688e-07,1.918690e-07,1.918693e-07,1.918695e-07,1.918697e-07,1.918700e-07,1.918702e-07,1.918704e-07,1.918707e-07,1.918709e-07,1.918711e-07,1.918714e-07,1.918716e-07,1.918718e-07,1.918721e-07,1.918723e-07,1.918725e-07,1.918728e-07,1.918730e-07,1.918732e-07,1.918735e-07,1.918737e-07,1.918739e-07,1.918742e-07,1.918744e-07,1.918746e-07,1.918749e-07,1.918751e-07,1.918753e-07,1.918756e-07,1.918758e-07,1.918760e-07,1.918763e-07,1.918765e-07,1.918767e-07,1.918770e-07,1.918772e-07,1.918774e-07,1.918777e-07,1.918779e-07,1.918781e-07,1.918784e-07,1.918786e-07,1.918788e-07,1.918791e-07,1.918793e-07,1.918795e-07,1.918798e-07,1.918800e-07,1.918802e-07,1.918805e-07,1.918807e-07,1.918809e-07,1.918812e-07,1.918814e-07,1.918816e-07,1.918819e-07,1.918821e-07,1.918823e-07,1.918826e-07,1.918828e-07,1.918831e-07,1.918833e-07,1.918835e-07,1.918838e-07,1.918840e-07,1.918842e-07,1.918845e-07,1.918847e-07,1.918849e-07,1.918852e-07,1.918854e-07,1.918856e-07,1.918859e-07,1.918861e-07,1.918863e-07,1.918866e-07,1.918868e-07,1.918870e-07,1.918873e-07,1.918875e-07,1.918877e-07,1.918880e-07,1.918882e-07,1.918884e-07,1.918887e-07,1.918889e-07,1.918891e-07,1.918894e-07,1.918896e-07,1.918898e-07,1.918901e-07,1.918903e-07,1.918905e-07,1.918908e-07,1.918910e-07,1.918912e-07,1.918915e-07,1.918917e-07,1.918919e-07,1.918922e-07,1.918924e-07,1.918926e-07,1.918929e-07,1.918931e-07,1.918933e-07,1.918936e-07,1.918938e-07,1.918940e-07,1.918943e-07,1.918945e-07,1.918947e-07,1.918950e-07,1.918952e-07,1.918954e-07,1.918957e-07,1.918959e-07,1.918961e-07,1.918964e-07,1.918966e-07,1.918968e-07,1.918971e-07,1.918973e-07,1.918975e-07,1.918978e-07,1.918980e-07,1.918982e-07,1.918985e-07,1.918987e-07,1.918989e-07,1.918992e-07,1.918994e-07,1.918996e-07,1.918999e-07,1.919001e-07,1.919003e-07,1.919006e-07,1.919008e-07,1.919010e-07,1.919013e-07,1.919015e-07,1.919017e-07,1.919020e-07,1.919022e-07,1.919024e-07,1.919027e-07,1.919029e-07,1.919031e-07,1.919034e-07,1.919036e-07,1.919038e-07,1.919041e-07,1.919043e-07,1.919045e-07,1.919048e-07,1.919050e-07,1.919052e-07,1.919055e-07,1.919057e-07,1.919059e-07,1.919062e-07,1.919064e-07,1.919066e-07,1.919069e-07,1.919071e-07,1.919073e-07,1.919076e-07,1.919078e-07,1.919080e-07,1.919083e-07,1.919085e-07,1.919087e-07,1.919090e-07,1.919092e-07,1.919094e-07,1.919097e-07,1.919099e-07,1.919101e-07,1.919104e-07,1.919106e-07,1.919108e-07,1.919111e-07,1.919113e-07,1.919115e-07,1.919118e-07,1.919120e-07,1.919122e-07,1.919125e-07,1.919127e-07,1.919129e-07,1.919132e-07,1.919134e-07,1.919136e-07,1.919139e-07,1.919141e-07,1.919143e-07,1.919146e-07,1.919148e-07,1.919150e-07,1.919153e-07,1.919155e-07,1.919157e-07,1.919160e-07,1.919162e-07,1.919164e-07,1.919166e-07,1.919169e-07,1.919171e-07,1.919173e-07,1.919176e-07,1.919178e-07,1.919180e-07,1.919183e-07,1.919185e-07,1.919187e-07,1.919190e-07,1.919192e-07,1.919194e-07,1.919197e-07,1.919199e-07,1.919201e-07,1.919204e-07,1.919206e-07,1.919208e-07,1.919211e-07,1.919213e-07,1.919215e-07,1.919218e-07,1.919220e-07,1.919222e-07,1.919225e-07,1.919227e-07,1.919229e-07,1.919232e-07,1.919234e-07,1.919236e-07,1.919239e-07,1.919241e-07,1.919243e-07,1.919246e-07,1.919248e-07,1.919250e-07,1.919253e-07,1.919255e-07,1.919257e-07,1.919260e-07,1.919262e-07,1.919264e-07,1.919267e-07,1.919269e-07,1.919271e-07,1.919274e-07,1.919276e-07,1.919278e-07,1.919281e-07,1.919283e-07,1.919285e-07,1.919288e-07,1.919290e-07,1.919292e-07,1.919295e-07,1.919297e-07,1.919299e-07,1.919302e-07,1.919304e-07,1.919306e-07,1.919309e-07,1.919311e-07,1.919313e-07,1.919316e-07,1.919318e-07,1.919320e-07,1.919322e-07,1.919325e-07,1.919327e-07,1.919329e-07,1.919332e-07,1.919334e-07,1.919336e-07,1.919339e-07,1.919341e-07,1.919343e-07,1.919346e-07,1.919348e-07,1.919350e-07,1.919353e-07,1.919355e-07,1.919357e-07,1.919360e-07,1.919362e-07,1.919364e-07,1.919367e-07,1.919369e-07,1.919371e-07,1.919374e-07,1.919376e-07,1.919378e-07,1.919381e-07,1.919383e-07,1.919385e-07,1.919388e-07,1.919390e-07,1.919392e-07,1.919395e-07,1.919397e-07,1.919399e-07,1.919402e-07,1.919404e-07,1.919406e-07,1.919409e-07,1.919411e-07,1.919413e-07,1.919416e-07,1.919418e-07,1.919420e-07,1.919423e-07,1.919425e-07,1.919427e-07,1.919429e-07,1.919432e-07,1.919434e-07,1.919436e-07,1.919439e-07,1.919441e-07,1.919443e-07,1.919446e-07,1.919448e-07,1.919450e-07,1.919453e-07,1.919455e-07,1.919457e-07,1.919460e-07,1.919462e-07,1.919464e-07,1.919467e-07,1.919469e-07,1.919471e-07,1.919474e-07,1.919476e-07,1.919478e-07,1.919481e-07,1.919483e-07,1.919485e-07,1.919488e-07,1.919490e-07,1.919492e-07,1.919495e-07,1.919497e-07,1.919499e-07,1.919502e-07,1.919504e-07,1.919506e-07,1.919508e-07,1.919511e-07,1.919513e-07,1.919515e-07,1.919518e-07,1.919520e-07,1.919522e-07,1.919525e-07,1.919527e-07,1.919529e-07,1.919532e-07,1.919534e-07,1.919536e-07,1.919539e-07,1.919541e-07,1.919543e-07,1.919546e-07,1.919548e-07,1.919550e-07,1.919553e-07,1.919555e-07,1.919557e-07,1.919560e-07,1.919562e-07,1.919564e-07,1.919567e-07,1.919569e-07,1.919571e-07,1.919574e-07,1.919576e-07,1.919578e-07,1.919580e-07,1.919583e-07,1.919585e-07,1.919587e-07,1.919590e-07,1.919592e-07,1.919594e-07,1.919597e-07,1.919599e-07,1.919601e-07,1.919604e-07,1.919606e-07,1.919608e-07,1.919611e-07,1.919613e-07,1.919615e-07,1.919618e-07,1.919620e-07,1.919622e-07,1.919625e-07,1.919627e-07,1.919629e-07,1.919632e-07,1.919634e-07,1.919636e-07,1.919639e-07,1.919641e-07,1.919643e-07,1.919645e-07,1.919648e-07,1.919650e-07,1.919652e-07,1.919655e-07,1.919657e-07,1.919659e-07,1.919662e-07,1.919664e-07,1.919666e-07,1.919669e-07,1.919671e-07,1.919673e-07,1.919676e-07,1.919678e-07,1.919680e-07,1.919683e-07,1.919685e-07,1.919687e-07,1.919690e-07,1.919692e-07,1.919694e-07,1.919697e-07,1.919699e-07,1.919701e-07,1.919703e-07,1.919706e-07,1.919708e-07,1.919710e-07,1.919713e-07,1.919715e-07,1.919717e-07,1.919720e-07,1.919722e-07,1.919724e-07,1.919727e-07,1.919729e-07,1.919731e-07,1.919734e-07,1.919736e-07,1.919738e-07,1.919741e-07,1.919743e-07,1.919745e-07,1.919748e-07,1.919750e-07,1.919752e-07,1.919754e-07,1.919757e-07,1.919759e-07,1.919761e-07,1.919764e-07,1.919766e-07,1.919768e-07,1.919771e-07,1.919773e-07,1.919775e-07,1.919778e-07,1.919780e-07,1.919782e-07,1.919785e-07,1.919787e-07,1.919789e-07,1.919792e-07,1.919794e-07,1.919796e-07,1.919799e-07,1.919801e-07,1.919803e-07,1.919805e-07,1.919808e-07,1.919810e-07,1.919812e-07,1.919815e-07,1.919817e-07,1.919819e-07,1.919822e-07,1.919824e-07,1.919826e-07,1.919829e-07,1.919831e-07,1.919833e-07,1.919836e-07,1.919838e-07,1.919840e-07,1.919843e-07,1.919845e-07,1.919847e-07,1.919850e-07,1.919852e-07,1.919854e-07,1.919856e-07,1.919859e-07,1.919861e-07,1.919863e-07,1.919866e-07,1.919868e-07,1.919870e-07,1.919873e-07,1.919875e-07,1.919877e-07,1.919880e-07,1.919882e-07,1.919884e-07,1.919887e-07,1.919889e-07,1.919891e-07,1.919894e-07,1.919896e-07,1.919898e-07,1.919900e-07,1.919903e-07,1.919905e-07,1.919907e-07,1.919910e-07,1.919912e-07,1.919914e-07,1.919917e-07,1.919919e-07,1.919921e-07,1.919924e-07,1.919926e-07,1.919928e-07,1.919931e-07,1.919933e-07,1.919935e-07,1.919937e-07,1.919940e-07,1.919942e-07,1.919944e-07,1.919947e-07,1.919949e-07,1.919951e-07,1.919954e-07,1.919956e-07,1.919958e-07,1.919961e-07,1.919963e-07,1.919965e-07,1.919968e-07,1.919970e-07,1.919972e-07,1.919975e-07,1.919977e-07,1.919979e-07,1.919981e-07,1.919984e-07,1.919986e-07,1.919988e-07,1.919991e-07,1.919993e-07,1.919995e-07,1.919998e-07,1.920000e-07,1.920002e-07,1.920005e-07,1.920007e-07,1.920009e-07,1.920012e-07,1.920014e-07,1.920016e-07,1.920018e-07,1.920021e-07,1.920023e-07,1.920025e-07,1.920028e-07,1.920030e-07,1.920032e-07,1.920035e-07,1.920037e-07,1.920039e-07,1.920042e-07,1.920044e-07,1.920046e-07,1.920049e-07,1.920051e-07,1.920053e-07,1.920055e-07,1.920058e-07,1.920060e-07,1.920062e-07,1.920065e-07,1.920067e-07,1.920069e-07,1.920072e-07,1.920074e-07,1.920076e-07,1.920079e-07,1.920081e-07,1.920083e-07,1.920086e-07,1.920088e-07,1.920090e-07,1.920092e-07,1.920095e-07,1.920097e-07,1.920099e-07,1.920102e-07,1.920104e-07,1.920106e-07,1.920109e-07,1.920111e-07,1.920113e-07,1.920116e-07,1.920118e-07,1.920120e-07,1.920123e-07,1.920125e-07,1.920127e-07,1.920129e-07,1.920132e-07,1.920134e-07,1.920136e-07,1.920139e-07,1.920141e-07,1.920143e-07,1.920146e-07,1.920148e-07,1.920150e-07,1.920153e-07,1.920155e-07,1.920157e-07,1.920159e-07,1.920162e-07,1.920164e-07,1.920166e-07,1.920169e-07,1.920171e-07,1.920173e-07,1.920176e-07,1.920178e-07,1.920180e-07,1.920183e-07,1.920185e-07,1.920187e-07,1.920190e-07,1.920192e-07,1.920194e-07,1.920196e-07,1.920199e-07,1.920201e-07,1.920203e-07,1.920206e-07,1.920208e-07,1.920210e-07,1.920213e-07,1.920215e-07,1.920217e-07,1.920220e-07,1.920222e-07,1.920224e-07,1.920226e-07,1.920229e-07,1.920231e-07,1.920233e-07,1.920236e-07,1.920238e-07,1.920240e-07,1.920243e-07,1.920245e-07,1.920247e-07,1.920250e-07,1.920252e-07,1.920254e-07,1.920256e-07,1.920259e-07,1.920261e-07,1.920263e-07,1.920266e-07,1.920268e-07,1.920270e-07,1.920273e-07,1.920275e-07,1.920277e-07,1.920280e-07,1.920282e-07,1.920284e-07,1.920286e-07,1.920289e-07,1.920291e-07,1.920293e-07,1.920296e-07,1.920298e-07,1.920300e-07,1.920303e-07,1.920305e-07,1.920307e-07,1.920310e-07,1.920312e-07,1.920314e-07,1.920316e-07,1.920319e-07,1.920321e-07,1.920323e-07,1.920326e-07,1.920328e-07,1.920330e-07,1.920333e-07,1.920335e-07,1.920337e-07,1.920340e-07,1.920342e-07,1.920344e-07,1.920346e-07,1.920349e-07,1.920351e-07,1.920353e-07,1.920356e-07,1.920358e-07,1.920360e-07,1.920363e-07,1.920365e-07,1.920367e-07,1.920370e-07,1.920372e-07,1.920374e-07,1.920376e-07,1.920379e-07,1.920381e-07,1.920383e-07,1.920386e-07,1.920388e-07,1.920390e-07,1.920393e-07,1.920395e-07,1.920397e-07,1.920400e-07,1.920402e-07,1.920404e-07,1.920406e-07,1.920409e-07,1.920411e-07,1.920413e-07,1.920416e-07,1.920418e-07,1.920420e-07,1.920423e-07,1.920425e-07,1.920427e-07,1.920429e-07,1.920432e-07,1.920434e-07,1.920436e-07,1.920439e-07,1.920441e-07,1.920443e-07,1.920446e-07,1.920448e-07,1.920450e-07,1.920453e-07,1.920455e-07,1.920457e-07,1.920459e-07,1.920462e-07,1.920464e-07,1.920466e-07,1.920469e-07,1.920471e-07,1.920473e-07,1.920476e-07,1.920478e-07,1.920480e-07,1.920482e-07,1.920485e-07,1.920487e-07,1.920489e-07,1.920492e-07,1.920494e-07,1.920496e-07,1.920499e-07,1.920501e-07,1.920503e-07,1.920506e-07,1.920508e-07,1.920510e-07,1.920512e-07,1.920515e-07,1.920517e-07,1.920519e-07,1.920522e-07,1.920524e-07,1.920526e-07,1.920529e-07,1.920531e-07,1.920533e-07,1.920535e-07,1.920538e-07,1.920540e-07,1.920542e-07,1.920545e-07,1.920547e-07,1.920549e-07,1.920552e-07,1.920554e-07,1.920556e-07,1.920558e-07,1.920561e-07,1.920563e-07,1.920565e-07,1.920568e-07,1.920570e-07,1.920572e-07,1.920575e-07,1.920577e-07,1.920579e-07,1.920582e-07,1.920584e-07,1.920586e-07,1.920588e-07,1.920591e-07,1.920593e-07,1.920595e-07,1.920598e-07,1.920600e-07,1.920602e-07,1.920605e-07,1.920607e-07,1.920609e-07,1.920611e-07,1.920614e-07,1.920616e-07,1.920618e-07,1.920621e-07,1.920623e-07,1.920625e-07,1.920628e-07,1.920630e-07,1.920632e-07,1.920634e-07,1.920637e-07,1.920639e-07,1.920641e-07,1.920644e-07,1.920646e-07,1.920648e-07,1.920651e-07,1.920653e-07,1.920655e-07,1.920657e-07,1.920660e-07,1.920662e-07,1.920664e-07,1.920667e-07,1.920669e-07,1.920671e-07,1.920674e-07,1.920676e-07,1.920678e-07,1.920680e-07,1.920683e-07,1.920685e-07,1.920687e-07,1.920690e-07,1.920692e-07,1.920694e-07,1.920697e-07,1.920699e-07,1.920701e-07,1.920703e-07,1.920706e-07,1.920708e-07,1.920710e-07,1.920713e-07,1.920715e-07,1.920717e-07,1.920720e-07,1.920722e-07,1.920724e-07,1.920726e-07,1.920729e-07,1.920731e-07,1.920733e-07,1.920736e-07,1.920738e-07,1.920740e-07,1.920743e-07,1.920745e-07,1.920747e-07,1.920749e-07,1.920752e-07,1.920754e-07,1.920756e-07,1.920759e-07,1.920761e-07,1.920763e-07,1.920766e-07,1.920768e-07,1.920770e-07,1.920772e-07,1.920775e-07,1.920777e-07,1.920779e-07,1.920782e-07,1.920784e-07,1.920786e-07,1.920788e-07,1.920791e-07,1.920793e-07,1.920795e-07,1.920798e-07,1.920800e-07,1.920802e-07,1.920805e-07,1.920807e-07,1.920809e-07,1.920811e-07,1.920814e-07,1.920816e-07,1.920818e-07,1.920821e-07,1.920823e-07,1.920825e-07,1.920828e-07,1.920830e-07,1.920832e-07,1.920834e-07,1.920837e-07,1.920839e-07,1.920841e-07,1.920844e-07,1.920846e-07,1.920848e-07,1.920851e-07,1.920853e-07,1.920855e-07,1.920857e-07,1.920860e-07,1.920862e-07,1.920864e-07,1.920867e-07,1.920869e-07,1.920871e-07,1.920873e-07,1.920876e-07,1.920878e-07,1.920880e-07,1.920883e-07,1.920885e-07,1.920887e-07,1.920890e-07,1.920892e-07,1.920894e-07,1.920896e-07,1.920899e-07,1.920901e-07,1.920903e-07,1.920906e-07,1.920908e-07,1.920910e-07,1.920913e-07,1.920915e-07,1.920917e-07,1.920919e-07,1.920922e-07,1.920924e-07,1.920926e-07,1.920929e-07,1.920931e-07,1.920933e-07,1.920935e-07,1.920938e-07,1.920940e-07,1.920942e-07,1.920945e-07,1.920947e-07,1.920949e-07,1.920952e-07,1.920954e-07,1.920956e-07,1.920958e-07,1.920961e-07,1.920963e-07,1.920965e-07,1.920968e-07,1.920970e-07,1.920972e-07,1.920974e-07,1.920977e-07,1.920979e-07,1.920981e-07,1.920984e-07,1.920986e-07,1.920988e-07,1.920991e-07,1.920993e-07,1.920995e-07,1.920997e-07,1.921000e-07,1.921002e-07,1.921004e-07,1.921007e-07,1.921009e-07,1.921011e-07,1.921013e-07,1.921016e-07,1.921018e-07,1.921020e-07,1.921023e-07,1.921025e-07,1.921027e-07,1.921030e-07,1.921032e-07,1.921034e-07,1.921036e-07,1.921039e-07,1.921041e-07,1.921043e-07,1.921046e-07,1.921048e-07,1.921050e-07,1.921052e-07,1.921055e-07,1.921057e-07,1.921059e-07,1.921062e-07,1.921064e-07,1.921066e-07,1.921068e-07,1.921071e-07,1.921073e-07,1.921075e-07,1.921078e-07,1.921080e-07,1.921082e-07,1.921085e-07,1.921087e-07,1.921089e-07,1.921091e-07,1.921094e-07,1.921096e-07,1.921098e-07,1.921101e-07,1.921103e-07,1.921105e-07,1.921107e-07,1.921110e-07,1.921112e-07,1.921114e-07,1.921117e-07,1.921119e-07,1.921121e-07,1.921124e-07,1.921126e-07,1.921128e-07,1.921130e-07,1.921133e-07,1.921135e-07,1.921137e-07,1.921140e-07,1.921142e-07,1.921144e-07,1.921146e-07,1.921149e-07,1.921151e-07,1.921153e-07,1.921156e-07,1.921158e-07,1.921160e-07,1.921162e-07,1.921165e-07,1.921167e-07,1.921169e-07,1.921172e-07,1.921174e-07,1.921176e-07,1.921178e-07,1.921181e-07,1.921183e-07,1.921185e-07,1.921188e-07,1.921190e-07,1.921192e-07,1.921195e-07,1.921197e-07,1.921199e-07,1.921201e-07,1.921204e-07,1.921206e-07,1.921208e-07,1.921211e-07,1.921213e-07,1.921215e-07,1.921217e-07,1.921220e-07,1.921222e-07,1.921224e-07,1.921227e-07,1.921229e-07,1.921231e-07,1.921233e-07,1.921236e-07,1.921238e-07,1.921240e-07,1.921243e-07,1.921245e-07,1.921247e-07,1.921249e-07,1.921252e-07,1.921254e-07,1.921256e-07,1.921259e-07,1.921261e-07,1.921263e-07,1.921265e-07,1.921268e-07,1.921270e-07,1.921272e-07,1.921275e-07,1.921277e-07,1.921279e-07,1.921281e-07,1.921284e-07,1.921286e-07,1.921288e-07,1.921291e-07,1.921293e-07,1.921295e-07,1.921298e-07,1.921300e-07,1.921302e-07,1.921304e-07,1.921307e-07,1.921309e-07,1.921311e-07,1.921314e-07,1.921316e-07,1.921318e-07,1.921320e-07,1.921323e-07,1.921325e-07,1.921327e-07,1.921330e-07,1.921332e-07,1.921334e-07,1.921336e-07,1.921339e-07,1.921341e-07,1.921343e-07,1.921346e-07,1.921348e-07,1.921350e-07,1.921352e-07,1.921355e-07,1.921357e-07,1.921359e-07,1.921362e-07,1.921364e-07,1.921366e-07,1.921368e-07,1.921371e-07,1.921373e-07,1.921375e-07,1.921378e-07,1.921380e-07,1.921382e-07,1.921384e-07,1.921387e-07,1.921389e-07,1.921391e-07,1.921394e-07,1.921396e-07,1.921398e-07,1.921400e-07,1.921403e-07,1.921405e-07,1.921407e-07,1.921410e-07,1.921412e-07,1.921414e-07,1.921416e-07,1.921419e-07,1.921421e-07,1.921423e-07,1.921426e-07,1.921428e-07,1.921430e-07,1.921432e-07,1.921435e-07,1.921437e-07,1.921439e-07,1.921442e-07,1.921444e-07,1.921446e-07,1.921448e-07,1.921451e-07,1.921453e-07,1.921455e-07,1.921458e-07,1.921460e-07,1.921462e-07,1.921464e-07,1.921467e-07,1.921469e-07,1.921471e-07,1.921474e-07,1.921476e-07,1.921478e-07,1.921480e-07,1.921483e-07,1.921485e-07,1.921487e-07,1.921490e-07,1.921492e-07,1.921494e-07,1.921496e-07,1.921499e-07,1.921501e-07,1.921503e-07,1.921506e-07,1.921508e-07,1.921510e-07,1.921512e-07,1.921515e-07,1.921517e-07,1.921519e-07,1.921522e-07,1.921524e-07,1.921526e-07,1.921528e-07,1.921531e-07,1.921533e-07,1.921535e-07,1.921537e-07,1.921540e-07,1.921542e-07,1.921544e-07,1.921547e-07,1.921549e-07,1.921551e-07,1.921553e-07,1.921556e-07,1.921558e-07,1.921560e-07,1.921563e-07,1.921565e-07,1.921567e-07,1.921569e-07,1.921572e-07,1.921574e-07,1.921576e-07,1.921579e-07,1.921581e-07,1.921583e-07,1.921585e-07,1.921588e-07,1.921590e-07,1.921592e-07,1.921595e-07,1.921597e-07,1.921599e-07,1.921601e-07,1.921604e-07,1.921606e-07,1.921608e-07,1.921611e-07,1.921613e-07,1.921615e-07,1.921617e-07,1.921620e-07,1.921622e-07,1.921624e-07,1.921627e-07,1.921629e-07,1.921631e-07,1.921633e-07,1.921636e-07,1.921638e-07,1.921640e-07,1.921642e-07,1.921645e-07,1.921647e-07,1.921649e-07,1.921652e-07,1.921654e-07,1.921656e-07,1.921658e-07,1.921661e-07,1.921663e-07,1.921665e-07,1.921668e-07,1.921670e-07,1.921672e-07,1.921674e-07,1.921677e-07,1.921679e-07,1.921681e-07,1.921684e-07,1.921686e-07,1.921688e-07,1.921690e-07,1.921693e-07,1.921695e-07,1.921697e-07,1.921699e-07,1.921702e-07,1.921704e-07,1.921706e-07,1.921709e-07,1.921711e-07,1.921713e-07,1.921715e-07,1.921718e-07,1.921720e-07,1.921722e-07,1.921725e-07,1.921727e-07,1.921729e-07,1.921731e-07,1.921734e-07,1.921736e-07,1.921738e-07,1.921741e-07,1.921743e-07,1.921745e-07,1.921747e-07,1.921750e-07,1.921752e-07,1.921754e-07,1.921756e-07,1.921759e-07,1.921761e-07,1.921763e-07,1.921766e-07,1.921768e-07,1.921770e-07,1.921772e-07,1.921775e-07,1.921777e-07,1.921779e-07,1.921782e-07,1.921784e-07,1.921786e-07,1.921788e-07,1.921791e-07,1.921793e-07,1.921795e-07,1.921797e-07,1.921800e-07,1.921802e-07,1.921804e-07,1.921807e-07,1.921809e-07,1.921811e-07,1.921813e-07,1.921816e-07,1.921818e-07,1.921820e-07,1.921823e-07,1.921825e-07,1.921827e-07,1.921829e-07,1.921832e-07,1.921834e-07,1.921836e-07,1.921838e-07,1.921841e-07,1.921843e-07,1.921845e-07,1.921848e-07,1.921850e-07,1.921852e-07,1.921854e-07,1.921857e-07,1.921859e-07,1.921861e-07,1.921864e-07,1.921866e-07,1.921868e-07,1.921870e-07,1.921873e-07,1.921875e-07,1.921877e-07,1.921879e-07,1.921882e-07,1.921884e-07,1.921886e-07,1.921889e-07,1.921891e-07,1.921893e-07,1.921895e-07,1.921898e-07,1.921900e-07,1.921902e-07,1.921905e-07,1.921907e-07,1.921909e-07,1.921911e-07,1.921914e-07,1.921916e-07,1.921918e-07,1.921920e-07,1.921923e-07,1.921925e-07,1.921927e-07,1.921930e-07,1.921932e-07,1.921934e-07,1.921936e-07,1.921939e-07,1.921941e-07,1.921943e-07,1.921945e-07,1.921948e-07,1.921950e-07,1.921952e-07,1.921955e-07,1.921957e-07,1.921959e-07,1.921961e-07,1.921964e-07,1.921966e-07,1.921968e-07,1.921970e-07,1.921973e-07,1.921975e-07,1.921977e-07,1.921980e-07,1.921982e-07,1.921984e-07,1.921986e-07,1.921989e-07,1.921991e-07,1.921993e-07,1.921996e-07,1.921998e-07,1.922000e-07,1.922002e-07,1.922005e-07,1.922007e-07,1.922009e-07,1.922011e-07,1.922014e-07,1.922016e-07,1.922018e-07,1.922021e-07,1.922023e-07,1.922025e-07,1.922027e-07,1.922030e-07,1.922032e-07,1.922034e-07,1.922036e-07,1.922039e-07,1.922041e-07,1.922043e-07,1.922046e-07,1.922048e-07,1.922050e-07,1.922052e-07,1.922055e-07,1.922057e-07,1.922059e-07,1.922061e-07,1.922064e-07,1.922066e-07,1.922068e-07,1.922071e-07,1.922073e-07,1.922075e-07,1.922077e-07,1.922080e-07,1.922082e-07,1.922084e-07,1.922086e-07,1.922089e-07,1.922091e-07,1.922093e-07,1.922096e-07,1.922098e-07,1.922100e-07,1.922102e-07,1.922105e-07,1.922107e-07,1.922109e-07,1.922111e-07,1.922114e-07,1.922116e-07,1.922118e-07,1.922121e-07,1.922123e-07,1.922125e-07,1.922127e-07,1.922130e-07,1.922132e-07,1.922134e-07,1.922136e-07,1.922139e-07,1.922141e-07,1.922143e-07,1.922146e-07,1.922148e-07,1.922150e-07,1.922152e-07,1.922155e-07,1.922157e-07,1.922159e-07,1.922161e-07,1.922164e-07,1.922166e-07,1.922168e-07,1.922171e-07,1.922173e-07,1.922175e-07,1.922177e-07,1.922180e-07,1.922182e-07,1.922184e-07,1.922186e-07,1.922189e-07,1.922191e-07,1.922193e-07,1.922195e-07,1.922198e-07,1.922200e-07,1.922202e-07,1.922205e-07,1.922207e-07,1.922209e-07,1.922211e-07,1.922214e-07,1.922216e-07,1.922218e-07,1.922220e-07,1.922223e-07,1.922225e-07,1.922227e-07,1.922230e-07,1.922232e-07,1.922234e-07,1.922236e-07,1.922239e-07,1.922241e-07,1.922243e-07,1.922245e-07,1.922248e-07,1.922250e-07,1.922252e-07,1.922254e-07,1.922257e-07,1.922259e-07,1.922261e-07,1.922264e-07,1.922266e-07,1.922268e-07,1.922270e-07,1.922273e-07,1.922275e-07,1.922277e-07,1.922279e-07,1.922282e-07,1.922284e-07,1.922286e-07,1.922289e-07,1.922291e-07,1.922293e-07,1.922295e-07,1.922298e-07,1.922300e-07,1.922302e-07,1.922304e-07,1.922307e-07,1.922309e-07,1.922311e-07,1.922313e-07,1.922316e-07,1.922318e-07,1.922320e-07,1.922323e-07,1.922325e-07,1.922327e-07,1.922329e-07,1.922332e-07,1.922334e-07,1.922336e-07,1.922338e-07,1.922341e-07,1.922343e-07,1.922345e-07,1.922348e-07,1.922350e-07,1.922352e-07,1.922354e-07,1.922357e-07,1.922359e-07,1.922361e-07,1.922363e-07,1.922366e-07,1.922368e-07,1.922370e-07,1.922372e-07,1.922375e-07,1.922377e-07,1.922379e-07,1.922382e-07,1.922384e-07,1.922386e-07,1.922388e-07,1.922391e-07,1.922393e-07,1.922395e-07,1.922397e-07,1.922400e-07,1.922402e-07,1.922404e-07,1.922406e-07,1.922409e-07,1.922411e-07,1.922413e-07,1.922416e-07,1.922418e-07,1.922420e-07,1.922422e-07,1.922425e-07,1.922427e-07,1.922429e-07,1.922431e-07,1.922434e-07,1.922436e-07,1.922438e-07,1.922440e-07,1.922443e-07,1.922445e-07,1.922447e-07,1.922449e-07,1.922452e-07,1.922454e-07,1.922456e-07,1.922459e-07,1.922461e-07,1.922463e-07,1.922465e-07,1.922468e-07,1.922470e-07,1.922472e-07,1.922474e-07,1.922477e-07,1.922479e-07,1.922481e-07,1.922483e-07,1.922486e-07,1.922488e-07,1.922490e-07,1.922493e-07,1.922495e-07,1.922497e-07,1.922499e-07,1.922502e-07,1.922504e-07,1.922506e-07,1.922508e-07,1.922511e-07,1.922513e-07,1.922515e-07,1.922517e-07,1.922520e-07,1.922522e-07,1.922524e-07,1.922526e-07,1.922529e-07,1.922531e-07,1.922533e-07,1.922536e-07,1.922538e-07,1.922540e-07,1.922542e-07,1.922545e-07,1.922547e-07,1.922549e-07,1.922551e-07,1.922554e-07,1.922556e-07,1.922558e-07,1.922560e-07,1.922563e-07,1.922565e-07,1.922567e-07,1.922569e-07,1.922572e-07,1.922574e-07,1.922576e-07,1.922579e-07,1.922581e-07,1.922583e-07,1.922585e-07,1.922588e-07,1.922590e-07,1.922592e-07,1.922594e-07,1.922597e-07,1.922599e-07,1.922601e-07,1.922603e-07,1.922606e-07,1.922608e-07,1.922610e-07,1.922612e-07,1.922615e-07,1.922617e-07,1.922619e-07,1.922622e-07,1.922624e-07,1.922626e-07,1.922628e-07,1.922631e-07,1.922633e-07,1.922635e-07,1.922637e-07,1.922640e-07,1.922642e-07,1.922644e-07,1.922646e-07,1.922649e-07,1.922651e-07,1.922653e-07,1.922655e-07,1.922658e-07,1.922660e-07,1.922662e-07,1.922665e-07,1.922667e-07,1.922669e-07,1.922671e-07,1.922674e-07,1.922676e-07,1.922678e-07,1.922680e-07,1.922683e-07,1.922685e-07,1.922687e-07,1.922689e-07,1.922692e-07,1.922694e-07,1.922696e-07,1.922698e-07,1.922701e-07,1.922703e-07,1.922705e-07,1.922707e-07,1.922710e-07,1.922712e-07,1.922714e-07,1.922717e-07,1.922719e-07,1.922721e-07,1.922723e-07,1.922726e-07,1.922728e-07,1.922730e-07,1.922732e-07,1.922735e-07,1.922737e-07,1.922739e-07,1.922741e-07,1.922744e-07,1.922746e-07,1.922748e-07,1.922750e-07,1.922753e-07,1.922755e-07,1.922757e-07,1.922759e-07,1.922762e-07,1.922764e-07,1.922766e-07,1.922768e-07,1.922771e-07,1.922773e-07,1.922775e-07,1.922778e-07,1.922780e-07,1.922782e-07,1.922784e-07,1.922787e-07,1.922789e-07,1.922791e-07,1.922793e-07,1.922796e-07,1.922798e-07,1.922800e-07,1.922802e-07,1.922805e-07,1.922807e-07,1.922809e-07,1.922811e-07,1.922814e-07,1.922816e-07,1.922818e-07,1.922820e-07,1.922823e-07,1.922825e-07,1.922827e-07,1.922829e-07,1.922832e-07,1.922834e-07,1.922836e-07,1.922839e-07,1.922841e-07,1.922843e-07,1.922845e-07,1.922848e-07,1.922850e-07,1.922852e-07,1.922854e-07,1.922857e-07,1.922859e-07,1.922861e-07,1.922863e-07,1.922866e-07,1.922868e-07,1.922870e-07,1.922872e-07,1.922875e-07,1.922877e-07,1.922879e-07,1.922881e-07,1.922884e-07,1.922886e-07,1.922888e-07,1.922890e-07,1.922893e-07,1.922895e-07,1.922897e-07,1.922899e-07,1.922902e-07,1.922904e-07,1.922906e-07,1.922908e-07,1.922911e-07,1.922913e-07,1.922915e-07,1.922918e-07,1.922920e-07,1.922922e-07,1.922924e-07,1.922927e-07,1.922929e-07,1.922931e-07,1.922933e-07,1.922936e-07,1.922938e-07,1.922940e-07,1.922942e-07,1.922945e-07,1.922947e-07,1.922949e-07,1.922951e-07,1.922954e-07,1.922956e-07,1.922958e-07,1.922960e-07,1.922963e-07,1.922965e-07,1.922967e-07,1.922969e-07,1.922972e-07,1.922974e-07,1.922976e-07,1.922978e-07,1.922981e-07,1.922983e-07,1.922985e-07,1.922987e-07,1.922990e-07,1.922992e-07,1.922994e-07,1.922996e-07,1.922999e-07,1.923001e-07,1.923003e-07,1.923005e-07,1.923008e-07,1.923010e-07,1.923012e-07,1.923014e-07,1.923017e-07,1.923019e-07,1.923021e-07,1.923024e-07,1.923026e-07,1.923028e-07,1.923030e-07,1.923033e-07,1.923035e-07,1.923037e-07,1.923039e-07,1.923042e-07,1.923044e-07,1.923046e-07,1.923048e-07,1.923051e-07,1.923053e-07,1.923055e-07,1.923057e-07,1.923060e-07,1.923062e-07,1.923064e-07,1.923066e-07,1.923069e-07,1.923071e-07,1.923073e-07,1.923075e-07,1.923078e-07,1.923080e-07,1.923082e-07,1.923084e-07,1.923087e-07,1.923089e-07,1.923091e-07,1.923093e-07,1.923096e-07,1.923098e-07,1.923100e-07,1.923102e-07,1.923105e-07,1.923107e-07,1.923109e-07,1.923111e-07,1.923114e-07,1.923116e-07,1.923118e-07,1.923120e-07,1.923123e-07,1.923125e-07,1.923127e-07,1.923129e-07,1.923132e-07,1.923134e-07,1.923136e-07,1.923138e-07,1.923141e-07,1.923143e-07,1.923145e-07,1.923147e-07,1.923150e-07,1.923152e-07,1.923154e-07,1.923156e-07,1.923159e-07,1.923161e-07,1.923163e-07,1.923165e-07,1.923168e-07,1.923170e-07,1.923172e-07,1.923174e-07,1.923177e-07,1.923179e-07,1.923181e-07,1.923183e-07,1.923186e-07,1.923188e-07,1.923190e-07,1.923192e-07,1.923195e-07,1.923197e-07,1.923199e-07,1.923201e-07,1.923204e-07,1.923206e-07,1.923208e-07,1.923210e-07,1.923213e-07,1.923215e-07,1.923217e-07,1.923219e-07,1.923222e-07,1.923224e-07,1.923226e-07,1.923228e-07,1.923231e-07,1.923233e-07,1.923235e-07,1.923237e-07,1.923240e-07,1.923242e-07,1.923244e-07,1.923246e-07,1.923249e-07,1.923251e-07,1.923253e-07,1.923255e-07,1.923258e-07,1.923260e-07,1.923262e-07,1.923264e-07,1.923267e-07,1.923269e-07,1.923271e-07,1.923273e-07,1.923276e-07,1.923278e-07,1.923280e-07,1.923282e-07,1.923285e-07,1.923287e-07,1.923289e-07,1.923291e-07,1.923294e-07,1.923296e-07,1.923298e-07,1.923300e-07,1.923303e-07,1.923305e-07,1.923307e-07,1.923309e-07,1.923312e-07,1.923314e-07,1.923316e-07,1.923318e-07,1.923321e-07,1.923323e-07,1.923325e-07,1.923327e-07,1.923330e-07,1.923332e-07,1.923334e-07,1.923336e-07,1.923339e-07,1.923341e-07,1.923343e-07,1.923345e-07,1.923348e-07,1.923350e-07,1.923352e-07,1.923354e-07,1.923357e-07,1.923359e-07,1.923361e-07,1.923363e-07,1.923366e-07,1.923368e-07,1.923370e-07,1.923372e-07,1.923375e-07,1.923377e-07,1.923379e-07,1.923381e-07,1.923384e-07,1.923386e-07,1.923388e-07,1.923390e-07,1.923393e-07,1.923395e-07,1.923397e-07,1.923399e-07,1.923402e-07,1.923404e-07,1.923406e-07,1.923408e-07,1.923411e-07,1.923413e-07,1.923415e-07,1.923417e-07,1.923420e-07,1.923422e-07,1.923424e-07,1.923426e-07,1.923429e-07,1.923431e-07,1.923433e-07,1.923435e-07,1.923438e-07,1.923440e-07,1.923442e-07,1.923444e-07,1.923447e-07,1.923449e-07,1.923451e-07,1.923453e-07,1.923456e-07,1.923458e-07,1.923460e-07,1.923462e-07,1.923465e-07,1.923467e-07,1.923469e-07,1.923471e-07,1.923474e-07,1.923476e-07,1.923478e-07,1.923480e-07,1.923483e-07,1.923485e-07,1.923487e-07,1.923489e-07,1.923491e-07,1.923494e-07,1.923496e-07,1.923498e-07,1.923500e-07,1.923503e-07,1.923505e-07,1.923507e-07,1.923509e-07,1.923512e-07,1.923514e-07,1.923516e-07,1.923518e-07,1.923521e-07,1.923523e-07,1.923525e-07,1.923527e-07,1.923530e-07,1.923532e-07,1.923534e-07,1.923536e-07,1.923539e-07,1.923541e-07,1.923543e-07,1.923545e-07,1.923548e-07,1.923550e-07,1.923552e-07,1.923554e-07,1.923557e-07,1.923559e-07,1.923561e-07,1.923563e-07,1.923566e-07,1.923568e-07,1.923570e-07,1.923572e-07,1.923575e-07,1.923577e-07,1.923579e-07,1.923581e-07,1.923584e-07,1.923586e-07,1.923588e-07,1.923590e-07,1.923592e-07,1.923595e-07,1.923597e-07,1.923599e-07,1.923601e-07,1.923604e-07,1.923606e-07,1.923608e-07,1.923610e-07,1.923613e-07,1.923615e-07,1.923617e-07,1.923619e-07,1.923622e-07,1.923624e-07,1.923626e-07,1.923628e-07,1.923631e-07,1.923633e-07,1.923635e-07,1.923637e-07,1.923640e-07,1.923642e-07,1.923644e-07,1.923646e-07,1.923649e-07,1.923651e-07,1.923653e-07,1.923655e-07,1.923658e-07,1.923660e-07,1.923662e-07,1.923664e-07,1.923666e-07,1.923669e-07,1.923671e-07,1.923673e-07,1.923675e-07,1.923678e-07,1.923680e-07,1.923682e-07,1.923684e-07,1.923687e-07,1.923689e-07,1.923691e-07,1.923693e-07,1.923696e-07,1.923698e-07,1.923700e-07,1.923702e-07,1.923705e-07,1.923707e-07,1.923709e-07,1.923711e-07,1.923714e-07,1.923716e-07,1.923718e-07,1.923720e-07,1.923723e-07,1.923725e-07,1.923727e-07,1.923729e-07,1.923731e-07,1.923734e-07,1.923736e-07,1.923738e-07,1.923740e-07,1.923743e-07,1.923745e-07,1.923747e-07,1.923749e-07,1.923752e-07,1.923754e-07,1.923756e-07,1.923758e-07,1.923761e-07,1.923763e-07,1.923765e-07,1.923767e-07,1.923770e-07,1.923772e-07,1.923774e-07,1.923776e-07,1.923779e-07,1.923781e-07,1.923783e-07,1.923785e-07,1.923788e-07,1.923790e-07,1.923792e-07,1.923794e-07,1.923796e-07,1.923799e-07,1.923801e-07,1.923803e-07,1.923805e-07,1.923808e-07,1.923810e-07,1.923812e-07,1.923814e-07,1.923817e-07,1.923819e-07,1.923821e-07,1.923823e-07,1.923826e-07,1.923828e-07,1.923830e-07,1.923832e-07,1.923835e-07,1.923837e-07,1.923839e-07,1.923841e-07,1.923843e-07,1.923846e-07,1.923848e-07,1.923850e-07,1.923852e-07,1.923855e-07,1.923857e-07,1.923859e-07,1.923861e-07,1.923864e-07,1.923866e-07,1.923868e-07,1.923870e-07,1.923873e-07,1.923875e-07,1.923877e-07,1.923879e-07,1.923882e-07,1.923884e-07,1.923886e-07,1.923888e-07,1.923890e-07,1.923893e-07,1.923895e-07,1.923897e-07,1.923899e-07,1.923902e-07,1.923904e-07,1.923906e-07,1.923908e-07,1.923911e-07,1.923913e-07,1.923915e-07,1.923917e-07,1.923920e-07,1.923922e-07,1.923924e-07,1.923926e-07,1.923929e-07,1.923931e-07,1.923933e-07,1.923935e-07,1.923937e-07,1.923940e-07,1.923942e-07,1.923944e-07,1.923946e-07,1.923949e-07,1.923951e-07,1.923953e-07,1.923955e-07,1.923958e-07,1.923960e-07,1.923962e-07,1.923964e-07,1.923967e-07,1.923969e-07,1.923971e-07,1.923973e-07,1.923975e-07,1.923978e-07,1.923980e-07,1.923982e-07,1.923984e-07,1.923987e-07,1.923989e-07,1.923991e-07,1.923993e-07,1.923996e-07,1.923998e-07,1.924000e-07,1.924002e-07,1.924005e-07,1.924007e-07,1.924009e-07,1.924011e-07,1.924013e-07,1.924016e-07,1.924018e-07,1.924020e-07,1.924022e-07,1.924025e-07,1.924027e-07,1.924029e-07,1.924031e-07,1.924034e-07,1.924036e-07,1.924038e-07,1.924040e-07,1.924043e-07,1.924045e-07,1.924047e-07,1.924049e-07,1.924051e-07,1.924054e-07,1.924056e-07,1.924058e-07,1.924060e-07,1.924063e-07,1.924065e-07,1.924067e-07,1.924069e-07,1.924072e-07,1.924074e-07,1.924076e-07,1.924078e-07,1.924081e-07,1.924083e-07,1.924085e-07,1.924087e-07,1.924089e-07,1.924092e-07,1.924094e-07,1.924096e-07,1.924098e-07,1.924101e-07,1.924103e-07,1.924105e-07,1.924107e-07,1.924110e-07,1.924112e-07,1.924114e-07,1.924116e-07,1.924119e-07,1.924121e-07,1.924123e-07,1.924125e-07,1.924127e-07,1.924130e-07,1.924132e-07,1.924134e-07,1.924136e-07,1.924139e-07,1.924141e-07,1.924143e-07,1.924145e-07,1.924148e-07,1.924150e-07,1.924152e-07,1.924154e-07,1.924156e-07,1.924159e-07,1.924161e-07,1.924163e-07,1.924165e-07,1.924168e-07,1.924170e-07,1.924172e-07,1.924174e-07,1.924177e-07,1.924179e-07,1.924181e-07,1.924183e-07,1.924185e-07,1.924188e-07,1.924190e-07,1.924192e-07,1.924194e-07,1.924197e-07,1.924199e-07,1.924201e-07,1.924203e-07,1.924206e-07,1.924208e-07,1.924210e-07,1.924212e-07,1.924215e-07,1.924217e-07,1.924219e-07,1.924221e-07,1.924223e-07,1.924226e-07,1.924228e-07,1.924230e-07,1.924232e-07,1.924235e-07,1.924237e-07,1.924239e-07,1.924241e-07,1.924244e-07,1.924246e-07,1.924248e-07,1.924250e-07,1.924252e-07,1.924255e-07,1.924257e-07,1.924259e-07,1.924261e-07,1.924264e-07,1.924266e-07,1.924268e-07,1.924270e-07,1.924273e-07,1.924275e-07,1.924277e-07,1.924279e-07,1.924281e-07,1.924284e-07,1.924286e-07,1.924288e-07,1.924290e-07,1.924293e-07,1.924295e-07,1.924297e-07,1.924299e-07,1.924302e-07,1.924304e-07,1.924306e-07,1.924308e-07,1.924310e-07,1.924313e-07,1.924315e-07,1.924317e-07,1.924319e-07,1.924322e-07,1.924324e-07,1.924326e-07,1.924328e-07,1.924330e-07,1.924333e-07,1.924335e-07,1.924337e-07,1.924339e-07,1.924342e-07,1.924344e-07,1.924346e-07,1.924348e-07,1.924351e-07,1.924353e-07,1.924355e-07,1.924357e-07,1.924359e-07,1.924362e-07,1.924364e-07,1.924366e-07,1.924368e-07,1.924371e-07,1.924373e-07,1.924375e-07,1.924377e-07,1.924380e-07,1.924382e-07,1.924384e-07,1.924386e-07,1.924388e-07,1.924391e-07,1.924393e-07,1.924395e-07,1.924397e-07,1.924400e-07,1.924402e-07,1.924404e-07,1.924406e-07,1.924408e-07,1.924411e-07,1.924413e-07,1.924415e-07,1.924417e-07,1.924420e-07,1.924422e-07,1.924424e-07,1.924426e-07,1.924429e-07,1.924431e-07,1.924433e-07,1.924435e-07,1.924437e-07,1.924440e-07,1.924442e-07,1.924444e-07,1.924446e-07,1.924449e-07,1.924451e-07,1.924453e-07,1.924455e-07,1.924457e-07,1.924460e-07,1.924462e-07,1.924464e-07,1.924466e-07,1.924469e-07,1.924471e-07,1.924473e-07,1.924475e-07,1.924478e-07,1.924480e-07,1.924482e-07,1.924484e-07,1.924486e-07,1.924489e-07,1.924491e-07,1.924493e-07,1.924495e-07,1.924498e-07,1.924500e-07,1.924502e-07,1.924504e-07,1.924506e-07,1.924509e-07,1.924511e-07,1.924513e-07,1.924515e-07,1.924518e-07,1.924520e-07,1.924522e-07,1.924524e-07,1.924527e-07,1.924529e-07,1.924531e-07,1.924533e-07,1.924535e-07,1.924538e-07,1.924540e-07,1.924542e-07,1.924544e-07,1.924547e-07,1.924549e-07,1.924551e-07,1.924553e-07,1.924555e-07,1.924558e-07,1.924560e-07,1.924562e-07,1.924564e-07,1.924567e-07,1.924569e-07,1.924571e-07,1.924573e-07,1.924575e-07,1.924578e-07,1.924580e-07,1.924582e-07,1.924584e-07,1.924587e-07,1.924589e-07,1.924591e-07,1.924593e-07,1.924595e-07,1.924598e-07,1.924600e-07,1.924602e-07,1.924604e-07,1.924607e-07,1.924609e-07,1.924611e-07,1.924613e-07,1.924615e-07,1.924618e-07,1.924620e-07,1.924622e-07,1.924624e-07,1.924627e-07,1.924629e-07,1.924631e-07,1.924633e-07,1.924636e-07,1.924638e-07,1.924640e-07,1.924642e-07,1.924644e-07,1.924647e-07,1.924649e-07,1.924651e-07,1.924653e-07,1.924656e-07,1.924658e-07,1.924660e-07,1.924662e-07,1.924664e-07,1.924667e-07,1.924669e-07,1.924671e-07,1.924673e-07,1.924676e-07,1.924678e-07,1.924680e-07,1.924682e-07,1.924684e-07,1.924687e-07,1.924689e-07,1.924691e-07,1.924693e-07,1.924696e-07,1.924698e-07,1.924700e-07,1.924702e-07,1.924704e-07,1.924707e-07,1.924709e-07,1.924711e-07,1.924713e-07,1.924716e-07,1.924718e-07,1.924720e-07,1.924722e-07,1.924724e-07,1.924727e-07,1.924729e-07,1.924731e-07,1.924733e-07,1.924736e-07,1.924738e-07,1.924740e-07,1.924742e-07,1.924744e-07,1.924747e-07,1.924749e-07,1.924751e-07,1.924753e-07,1.924756e-07,1.924758e-07,1.924760e-07,1.924762e-07,1.924764e-07,1.924767e-07,1.924769e-07,1.924771e-07,1.924773e-07,1.924776e-07,1.924778e-07,1.924780e-07,1.924782e-07,1.924784e-07,1.924787e-07,1.924789e-07,1.924791e-07,1.924793e-07,1.924795e-07,1.924798e-07,1.924800e-07,1.924802e-07,1.924804e-07,1.924807e-07,1.924809e-07,1.924811e-07,1.924813e-07,1.924815e-07,1.924818e-07,1.924820e-07,1.924822e-07,1.924824e-07,1.924827e-07,1.924829e-07,1.924831e-07,1.924833e-07,1.924835e-07,1.924838e-07,1.924840e-07,1.924842e-07,1.924844e-07,1.924847e-07,1.924849e-07,1.924851e-07,1.924853e-07,1.924855e-07,1.924858e-07,1.924860e-07,1.924862e-07,1.924864e-07,1.924867e-07,1.924869e-07,1.924871e-07,1.924873e-07,1.924875e-07,1.924878e-07,1.924880e-07,1.924882e-07,1.924884e-07,1.924886e-07,1.924889e-07,1.924891e-07,1.924893e-07,1.924895e-07,1.924898e-07,1.924900e-07,1.924902e-07,1.924904e-07,1.924906e-07,1.924909e-07,1.924911e-07,1.924913e-07,1.924915e-07,1.924918e-07,1.924920e-07,1.924922e-07,1.924924e-07,1.924926e-07,1.924929e-07,1.924931e-07,1.924933e-07,1.924935e-07,1.924938e-07,1.924940e-07,1.924942e-07,1.924944e-07,1.924946e-07,1.924949e-07,1.924951e-07,1.924953e-07,1.924955e-07,1.924957e-07,1.924960e-07,1.924962e-07,1.924964e-07,1.924966e-07,1.924969e-07,1.924971e-07,1.924973e-07,1.924975e-07,1.924977e-07,1.924980e-07,1.924982e-07,1.924984e-07,1.924986e-07,1.924989e-07,1.924991e-07,1.924993e-07,1.924995e-07,1.924997e-07,1.925000e-07,1.925002e-07,1.925004e-07,1.925006e-07,1.925008e-07,1.925011e-07,1.925013e-07,1.925015e-07,1.925017e-07,1.925020e-07,1.925022e-07,1.925024e-07,1.925026e-07,1.925028e-07,1.925031e-07,1.925033e-07,1.925035e-07,1.925037e-07,1.925039e-07,1.925042e-07,1.925044e-07,1.925046e-07,1.925048e-07,1.925051e-07,1.925053e-07,1.925055e-07,1.925057e-07,1.925059e-07,1.925062e-07,1.925064e-07,1.925066e-07,1.925068e-07,1.925071e-07,1.925073e-07,1.925075e-07,1.925077e-07,1.925079e-07,1.925082e-07,1.925084e-07,1.925086e-07,1.925088e-07,1.925090e-07,1.925093e-07,1.925095e-07,1.925097e-07,1.925099e-07,1.925102e-07,1.925104e-07,1.925106e-07,1.925108e-07,1.925110e-07,1.925113e-07,1.925115e-07,1.925117e-07,1.925119e-07,1.925121e-07,1.925124e-07,1.925126e-07,1.925128e-07,1.925130e-07,1.925133e-07,1.925135e-07,1.925137e-07,1.925139e-07,1.925141e-07,1.925144e-07,1.925146e-07,1.925148e-07,1.925150e-07,1.925152e-07,1.925155e-07,1.925157e-07,1.925159e-07,1.925161e-07,1.925164e-07,1.925166e-07,1.925168e-07,1.925170e-07,1.925172e-07,1.925175e-07,1.925177e-07,1.925179e-07,1.925181e-07,1.925183e-07,1.925186e-07,1.925188e-07,1.925190e-07,1.925192e-07,1.925195e-07,1.925197e-07,1.925199e-07,1.925201e-07,1.925203e-07,1.925206e-07,1.925208e-07,1.925210e-07,1.925212e-07,1.925214e-07,1.925217e-07,1.925219e-07,1.925221e-07,1.925223e-07,1.925225e-07,1.925228e-07,1.925230e-07,1.925232e-07,1.925234e-07,1.925237e-07,1.925239e-07,1.925241e-07,1.925243e-07,1.925245e-07,1.925248e-07,1.925250e-07,1.925252e-07,1.925254e-07,1.925256e-07,1.925259e-07,1.925261e-07,1.925263e-07,1.925265e-07,1.925268e-07,1.925270e-07,1.925272e-07,1.925274e-07,1.925276e-07,1.925279e-07,1.925281e-07,1.925283e-07,1.925285e-07,1.925287e-07,1.925290e-07,1.925292e-07,1.925294e-07,1.925296e-07,1.925298e-07,1.925301e-07,1.925303e-07,1.925305e-07,1.925307e-07,1.925310e-07,1.925312e-07,1.925314e-07,1.925316e-07,1.925318e-07,1.925321e-07,1.925323e-07,1.925325e-07,1.925327e-07,1.925329e-07,1.925332e-07,1.925334e-07,1.925336e-07,1.925338e-07,1.925340e-07,1.925343e-07,1.925345e-07,1.925347e-07,1.925349e-07,1.925352e-07,1.925354e-07,1.925356e-07,1.925358e-07,1.925360e-07,1.925363e-07,1.925365e-07,1.925367e-07,1.925369e-07,1.925371e-07,1.925374e-07,1.925376e-07,1.925378e-07,1.925380e-07,1.925382e-07,1.925385e-07,1.925387e-07,1.925389e-07,1.925391e-07,1.925393e-07,1.925396e-07,1.925398e-07,1.925400e-07,1.925402e-07,1.925405e-07,1.925407e-07,1.925409e-07,1.925411e-07,1.925413e-07,1.925416e-07,1.925418e-07,1.925420e-07,1.925422e-07,1.925424e-07,1.925427e-07,1.925429e-07,1.925431e-07,1.925433e-07,1.925435e-07,1.925438e-07,1.925440e-07,1.925442e-07,1.925444e-07,1.925447e-07,1.925449e-07,1.925451e-07,1.925453e-07,1.925455e-07,1.925458e-07,1.925460e-07,1.925462e-07,1.925464e-07,1.925466e-07,1.925469e-07,1.925471e-07,1.925473e-07,1.925475e-07,1.925477e-07,1.925480e-07,1.925482e-07,1.925484e-07,1.925486e-07,1.925488e-07,1.925491e-07,1.925493e-07,1.925495e-07,1.925497e-07,1.925499e-07,1.925502e-07,1.925504e-07,1.925506e-07,1.925508e-07,1.925511e-07,1.925513e-07,1.925515e-07,1.925517e-07,1.925519e-07,1.925522e-07,1.925524e-07,1.925526e-07,1.925528e-07,1.925530e-07,1.925533e-07,1.925535e-07,1.925537e-07,1.925539e-07,1.925541e-07,1.925544e-07,1.925546e-07,1.925548e-07,1.925550e-07,1.925552e-07,1.925555e-07,1.925557e-07,1.925559e-07,1.925561e-07,1.925563e-07,1.925566e-07,1.925568e-07,1.925570e-07,1.925572e-07,1.925575e-07,1.925577e-07,1.925579e-07,1.925581e-07,1.925583e-07,1.925586e-07,1.925588e-07,1.925590e-07,1.925592e-07,1.925594e-07,1.925597e-07,1.925599e-07,1.925601e-07,1.925603e-07,1.925605e-07,1.925608e-07,1.925610e-07,1.925612e-07,1.925614e-07,1.925616e-07,1.925619e-07,1.925621e-07,1.925623e-07,1.925625e-07,1.925627e-07,1.925630e-07,1.925632e-07,1.925634e-07,1.925636e-07,1.925638e-07,1.925641e-07,1.925643e-07,1.925645e-07,1.925647e-07,1.925649e-07,1.925652e-07,1.925654e-07,1.925656e-07,1.925658e-07,1.925661e-07,1.925663e-07,1.925665e-07,1.925667e-07,1.925669e-07,1.925672e-07,1.925674e-07,1.925676e-07,1.925678e-07,1.925680e-07,1.925683e-07,1.925685e-07,1.925687e-07,1.925689e-07,1.925691e-07,1.925694e-07,1.925696e-07,1.925698e-07,1.925700e-07,1.925702e-07,1.925705e-07,1.925707e-07,1.925709e-07,1.925711e-07,1.925713e-07,1.925716e-07,1.925718e-07,1.925720e-07,1.925722e-07,1.925724e-07,1.925727e-07,1.925729e-07,1.925731e-07,1.925733e-07,1.925735e-07,1.925738e-07,1.925740e-07,1.925742e-07,1.925744e-07,1.925746e-07,1.925749e-07,1.925751e-07,1.925753e-07,1.925755e-07,1.925757e-07,1.925760e-07,1.925762e-07,1.925764e-07,1.925766e-07,1.925768e-07,1.925771e-07,1.925773e-07,1.925775e-07,1.925777e-07,1.925779e-07,1.925782e-07,1.925784e-07,1.925786e-07,1.925788e-07,1.925790e-07,1.925793e-07,1.925795e-07,1.925797e-07,1.925799e-07,1.925801e-07,1.925804e-07,1.925806e-07,1.925808e-07,1.925810e-07,1.925812e-07,1.925815e-07,1.925817e-07,1.925819e-07,1.925821e-07,1.925823e-07,1.925826e-07,1.925828e-07,1.925830e-07,1.925832e-07,1.925835e-07,1.925837e-07,1.925839e-07,1.925841e-07,1.925843e-07,1.925846e-07,1.925848e-07,1.925850e-07,1.925852e-07,1.925854e-07,1.925857e-07,1.925859e-07,1.925861e-07,1.925863e-07,1.925865e-07,1.925868e-07,1.925870e-07,1.925872e-07,1.925874e-07,1.925876e-07,1.925879e-07,1.925881e-07,1.925883e-07,1.925885e-07,1.925887e-07,1.925890e-07,1.925892e-07,1.925894e-07,1.925896e-07,1.925898e-07,1.925901e-07,1.925903e-07,1.925905e-07,1.925907e-07,1.925909e-07,1.925912e-07,1.925914e-07,1.925916e-07,1.925918e-07,1.925920e-07,1.925923e-07,1.925925e-07,1.925927e-07,1.925929e-07,1.925931e-07,1.925933e-07,1.925936e-07,1.925938e-07,1.925940e-07,1.925942e-07,1.925944e-07,1.925947e-07,1.925949e-07,1.925951e-07,1.925953e-07,1.925955e-07,1.925958e-07,1.925960e-07,1.925962e-07,1.925964e-07,1.925966e-07,1.925969e-07,1.925971e-07,1.925973e-07,1.925975e-07,1.925977e-07,1.925980e-07,1.925982e-07,1.925984e-07,1.925986e-07,1.925988e-07,1.925991e-07,1.925993e-07,1.925995e-07,1.925997e-07,1.925999e-07,1.926002e-07,1.926004e-07,1.926006e-07,1.926008e-07,1.926010e-07,1.926013e-07,1.926015e-07,1.926017e-07,1.926019e-07,1.926021e-07,1.926024e-07,1.926026e-07,1.926028e-07,1.926030e-07,1.926032e-07,1.926035e-07,1.926037e-07,1.926039e-07,1.926041e-07,1.926043e-07,1.926046e-07,1.926048e-07,1.926050e-07,1.926052e-07,1.926054e-07,1.926057e-07,1.926059e-07,1.926061e-07,1.926063e-07,1.926065e-07,1.926068e-07,1.926070e-07,1.926072e-07,1.926074e-07,1.926076e-07,1.926079e-07,1.926081e-07,1.926083e-07,1.926085e-07,1.926087e-07,1.926090e-07,1.926092e-07,1.926094e-07,1.926096e-07,1.926098e-07,1.926101e-07,1.926103e-07,1.926105e-07,1.926107e-07,1.926109e-07,1.926111e-07,1.926114e-07,1.926116e-07,1.926118e-07,1.926120e-07,1.926122e-07,1.926125e-07,1.926127e-07,1.926129e-07,1.926131e-07,1.926133e-07,1.926136e-07,1.926138e-07,1.926140e-07,1.926142e-07,1.926144e-07,1.926147e-07,1.926149e-07,1.926151e-07,1.926153e-07,1.926155e-07,1.926158e-07,1.926160e-07,1.926162e-07,1.926164e-07,1.926166e-07,1.926169e-07,1.926171e-07,1.926173e-07,1.926175e-07,1.926177e-07,1.926180e-07,1.926182e-07,1.926184e-07,1.926186e-07,1.926188e-07,1.926190e-07,1.926193e-07,1.926195e-07,1.926197e-07,1.926199e-07,1.926201e-07,1.926204e-07,1.926206e-07,1.926208e-07,1.926210e-07,1.926212e-07,1.926215e-07,1.926217e-07,1.926219e-07,1.926221e-07,1.926223e-07,1.926226e-07,1.926228e-07,1.926230e-07,1.926232e-07,1.926234e-07,1.926237e-07,1.926239e-07,1.926241e-07,1.926243e-07,1.926245e-07,1.926248e-07,1.926250e-07,1.926252e-07,1.926254e-07,1.926256e-07,1.926258e-07,1.926261e-07,1.926263e-07,1.926265e-07,1.926267e-07,1.926269e-07,1.926272e-07,1.926274e-07,1.926276e-07,1.926278e-07,1.926280e-07,1.926283e-07,1.926285e-07,1.926287e-07,1.926289e-07,1.926291e-07,1.926294e-07,1.926296e-07,1.926298e-07,1.926300e-07,1.926302e-07,1.926305e-07,1.926307e-07,1.926309e-07,1.926311e-07,1.926313e-07,1.926315e-07,1.926318e-07,1.926320e-07,1.926322e-07,1.926324e-07,1.926326e-07,1.926329e-07,1.926331e-07,1.926333e-07,1.926335e-07,1.926337e-07,1.926340e-07,1.926342e-07,1.926344e-07,1.926346e-07,1.926348e-07,1.926351e-07,1.926353e-07,1.926355e-07,1.926357e-07,1.926359e-07,1.926362e-07,1.926364e-07,1.926366e-07,1.926368e-07,1.926370e-07,1.926372e-07,1.926375e-07,1.926377e-07,1.926379e-07,1.926381e-07,1.926383e-07,1.926386e-07,1.926388e-07,1.926390e-07,1.926392e-07,1.926394e-07,1.926397e-07,1.926399e-07,1.926401e-07,1.926403e-07,1.926405e-07,1.926408e-07,1.926410e-07,1.926412e-07,1.926414e-07,1.926416e-07,1.926418e-07,1.926421e-07,1.926423e-07,1.926425e-07,1.926427e-07,1.926429e-07,1.926432e-07,1.926434e-07,1.926436e-07,1.926438e-07,1.926440e-07,1.926443e-07,1.926445e-07,1.926447e-07,1.926449e-07,1.926451e-07,1.926454e-07,1.926456e-07,1.926458e-07,1.926460e-07,1.926462e-07,1.926464e-07,1.926467e-07,1.926469e-07,1.926471e-07,1.926473e-07,1.926475e-07,1.926478e-07,1.926480e-07,1.926482e-07,1.926484e-07,1.926486e-07,1.926489e-07,1.926491e-07,1.926493e-07,1.926495e-07,1.926497e-07,1.926499e-07,1.926502e-07,1.926504e-07,1.926506e-07,1.926508e-07,1.926510e-07,1.926513e-07,1.926515e-07,1.926517e-07,1.926519e-07,1.926521e-07,1.926524e-07,1.926526e-07,1.926528e-07,1.926530e-07,1.926532e-07,1.926534e-07,1.926537e-07,1.926539e-07,1.926541e-07,1.926543e-07,1.926545e-07,1.926548e-07,1.926550e-07,1.926552e-07,1.926554e-07,1.926556e-07,1.926559e-07,1.926561e-07,1.926563e-07,1.926565e-07,1.926567e-07,1.926569e-07,1.926572e-07,1.926574e-07,1.926576e-07,1.926578e-07,1.926580e-07,1.926583e-07,1.926585e-07,1.926587e-07,1.926589e-07,1.926591e-07,1.926594e-07,1.926596e-07,1.926598e-07,1.926600e-07,1.926602e-07,1.926604e-07,1.926607e-07,1.926609e-07,1.926611e-07,1.926613e-07,1.926615e-07,1.926618e-07,1.926620e-07,1.926622e-07,1.926624e-07,1.926626e-07,1.926629e-07,1.926631e-07,1.926633e-07,1.926635e-07,1.926637e-07,1.926639e-07,1.926642e-07,1.926644e-07,1.926646e-07,1.926648e-07,1.926650e-07,1.926653e-07,1.926655e-07,1.926657e-07,1.926659e-07,1.926661e-07,1.926663e-07,1.926666e-07,1.926668e-07,1.926670e-07,1.926672e-07,1.926674e-07,1.926677e-07,1.926679e-07,1.926681e-07,1.926683e-07,1.926685e-07,1.926688e-07,1.926690e-07,1.926692e-07,1.926694e-07,1.926696e-07,1.926698e-07,1.926701e-07,1.926703e-07,1.926705e-07,1.926707e-07,1.926709e-07,1.926712e-07,1.926714e-07,1.926716e-07,1.926718e-07,1.926720e-07,1.926722e-07,1.926725e-07,1.926727e-07,1.926729e-07,1.926731e-07,1.926733e-07,1.926736e-07,1.926738e-07,1.926740e-07,1.926742e-07,1.926744e-07,1.926746e-07,1.926749e-07,1.926751e-07,1.926753e-07,1.926755e-07,1.926757e-07,1.926760e-07,1.926762e-07,1.926764e-07,1.926766e-07,1.926768e-07,1.926771e-07,1.926773e-07,1.926775e-07,1.926777e-07,1.926779e-07,1.926781e-07,1.926784e-07,1.926786e-07,1.926788e-07,1.926790e-07,1.926792e-07,1.926795e-07,1.926797e-07,1.926799e-07,1.926801e-07,1.926803e-07,1.926805e-07,1.926808e-07,1.926810e-07,1.926812e-07,1.926814e-07,1.926816e-07,1.926819e-07,1.926821e-07,1.926823e-07,1.926825e-07,1.926827e-07,1.926829e-07,1.926832e-07,1.926834e-07,1.926836e-07,1.926838e-07,1.926840e-07,1.926843e-07,1.926845e-07,1.926847e-07,1.926849e-07,1.926851e-07,1.926853e-07,1.926856e-07,1.926858e-07,1.926860e-07,1.926862e-07,1.926864e-07,1.926867e-07,1.926869e-07,1.926871e-07,1.926873e-07,1.926875e-07,1.926877e-07,1.926880e-07,1.926882e-07,1.926884e-07,1.926886e-07,1.926888e-07,1.926891e-07,1.926893e-07,1.926895e-07,1.926897e-07,1.926899e-07,1.926901e-07,1.926904e-07,1.926906e-07,1.926908e-07,1.926910e-07,1.926912e-07,1.926915e-07,1.926917e-07,1.926919e-07,1.926921e-07,1.926923e-07,1.926925e-07,1.926928e-07,1.926930e-07,1.926932e-07,1.926934e-07,1.926936e-07,1.926939e-07,1.926941e-07,1.926943e-07,1.926945e-07,1.926947e-07,1.926949e-07,1.926952e-07,1.926954e-07,1.926956e-07,1.926958e-07,1.926960e-07,1.926962e-07,1.926965e-07,1.926967e-07,1.926969e-07,1.926971e-07,1.926973e-07,1.926976e-07,1.926978e-07,1.926980e-07,1.926982e-07,1.926984e-07,1.926986e-07,1.926989e-07,1.926991e-07,1.926993e-07,1.926995e-07,1.926997e-07,1.927000e-07,1.927002e-07,1.927004e-07,1.927006e-07,1.927008e-07,1.927010e-07,1.927013e-07,1.927015e-07,1.927017e-07,1.927019e-07,1.927021e-07,1.927024e-07,1.927026e-07,1.927028e-07,1.927030e-07,1.927032e-07,1.927034e-07,1.927037e-07,1.927039e-07,1.927041e-07,1.927043e-07,1.927045e-07,1.927047e-07,1.927050e-07,1.927052e-07,1.927054e-07,1.927056e-07,1.927058e-07,1.927061e-07,1.927063e-07,1.927065e-07,1.927067e-07,1.927069e-07,1.927071e-07,1.927074e-07,1.927076e-07,1.927078e-07,1.927080e-07,1.927082e-07,1.927084e-07,1.927087e-07,1.927089e-07,1.927091e-07,1.927093e-07,1.927095e-07,1.927098e-07,1.927100e-07,1.927102e-07,1.927104e-07,1.927106e-07,1.927108e-07,1.927111e-07,1.927113e-07,1.927115e-07,1.927117e-07,1.927119e-07,1.927122e-07,1.927124e-07,1.927126e-07,1.927128e-07,1.927130e-07,1.927132e-07,1.927135e-07,1.927137e-07,1.927139e-07,1.927141e-07,1.927143e-07,1.927145e-07,1.927148e-07,1.927150e-07,1.927152e-07,1.927154e-07,1.927156e-07,1.927159e-07,1.927161e-07,1.927163e-07,1.927165e-07,1.927167e-07,1.927169e-07,1.927172e-07,1.927174e-07,1.927176e-07,1.927178e-07,1.927180e-07,1.927182e-07,1.927185e-07,1.927187e-07,1.927189e-07,1.927191e-07,1.927193e-07,1.927195e-07,1.927198e-07,1.927200e-07,1.927202e-07,1.927204e-07,1.927206e-07,1.927209e-07,1.927211e-07,1.927213e-07,1.927215e-07,1.927217e-07,1.927219e-07,1.927222e-07,1.927224e-07,1.927226e-07,1.927228e-07,1.927230e-07,1.927232e-07,1.927235e-07,1.927237e-07,1.927239e-07,1.927241e-07,1.927243e-07,1.927246e-07,1.927248e-07,1.927250e-07,1.927252e-07,1.927254e-07,1.927256e-07,1.927259e-07,1.927261e-07,1.927263e-07,1.927265e-07,1.927267e-07,1.927269e-07,1.927272e-07,1.927274e-07,1.927276e-07,1.927278e-07,1.927280e-07,1.927282e-07,1.927285e-07,1.927287e-07,1.927289e-07,1.927291e-07,1.927293e-07,1.927296e-07,1.927298e-07,1.927300e-07,1.927302e-07,1.927304e-07,1.927306e-07,1.927309e-07,1.927311e-07,1.927313e-07,1.927315e-07,1.927317e-07,1.927319e-07,1.927322e-07,1.927324e-07,1.927326e-07,1.927328e-07,1.927330e-07,1.927332e-07,1.927335e-07,1.927337e-07,1.927339e-07,1.927341e-07,1.927343e-07,1.927345e-07,1.927348e-07,1.927350e-07,1.927352e-07,1.927354e-07,1.927356e-07,1.927359e-07,1.927361e-07,1.927363e-07,1.927365e-07,1.927367e-07,1.927369e-07,1.927372e-07,1.927374e-07,1.927376e-07,1.927378e-07,1.927380e-07,1.927382e-07,1.927385e-07,1.927387e-07,1.927389e-07,1.927391e-07,1.927393e-07,1.927395e-07,1.927398e-07,1.927400e-07,1.927402e-07,1.927404e-07,1.927406e-07,1.927408e-07,1.927411e-07,1.927413e-07,1.927415e-07,1.927417e-07,1.927419e-07,1.927422e-07,1.927424e-07,1.927426e-07,1.927428e-07,1.927430e-07,1.927432e-07,1.927435e-07,1.927437e-07,1.927439e-07,1.927441e-07,1.927443e-07,1.927445e-07,1.927448e-07,1.927450e-07,1.927452e-07,1.927454e-07,1.927456e-07,1.927458e-07,1.927461e-07,1.927463e-07,1.927465e-07,1.927467e-07,1.927469e-07,1.927471e-07,1.927474e-07,1.927476e-07,1.927478e-07,1.927480e-07,1.927482e-07,1.927484e-07,1.927487e-07,1.927489e-07,1.927491e-07,1.927493e-07,1.927495e-07,1.927497e-07,1.927500e-07,1.927502e-07,1.927504e-07,1.927506e-07,1.927508e-07,1.927511e-07,1.927513e-07,1.927515e-07,1.927517e-07,1.927519e-07,1.927521e-07,1.927524e-07,1.927526e-07,1.927528e-07,1.927530e-07,1.927532e-07,1.927534e-07,1.927537e-07,1.927539e-07,1.927541e-07,1.927543e-07,1.927545e-07,1.927547e-07,1.927550e-07,1.927552e-07,1.927554e-07,1.927556e-07,1.927558e-07,1.927560e-07,1.927563e-07,1.927565e-07,1.927567e-07,1.927569e-07,1.927571e-07,1.927573e-07,1.927576e-07,1.927578e-07,1.927580e-07,1.927582e-07,1.927584e-07,1.927586e-07,1.927589e-07,1.927591e-07,1.927593e-07,1.927595e-07,1.927597e-07,1.927599e-07,1.927602e-07,1.927604e-07,1.927606e-07,1.927608e-07,1.927610e-07,1.927612e-07,1.927615e-07,1.927617e-07,1.927619e-07,1.927621e-07,1.927623e-07,1.927625e-07,1.927628e-07,1.927630e-07,1.927632e-07,1.927634e-07,1.927636e-07,1.927638e-07,1.927641e-07,1.927643e-07,1.927645e-07,1.927647e-07,1.927649e-07,1.927651e-07,1.927654e-07,1.927656e-07,1.927658e-07,1.927660e-07,1.927662e-07,1.927664e-07,1.927667e-07,1.927669e-07,1.927671e-07,1.927673e-07,1.927675e-07,1.927677e-07,1.927680e-07,1.927682e-07,1.927684e-07,1.927686e-07,1.927688e-07,1.927690e-07,1.927693e-07,1.927695e-07,1.927697e-07,1.927699e-07,1.927701e-07,1.927703e-07,1.927706e-07,1.927708e-07,1.927710e-07,1.927712e-07,1.927714e-07,1.927716e-07,1.927719e-07,1.927721e-07,1.927723e-07,1.927725e-07,1.927727e-07,1.927729e-07,1.927732e-07,1.927734e-07,1.927736e-07,1.927738e-07,1.927740e-07,1.927742e-07,1.927745e-07,1.927747e-07,1.927749e-07,1.927751e-07,1.927753e-07,1.927755e-07,1.927758e-07,1.927760e-07,1.927762e-07,1.927764e-07,1.927766e-07,1.927768e-07,1.927771e-07,1.927773e-07,1.927775e-07,1.927777e-07,1.927779e-07,1.927781e-07,1.927784e-07,1.927786e-07,1.927788e-07,1.927790e-07,1.927792e-07,1.927794e-07,1.927797e-07,1.927799e-07,1.927801e-07,1.927803e-07,1.927805e-07,1.927807e-07,1.927810e-07,1.927812e-07,1.927814e-07,1.927816e-07,1.927818e-07,1.927820e-07,1.927823e-07,1.927825e-07,1.927827e-07,1.927829e-07,1.927831e-07,1.927833e-07,1.927835e-07,1.927838e-07,1.927840e-07,1.927842e-07,1.927844e-07,1.927846e-07,1.927848e-07,1.927851e-07,1.927853e-07,1.927855e-07,1.927857e-07,1.927859e-07,1.927861e-07,1.927864e-07,1.927866e-07,1.927868e-07,1.927870e-07,1.927872e-07,1.927874e-07,1.927877e-07,1.927879e-07,1.927881e-07,1.927883e-07,1.927885e-07,1.927887e-07,1.927890e-07,1.927892e-07,1.927894e-07,1.927896e-07,1.927898e-07,1.927900e-07,1.927903e-07,1.927905e-07,1.927907e-07,1.927909e-07,1.927911e-07,1.927913e-07,1.927916e-07,1.927918e-07,1.927920e-07,1.927922e-07,1.927924e-07,1.927926e-07,1.927928e-07,1.927931e-07,1.927933e-07,1.927935e-07,1.927937e-07,1.927939e-07,1.927941e-07,1.927944e-07,1.927946e-07,1.927948e-07,1.927950e-07,1.927952e-07,1.927954e-07,1.927957e-07,1.927959e-07,1.927961e-07,1.927963e-07,1.927965e-07,1.927967e-07,1.927970e-07,1.927972e-07,1.927974e-07,1.927976e-07,1.927978e-07,1.927980e-07,1.927983e-07,1.927985e-07,1.927987e-07,1.927989e-07,1.927991e-07,1.927993e-07,1.927995e-07,1.927998e-07,1.928000e-07,1.928002e-07,1.928004e-07,1.928006e-07,1.928008e-07,1.928011e-07,1.928013e-07,1.928015e-07,1.928017e-07,1.928019e-07,1.928021e-07,1.928024e-07,1.928026e-07,1.928028e-07,1.928030e-07,1.928032e-07,1.928034e-07,1.928037e-07,1.928039e-07,1.928041e-07,1.928043e-07,1.928045e-07,1.928047e-07,1.928049e-07,1.928052e-07,1.928054e-07,1.928056e-07,1.928058e-07,1.928060e-07,1.928062e-07,1.928065e-07,1.928067e-07,1.928069e-07,1.928071e-07,1.928073e-07,1.928075e-07,1.928078e-07,1.928080e-07,1.928082e-07,1.928084e-07,1.928086e-07,1.928088e-07,1.928091e-07,1.928093e-07,1.928095e-07,1.928097e-07,1.928099e-07,1.928101e-07,1.928103e-07,1.928106e-07,1.928108e-07,1.928110e-07,1.928112e-07,1.928114e-07,1.928116e-07,1.928119e-07,1.928121e-07,1.928123e-07,1.928125e-07,1.928127e-07,1.928129e-07,1.928132e-07,1.928134e-07,1.928136e-07,1.928138e-07,1.928140e-07,1.928142e-07,1.928144e-07,1.928147e-07,1.928149e-07,1.928151e-07,1.928153e-07,1.928155e-07,1.928157e-07,1.928160e-07,1.928162e-07,1.928164e-07,1.928166e-07,1.928168e-07,1.928170e-07,1.928173e-07,1.928175e-07,1.928177e-07,1.928179e-07,1.928181e-07,1.928183e-07,1.928185e-07,1.928188e-07,1.928190e-07,1.928192e-07,1.928194e-07,1.928196e-07,1.928198e-07,1.928201e-07,1.928203e-07,1.928205e-07,1.928207e-07,1.928209e-07,1.928211e-07,1.928213e-07,1.928216e-07,1.928218e-07,1.928220e-07,1.928222e-07,1.928224e-07,1.928226e-07,1.928229e-07,1.928231e-07,1.928233e-07,1.928235e-07,1.928237e-07,1.928239e-07,1.928242e-07,1.928244e-07,1.928246e-07,1.928248e-07,1.928250e-07,1.928252e-07,1.928254e-07,1.928257e-07,1.928259e-07,1.928261e-07,1.928263e-07,1.928265e-07,1.928267e-07,1.928270e-07,1.928272e-07,1.928274e-07,1.928276e-07,1.928278e-07,1.928280e-07,1.928282e-07,1.928285e-07,1.928287e-07,1.928289e-07,1.928291e-07,1.928293e-07,1.928295e-07,1.928298e-07,1.928300e-07,1.928302e-07,1.928304e-07,1.928306e-07,1.928308e-07,1.928310e-07,1.928313e-07,1.928315e-07,1.928317e-07,1.928319e-07,1.928321e-07,1.928323e-07,1.928326e-07,1.928328e-07,1.928330e-07,1.928332e-07,1.928334e-07,1.928336e-07,1.928339e-07,1.928341e-07,1.928343e-07,1.928345e-07,1.928347e-07,1.928349e-07,1.928351e-07,1.928354e-07,1.928356e-07,1.928358e-07,1.928360e-07,1.928362e-07,1.928364e-07,1.928367e-07,1.928369e-07,1.928371e-07,1.928373e-07,1.928375e-07,1.928377e-07,1.928379e-07,1.928382e-07,1.928384e-07,1.928386e-07,1.928388e-07,1.928390e-07,1.928392e-07,1.928395e-07,1.928397e-07,1.928399e-07,1.928401e-07,1.928403e-07,1.928405e-07,1.928407e-07,1.928410e-07,1.928412e-07,1.928414e-07,1.928416e-07,1.928418e-07,1.928420e-07,1.928422e-07,1.928425e-07,1.928427e-07,1.928429e-07,1.928431e-07,1.928433e-07,1.928435e-07,1.928438e-07,1.928440e-07,1.928442e-07,1.928444e-07,1.928446e-07,1.928448e-07,1.928450e-07,1.928453e-07,1.928455e-07,1.928457e-07,1.928459e-07,1.928461e-07,1.928463e-07,1.928466e-07,1.928468e-07,1.928470e-07,1.928472e-07,1.928474e-07,1.928476e-07,1.928478e-07,1.928481e-07,1.928483e-07,1.928485e-07,1.928487e-07,1.928489e-07,1.928491e-07,1.928494e-07,1.928496e-07,1.928498e-07,1.928500e-07,1.928502e-07,1.928504e-07,1.928506e-07,1.928509e-07,1.928511e-07,1.928513e-07,1.928515e-07,1.928517e-07,1.928519e-07,1.928521e-07,1.928524e-07,1.928526e-07,1.928528e-07,1.928530e-07,1.928532e-07,1.928534e-07,1.928537e-07,1.928539e-07,1.928541e-07,1.928543e-07,1.928545e-07,1.928547e-07,1.928549e-07,1.928552e-07,1.928554e-07,1.928556e-07,1.928558e-07,1.928560e-07,1.928562e-07,1.928564e-07,1.928567e-07,1.928569e-07,1.928571e-07,1.928573e-07,1.928575e-07,1.928577e-07,1.928580e-07,1.928582e-07,1.928584e-07,1.928586e-07,1.928588e-07,1.928590e-07,1.928592e-07,1.928595e-07,1.928597e-07,1.928599e-07,1.928601e-07,1.928603e-07,1.928605e-07,1.928607e-07,1.928610e-07,1.928612e-07,1.928614e-07,1.928616e-07,1.928618e-07,1.928620e-07,1.928623e-07,1.928625e-07,1.928627e-07,1.928629e-07,1.928631e-07,1.928633e-07,1.928635e-07,1.928638e-07,1.928640e-07,1.928642e-07,1.928644e-07,1.928646e-07,1.928648e-07,1.928650e-07,1.928653e-07,1.928655e-07,1.928657e-07,1.928659e-07,1.928661e-07,1.928663e-07,1.928665e-07,1.928668e-07,1.928670e-07,1.928672e-07,1.928674e-07,1.928676e-07,1.928678e-07,1.928681e-07,1.928683e-07,1.928685e-07,1.928687e-07,1.928689e-07,1.928691e-07,1.928693e-07,1.928696e-07,1.928698e-07,1.928700e-07,1.928702e-07,1.928704e-07,1.928706e-07,1.928708e-07,1.928711e-07,1.928713e-07,1.928715e-07,1.928717e-07,1.928719e-07,1.928721e-07,1.928723e-07,1.928726e-07,1.928728e-07,1.928730e-07,1.928732e-07,1.928734e-07,1.928736e-07,1.928739e-07,1.928741e-07,1.928743e-07,1.928745e-07,1.928747e-07,1.928749e-07,1.928751e-07,1.928754e-07,1.928756e-07,1.928758e-07,1.928760e-07,1.928762e-07,1.928764e-07,1.928766e-07,1.928769e-07,1.928771e-07,1.928773e-07,1.928775e-07,1.928777e-07,1.928779e-07,1.928781e-07,1.928784e-07,1.928786e-07,1.928788e-07,1.928790e-07,1.928792e-07,1.928794e-07,1.928796e-07,1.928799e-07,1.928801e-07,1.928803e-07,1.928805e-07,1.928807e-07,1.928809e-07,1.928811e-07,1.928814e-07,1.928816e-07,1.928818e-07,1.928820e-07,1.928822e-07,1.928824e-07,1.928827e-07,1.928829e-07,1.928831e-07,1.928833e-07,1.928835e-07,1.928837e-07,1.928839e-07,1.928842e-07,1.928844e-07,1.928846e-07,1.928848e-07,1.928850e-07,1.928852e-07,1.928854e-07,1.928857e-07,1.928859e-07,1.928861e-07,1.928863e-07,1.928865e-07,1.928867e-07,1.928869e-07,1.928872e-07,1.928874e-07,1.928876e-07,1.928878e-07,1.928880e-07,1.928882e-07,1.928884e-07,1.928887e-07,1.928889e-07,1.928891e-07,1.928893e-07,1.928895e-07,1.928897e-07,1.928899e-07,1.928902e-07,1.928904e-07,1.928906e-07,1.928908e-07,1.928910e-07,1.928912e-07,1.928914e-07,1.928917e-07,1.928919e-07,1.928921e-07,1.928923e-07,1.928925e-07,1.928927e-07,1.928929e-07,1.928932e-07,1.928934e-07,1.928936e-07,1.928938e-07,1.928940e-07,1.928942e-07,1.928944e-07,1.928947e-07,1.928949e-07,1.928951e-07,1.928953e-07,1.928955e-07,1.928957e-07,1.928959e-07,1.928962e-07,1.928964e-07,1.928966e-07,1.928968e-07,1.928970e-07,1.928972e-07,1.928974e-07,1.928977e-07,1.928979e-07,1.928981e-07,1.928983e-07,1.928985e-07,1.928987e-07,1.928989e-07,1.928992e-07,1.928994e-07,1.928996e-07,1.928998e-07,1.929000e-07,1.929002e-07,1.929004e-07,1.929007e-07,1.929009e-07,1.929011e-07,1.929013e-07,1.929015e-07,1.929017e-07,1.929019e-07,1.929022e-07,1.929024e-07,1.929026e-07,1.929028e-07,1.929030e-07,1.929032e-07,1.929034e-07,1.929037e-07,1.929039e-07,1.929041e-07,1.929043e-07,1.929045e-07,1.929047e-07,1.929049e-07,1.929052e-07,1.929054e-07,1.929056e-07,1.929058e-07,1.929060e-07,1.929062e-07,1.929064e-07,1.929067e-07,1.929069e-07,1.929071e-07,1.929073e-07,1.929075e-07,1.929077e-07,1.929079e-07,1.929082e-07,1.929084e-07,1.929086e-07,1.929088e-07,1.929090e-07,1.929092e-07,1.929094e-07,1.929097e-07,1.929099e-07,1.929101e-07,1.929103e-07,1.929105e-07,1.929107e-07,1.929109e-07,1.929111e-07,1.929114e-07,1.929116e-07,1.929118e-07,1.929120e-07,1.929122e-07,1.929124e-07,1.929126e-07,1.929129e-07,1.929131e-07,1.929133e-07,1.929135e-07,1.929137e-07,1.929139e-07,1.929141e-07,1.929144e-07,1.929146e-07,1.929148e-07,1.929150e-07,1.929152e-07,1.929154e-07,1.929156e-07,1.929159e-07,1.929161e-07,1.929163e-07,1.929165e-07,1.929167e-07,1.929169e-07,1.929171e-07,1.929174e-07,1.929176e-07,1.929178e-07,1.929180e-07,1.929182e-07,1.929184e-07,1.929186e-07,1.929189e-07,1.929191e-07,1.929193e-07,1.929195e-07,1.929197e-07,1.929199e-07,1.929201e-07,1.929203e-07,1.929206e-07,1.929208e-07,1.929210e-07,1.929212e-07,1.929214e-07,1.929216e-07,1.929218e-07,1.929221e-07,1.929223e-07,1.929225e-07,1.929227e-07,1.929229e-07,1.929231e-07,1.929233e-07,1.929236e-07,1.929238e-07,1.929240e-07,1.929242e-07,1.929244e-07,1.929246e-07,1.929248e-07,1.929251e-07,1.929253e-07,1.929255e-07,1.929257e-07,1.929259e-07,1.929261e-07,1.929263e-07,1.929265e-07,1.929268e-07,1.929270e-07,1.929272e-07,1.929274e-07,1.929276e-07,1.929278e-07,1.929280e-07,1.929283e-07,1.929285e-07,1.929287e-07,1.929289e-07,1.929291e-07,1.929293e-07,1.929295e-07,1.929298e-07,1.929300e-07,1.929302e-07,1.929304e-07,1.929306e-07,1.929308e-07,1.929310e-07,1.929312e-07,1.929315e-07,1.929317e-07,1.929319e-07,1.929321e-07,1.929323e-07,1.929325e-07,1.929327e-07,1.929330e-07,1.929332e-07,1.929334e-07,1.929336e-07,1.929338e-07,1.929340e-07,1.929342e-07,1.929345e-07,1.929347e-07,1.929349e-07,1.929351e-07,1.929353e-07,1.929355e-07,1.929357e-07,1.929359e-07,1.929362e-07,1.929364e-07,1.929366e-07,1.929368e-07,1.929370e-07,1.929372e-07,1.929374e-07,1.929377e-07,1.929379e-07,1.929381e-07,1.929383e-07,1.929385e-07,1.929387e-07,1.929389e-07,1.929391e-07,1.929394e-07,1.929396e-07,1.929398e-07,1.929400e-07,1.929402e-07,1.929404e-07,1.929406e-07,1.929409e-07,1.929411e-07,1.929413e-07,1.929415e-07,1.929417e-07,1.929419e-07,1.929421e-07,1.929424e-07,1.929426e-07,1.929428e-07,1.929430e-07,1.929432e-07,1.929434e-07,1.929436e-07,1.929438e-07,1.929441e-07,1.929443e-07,1.929445e-07,1.929447e-07,1.929449e-07,1.929451e-07,1.929453e-07,1.929456e-07,1.929458e-07,1.929460e-07,1.929462e-07,1.929464e-07,1.929466e-07,1.929468e-07,1.929470e-07,1.929473e-07,1.929475e-07,1.929477e-07,1.929479e-07,1.929481e-07,1.929483e-07,1.929485e-07,1.929488e-07,1.929490e-07,1.929492e-07,1.929494e-07,1.929496e-07,1.929498e-07,1.929500e-07,1.929502e-07,1.929505e-07,1.929507e-07,1.929509e-07,1.929511e-07,1.929513e-07,1.929515e-07,1.929517e-07,1.929520e-07,1.929522e-07,1.929524e-07,1.929526e-07,1.929528e-07,1.929530e-07,1.929532e-07,1.929534e-07,1.929537e-07,1.929539e-07,1.929541e-07,1.929543e-07,1.929545e-07,1.929547e-07,1.929549e-07,1.929552e-07,1.929554e-07,1.929556e-07,1.929558e-07,1.929560e-07,1.929562e-07,1.929564e-07,1.929566e-07,1.929569e-07,1.929571e-07,1.929573e-07,1.929575e-07,1.929577e-07,1.929579e-07,1.929581e-07,1.929583e-07,1.929586e-07,1.929588e-07,1.929590e-07,1.929592e-07,1.929594e-07,1.929596e-07,1.929598e-07,1.929601e-07,1.929603e-07,1.929605e-07,1.929607e-07,1.929609e-07,1.929611e-07,1.929613e-07,1.929615e-07,1.929618e-07,1.929620e-07,1.929622e-07,1.929624e-07,1.929626e-07,1.929628e-07,1.929630e-07,1.929633e-07,1.929635e-07,1.929637e-07,1.929639e-07,1.929641e-07,1.929643e-07,1.929645e-07,1.929647e-07,1.929650e-07,1.929652e-07,1.929654e-07,1.929656e-07,1.929658e-07,1.929660e-07,1.929662e-07,1.929664e-07,1.929667e-07,1.929669e-07,1.929671e-07,1.929673e-07,1.929675e-07,1.929677e-07,1.929679e-07,1.929681e-07,1.929684e-07,1.929686e-07,1.929688e-07,1.929690e-07,1.929692e-07,1.929694e-07,1.929696e-07,1.929699e-07,1.929701e-07,1.929703e-07,1.929705e-07,1.929707e-07,1.929709e-07,1.929711e-07,1.929713e-07,1.929716e-07,1.929718e-07,1.929720e-07,1.929722e-07,1.929724e-07,1.929726e-07,1.929728e-07,1.929730e-07,1.929733e-07,1.929735e-07,1.929737e-07,1.929739e-07,1.929741e-07,1.929743e-07,1.929745e-07,1.929747e-07,1.929750e-07,1.929752e-07,1.929754e-07,1.929756e-07,1.929758e-07,1.929760e-07,1.929762e-07,1.929765e-07,1.929767e-07,1.929769e-07,1.929771e-07,1.929773e-07,1.929775e-07,1.929777e-07,1.929779e-07,1.929782e-07,1.929784e-07,1.929786e-07,1.929788e-07,1.929790e-07,1.929792e-07,1.929794e-07,1.929796e-07,1.929799e-07,1.929801e-07,1.929803e-07,1.929805e-07,1.929807e-07,1.929809e-07,1.929811e-07,1.929813e-07,1.929816e-07,1.929818e-07,1.929820e-07,1.929822e-07,1.929824e-07,1.929826e-07,1.929828e-07,1.929830e-07,1.929833e-07,1.929835e-07,1.929837e-07,1.929839e-07,1.929841e-07,1.929843e-07,1.929845e-07,1.929847e-07,1.929850e-07,1.929852e-07,1.929854e-07,1.929856e-07,1.929858e-07,1.929860e-07,1.929862e-07,1.929865e-07,1.929867e-07,1.929869e-07,1.929871e-07,1.929873e-07,1.929875e-07,1.929877e-07,1.929879e-07,1.929882e-07,1.929884e-07,1.929886e-07,1.929888e-07,1.929890e-07,1.929892e-07,1.929894e-07,1.929896e-07,1.929899e-07,1.929901e-07,1.929903e-07,1.929905e-07,1.929907e-07,1.929909e-07,1.929911e-07,1.929913e-07,1.929916e-07,1.929918e-07,1.929920e-07,1.929922e-07,1.929924e-07,1.929926e-07,1.929928e-07,1.929930e-07,1.929933e-07,1.929935e-07,1.929937e-07,1.929939e-07,1.929941e-07,1.929943e-07,1.929945e-07,1.929947e-07,1.929950e-07,1.929952e-07,1.929954e-07,1.929956e-07,1.929958e-07,1.929960e-07,1.929962e-07,1.929964e-07,1.929967e-07,1.929969e-07,1.929971e-07,1.929973e-07,1.929975e-07,1.929977e-07,1.929979e-07,1.929981e-07,1.929984e-07,1.929986e-07,1.929988e-07,1.929990e-07,1.929992e-07,1.929994e-07,1.929996e-07,1.929998e-07,1.930001e-07,1.930003e-07,1.930005e-07,1.930007e-07,1.930009e-07,1.930011e-07,1.930013e-07,1.930015e-07,1.930018e-07,1.930020e-07,1.930022e-07,1.930024e-07,1.930026e-07,1.930028e-07,1.930030e-07,1.930032e-07,1.930034e-07,1.930037e-07,1.930039e-07,1.930041e-07,1.930043e-07,1.930045e-07,1.930047e-07,1.930049e-07,1.930051e-07,1.930054e-07,1.930056e-07,1.930058e-07,1.930060e-07,1.930062e-07,1.930064e-07,1.930066e-07,1.930068e-07,1.930071e-07,1.930073e-07,1.930075e-07,1.930077e-07,1.930079e-07,1.930081e-07,1.930083e-07,1.930085e-07,1.930088e-07,1.930090e-07,1.930092e-07,1.930094e-07,1.930096e-07,1.930098e-07,1.930100e-07,1.930102e-07,1.930105e-07,1.930107e-07,1.930109e-07,1.930111e-07,1.930113e-07,1.930115e-07,1.930117e-07,1.930119e-07,1.930122e-07,1.930124e-07,1.930126e-07,1.930128e-07,1.930130e-07,1.930132e-07,1.930134e-07,1.930136e-07,1.930138e-07,1.930141e-07,1.930143e-07,1.930145e-07,1.930147e-07,1.930149e-07,1.930151e-07,1.930153e-07,1.930155e-07,1.930158e-07,1.930160e-07,1.930162e-07,1.930164e-07,1.930166e-07,1.930168e-07,1.930170e-07,1.930172e-07,1.930175e-07,1.930177e-07,1.930179e-07,1.930181e-07,1.930183e-07,1.930185e-07,1.930187e-07,1.930189e-07,1.930192e-07,1.930194e-07,1.930196e-07,1.930198e-07,1.930200e-07,1.930202e-07,1.930204e-07,1.930206e-07,1.930208e-07,1.930211e-07,1.930213e-07,1.930215e-07,1.930217e-07,1.930219e-07,1.930221e-07,1.930223e-07,1.930225e-07,1.930228e-07,1.930230e-07,1.930232e-07,1.930234e-07,1.930236e-07,1.930238e-07,1.930240e-07,1.930242e-07,1.930245e-07,1.930247e-07,1.930249e-07,1.930251e-07,1.930253e-07,1.930255e-07,1.930257e-07,1.930259e-07,1.930261e-07,1.930264e-07,1.930266e-07,1.930268e-07,1.930270e-07,1.930272e-07,1.930274e-07,1.930276e-07,1.930278e-07,1.930281e-07,1.930283e-07,1.930285e-07,1.930287e-07,1.930289e-07,1.930291e-07,1.930293e-07,1.930295e-07,1.930297e-07,1.930300e-07,1.930302e-07,1.930304e-07,1.930306e-07,1.930308e-07,1.930310e-07,1.930312e-07,1.930314e-07,1.930317e-07,1.930319e-07,1.930321e-07,1.930323e-07,1.930325e-07,1.930327e-07,1.930329e-07,1.930331e-07,1.930333e-07,1.930336e-07,1.930338e-07,1.930340e-07,1.930342e-07,1.930344e-07,1.930346e-07,1.930348e-07,1.930350e-07,1.930353e-07,1.930355e-07,1.930357e-07,1.930359e-07,1.930361e-07,1.930363e-07,1.930365e-07,1.930367e-07,1.930369e-07,1.930372e-07,1.930374e-07,1.930376e-07,1.930378e-07,1.930380e-07,1.930382e-07,1.930384e-07,1.930386e-07,1.930389e-07,1.930391e-07,1.930393e-07,1.930395e-07,1.930397e-07,1.930399e-07,1.930401e-07,1.930403e-07,1.930405e-07,1.930408e-07,1.930410e-07,1.930412e-07,1.930414e-07,1.930416e-07,1.930418e-07,1.930420e-07,1.930422e-07,1.930425e-07,1.930427e-07,1.930429e-07,1.930431e-07,1.930433e-07,1.930435e-07,1.930437e-07,1.930439e-07,1.930441e-07,1.930444e-07,1.930446e-07,1.930448e-07,1.930450e-07,1.930452e-07,1.930454e-07,1.930456e-07,1.930458e-07,1.930460e-07,1.930463e-07,1.930465e-07,1.930467e-07,1.930469e-07,1.930471e-07,1.930473e-07,1.930475e-07,1.930477e-07,1.930480e-07,1.930482e-07,1.930484e-07,1.930486e-07,1.930488e-07,1.930490e-07,1.930492e-07,1.930494e-07,1.930496e-07,1.930499e-07,1.930501e-07,1.930503e-07,1.930505e-07,1.930507e-07,1.930509e-07,1.930511e-07,1.930513e-07,1.930515e-07,1.930518e-07,1.930520e-07,1.930522e-07,1.930524e-07,1.930526e-07,1.930528e-07,1.930530e-07,1.930532e-07,1.930535e-07,1.930537e-07,1.930539e-07,1.930541e-07,1.930543e-07,1.930545e-07,1.930547e-07,1.930549e-07,1.930551e-07,1.930554e-07,1.930556e-07,1.930558e-07,1.930560e-07,1.930562e-07,1.930564e-07,1.930566e-07,1.930568e-07,1.930570e-07,1.930573e-07,1.930575e-07,1.930577e-07,1.930579e-07,1.930581e-07,1.930583e-07,1.930585e-07,1.930587e-07,1.930589e-07,1.930592e-07,1.930594e-07,1.930596e-07,1.930598e-07,1.930600e-07,1.930602e-07,1.930604e-07,1.930606e-07,1.930608e-07,1.930611e-07,1.930613e-07,1.930615e-07,1.930617e-07,1.930619e-07,1.930621e-07,1.930623e-07,1.930625e-07,1.930627e-07,1.930630e-07,1.930632e-07,1.930634e-07,1.930636e-07,1.930638e-07,1.930640e-07,1.930642e-07,1.930644e-07,1.930647e-07,1.930649e-07,1.930651e-07,1.930653e-07,1.930655e-07,1.930657e-07,1.930659e-07,1.930661e-07,1.930663e-07,1.930666e-07,1.930668e-07,1.930670e-07,1.930672e-07,1.930674e-07,1.930676e-07,1.930678e-07,1.930680e-07,1.930682e-07,1.930685e-07,1.930687e-07,1.930689e-07,1.930691e-07,1.930693e-07,1.930695e-07,1.930697e-07,1.930699e-07,1.930701e-07,1.930704e-07,1.930706e-07,1.930708e-07,1.930710e-07,1.930712e-07,1.930714e-07,1.930716e-07,1.930718e-07,1.930720e-07,1.930723e-07,1.930725e-07,1.930727e-07,1.930729e-07,1.930731e-07,1.930733e-07,1.930735e-07,1.930737e-07,1.930739e-07,1.930742e-07,1.930744e-07,1.930746e-07,1.930748e-07,1.930750e-07,1.930752e-07,1.930754e-07,1.930756e-07,1.930758e-07,1.930761e-07,1.930763e-07,1.930765e-07,1.930767e-07,1.930769e-07,1.930771e-07,1.930773e-07,1.930775e-07,1.930777e-07,1.930780e-07,1.930782e-07,1.930784e-07,1.930786e-07,1.930788e-07,1.930790e-07,1.930792e-07,1.930794e-07,1.930796e-07,1.930798e-07,1.930801e-07,1.930803e-07,1.930805e-07,1.930807e-07,1.930809e-07,1.930811e-07,1.930813e-07,1.930815e-07,1.930817e-07,1.930820e-07,1.930822e-07,1.930824e-07,1.930826e-07,1.930828e-07,1.930830e-07,1.930832e-07,1.930834e-07,1.930836e-07,1.930839e-07,1.930841e-07,1.930843e-07,1.930845e-07,1.930847e-07,1.930849e-07,1.930851e-07,1.930853e-07,1.930855e-07,1.930858e-07,1.930860e-07,1.930862e-07,1.930864e-07,1.930866e-07,1.930868e-07,1.930870e-07,1.930872e-07,1.930874e-07,1.930877e-07,1.930879e-07,1.930881e-07,1.930883e-07,1.930885e-07,1.930887e-07,1.930889e-07,1.930891e-07,1.930893e-07,1.930895e-07,1.930898e-07,1.930900e-07,1.930902e-07,1.930904e-07,1.930906e-07,1.930908e-07,1.930910e-07,1.930912e-07,1.930914e-07,1.930917e-07,1.930919e-07,1.930921e-07,1.930923e-07,1.930925e-07,1.930927e-07,1.930929e-07,1.930931e-07,1.930933e-07,1.930936e-07,1.930938e-07,1.930940e-07,1.930942e-07,1.930944e-07,1.930946e-07,1.930948e-07,1.930950e-07,1.930952e-07,1.930954e-07,1.930957e-07,1.930959e-07,1.930961e-07,1.930963e-07,1.930965e-07,1.930967e-07,1.930969e-07,1.930971e-07,1.930973e-07,1.930976e-07,1.930978e-07,1.930980e-07,1.930982e-07,1.930984e-07,1.930986e-07,1.930988e-07,1.930990e-07,1.930992e-07,1.930995e-07,1.930997e-07,1.930999e-07,1.931001e-07,1.931003e-07,1.931005e-07,1.931007e-07,1.931009e-07,1.931011e-07,1.931013e-07,1.931016e-07,1.931018e-07,1.931020e-07,1.931022e-07,1.931024e-07,1.931026e-07,1.931028e-07,1.931030e-07,1.931032e-07,1.931035e-07,1.931037e-07,1.931039e-07,1.931041e-07,1.931043e-07,1.931045e-07,1.931047e-07,1.931049e-07,1.931051e-07,1.931053e-07,1.931056e-07,1.931058e-07,1.931060e-07,1.931062e-07,1.931064e-07,1.931066e-07,1.931068e-07,1.931070e-07,1.931072e-07,1.931075e-07,1.931077e-07,1.931079e-07,1.931081e-07,1.931083e-07,1.931085e-07,1.931087e-07,1.931089e-07,1.931091e-07,1.931093e-07,1.931096e-07,1.931098e-07,1.931100e-07,1.931102e-07,1.931104e-07,1.931106e-07,1.931108e-07,1.931110e-07,1.931112e-07,1.931114e-07,1.931117e-07,1.931119e-07,1.931121e-07,1.931123e-07,1.931125e-07,1.931127e-07,1.931129e-07,1.931131e-07,1.931133e-07,1.931136e-07,1.931138e-07,1.931140e-07,1.931142e-07,1.931144e-07,1.931146e-07,1.931148e-07,1.931150e-07,1.931152e-07,1.931154e-07,1.931157e-07,1.931159e-07,1.931161e-07,1.931163e-07,1.931165e-07,1.931167e-07,1.931169e-07,1.931171e-07,1.931173e-07,1.931175e-07,1.931178e-07,1.931180e-07,1.931182e-07,1.931184e-07,1.931186e-07,1.931188e-07,1.931190e-07,1.931192e-07,1.931194e-07,1.931196e-07,1.931199e-07,1.931201e-07,1.931203e-07,1.931205e-07,1.931207e-07,1.931209e-07,1.931211e-07,1.931213e-07,1.931215e-07,1.931218e-07,1.931220e-07,1.931222e-07,1.931224e-07,1.931226e-07,1.931228e-07,1.931230e-07,1.931232e-07,1.931234e-07,1.931236e-07,1.931239e-07,1.931241e-07,1.931243e-07,1.931245e-07,1.931247e-07,1.931249e-07,1.931251e-07,1.931253e-07,1.931255e-07,1.931257e-07,1.931260e-07,1.931262e-07,1.931264e-07,1.931266e-07,1.931268e-07,1.931270e-07,1.931272e-07,1.931274e-07,1.931276e-07,1.931278e-07,1.931281e-07,1.931283e-07,1.931285e-07,1.931287e-07,1.931289e-07,1.931291e-07,1.931293e-07,1.931295e-07,1.931297e-07,1.931299e-07,1.931302e-07,1.931304e-07,1.931306e-07,1.931308e-07,1.931310e-07,1.931312e-07,1.931314e-07,1.931316e-07,1.931318e-07,1.931320e-07,1.931323e-07,1.931325e-07,1.931327e-07,1.931329e-07,1.931331e-07,1.931333e-07,1.931335e-07,1.931337e-07,1.931339e-07,1.931341e-07,1.931344e-07,1.931346e-07,1.931348e-07,1.931350e-07,1.931352e-07,1.931354e-07,1.931356e-07,1.931358e-07,1.931360e-07,1.931362e-07,1.931365e-07,1.931367e-07,1.931369e-07,1.931371e-07,1.931373e-07,1.931375e-07,1.931377e-07,1.931379e-07,1.931381e-07,1.931383e-07,1.931386e-07,1.931388e-07,1.931390e-07,1.931392e-07,1.931394e-07,1.931396e-07,1.931398e-07,1.931400e-07,1.931402e-07,1.931404e-07,1.931407e-07,1.931409e-07,1.931411e-07,1.931413e-07,1.931415e-07,1.931417e-07,1.931419e-07,1.931421e-07,1.931423e-07,1.931425e-07,1.931428e-07,1.931430e-07,1.931432e-07,1.931434e-07,1.931436e-07,1.931438e-07,1.931440e-07,1.931442e-07,1.931444e-07,1.931446e-07,1.931448e-07,1.931451e-07,1.931453e-07,1.931455e-07,1.931457e-07,1.931459e-07,1.931461e-07,1.931463e-07,1.931465e-07,1.931467e-07,1.931469e-07,1.931472e-07,1.931474e-07,1.931476e-07,1.931478e-07,1.931480e-07,1.931482e-07,1.931484e-07,1.931486e-07,1.931488e-07,1.931490e-07,1.931493e-07,1.931495e-07,1.931497e-07,1.931499e-07,1.931501e-07,1.931503e-07,1.931505e-07,1.931507e-07,1.931509e-07,1.931511e-07,1.931514e-07,1.931516e-07,1.931518e-07,1.931520e-07,1.931522e-07,1.931524e-07,1.931526e-07,1.931528e-07,1.931530e-07,1.931532e-07,1.931534e-07,1.931537e-07,1.931539e-07,1.931541e-07,1.931543e-07,1.931545e-07,1.931547e-07,1.931549e-07,1.931551e-07,1.931553e-07,1.931555e-07,1.931558e-07,1.931560e-07,1.931562e-07,1.931564e-07,1.931566e-07,1.931568e-07,1.931570e-07,1.931572e-07,1.931574e-07,1.931576e-07,1.931578e-07,1.931581e-07,1.931583e-07,1.931585e-07,1.931587e-07,1.931589e-07,1.931591e-07,1.931593e-07,1.931595e-07,1.931597e-07,1.931599e-07,1.931602e-07,1.931604e-07,1.931606e-07,1.931608e-07,1.931610e-07,1.931612e-07,1.931614e-07,1.931616e-07,1.931618e-07,1.931620e-07,1.931622e-07,1.931625e-07,1.931627e-07,1.931629e-07,1.931631e-07,1.931633e-07,1.931635e-07,1.931637e-07,1.931639e-07,1.931641e-07,1.931643e-07,1.931646e-07,1.931648e-07,1.931650e-07,1.931652e-07,1.931654e-07,1.931656e-07,1.931658e-07,1.931660e-07,1.931662e-07,1.931664e-07,1.931666e-07,1.931669e-07,1.931671e-07,1.931673e-07,1.931675e-07,1.931677e-07,1.931679e-07,1.931681e-07,1.931683e-07,1.931685e-07,1.931687e-07,1.931689e-07,1.931692e-07,1.931694e-07,1.931696e-07,1.931698e-07,1.931700e-07,1.931702e-07,1.931704e-07,1.931706e-07,1.931708e-07,1.931710e-07,1.931713e-07,1.931715e-07,1.931717e-07,1.931719e-07,1.931721e-07,1.931723e-07,1.931725e-07,1.931727e-07,1.931729e-07,1.931731e-07,1.931733e-07,1.931736e-07,1.931738e-07,1.931740e-07,1.931742e-07,1.931744e-07,1.931746e-07,1.931748e-07,1.931750e-07,1.931752e-07,1.931754e-07,1.931756e-07,1.931759e-07,1.931761e-07,1.931763e-07,1.931765e-07,1.931767e-07,1.931769e-07,1.931771e-07,1.931773e-07,1.931775e-07,1.931777e-07,1.931779e-07,1.931782e-07,1.931784e-07,1.931786e-07,1.931788e-07,1.931790e-07,1.931792e-07,1.931794e-07,1.931796e-07,1.931798e-07,1.931800e-07,1.931802e-07,1.931805e-07,1.931807e-07,1.931809e-07,1.931811e-07,1.931813e-07,1.931815e-07,1.931817e-07,1.931819e-07,1.931821e-07,1.931823e-07,1.931825e-07,1.931828e-07,1.931830e-07,1.931832e-07,1.931834e-07,1.931836e-07,1.931838e-07,1.931840e-07,1.931842e-07,1.931844e-07,1.931846e-07,1.931848e-07,1.931851e-07,1.931853e-07,1.931855e-07,1.931857e-07,1.931859e-07,1.931861e-07,1.931863e-07,1.931865e-07,1.931867e-07,1.931869e-07,1.931871e-07,1.931874e-07,1.931876e-07,1.931878e-07,1.931880e-07,1.931882e-07,1.931884e-07,1.931886e-07,1.931888e-07,1.931890e-07,1.931892e-07,1.931894e-07,1.931897e-07,1.931899e-07,1.931901e-07,1.931903e-07,1.931905e-07,1.931907e-07,1.931909e-07,1.931911e-07,1.931913e-07,1.931915e-07,1.931917e-07,1.931920e-07,1.931922e-07,1.931924e-07,1.931926e-07,1.931928e-07,1.931930e-07,1.931932e-07,1.931934e-07,1.931936e-07,1.931938e-07,1.931940e-07,1.931943e-07,1.931945e-07,1.931947e-07,1.931949e-07,1.931951e-07,1.931953e-07,1.931955e-07,1.931957e-07,1.931959e-07,1.931961e-07,1.931963e-07,1.931966e-07,1.931968e-07,1.931970e-07,1.931972e-07,1.931974e-07,1.931976e-07,1.931978e-07,1.931980e-07,1.931982e-07,1.931984e-07,1.931986e-07,1.931988e-07,1.931991e-07,1.931993e-07,1.931995e-07,1.931997e-07,1.931999e-07,1.932001e-07,1.932003e-07,1.932005e-07,1.932007e-07,1.932009e-07,1.932011e-07,1.932014e-07,1.932016e-07,1.932018e-07,1.932020e-07,1.932022e-07,1.932024e-07,1.932026e-07,1.932028e-07,1.932030e-07,1.932032e-07,1.932034e-07,1.932036e-07,1.932039e-07,1.932041e-07,1.932043e-07,1.932045e-07,1.932047e-07,1.932049e-07,1.932051e-07,1.932053e-07,1.932055e-07,1.932057e-07,1.932059e-07,1.932062e-07,1.932064e-07,1.932066e-07,1.932068e-07,1.932070e-07,1.932072e-07,1.932074e-07,1.932076e-07,1.932078e-07,1.932080e-07,1.932082e-07,1.932084e-07,1.932087e-07,1.932089e-07,1.932091e-07,1.932093e-07,1.932095e-07,1.932097e-07,1.932099e-07,1.932101e-07,1.932103e-07,1.932105e-07,1.932107e-07,1.932110e-07,1.932112e-07,1.932114e-07,1.932116e-07,1.932118e-07,1.932120e-07,1.932122e-07,1.932124e-07,1.932126e-07,1.932128e-07,1.932130e-07,1.932132e-07,1.932135e-07,1.932137e-07,1.932139e-07,1.932141e-07,1.932143e-07,1.932145e-07,1.932147e-07,1.932149e-07,1.932151e-07,1.932153e-07,1.932155e-07,1.932157e-07,1.932160e-07,1.932162e-07,1.932164e-07,1.932166e-07,1.932168e-07,1.932170e-07,1.932172e-07,1.932174e-07,1.932176e-07,1.932178e-07,1.932180e-07,1.932183e-07,1.932185e-07,1.932187e-07,1.932189e-07,1.932191e-07,1.932193e-07,1.932195e-07,1.932197e-07,1.932199e-07,1.932201e-07,1.932203e-07,1.932205e-07,1.932208e-07,1.932210e-07,1.932212e-07,1.932214e-07,1.932216e-07,1.932218e-07,1.932220e-07,1.932222e-07,1.932224e-07,1.932226e-07,1.932228e-07,1.932230e-07,1.932233e-07,1.932235e-07,1.932237e-07,1.932239e-07,1.932241e-07,1.932243e-07,1.932245e-07,1.932247e-07,1.932249e-07,1.932251e-07,1.932253e-07,1.932255e-07,1.932258e-07,1.932260e-07,1.932262e-07,1.932264e-07,1.932266e-07,1.932268e-07,1.932270e-07,1.932272e-07,1.932274e-07,1.932276e-07,1.932278e-07,1.932280e-07,1.932283e-07,1.932285e-07,1.932287e-07,1.932289e-07,1.932291e-07,1.932293e-07,1.932295e-07,1.932297e-07,1.932299e-07,1.932301e-07,1.932303e-07,1.932305e-07,1.932308e-07,1.932310e-07,1.932312e-07,1.932314e-07,1.932316e-07,1.932318e-07,1.932320e-07,1.932322e-07,1.932324e-07,1.932326e-07,1.932328e-07,1.932330e-07,1.932333e-07,1.932335e-07,1.932337e-07,1.932339e-07,1.932341e-07,1.932343e-07,1.932345e-07,1.932347e-07,1.932349e-07,1.932351e-07,1.932353e-07,1.932355e-07,1.932357e-07,1.932360e-07,1.932362e-07,1.932364e-07,1.932366e-07,1.932368e-07,1.932370e-07,1.932372e-07,1.932374e-07,1.932376e-07,1.932378e-07,1.932380e-07,1.932382e-07,1.932385e-07,1.932387e-07,1.932389e-07,1.932391e-07,1.932393e-07,1.932395e-07,1.932397e-07,1.932399e-07,1.932401e-07,1.932403e-07,1.932405e-07,1.932407e-07,1.932410e-07,1.932412e-07,1.932414e-07,1.932416e-07,1.932418e-07,1.932420e-07,1.932422e-07,1.932424e-07,1.932426e-07,1.932428e-07,1.932430e-07,1.932432e-07,1.932434e-07,1.932437e-07,1.932439e-07,1.932441e-07,1.932443e-07,1.932445e-07,1.932447e-07,1.932449e-07,1.932451e-07,1.932453e-07,1.932455e-07,1.932457e-07,1.932459e-07,1.932462e-07,1.932464e-07,1.932466e-07,1.932468e-07,1.932470e-07,1.932472e-07,1.932474e-07,1.932476e-07,1.932478e-07,1.932480e-07,1.932482e-07,1.932484e-07,1.932486e-07,1.932489e-07,1.932491e-07,1.932493e-07,1.932495e-07,1.932497e-07,1.932499e-07,1.932501e-07,1.932503e-07,1.932505e-07,1.932507e-07,1.932509e-07,1.932511e-07,1.932513e-07,1.932516e-07,1.932518e-07,1.932520e-07,1.932522e-07,1.932524e-07,1.932526e-07,1.932528e-07,1.932530e-07,1.932532e-07,1.932534e-07,1.932536e-07,1.932538e-07,1.932541e-07,1.932543e-07,1.932545e-07,1.932547e-07,1.932549e-07,1.932551e-07,1.932553e-07,1.932555e-07,1.932557e-07,1.932559e-07,1.932561e-07,1.932563e-07,1.932565e-07,1.932568e-07,1.932570e-07,1.932572e-07,1.932574e-07,1.932576e-07,1.932578e-07,1.932580e-07,1.932582e-07,1.932584e-07,1.932586e-07,1.932588e-07,1.932590e-07,1.932592e-07,1.932595e-07,1.932597e-07,1.932599e-07,1.932601e-07,1.932603e-07,1.932605e-07,1.932607e-07,1.932609e-07,1.932611e-07,1.932613e-07,1.932615e-07,1.932617e-07,1.932619e-07,1.932622e-07,1.932624e-07,1.932626e-07,1.932628e-07,1.932630e-07,1.932632e-07,1.932634e-07,1.932636e-07,1.932638e-07,1.932640e-07,1.932642e-07,1.932644e-07,1.932646e-07,1.932649e-07,1.932651e-07,1.932653e-07,1.932655e-07,1.932657e-07,1.932659e-07,1.932661e-07,1.932663e-07,1.932665e-07,1.932667e-07,1.932669e-07,1.932671e-07,1.932673e-07,1.932676e-07,1.932678e-07,1.932680e-07,1.932682e-07,1.932684e-07,1.932686e-07,1.932688e-07,1.932690e-07,1.932692e-07,1.932694e-07,1.932696e-07,1.932698e-07,1.932700e-07,1.932703e-07,1.932705e-07,1.932707e-07,1.932709e-07,1.932711e-07,1.932713e-07,1.932715e-07,1.932717e-07,1.932719e-07,1.932721e-07,1.932723e-07,1.932725e-07,1.932727e-07,1.932729e-07,1.932732e-07,1.932734e-07,1.932736e-07,1.932738e-07,1.932740e-07,1.932742e-07,1.932744e-07,1.932746e-07,1.932748e-07,1.932750e-07,1.932752e-07,1.932754e-07,1.932756e-07,1.932759e-07,1.932761e-07,1.932763e-07,1.932765e-07,1.932767e-07,1.932769e-07,1.932771e-07,1.932773e-07,1.932775e-07,1.932777e-07,1.932779e-07,1.932781e-07,1.932783e-07,1.932785e-07,1.932788e-07,1.932790e-07,1.932792e-07,1.932794e-07,1.932796e-07,1.932798e-07,1.932800e-07,1.932802e-07,1.932804e-07,1.932806e-07,1.932808e-07,1.932810e-07,1.932812e-07,1.932815e-07,1.932817e-07,1.932819e-07,1.932821e-07,1.932823e-07,1.932825e-07,1.932827e-07,1.932829e-07,1.932831e-07,1.932833e-07,1.932835e-07,1.932837e-07,1.932839e-07,1.932841e-07,1.932844e-07,1.932846e-07,1.932848e-07,1.932850e-07,1.932852e-07,1.932854e-07,1.932856e-07,1.932858e-07,1.932860e-07,1.932862e-07,1.932864e-07,1.932866e-07,1.932868e-07,1.932870e-07,1.932873e-07,1.932875e-07,1.932877e-07,1.932879e-07,1.932881e-07,1.932883e-07,1.932885e-07,1.932887e-07,1.932889e-07,1.932891e-07,1.932893e-07,1.932895e-07,1.932897e-07,1.932900e-07,1.932902e-07,1.932904e-07,1.932906e-07,1.932908e-07,1.932910e-07,1.932912e-07,1.932914e-07,1.932916e-07,1.932918e-07,1.932920e-07,1.932922e-07,1.932924e-07,1.932926e-07,1.932929e-07,1.932931e-07,1.932933e-07,1.932935e-07,1.932937e-07,1.932939e-07,1.932941e-07,1.932943e-07,1.932945e-07,1.932947e-07,1.932949e-07,1.932951e-07,1.932953e-07,1.932955e-07,1.932958e-07,1.932960e-07,1.932962e-07,1.932964e-07,1.932966e-07,1.932968e-07,1.932970e-07,1.932972e-07,1.932974e-07,1.932976e-07,1.932978e-07,1.932980e-07,1.932982e-07,1.932984e-07,1.932986e-07,1.932989e-07,1.932991e-07,1.932993e-07,1.932995e-07,1.932997e-07,1.932999e-07,1.933001e-07,1.933003e-07,1.933005e-07,1.933007e-07,1.933009e-07,1.933011e-07,1.933013e-07,1.933015e-07,1.933018e-07,1.933020e-07,1.933022e-07,1.933024e-07,1.933026e-07,1.933028e-07,1.933030e-07,1.933032e-07,1.933034e-07,1.933036e-07,1.933038e-07,1.933040e-07,1.933042e-07,1.933044e-07,1.933047e-07,1.933049e-07,1.933051e-07,1.933053e-07,1.933055e-07,1.933057e-07,1.933059e-07,1.933061e-07,1.933063e-07,1.933065e-07,1.933067e-07,1.933069e-07,1.933071e-07,1.933073e-07,1.933075e-07,1.933078e-07,1.933080e-07,1.933082e-07,1.933084e-07,1.933086e-07,1.933088e-07,1.933090e-07,1.933092e-07,1.933094e-07,1.933096e-07,1.933098e-07,1.933100e-07,1.933102e-07,1.933104e-07,1.933107e-07,1.933109e-07,1.933111e-07,1.933113e-07,1.933115e-07,1.933117e-07,1.933119e-07,1.933121e-07,1.933123e-07,1.933125e-07,1.933127e-07,1.933129e-07,1.933131e-07,1.933133e-07,1.933135e-07,1.933138e-07,1.933140e-07,1.933142e-07,1.933144e-07,1.933146e-07,1.933148e-07,1.933150e-07,1.933152e-07,1.933154e-07,1.933156e-07,1.933158e-07,1.933160e-07,1.933162e-07,1.933164e-07,1.933166e-07,1.933169e-07,1.933171e-07,1.933173e-07,1.933175e-07,1.933177e-07,1.933179e-07,1.933181e-07,1.933183e-07,1.933185e-07,1.933187e-07,1.933189e-07,1.933191e-07,1.933193e-07,1.933195e-07,1.933197e-07,1.933200e-07,1.933202e-07,1.933204e-07,1.933206e-07,1.933208e-07,1.933210e-07,1.933212e-07,1.933214e-07,1.933216e-07,1.933218e-07,1.933220e-07,1.933222e-07,1.933224e-07,1.933226e-07,1.933228e-07,1.933231e-07,1.933233e-07,1.933235e-07,1.933237e-07,1.933239e-07,1.933241e-07,1.933243e-07,1.933245e-07,1.933247e-07,1.933249e-07,1.933251e-07,1.933253e-07,1.933255e-07,1.933257e-07,1.933259e-07,1.933262e-07,1.933264e-07,1.933266e-07,1.933268e-07,1.933270e-07,1.933272e-07,1.933274e-07,1.933276e-07,1.933278e-07,1.933280e-07,1.933282e-07,1.933284e-07,1.933286e-07,1.933288e-07,1.933290e-07,1.933293e-07,1.933295e-07,1.933297e-07,1.933299e-07,1.933301e-07,1.933303e-07,1.933305e-07,1.933307e-07,1.933309e-07,1.933311e-07,1.933313e-07,1.933315e-07,1.933317e-07,1.933319e-07,1.933321e-07,1.933323e-07,1.933326e-07,1.933328e-07,1.933330e-07,1.933332e-07,1.933334e-07,1.933336e-07,1.933338e-07,1.933340e-07,1.933342e-07,1.933344e-07,1.933346e-07,1.933348e-07,1.933350e-07,1.933352e-07,1.933354e-07,1.933357e-07,1.933359e-07,1.933361e-07,1.933363e-07,1.933365e-07,1.933367e-07,1.933369e-07,1.933371e-07,1.933373e-07,1.933375e-07,1.933377e-07,1.933379e-07,1.933381e-07,1.933383e-07,1.933385e-07,1.933387e-07,1.933390e-07,1.933392e-07,1.933394e-07,1.933396e-07,1.933398e-07,1.933400e-07,1.933402e-07,1.933404e-07,1.933406e-07,1.933408e-07,1.933410e-07,1.933412e-07,1.933414e-07,1.933416e-07,1.933418e-07,1.933420e-07,1.933423e-07,1.933425e-07,1.933427e-07,1.933429e-07,1.933431e-07,1.933433e-07,1.933435e-07,1.933437e-07,1.933439e-07,1.933441e-07,1.933443e-07,1.933445e-07,1.933447e-07,1.933449e-07,1.933451e-07,1.933453e-07,1.933456e-07,1.933458e-07,1.933460e-07,1.933462e-07,1.933464e-07,1.933466e-07,1.933468e-07,1.933470e-07,1.933472e-07,1.933474e-07,1.933476e-07,1.933478e-07,1.933480e-07,1.933482e-07,1.933484e-07,1.933486e-07,1.933489e-07,1.933491e-07,1.933493e-07,1.933495e-07,1.933497e-07,1.933499e-07,1.933501e-07,1.933503e-07,1.933505e-07,1.933507e-07,1.933509e-07,1.933511e-07,1.933513e-07,1.933515e-07,1.933517e-07,1.933519e-07,1.933521e-07,1.933524e-07,1.933526e-07,1.933528e-07,1.933530e-07,1.933532e-07,1.933534e-07,1.933536e-07,1.933538e-07,1.933540e-07,1.933542e-07,1.933544e-07,1.933546e-07,1.933548e-07,1.933550e-07,1.933552e-07,1.933554e-07,1.933557e-07,1.933559e-07,1.933561e-07,1.933563e-07,1.933565e-07,1.933567e-07,1.933569e-07,1.933571e-07,1.933573e-07,1.933575e-07,1.933577e-07,1.933579e-07,1.933581e-07,1.933583e-07,1.933585e-07,1.933587e-07,1.933589e-07,1.933592e-07,1.933594e-07,1.933596e-07,1.933598e-07,1.933600e-07,1.933602e-07,1.933604e-07,1.933606e-07,1.933608e-07,1.933610e-07,1.933612e-07,1.933614e-07,1.933616e-07,1.933618e-07,1.933620e-07,1.933622e-07,1.933625e-07,1.933627e-07,1.933629e-07,1.933631e-07,1.933633e-07,1.933635e-07,1.933637e-07,1.933639e-07,1.933641e-07,1.933643e-07,1.933645e-07,1.933647e-07,1.933649e-07,1.933651e-07,1.933653e-07,1.933655e-07,1.933657e-07,1.933660e-07,1.933662e-07,1.933664e-07,1.933666e-07,1.933668e-07,1.933670e-07,1.933672e-07,1.933674e-07,1.933676e-07,1.933678e-07,1.933680e-07,1.933682e-07,1.933684e-07,1.933686e-07,1.933688e-07,1.933690e-07,1.933692e-07,1.933694e-07,1.933697e-07,1.933699e-07,1.933701e-07,1.933703e-07,1.933705e-07,1.933707e-07,1.933709e-07,1.933711e-07,1.933713e-07,1.933715e-07,1.933717e-07,1.933719e-07,1.933721e-07,1.933723e-07,1.933725e-07,1.933727e-07,1.933729e-07,1.933732e-07,1.933734e-07,1.933736e-07,1.933738e-07,1.933740e-07,1.933742e-07,1.933744e-07,1.933746e-07,1.933748e-07,1.933750e-07,1.933752e-07,1.933754e-07,1.933756e-07,1.933758e-07,1.933760e-07,1.933762e-07,1.933764e-07,1.933766e-07,1.933769e-07,1.933771e-07,1.933773e-07,1.933775e-07,1.933777e-07,1.933779e-07,1.933781e-07,1.933783e-07,1.933785e-07,1.933787e-07,1.933789e-07,1.933791e-07,1.933793e-07,1.933795e-07,1.933797e-07,1.933799e-07,1.933801e-07,1.933804e-07,1.933806e-07,1.933808e-07,1.933810e-07,1.933812e-07,1.933814e-07,1.933816e-07,1.933818e-07,1.933820e-07,1.933822e-07,1.933824e-07,1.933826e-07,1.933828e-07,1.933830e-07,1.933832e-07,1.933834e-07,1.933836e-07,1.933838e-07,1.933841e-07,1.933843e-07,1.933845e-07,1.933847e-07,1.933849e-07,1.933851e-07,1.933853e-07,1.933855e-07,1.933857e-07,1.933859e-07,1.933861e-07,1.933863e-07,1.933865e-07,1.933867e-07,1.933869e-07,1.933871e-07,1.933873e-07,1.933875e-07,1.933877e-07,1.933880e-07,1.933882e-07,1.933884e-07,1.933886e-07,1.933888e-07,1.933890e-07,1.933892e-07,1.933894e-07,1.933896e-07,1.933898e-07,1.933900e-07,1.933902e-07,1.933904e-07,1.933906e-07,1.933908e-07,1.933910e-07,1.933912e-07,1.933914e-07,1.933917e-07,1.933919e-07,1.933921e-07,1.933923e-07,1.933925e-07,1.933927e-07,1.933929e-07,1.933931e-07,1.933933e-07,1.933935e-07,1.933937e-07,1.933939e-07,1.933941e-07,1.933943e-07,1.933945e-07,1.933947e-07,1.933949e-07,1.933951e-07,1.933953e-07,1.933956e-07,1.933958e-07,1.933960e-07,1.933962e-07,1.933964e-07,1.933966e-07,1.933968e-07,1.933970e-07,1.933972e-07,1.933974e-07,1.933976e-07,1.933978e-07,1.933980e-07,1.933982e-07,1.933984e-07,1.933986e-07,1.933988e-07,1.933990e-07,1.933993e-07,1.933995e-07,1.933997e-07,1.933999e-07,1.934001e-07,1.934003e-07,1.934005e-07,1.934007e-07,1.934009e-07,1.934011e-07,1.934013e-07,1.934015e-07,1.934017e-07,1.934019e-07,1.934021e-07,1.934023e-07,1.934025e-07,1.934027e-07,1.934029e-07,1.934031e-07,1.934034e-07,1.934036e-07,1.934038e-07,1.934040e-07,1.934042e-07,1.934044e-07,1.934046e-07,1.934048e-07,1.934050e-07,1.934052e-07,1.934054e-07,1.934056e-07,1.934058e-07,1.934060e-07,1.934062e-07,1.934064e-07,1.934066e-07,1.934068e-07,1.934070e-07,1.934073e-07,1.934075e-07,1.934077e-07,1.934079e-07,1.934081e-07,1.934083e-07,1.934085e-07,1.934087e-07,1.934089e-07,1.934091e-07,1.934093e-07,1.934095e-07,1.934097e-07,1.934099e-07,1.934101e-07,1.934103e-07,1.934105e-07,1.934107e-07,1.934109e-07,1.934111e-07,1.934114e-07,1.934116e-07,1.934118e-07,1.934120e-07,1.934122e-07,1.934124e-07,1.934126e-07,1.934128e-07,1.934130e-07,1.934132e-07,1.934134e-07,1.934136e-07,1.934138e-07,1.934140e-07,1.934142e-07,1.934144e-07,1.934146e-07,1.934148e-07,1.934150e-07,1.934153e-07,1.934155e-07,1.934157e-07,1.934159e-07,1.934161e-07,1.934163e-07,1.934165e-07,1.934167e-07,1.934169e-07,1.934171e-07,1.934173e-07,1.934175e-07,1.934177e-07,1.934179e-07,1.934181e-07,1.934183e-07,1.934185e-07,1.934187e-07,1.934189e-07,1.934191e-07,1.934193e-07,1.934196e-07,1.934198e-07,1.934200e-07,1.934202e-07,1.934204e-07,1.934206e-07,1.934208e-07,1.934210e-07,1.934212e-07,1.934214e-07,1.934216e-07,1.934218e-07,1.934220e-07,1.934222e-07,1.934224e-07,1.934226e-07,1.934228e-07,1.934230e-07,1.934232e-07,1.934234e-07,1.934237e-07,1.934239e-07,1.934241e-07,1.934243e-07,1.934245e-07,1.934247e-07,1.934249e-07,1.934251e-07,1.934253e-07,1.934255e-07,1.934257e-07,1.934259e-07,1.934261e-07,1.934263e-07,1.934265e-07,1.934267e-07,1.934269e-07,1.934271e-07,1.934273e-07,1.934275e-07,1.934277e-07,1.934280e-07,1.934282e-07,1.934284e-07,1.934286e-07,1.934288e-07,1.934290e-07,1.934292e-07,1.934294e-07,1.934296e-07,1.934298e-07,1.934300e-07,1.934302e-07,1.934304e-07,1.934306e-07,1.934308e-07,1.934310e-07,1.934312e-07,1.934314e-07,1.934316e-07,1.934318e-07,1.934320e-07,1.934323e-07,1.934325e-07,1.934327e-07,1.934329e-07,1.934331e-07,1.934333e-07,1.934335e-07,1.934337e-07,1.934339e-07,1.934341e-07,1.934343e-07,1.934345e-07,1.934347e-07,1.934349e-07,1.934351e-07,1.934353e-07,1.934355e-07,1.934357e-07,1.934359e-07,1.934361e-07,1.934363e-07,1.934365e-07,1.934368e-07,1.934370e-07,1.934372e-07,1.934374e-07,1.934376e-07,1.934378e-07,1.934380e-07,1.934382e-07,1.934384e-07,1.934386e-07,1.934388e-07,1.934390e-07,1.934392e-07,1.934394e-07,1.934396e-07,1.934398e-07,1.934400e-07,1.934402e-07,1.934404e-07,1.934406e-07,1.934408e-07,1.934410e-07,1.934413e-07,1.934415e-07,1.934417e-07,1.934419e-07,1.934421e-07,1.934423e-07,1.934425e-07,1.934427e-07,1.934429e-07,1.934431e-07,1.934433e-07,1.934435e-07,1.934437e-07,1.934439e-07,1.934441e-07,1.934443e-07,1.934445e-07,1.934447e-07,1.934449e-07,1.934451e-07,1.934453e-07,1.934455e-07,1.934458e-07,1.934460e-07,1.934462e-07,1.934464e-07,1.934466e-07,1.934468e-07,1.934470e-07,1.934472e-07,1.934474e-07,1.934476e-07,1.934478e-07,1.934480e-07,1.934482e-07,1.934484e-07,1.934486e-07,1.934488e-07,1.934490e-07,1.934492e-07,1.934494e-07,1.934496e-07,1.934498e-07,1.934500e-07,1.934503e-07,1.934505e-07,1.934507e-07,1.934509e-07,1.934511e-07,1.934513e-07,1.934515e-07,1.934517e-07,1.934519e-07,1.934521e-07,1.934523e-07,1.934525e-07,1.934527e-07,1.934529e-07,1.934531e-07,1.934533e-07,1.934535e-07,1.934537e-07,1.934539e-07,1.934541e-07,1.934543e-07,1.934545e-07,1.934547e-07,1.934549e-07,1.934552e-07,1.934554e-07,1.934556e-07,1.934558e-07,1.934560e-07,1.934562e-07,1.934564e-07,1.934566e-07,1.934568e-07,1.934570e-07,1.934572e-07,1.934574e-07,1.934576e-07,1.934578e-07,1.934580e-07,1.934582e-07,1.934584e-07,1.934586e-07,1.934588e-07,1.934590e-07,1.934592e-07,1.934594e-07,1.934596e-07,1.934599e-07,1.934601e-07,1.934603e-07,1.934605e-07,1.934607e-07,1.934609e-07,1.934611e-07,1.934613e-07,1.934615e-07,1.934617e-07,1.934619e-07,1.934621e-07,1.934623e-07,1.934625e-07,1.934627e-07,1.934629e-07,1.934631e-07,1.934633e-07,1.934635e-07,1.934637e-07,1.934639e-07,1.934641e-07,1.934643e-07,1.934645e-07,1.934648e-07,1.934650e-07,1.934652e-07,1.934654e-07,1.934656e-07,1.934658e-07,1.934660e-07,1.934662e-07,1.934664e-07,1.934666e-07,1.934668e-07,1.934670e-07,1.934672e-07,1.934674e-07,1.934676e-07,1.934678e-07,1.934680e-07,1.934682e-07,1.934684e-07,1.934686e-07,1.934688e-07,1.934690e-07,1.934692e-07,1.934694e-07,1.934696e-07,1.934699e-07,1.934701e-07,1.934703e-07,1.934705e-07,1.934707e-07,1.934709e-07,1.934711e-07,1.934713e-07,1.934715e-07,1.934717e-07,1.934719e-07,1.934721e-07,1.934723e-07,1.934725e-07,1.934727e-07,1.934729e-07,1.934731e-07,1.934733e-07,1.934735e-07,1.934737e-07,1.934739e-07,1.934741e-07,1.934743e-07,1.934745e-07,1.934747e-07,1.934750e-07,1.934752e-07,1.934754e-07,1.934756e-07,1.934758e-07,1.934760e-07,1.934762e-07,1.934764e-07,1.934766e-07,1.934768e-07,1.934770e-07,1.934772e-07,1.934774e-07,1.934776e-07,1.934778e-07,1.934780e-07,1.934782e-07,1.934784e-07,1.934786e-07,1.934788e-07,1.934790e-07,1.934792e-07,1.934794e-07,1.934796e-07,1.934798e-07,1.934801e-07,1.934803e-07,1.934805e-07,1.934807e-07,1.934809e-07,1.934811e-07,1.934813e-07,1.934815e-07,1.934817e-07,1.934819e-07,1.934821e-07,1.934823e-07,1.934825e-07,1.934827e-07,1.934829e-07,1.934831e-07,1.934833e-07,1.934835e-07,1.934837e-07,1.934839e-07,1.934841e-07,1.934843e-07,1.934845e-07,1.934847e-07,1.934849e-07,1.934851e-07,1.934853e-07,1.934856e-07,1.934858e-07,1.934860e-07,1.934862e-07,1.934864e-07,1.934866e-07,1.934868e-07,1.934870e-07,1.934872e-07,1.934874e-07,1.934876e-07,1.934878e-07,1.934880e-07,1.934882e-07,1.934884e-07,1.934886e-07,1.934888e-07,1.934890e-07,1.934892e-07,1.934894e-07,1.934896e-07,1.934898e-07,1.934900e-07,1.934902e-07,1.934904e-07,1.934906e-07,1.934908e-07,1.934911e-07,1.934913e-07,1.934915e-07,1.934917e-07,1.934919e-07,1.934921e-07,1.934923e-07,1.934925e-07,1.934927e-07,1.934929e-07,1.934931e-07,1.934933e-07,1.934935e-07,1.934937e-07,1.934939e-07,1.934941e-07,1.934943e-07,1.934945e-07,1.934947e-07,1.934949e-07,1.934951e-07,1.934953e-07,1.934955e-07,1.934957e-07,1.934959e-07,1.934961e-07,1.934963e-07,1.934966e-07,1.934968e-07,1.934970e-07,1.934972e-07,1.934974e-07,1.934976e-07,1.934978e-07,1.934980e-07,1.934982e-07,1.934984e-07,1.934986e-07,1.934988e-07,1.934990e-07,1.934992e-07,1.934994e-07,1.934996e-07,1.934998e-07,1.935000e-07,1.935002e-07,1.935004e-07,1.935006e-07,1.935008e-07,1.935010e-07,1.935012e-07,1.935014e-07,1.935016e-07,1.935018e-07,1.935020e-07,1.935022e-07,1.935025e-07,1.935027e-07,1.935029e-07,1.935031e-07,1.935033e-07,1.935035e-07,1.935037e-07,1.935039e-07,1.935041e-07,1.935043e-07,1.935045e-07,1.935047e-07,1.935049e-07,1.935051e-07,1.935053e-07,1.935055e-07,1.935057e-07,1.935059e-07,1.935061e-07,1.935063e-07,1.935065e-07,1.935067e-07,1.935069e-07,1.935071e-07,1.935073e-07,1.935075e-07,1.935077e-07,1.935079e-07,1.935081e-07,1.935084e-07,1.935086e-07,1.935088e-07,1.935090e-07,1.935092e-07,1.935094e-07,1.935096e-07,1.935098e-07,1.935100e-07,1.935102e-07,1.935104e-07,1.935106e-07,1.935108e-07,1.935110e-07,1.935112e-07,1.935114e-07,1.935116e-07,1.935118e-07,1.935120e-07,1.935122e-07,1.935124e-07,1.935126e-07,1.935128e-07,1.935130e-07,1.935132e-07,1.935134e-07,1.935136e-07,1.935138e-07,1.935140e-07,1.935142e-07,1.935145e-07,1.935147e-07,1.935149e-07,1.935151e-07,1.935153e-07,1.935155e-07,1.935157e-07,1.935159e-07,1.935161e-07,1.935163e-07,1.935165e-07,1.935167e-07,1.935169e-07,1.935171e-07,1.935173e-07,1.935175e-07,1.935177e-07,1.935179e-07,1.935181e-07,1.935183e-07,1.935185e-07,1.935187e-07,1.935189e-07,1.935191e-07,1.935193e-07,1.935195e-07,1.935197e-07,1.935199e-07,1.935201e-07,1.935203e-07,1.935205e-07,1.935208e-07,1.935210e-07,1.935212e-07,1.935214e-07,1.935216e-07,1.935218e-07,1.935220e-07,1.935222e-07,1.935224e-07,1.935226e-07,1.935228e-07,1.935230e-07,1.935232e-07,1.935234e-07,1.935236e-07,1.935238e-07,1.935240e-07,1.935242e-07,1.935244e-07,1.935246e-07,1.935248e-07,1.935250e-07,1.935252e-07,1.935254e-07,1.935256e-07,1.935258e-07,1.935260e-07,1.935262e-07,1.935264e-07,1.935266e-07,1.935268e-07,1.935270e-07,1.935272e-07,1.935275e-07,1.935277e-07,1.935279e-07,1.935281e-07,1.935283e-07,1.935285e-07,1.935287e-07,1.935289e-07,1.935291e-07,1.935293e-07,1.935295e-07,1.935297e-07,1.935299e-07,1.935301e-07,1.935303e-07,1.935305e-07,1.935307e-07,1.935309e-07,1.935311e-07,1.935313e-07,1.935315e-07,1.935317e-07,1.935319e-07,1.935321e-07,1.935323e-07,1.935325e-07,1.935327e-07,1.935329e-07,1.935331e-07,1.935333e-07,1.935335e-07,1.935337e-07,1.935339e-07,1.935342e-07,1.935344e-07,1.935346e-07,1.935348e-07,1.935350e-07,1.935352e-07,1.935354e-07,1.935356e-07,1.935358e-07,1.935360e-07,1.935362e-07,1.935364e-07,1.935366e-07,1.935368e-07,1.935370e-07,1.935372e-07,1.935374e-07,1.935376e-07,1.935378e-07,1.935380e-07,1.935382e-07,1.935384e-07,1.935386e-07,1.935388e-07,1.935390e-07,1.935392e-07,1.935394e-07,1.935396e-07,1.935398e-07,1.935400e-07,1.935402e-07,1.935404e-07,1.935406e-07,1.935408e-07,1.935410e-07,1.935412e-07,1.935415e-07,1.935417e-07,1.935419e-07,1.935421e-07,1.935423e-07,1.935425e-07,1.935427e-07,1.935429e-07,1.935431e-07,1.935433e-07,1.935435e-07,1.935437e-07,1.935439e-07,1.935441e-07,1.935443e-07,1.935445e-07,1.935447e-07,1.935449e-07,1.935451e-07,1.935453e-07,1.935455e-07,1.935457e-07,1.935459e-07,1.935461e-07,1.935463e-07,1.935465e-07,1.935467e-07,1.935469e-07,1.935471e-07,1.935473e-07,1.935475e-07,1.935477e-07,1.935479e-07,1.935481e-07,1.935483e-07,1.935485e-07,1.935488e-07,1.935490e-07,1.935492e-07,1.935494e-07,1.935496e-07,1.935498e-07,1.935500e-07,1.935502e-07,1.935504e-07,1.935506e-07,1.935508e-07,1.935510e-07,1.935512e-07,1.935514e-07,1.935516e-07,1.935518e-07,1.935520e-07,1.935522e-07,1.935524e-07,1.935526e-07,1.935528e-07,1.935530e-07,1.935532e-07,1.935534e-07,1.935536e-07,1.935538e-07,1.935540e-07,1.935542e-07,1.935544e-07,1.935546e-07,1.935548e-07,1.935550e-07,1.935552e-07,1.935554e-07,1.935556e-07,1.935558e-07,1.935560e-07,1.935562e-07,1.935564e-07,1.935567e-07,1.935569e-07,1.935571e-07,1.935573e-07,1.935575e-07,1.935577e-07,1.935579e-07,1.935581e-07,1.935583e-07,1.935585e-07,1.935587e-07,1.935589e-07,1.935591e-07,1.935593e-07,1.935595e-07,1.935597e-07,1.935599e-07,1.935601e-07,1.935603e-07,1.935605e-07,1.935607e-07,1.935609e-07,1.935611e-07,1.935613e-07,1.935615e-07,1.935617e-07,1.935619e-07,1.935621e-07,1.935623e-07,1.935625e-07,1.935627e-07,1.935629e-07,1.935631e-07,1.935633e-07,1.935635e-07,1.935637e-07,1.935639e-07,1.935641e-07,1.935643e-07,1.935645e-07,1.935647e-07,1.935650e-07,1.935652e-07,1.935654e-07,1.935656e-07,1.935658e-07,1.935660e-07,1.935662e-07,1.935664e-07,1.935666e-07,1.935668e-07,1.935670e-07,1.935672e-07,1.935674e-07,1.935676e-07,1.935678e-07,1.935680e-07,1.935682e-07,1.935684e-07,1.935686e-07,1.935688e-07,1.935690e-07,1.935692e-07,1.935694e-07,1.935696e-07,1.935698e-07,1.935700e-07,1.935702e-07,1.935704e-07,1.935706e-07,1.935708e-07,1.935710e-07,1.935712e-07,1.935714e-07,1.935716e-07,1.935718e-07,1.935720e-07,1.935722e-07,1.935724e-07,1.935726e-07,1.935728e-07,1.935730e-07,1.935732e-07,1.935734e-07,1.935737e-07,1.935739e-07,1.935741e-07,1.935743e-07,1.935745e-07,1.935747e-07,1.935749e-07,1.935751e-07,1.935753e-07,1.935755e-07,1.935757e-07,1.935759e-07,1.935761e-07,1.935763e-07,1.935765e-07,1.935767e-07,1.935769e-07,1.935771e-07,1.935773e-07,1.935775e-07,1.935777e-07,1.935779e-07,1.935781e-07,1.935783e-07,1.935785e-07,1.935787e-07,1.935789e-07,1.935791e-07,1.935793e-07,1.935795e-07,1.935797e-07,1.935799e-07,1.935801e-07,1.935803e-07,1.935805e-07,1.935807e-07,1.935809e-07,1.935811e-07,1.935813e-07,1.935815e-07,1.935817e-07,1.935819e-07,1.935821e-07,1.935823e-07,1.935825e-07,1.935827e-07,1.935830e-07,1.935832e-07,1.935834e-07,1.935836e-07,1.935838e-07,1.935840e-07,1.935842e-07,1.935844e-07,1.935846e-07,1.935848e-07,1.935850e-07,1.935852e-07,1.935854e-07,1.935856e-07,1.935858e-07,1.935860e-07,1.935862e-07,1.935864e-07,1.935866e-07,1.935868e-07,1.935870e-07,1.935872e-07,1.935874e-07,1.935876e-07,1.935878e-07,1.935880e-07,1.935882e-07,1.935884e-07,1.935886e-07,1.935888e-07,1.935890e-07,1.935892e-07,1.935894e-07,1.935896e-07,1.935898e-07,1.935900e-07,1.935902e-07,1.935904e-07,1.935906e-07,1.935908e-07,1.935910e-07,1.935912e-07,1.935914e-07,1.935916e-07,1.935918e-07,1.935920e-07,1.935922e-07,1.935924e-07,1.935926e-07,1.935928e-07,1.935930e-07,1.935933e-07,1.935935e-07,1.935937e-07,1.935939e-07,1.935941e-07,1.935943e-07,1.935945e-07,1.935947e-07,1.935949e-07,1.935951e-07,1.935953e-07,1.935955e-07,1.935957e-07,1.935959e-07,1.935961e-07,1.935963e-07,1.935965e-07,1.935967e-07,1.935969e-07,1.935971e-07,1.935973e-07,1.935975e-07,1.935977e-07,1.935979e-07,1.935981e-07,1.935983e-07,1.935985e-07,1.935987e-07,1.935989e-07,1.935991e-07,1.935993e-07,1.935995e-07,1.935997e-07,1.935999e-07,1.936001e-07,1.936003e-07,1.936005e-07,1.936007e-07,1.936009e-07,1.936011e-07,1.936013e-07,1.936015e-07,1.936017e-07,1.936019e-07,1.936021e-07,1.936023e-07,1.936025e-07,1.936027e-07,1.936029e-07,1.936031e-07,1.936033e-07,1.936035e-07,1.936037e-07,1.936039e-07,1.936041e-07,1.936043e-07,1.936046e-07,1.936048e-07,1.936050e-07,1.936052e-07,1.936054e-07,1.936056e-07,1.936058e-07,1.936060e-07,1.936062e-07,1.936064e-07,1.936066e-07,1.936068e-07,1.936070e-07,1.936072e-07,1.936074e-07,1.936076e-07,1.936078e-07,1.936080e-07,1.936082e-07,1.936084e-07,1.936086e-07,1.936088e-07,1.936090e-07,1.936092e-07,1.936094e-07,1.936096e-07,1.936098e-07,1.936100e-07,1.936102e-07,1.936104e-07,1.936106e-07,1.936108e-07,1.936110e-07,1.936112e-07,1.936114e-07,1.936116e-07,1.936118e-07,1.936120e-07,1.936122e-07,1.936124e-07,1.936126e-07,1.936128e-07,1.936130e-07,1.936132e-07,1.936134e-07,1.936136e-07,1.936138e-07,1.936140e-07,1.936142e-07,1.936144e-07,1.936146e-07,1.936148e-07,1.936150e-07,1.936152e-07,1.936154e-07,1.936156e-07,1.936158e-07,1.936160e-07,1.936162e-07,1.936164e-07,1.936166e-07,1.936168e-07,1.936171e-07,1.936173e-07,1.936175e-07,1.936177e-07,1.936179e-07,1.936181e-07,1.936183e-07,1.936185e-07,1.936187e-07,1.936189e-07,1.936191e-07,1.936193e-07,1.936195e-07,1.936197e-07,1.936199e-07,1.936201e-07,1.936203e-07,1.936205e-07,1.936207e-07,1.936209e-07,1.936211e-07,1.936213e-07,1.936215e-07,1.936217e-07,1.936219e-07,1.936221e-07,1.936223e-07,1.936225e-07,1.936227e-07,1.936229e-07,1.936231e-07,1.936233e-07,1.936235e-07,1.936237e-07,1.936239e-07,1.936241e-07,1.936243e-07,1.936245e-07,1.936247e-07,1.936249e-07,1.936251e-07,1.936253e-07,1.936255e-07,1.936257e-07,1.936259e-07,1.936261e-07,1.936263e-07,1.936265e-07,1.936267e-07,1.936269e-07,1.936271e-07,1.936273e-07,1.936275e-07,1.936277e-07,1.936279e-07,1.936281e-07,1.936283e-07,1.936285e-07,1.936287e-07,1.936289e-07,1.936291e-07,1.936293e-07,1.936295e-07,1.936297e-07,1.936299e-07,1.936301e-07,1.936303e-07,1.936305e-07,1.936307e-07,1.936309e-07,1.936311e-07,1.936313e-07,1.936315e-07,1.936317e-07,1.936320e-07,1.936322e-07,1.936324e-07,1.936326e-07,1.936328e-07,1.936330e-07,1.936332e-07,1.936334e-07,1.936336e-07,1.936338e-07,1.936340e-07,1.936342e-07,1.936344e-07,1.936346e-07,1.936348e-07,1.936350e-07,1.936352e-07,1.936354e-07,1.936356e-07,1.936358e-07,1.936360e-07,1.936362e-07,1.936364e-07,1.936366e-07,1.936368e-07,1.936370e-07,1.936372e-07,1.936374e-07,1.936376e-07,1.936378e-07,1.936380e-07,1.936382e-07,1.936384e-07,1.936386e-07,1.936388e-07,1.936390e-07,1.936392e-07,1.936394e-07,1.936396e-07,1.936398e-07,1.936400e-07,1.936402e-07,1.936404e-07,1.936406e-07,1.936408e-07,1.936410e-07,1.936412e-07,1.936414e-07,1.936416e-07,1.936418e-07,1.936420e-07,1.936422e-07,1.936424e-07,1.936426e-07,1.936428e-07,1.936430e-07,1.936432e-07,1.936434e-07,1.936436e-07,1.936438e-07,1.936440e-07,1.936442e-07,1.936444e-07,1.936446e-07,1.936448e-07,1.936450e-07,1.936452e-07,1.936454e-07,1.936456e-07,1.936458e-07,1.936460e-07,1.936462e-07,1.936464e-07,1.936466e-07,1.936468e-07,1.936470e-07,1.936472e-07,1.936474e-07,1.936476e-07,1.936478e-07,1.936480e-07,1.936482e-07,1.936484e-07,1.936486e-07,1.936488e-07,1.936490e-07,1.936492e-07,1.936494e-07,1.936496e-07,1.936498e-07,1.936500e-07,1.936502e-07,1.936504e-07,1.936506e-07,1.936508e-07,1.936511e-07,1.936513e-07,1.936515e-07,1.936517e-07,1.936519e-07,1.936521e-07,1.936523e-07,1.936525e-07,1.936527e-07,1.936529e-07,1.936531e-07,1.936533e-07,1.936535e-07,1.936537e-07,1.936539e-07,1.936541e-07,1.936543e-07,1.936545e-07,1.936547e-07,1.936549e-07,1.936551e-07,1.936553e-07,1.936555e-07,1.936557e-07,1.936559e-07,1.936561e-07,1.936563e-07,1.936565e-07,1.936567e-07,1.936569e-07,1.936571e-07,1.936573e-07,1.936575e-07,1.936577e-07,1.936579e-07,1.936581e-07,1.936583e-07,1.936585e-07,1.936587e-07,1.936589e-07,1.936591e-07,1.936593e-07,1.936595e-07,1.936597e-07,1.936599e-07,1.936601e-07,1.936603e-07,1.936605e-07,1.936607e-07,1.936609e-07,1.936611e-07,1.936613e-07,1.936615e-07,1.936617e-07,1.936619e-07,1.936621e-07,1.936623e-07,1.936625e-07,1.936627e-07,1.936629e-07,1.936631e-07,1.936633e-07,1.936635e-07,1.936637e-07,1.936639e-07,1.936641e-07,1.936643e-07,1.936645e-07,1.936647e-07,1.936649e-07,1.936651e-07,1.936653e-07,1.936655e-07,1.936657e-07,1.936659e-07,1.936661e-07,1.936663e-07,1.936665e-07,1.936667e-07,1.936669e-07,1.936671e-07,1.936673e-07,1.936675e-07,1.936677e-07,1.936679e-07,1.936681e-07,1.936683e-07,1.936685e-07,1.936687e-07,1.936689e-07,1.936691e-07,1.936693e-07,1.936695e-07,1.936697e-07,1.936699e-07,1.936701e-07,1.936703e-07,1.936705e-07,1.936707e-07,1.936709e-07,1.936711e-07,1.936713e-07,1.936715e-07,1.936717e-07,1.936719e-07,1.936721e-07,1.936723e-07,1.936725e-07,1.936727e-07,1.936729e-07,1.936731e-07,1.936733e-07,1.936735e-07,1.936737e-07,1.936739e-07,1.936741e-07,1.936743e-07,1.936745e-07,1.936747e-07,1.936749e-07,1.936751e-07,1.936753e-07,1.936755e-07,1.936757e-07,1.936759e-07,1.936761e-07,1.936763e-07,1.936765e-07,1.936767e-07,1.936769e-07,1.936771e-07,1.936773e-07,1.936775e-07,1.936777e-07,1.936779e-07,1.936781e-07,1.936783e-07,1.936785e-07,1.936787e-07,1.936789e-07,1.936791e-07,1.936793e-07,1.936795e-07,1.936797e-07,1.936799e-07,1.936801e-07,1.936803e-07,1.936805e-07,1.936807e-07,1.936809e-07,1.936811e-07,1.936813e-07,1.936815e-07,1.936817e-07,1.936819e-07,1.936821e-07,1.936823e-07,1.936825e-07,1.936827e-07,1.936829e-07,1.936832e-07,1.936834e-07,1.936836e-07,1.936838e-07,1.936840e-07,1.936842e-07,1.936844e-07,1.936846e-07,1.936848e-07,1.936850e-07,1.936852e-07,1.936854e-07,1.936856e-07,1.936858e-07,1.936860e-07,1.936862e-07,1.936864e-07,1.936866e-07,1.936868e-07,1.936870e-07,1.936872e-07,1.936874e-07,1.936876e-07,1.936878e-07,1.936880e-07,1.936882e-07,1.936884e-07,1.936886e-07,1.936888e-07,1.936890e-07,1.936892e-07,1.936894e-07,1.936896e-07,1.936898e-07,1.936900e-07,1.936902e-07,1.936904e-07,1.936906e-07,1.936908e-07,1.936910e-07,1.936912e-07,1.936914e-07,1.936916e-07,1.936918e-07,1.936920e-07,1.936922e-07,1.936924e-07,1.936926e-07,1.936928e-07,1.936930e-07,1.936932e-07,1.936934e-07,1.936936e-07,1.936938e-07,1.936940e-07,1.936942e-07,1.936944e-07,1.936946e-07,1.936948e-07,1.936950e-07,1.936952e-07,1.936954e-07,1.936956e-07,1.936958e-07,1.936960e-07,1.936962e-07,1.936964e-07,1.936966e-07,1.936968e-07,1.936970e-07,1.936972e-07,1.936974e-07,1.936976e-07,1.936978e-07,1.936980e-07,1.936982e-07,1.936984e-07,1.936986e-07,1.936988e-07,1.936990e-07,1.936992e-07,1.936994e-07,1.936996e-07,1.936998e-07,1.937000e-07,1.937002e-07,1.937004e-07,1.937006e-07,1.937008e-07,1.937010e-07,1.937012e-07,1.937014e-07,1.937016e-07,1.937018e-07,1.937020e-07,1.937022e-07,1.937024e-07,1.937026e-07,1.937028e-07,1.937030e-07,1.937032e-07,1.937034e-07,1.937036e-07,1.937038e-07,1.937040e-07,1.937042e-07,1.937044e-07,1.937046e-07,1.937048e-07,1.937050e-07,1.937052e-07,1.937054e-07,1.937056e-07,1.937058e-07,1.937060e-07,1.937062e-07,1.937064e-07,1.937066e-07,1.937068e-07,1.937070e-07,1.937072e-07,1.937074e-07,1.937076e-07,1.937078e-07,1.937080e-07,1.937082e-07,1.937084e-07,1.937086e-07,1.937088e-07,1.937090e-07,1.937092e-07,1.937094e-07,1.937096e-07,1.937098e-07,1.937100e-07,1.937102e-07,1.937104e-07,1.937106e-07,1.937108e-07,1.937110e-07,1.937112e-07,1.937114e-07,1.937116e-07,1.937118e-07,1.937120e-07,1.937122e-07,1.937124e-07,1.937126e-07,1.937128e-07,1.937130e-07,1.937132e-07,1.937134e-07,1.937136e-07,1.937138e-07,1.937140e-07,1.937142e-07,1.937144e-07,1.937146e-07,1.937148e-07,1.937150e-07,1.937152e-07,1.937154e-07,1.937156e-07,1.937158e-07,1.937160e-07,1.937162e-07,1.937164e-07,1.937166e-07,1.937168e-07,1.937170e-07,1.937172e-07,1.937174e-07,1.937176e-07,1.937178e-07,1.937180e-07,1.937182e-07,1.937184e-07,1.937186e-07,1.937188e-07,1.937190e-07,1.937192e-07,1.937194e-07,1.937196e-07,1.937198e-07,1.937200e-07,1.937202e-07,1.937204e-07,1.937206e-07,1.937208e-07,1.937210e-07,1.937212e-07,1.937214e-07,1.937216e-07,1.937218e-07,1.937220e-07,1.937222e-07,1.937224e-07,1.937226e-07,1.937228e-07,1.937230e-07,1.937232e-07,1.937234e-07,1.937236e-07,1.937237e-07,1.937239e-07,1.937241e-07,1.937243e-07,1.937245e-07,1.937247e-07,1.937249e-07,1.937251e-07,1.937253e-07,1.937255e-07,1.937257e-07,1.937259e-07,1.937261e-07,1.937263e-07,1.937265e-07,1.937267e-07,1.937269e-07,1.937271e-07,1.937273e-07,1.937275e-07,1.937277e-07,1.937279e-07,1.937281e-07,1.937283e-07,1.937285e-07,1.937287e-07,1.937289e-07,1.937291e-07,1.937293e-07,1.937295e-07,1.937297e-07,1.937299e-07,1.937301e-07,1.937303e-07,1.937305e-07,1.937307e-07,1.937309e-07,1.937311e-07,1.937313e-07,1.937315e-07,1.937317e-07,1.937319e-07,1.937321e-07,1.937323e-07,1.937325e-07,1.937327e-07,1.937329e-07,1.937331e-07,1.937333e-07,1.937335e-07,1.937337e-07,1.937339e-07,1.937341e-07,1.937343e-07,1.937345e-07,1.937347e-07,1.937349e-07,1.937351e-07,1.937353e-07,1.937355e-07,1.937357e-07,1.937359e-07,1.937361e-07,1.937363e-07,1.937365e-07,1.937367e-07,1.937369e-07,1.937371e-07,1.937373e-07,1.937375e-07,1.937377e-07,1.937379e-07,1.937381e-07,1.937383e-07,1.937385e-07,1.937387e-07,1.937389e-07,1.937391e-07,1.937393e-07,1.937395e-07,1.937397e-07,1.937399e-07,1.937401e-07,1.937403e-07,1.937405e-07,1.937407e-07,1.937409e-07,1.937411e-07,1.937413e-07,1.937415e-07,1.937417e-07,1.937419e-07,1.937421e-07,1.937423e-07,1.937425e-07,1.937427e-07,1.937429e-07,1.937431e-07,1.937433e-07,1.937435e-07,1.937437e-07,1.937439e-07,1.937441e-07,1.937443e-07,1.937445e-07,1.937447e-07,1.937449e-07,1.937451e-07,1.937453e-07,1.937455e-07,1.937457e-07,1.937459e-07,1.937461e-07,1.937463e-07,1.937465e-07,1.937467e-07,1.937469e-07,1.937471e-07,1.937473e-07,1.937475e-07,1.937477e-07,1.937479e-07,1.937481e-07,1.937483e-07,1.937485e-07,1.937487e-07,1.937489e-07,1.937491e-07,1.937493e-07,1.937495e-07,1.937497e-07,1.937499e-07,1.937501e-07,1.937503e-07,1.937505e-07,1.937507e-07,1.937509e-07,1.937511e-07,1.937513e-07,1.937515e-07,1.937517e-07,1.937519e-07,1.937521e-07,1.937523e-07,1.937525e-07,1.937527e-07,1.937529e-07,1.937531e-07,1.937533e-07,1.937535e-07,1.937537e-07,1.937539e-07,1.937541e-07,1.937543e-07,1.937545e-07,1.937547e-07,1.937549e-07,1.937551e-07,1.937553e-07,1.937555e-07,1.937557e-07,1.937558e-07,1.937560e-07,1.937562e-07,1.937564e-07,1.937566e-07,1.937568e-07,1.937570e-07,1.937572e-07,1.937574e-07,1.937576e-07,1.937578e-07,1.937580e-07,1.937582e-07,1.937584e-07,1.937586e-07,1.937588e-07,1.937590e-07,1.937592e-07,1.937594e-07,1.937596e-07,1.937598e-07,1.937600e-07,1.937602e-07,1.937604e-07,1.937606e-07,1.937608e-07,1.937610e-07,1.937612e-07,1.937614e-07,1.937616e-07,1.937618e-07,1.937620e-07,1.937622e-07,1.937624e-07,1.937626e-07,1.937628e-07,1.937630e-07,1.937632e-07,1.937634e-07,1.937636e-07,1.937638e-07,1.937640e-07,1.937642e-07,1.937644e-07,1.937646e-07,1.937648e-07,1.937650e-07,1.937652e-07,1.937654e-07,1.937656e-07,1.937658e-07,1.937660e-07,1.937662e-07,1.937664e-07,1.937666e-07,1.937668e-07,1.937670e-07,1.937672e-07,1.937674e-07,1.937676e-07,1.937678e-07,1.937680e-07,1.937682e-07,1.937684e-07,1.937686e-07,1.937688e-07,1.937690e-07,1.937692e-07,1.937694e-07,1.937696e-07,1.937698e-07,1.937700e-07,1.937702e-07,1.937704e-07,1.937706e-07,1.937708e-07,1.937710e-07,1.937712e-07,1.937714e-07,1.937716e-07,1.937718e-07,1.937720e-07,1.937722e-07,1.937724e-07,1.937726e-07,1.937728e-07,1.937730e-07,1.937732e-07,1.937734e-07,1.937736e-07,1.937738e-07,1.937740e-07,1.937742e-07,1.937744e-07,1.937746e-07,1.937747e-07,1.937749e-07,1.937751e-07,1.937753e-07,1.937755e-07,1.937757e-07,1.937759e-07,1.937761e-07,1.937763e-07,1.937765e-07,1.937767e-07,1.937769e-07,1.937771e-07,1.937773e-07,1.937775e-07,1.937777e-07,1.937779e-07,1.937781e-07,1.937783e-07,1.937785e-07,1.937787e-07,1.937789e-07,1.937791e-07,1.937793e-07,1.937795e-07,1.937797e-07,1.937799e-07,1.937801e-07,1.937803e-07,1.937805e-07,1.937807e-07,1.937809e-07,1.937811e-07,1.937813e-07,1.937815e-07,1.937817e-07,1.937819e-07,1.937821e-07,1.937823e-07,1.937825e-07,1.937827e-07,1.937829e-07,1.937831e-07,1.937833e-07,1.937835e-07,1.937837e-07,1.937839e-07,1.937841e-07,1.937843e-07,1.937845e-07,1.937847e-07,1.937849e-07,1.937851e-07,1.937853e-07,1.937855e-07,1.937857e-07,1.937859e-07,1.937861e-07,1.937863e-07,1.937865e-07,1.937867e-07,1.937869e-07,1.937871e-07,1.937873e-07,1.937875e-07,1.937877e-07,1.937879e-07,1.937881e-07,1.937883e-07,1.937885e-07,1.937887e-07,1.937889e-07,1.937891e-07,1.937893e-07,1.937895e-07,1.937896e-07,1.937898e-07,1.937900e-07,1.937902e-07,1.937904e-07,1.937906e-07,1.937908e-07,1.937910e-07,1.937912e-07,1.937914e-07,1.937916e-07,1.937918e-07,1.937920e-07,1.937922e-07,1.937924e-07,1.937926e-07,1.937928e-07,1.937930e-07,1.937932e-07,1.937934e-07,1.937936e-07,1.937938e-07,1.937940e-07,1.937942e-07,1.937944e-07,1.937946e-07,1.937948e-07,1.937950e-07,1.937952e-07,1.937954e-07,1.937956e-07,1.937958e-07,1.937960e-07,1.937962e-07,1.937964e-07,1.937966e-07,1.937968e-07,1.937970e-07,1.937972e-07,1.937974e-07,1.937976e-07,1.937978e-07,1.937980e-07,1.937982e-07,1.937984e-07,1.937986e-07,1.937988e-07,1.937990e-07,1.937992e-07,1.937994e-07,1.937996e-07,1.937998e-07,1.938000e-07,1.938002e-07,1.938004e-07,1.938006e-07,1.938008e-07,1.938010e-07,1.938012e-07,1.938014e-07,1.938016e-07,1.938018e-07,1.938020e-07,1.938021e-07,1.938023e-07,1.938025e-07,1.938027e-07,1.938029e-07,1.938031e-07,1.938033e-07,1.938035e-07,1.938037e-07,1.938039e-07,1.938041e-07,1.938043e-07,1.938045e-07,1.938047e-07,1.938049e-07,1.938051e-07,1.938053e-07,1.938055e-07,1.938057e-07,1.938059e-07,1.938061e-07,1.938063e-07,1.938065e-07,1.938067e-07,1.938069e-07,1.938071e-07,1.938073e-07,1.938075e-07,1.938077e-07,1.938079e-07,1.938081e-07,1.938083e-07,1.938085e-07,1.938087e-07,1.938089e-07,1.938091e-07,1.938093e-07,1.938095e-07,1.938097e-07,1.938099e-07,1.938101e-07,1.938103e-07,1.938105e-07,1.938107e-07,1.938109e-07,1.938111e-07,1.938113e-07,1.938115e-07,1.938117e-07,1.938119e-07,1.938121e-07,1.938123e-07,1.938125e-07,1.938127e-07,1.938129e-07,1.938131e-07,1.938133e-07,1.938134e-07,1.938136e-07,1.938138e-07,1.938140e-07,1.938142e-07,1.938144e-07,1.938146e-07,1.938148e-07,1.938150e-07,1.938152e-07,1.938154e-07,1.938156e-07,1.938158e-07,1.938160e-07,1.938162e-07,1.938164e-07,1.938166e-07,1.938168e-07,1.938170e-07,1.938172e-07,1.938174e-07,1.938176e-07,1.938178e-07,1.938180e-07,1.938182e-07,1.938184e-07,1.938186e-07,1.938188e-07,1.938190e-07,1.938192e-07,1.938194e-07,1.938196e-07,1.938198e-07,1.938200e-07,1.938202e-07,1.938204e-07,1.938206e-07,1.938208e-07,1.938210e-07,1.938212e-07,1.938214e-07,1.938216e-07,1.938218e-07,1.938220e-07,1.938222e-07,1.938224e-07,1.938226e-07,1.938228e-07,1.938230e-07,1.938232e-07,1.938234e-07,1.938235e-07,1.938237e-07,1.938239e-07,1.938241e-07,1.938243e-07,1.938245e-07,1.938247e-07,1.938249e-07,1.938251e-07,1.938253e-07,1.938255e-07,1.938257e-07,1.938259e-07,1.938261e-07,1.938263e-07,1.938265e-07,1.938267e-07,1.938269e-07,1.938271e-07,1.938273e-07,1.938275e-07,1.938277e-07,1.938279e-07,1.938281e-07,1.938283e-07,1.938285e-07,1.938287e-07,1.938289e-07,1.938291e-07,1.938293e-07,1.938295e-07,1.938297e-07,1.938299e-07,1.938301e-07,1.938303e-07,1.938305e-07,1.938307e-07,1.938309e-07,1.938311e-07,1.938313e-07,1.938315e-07,1.938317e-07,1.938319e-07,1.938321e-07,1.938323e-07,1.938325e-07,1.938327e-07,1.938328e-07,1.938330e-07,1.938332e-07,1.938334e-07,1.938336e-07,1.938338e-07,1.938340e-07,1.938342e-07,1.938344e-07,1.938346e-07,1.938348e-07,1.938350e-07,1.938352e-07,1.938354e-07,1.938356e-07,1.938358e-07,1.938360e-07,1.938362e-07,1.938364e-07,1.938366e-07,1.938368e-07,1.938370e-07,1.938372e-07,1.938374e-07,1.938376e-07,1.938378e-07,1.938380e-07,1.938382e-07,1.938384e-07,1.938386e-07,1.938388e-07,1.938390e-07,1.938392e-07,1.938394e-07,1.938396e-07,1.938398e-07,1.938400e-07,1.938402e-07,1.938404e-07,1.938406e-07,1.938408e-07,1.938410e-07,1.938412e-07,1.938414e-07,1.938415e-07,1.938417e-07,1.938419e-07,1.938421e-07,1.938423e-07,1.938425e-07,1.938427e-07,1.938429e-07,1.938431e-07,1.938433e-07,1.938435e-07,1.938437e-07,1.938439e-07,1.938441e-07,1.938443e-07,1.938445e-07,1.938447e-07,1.938449e-07,1.938451e-07,1.938453e-07,1.938455e-07,1.938457e-07,1.938459e-07,1.938461e-07,1.938463e-07,1.938465e-07,1.938467e-07,1.938469e-07,1.938471e-07,1.938473e-07,1.938475e-07,1.938477e-07,1.938479e-07,1.938481e-07,1.938483e-07,1.938485e-07,1.938487e-07,1.938489e-07,1.938491e-07,1.938493e-07,1.938495e-07,1.938496e-07,1.938498e-07,1.938500e-07,1.938502e-07,1.938504e-07,1.938506e-07,1.938508e-07,1.938510e-07,1.938512e-07,1.938514e-07,1.938516e-07,1.938518e-07,1.938520e-07,1.938522e-07,1.938524e-07,1.938526e-07,1.938528e-07,1.938530e-07,1.938532e-07,1.938534e-07,1.938536e-07,1.938538e-07,1.938540e-07,1.938542e-07,1.938544e-07,1.938546e-07,1.938548e-07,1.938550e-07,1.938552e-07,1.938554e-07,1.938556e-07,1.938558e-07,1.938560e-07,1.938562e-07,1.938564e-07,1.938566e-07,1.938568e-07,1.938570e-07,1.938572e-07,1.938574e-07,1.938575e-07,1.938577e-07,1.938579e-07,1.938581e-07,1.938583e-07,1.938585e-07,1.938587e-07,1.938589e-07,1.938591e-07,1.938593e-07,1.938595e-07,1.938597e-07,1.938599e-07,1.938601e-07,1.938603e-07,1.938605e-07,1.938607e-07,1.938609e-07,1.938611e-07,1.938613e-07,1.938615e-07,1.938617e-07,1.938619e-07,1.938621e-07,1.938623e-07,1.938625e-07,1.938627e-07,1.938629e-07,1.938631e-07,1.938633e-07,1.938635e-07,1.938637e-07,1.938639e-07,1.938641e-07,1.938643e-07,1.938645e-07,1.938647e-07,1.938648e-07,1.938650e-07,1.938652e-07,1.938654e-07,1.938656e-07,1.938658e-07,1.938660e-07,1.938662e-07,1.938664e-07,1.938666e-07,1.938668e-07,1.938670e-07,1.938672e-07,1.938674e-07,1.938676e-07,1.938678e-07,1.938680e-07,1.938682e-07,1.938684e-07,1.938686e-07,1.938688e-07,1.938690e-07,1.938692e-07,1.938694e-07,1.938696e-07,1.938698e-07,1.938700e-07,1.938702e-07,1.938704e-07,1.938706e-07,1.938708e-07,1.938710e-07,1.938712e-07,1.938714e-07,1.938716e-07,1.938718e-07,1.938719e-07,1.938721e-07,1.938723e-07,1.938725e-07,1.938727e-07,1.938729e-07,1.938731e-07,1.938733e-07,1.938735e-07,1.938737e-07,1.938739e-07,1.938741e-07,1.938743e-07,1.938745e-07,1.938747e-07,1.938749e-07,1.938751e-07,1.938753e-07,1.938755e-07,1.938757e-07,1.938759e-07,1.938761e-07,1.938763e-07,1.938765e-07,1.938767e-07,1.938769e-07,1.938771e-07,1.938773e-07,1.938775e-07,1.938777e-07,1.938779e-07,1.938781e-07,1.938783e-07,1.938785e-07,1.938786e-07,1.938788e-07,1.938790e-07,1.938792e-07,1.938794e-07,1.938796e-07,1.938798e-07,1.938800e-07,1.938802e-07,1.938804e-07,1.938806e-07,1.938808e-07,1.938810e-07,1.938812e-07,1.938814e-07,1.938816e-07,1.938818e-07,1.938820e-07,1.938822e-07,1.938824e-07,1.938826e-07,1.938828e-07,1.938830e-07,1.938832e-07,1.938834e-07,1.938836e-07,1.938838e-07,1.938840e-07,1.938842e-07,1.938844e-07,1.938846e-07,1.938848e-07,1.938850e-07,1.938851e-07,1.938853e-07,1.938855e-07,1.938857e-07,1.938859e-07,1.938861e-07,1.938863e-07,1.938865e-07,1.938867e-07,1.938869e-07,1.938871e-07,1.938873e-07,1.938875e-07,1.938877e-07,1.938879e-07,1.938881e-07,1.938883e-07,1.938885e-07,1.938887e-07,1.938889e-07,1.938891e-07,1.938893e-07,1.938895e-07,1.938897e-07,1.938899e-07,1.938901e-07,1.938903e-07,1.938905e-07,1.938907e-07,1.938909e-07,1.938911e-07,1.938913e-07,1.938914e-07,1.938916e-07,1.938918e-07,1.938920e-07,1.938922e-07,1.938924e-07,1.938926e-07,1.938928e-07,1.938930e-07,1.938932e-07,1.938934e-07,1.938936e-07,1.938938e-07,1.938940e-07,1.938942e-07,1.938944e-07,1.938946e-07,1.938948e-07,1.938950e-07,1.938952e-07,1.938954e-07,1.938956e-07,1.938958e-07,1.938960e-07,1.938962e-07,1.938964e-07,1.938966e-07,1.938968e-07,1.938970e-07,1.938972e-07,1.938974e-07,1.938975e-07,1.938977e-07,1.938979e-07,1.938981e-07,1.938983e-07,1.938985e-07,1.938987e-07,1.938989e-07,1.938991e-07,1.938993e-07,1.938995e-07,1.938997e-07,1.938999e-07,1.939001e-07,1.939003e-07,1.939005e-07,1.939007e-07,1.939009e-07,1.939011e-07,1.939013e-07,1.939015e-07,1.939017e-07,1.939019e-07,1.939021e-07,1.939023e-07,1.939025e-07,1.939027e-07,1.939029e-07,1.939031e-07,1.939033e-07,1.939034e-07,1.939036e-07,1.939038e-07,1.939040e-07,1.939042e-07,1.939044e-07,1.939046e-07,1.939048e-07,1.939050e-07,1.939052e-07,1.939054e-07,1.939056e-07,1.939058e-07,1.939060e-07,1.939062e-07,1.939064e-07,1.939066e-07,1.939068e-07,1.939070e-07,1.939072e-07,1.939074e-07,1.939076e-07,1.939078e-07,1.939080e-07,1.939082e-07,1.939084e-07,1.939086e-07,1.939088e-07,1.939090e-07,1.939091e-07,1.939093e-07,1.939095e-07,1.939097e-07,1.939099e-07,1.939101e-07,1.939103e-07,1.939105e-07,1.939107e-07,1.939109e-07,1.939111e-07,1.939113e-07,1.939115e-07,1.939117e-07,1.939119e-07,1.939121e-07,1.939123e-07,1.939125e-07,1.939127e-07,1.939129e-07,1.939131e-07,1.939133e-07,1.939135e-07,1.939137e-07,1.939139e-07,1.939141e-07,1.939143e-07,1.939145e-07,1.939146e-07,1.939148e-07,1.939150e-07,1.939152e-07,1.939154e-07,1.939156e-07,1.939158e-07,1.939160e-07,1.939162e-07,1.939164e-07,1.939166e-07,1.939168e-07,1.939170e-07,1.939172e-07,1.939174e-07,1.939176e-07,1.939178e-07,1.939180e-07,1.939182e-07,1.939184e-07,1.939186e-07,1.939188e-07,1.939190e-07,1.939192e-07,1.939194e-07,1.939196e-07,1.939198e-07,1.939200e-07,1.939201e-07,1.939203e-07,1.939205e-07,1.939207e-07,1.939209e-07,1.939211e-07,1.939213e-07,1.939215e-07,1.939217e-07,1.939219e-07,1.939221e-07,1.939223e-07,1.939225e-07,1.939227e-07,1.939229e-07,1.939231e-07,1.939233e-07,1.939235e-07,1.939237e-07,1.939239e-07,1.939241e-07,1.939243e-07,1.939245e-07,1.939247e-07,1.939249e-07,1.939251e-07,1.939253e-07,1.939254e-07,1.939256e-07,1.939258e-07,1.939260e-07,1.939262e-07,1.939264e-07,1.939266e-07,1.939268e-07,1.939270e-07,1.939272e-07,1.939274e-07,1.939276e-07,1.939278e-07,1.939280e-07,1.939282e-07,1.939284e-07,1.939286e-07,1.939288e-07,1.939290e-07,1.939292e-07,1.939294e-07,1.939296e-07,1.939298e-07,1.939300e-07,1.939302e-07,1.939304e-07,1.939305e-07,1.939307e-07,1.939309e-07,1.939311e-07,1.939313e-07,1.939315e-07,1.939317e-07,1.939319e-07,1.939321e-07,1.939323e-07,1.939325e-07,1.939327e-07,1.939329e-07,1.939331e-07,1.939333e-07,1.939335e-07,1.939337e-07,1.939339e-07,1.939341e-07,1.939343e-07,1.939345e-07,1.939347e-07,1.939349e-07,1.939351e-07,1.939353e-07,1.939355e-07,1.939356e-07,1.939358e-07,1.939360e-07,1.939362e-07,1.939364e-07,1.939366e-07,1.939368e-07,1.939370e-07,1.939372e-07,1.939374e-07,1.939376e-07,1.939378e-07,1.939380e-07,1.939382e-07,1.939384e-07,1.939386e-07,1.939388e-07,1.939390e-07,1.939392e-07,1.939394e-07,1.939396e-07,1.939398e-07,1.939400e-07,1.939402e-07,1.939404e-07,1.939405e-07,1.939407e-07,1.939409e-07,1.939411e-07,1.939413e-07,1.939415e-07,1.939417e-07,1.939419e-07,1.939421e-07,1.939423e-07,1.939425e-07,1.939427e-07,1.939429e-07,1.939431e-07,1.939433e-07,1.939435e-07,1.939437e-07,1.939439e-07,1.939441e-07,1.939443e-07,1.939445e-07,1.939447e-07,1.939449e-07,1.939451e-07,1.939453e-07,1.939454e-07,1.939456e-07,1.939458e-07,1.939460e-07,1.939462e-07,1.939464e-07,1.939466e-07,1.939468e-07,1.939470e-07,1.939472e-07,1.939474e-07,1.939476e-07,1.939478e-07,1.939480e-07,1.939482e-07,1.939484e-07,1.939486e-07,1.939488e-07,1.939490e-07,1.939492e-07,1.939494e-07,1.939496e-07,1.939498e-07,1.939500e-07,1.939501e-07,1.939503e-07,1.939505e-07,1.939507e-07,1.939509e-07,1.939511e-07,1.939513e-07,1.939515e-07,1.939517e-07,1.939519e-07,1.939521e-07,1.939523e-07,1.939525e-07,1.939527e-07,1.939529e-07,1.939531e-07,1.939533e-07,1.939535e-07,1.939537e-07,1.939539e-07,1.939541e-07,1.939543e-07,1.939545e-07,1.939547e-07,1.939548e-07,1.939550e-07,1.939552e-07,1.939554e-07,1.939556e-07,1.939558e-07,1.939560e-07,1.939562e-07,1.939564e-07,1.939566e-07,1.939568e-07,1.939570e-07,1.939572e-07,1.939574e-07,1.939576e-07,1.939578e-07,1.939580e-07,1.939582e-07,1.939584e-07,1.939586e-07,1.939588e-07,1.939590e-07,1.939592e-07,1.939593e-07,1.939595e-07,1.939597e-07,1.939599e-07,1.939601e-07,1.939603e-07,1.939605e-07,1.939607e-07,1.939609e-07,1.939611e-07,1.939613e-07,1.939615e-07,1.939617e-07,1.939619e-07,1.939621e-07,1.939623e-07,1.939625e-07,1.939627e-07,1.939629e-07,1.939631e-07,1.939633e-07,1.939635e-07,1.939637e-07,1.939638e-07,1.939640e-07,1.939642e-07,1.939644e-07,1.939646e-07,1.939648e-07,1.939650e-07,1.939652e-07,1.939654e-07,1.939656e-07,1.939658e-07,1.939660e-07,1.939662e-07,1.939664e-07,1.939666e-07,1.939668e-07,1.939670e-07,1.939672e-07,1.939674e-07,1.939676e-07,1.939678e-07,1.939680e-07,1.939681e-07,1.939683e-07,1.939685e-07,1.939687e-07,1.939689e-07,1.939691e-07,1.939693e-07,1.939695e-07,1.939697e-07,1.939699e-07,1.939701e-07,1.939703e-07,1.939705e-07,1.939707e-07,1.939709e-07,1.939711e-07,1.939713e-07,1.939715e-07,1.939717e-07,1.939719e-07,1.939721e-07,1.939723e-07,1.939725e-07,1.939726e-07,1.939728e-07,1.939730e-07,1.939732e-07,1.939734e-07,1.939736e-07,1.939738e-07,1.939740e-07,1.939742e-07,1.939744e-07,1.939746e-07,1.939748e-07,1.939750e-07,1.939752e-07,1.939754e-07,1.939756e-07,1.939758e-07,1.939760e-07,1.939762e-07,1.939764e-07,1.939766e-07,1.939767e-07,1.939769e-07,1.939771e-07,1.939773e-07,1.939775e-07,1.939777e-07,1.939779e-07,1.939781e-07,1.939783e-07,1.939785e-07,1.939787e-07,1.939789e-07,1.939791e-07,1.939793e-07,1.939795e-07,1.939797e-07,1.939799e-07,1.939801e-07,1.939803e-07,1.939805e-07,1.939807e-07,1.939809e-07,1.939810e-07,1.939812e-07,1.939814e-07,1.939816e-07,1.939818e-07,1.939820e-07,1.939822e-07,1.939824e-07,1.939826e-07,1.939828e-07,1.939830e-07,1.939832e-07,1.939834e-07,1.939836e-07,1.939838e-07,1.939840e-07,1.939842e-07,1.939844e-07,1.939846e-07,1.939848e-07,1.939850e-07,1.939851e-07,1.939853e-07,1.939855e-07,1.939857e-07,1.939859e-07,1.939861e-07,1.939863e-07,1.939865e-07,1.939867e-07,1.939869e-07,1.939871e-07,1.939873e-07,1.939875e-07,1.939877e-07,1.939879e-07,1.939881e-07,1.939883e-07,1.939885e-07,1.939887e-07,1.939889e-07,1.939891e-07,1.939892e-07,1.939894e-07,1.939896e-07,1.939898e-07,1.939900e-07,1.939902e-07,1.939904e-07,1.939906e-07,1.939908e-07,1.939910e-07,1.939912e-07,1.939914e-07,1.939916e-07,1.939918e-07,1.939920e-07,1.939922e-07,1.939924e-07,1.939926e-07,1.939928e-07,1.939930e-07,1.939932e-07,1.939933e-07,1.939935e-07,1.939937e-07,1.939939e-07,1.939941e-07,1.939943e-07,1.939945e-07,1.939947e-07,1.939949e-07,1.939951e-07,1.939953e-07,1.939955e-07,1.939957e-07,1.939959e-07,1.939961e-07,1.939963e-07,1.939965e-07,1.939967e-07,1.939969e-07,1.939971e-07,1.939972e-07,1.939974e-07,1.939976e-07,1.939978e-07,1.939980e-07,1.939982e-07,1.939984e-07,1.939986e-07,1.939988e-07,1.939990e-07,1.939992e-07,1.939994e-07,1.939996e-07,1.939998e-07,1.940000e-07,1.940002e-07,1.940004e-07,1.940006e-07,1.940008e-07,1.940010e-07,1.940011e-07,1.940013e-07,1.940015e-07,1.940017e-07,1.940019e-07,1.940021e-07,1.940023e-07,1.940025e-07,1.940027e-07,1.940029e-07,1.940031e-07,1.940033e-07,1.940035e-07,1.940037e-07,1.940039e-07,1.940041e-07,1.940043e-07,1.940045e-07,1.940047e-07,1.940049e-07,1.940050e-07,1.940052e-07,1.940054e-07,1.940056e-07,1.940058e-07,1.940060e-07,1.940062e-07,1.940064e-07,1.940066e-07,1.940068e-07,1.940070e-07,1.940072e-07,1.940074e-07,1.940076e-07,1.940078e-07,1.940080e-07,1.940082e-07,1.940084e-07,1.940086e-07,1.940087e-07,1.940089e-07,1.940091e-07,1.940093e-07,1.940095e-07,1.940097e-07,1.940099e-07,1.940101e-07,1.940103e-07,1.940105e-07,1.940107e-07,1.940109e-07,1.940111e-07,1.940113e-07,1.940115e-07,1.940117e-07,1.940119e-07,1.940121e-07,1.940123e-07,1.940125e-07,1.940126e-07,1.940128e-07,1.940130e-07,1.940132e-07,1.940134e-07,1.940136e-07,1.940138e-07,1.940140e-07,1.940142e-07,1.940144e-07,1.940146e-07,1.940148e-07,1.940150e-07,1.940152e-07,1.940154e-07,1.940156e-07,1.940158e-07,1.940160e-07,1.940162e-07,1.940163e-07,1.940165e-07,1.940167e-07,1.940169e-07,1.940171e-07,1.940173e-07,1.940175e-07,1.940177e-07,1.940179e-07,1.940181e-07,1.940183e-07,1.940185e-07,1.940187e-07,1.940189e-07,1.940191e-07,1.940193e-07,1.940195e-07,1.940197e-07,1.940198e-07,1.940200e-07,1.940202e-07,1.940204e-07,1.940206e-07,1.940208e-07,1.940210e-07,1.940212e-07,1.940214e-07,1.940216e-07,1.940218e-07,1.940220e-07,1.940222e-07,1.940224e-07,1.940226e-07,1.940228e-07,1.940230e-07,1.940232e-07,1.940234e-07,1.940235e-07,1.940237e-07,1.940239e-07,1.940241e-07,1.940243e-07,1.940245e-07,1.940247e-07,1.940249e-07,1.940251e-07,1.940253e-07,1.940255e-07,1.940257e-07,1.940259e-07,1.940261e-07,1.940263e-07,1.940265e-07,1.940267e-07,1.940269e-07,1.940271e-07,1.940272e-07,1.940274e-07,1.940276e-07,1.940278e-07,1.940280e-07,1.940282e-07,1.940284e-07,1.940286e-07,1.940288e-07,1.940290e-07,1.940292e-07,1.940294e-07,1.940296e-07,1.940298e-07,1.940300e-07,1.940302e-07,1.940304e-07,1.940306e-07,1.940307e-07,1.940309e-07,1.940311e-07,1.940313e-07,1.940315e-07,1.940317e-07,1.940319e-07,1.940321e-07,1.940323e-07,1.940325e-07,1.940327e-07,1.940329e-07,1.940331e-07,1.940333e-07,1.940335e-07,1.940337e-07,1.940339e-07,1.940341e-07,1.940342e-07,1.940344e-07,1.940346e-07,1.940348e-07,1.940350e-07,1.940352e-07,1.940354e-07,1.940356e-07,1.940358e-07,1.940360e-07,1.940362e-07,1.940364e-07,1.940366e-07,1.940368e-07,1.940370e-07,1.940372e-07,1.940374e-07,1.940376e-07,1.940377e-07,1.940379e-07,1.940381e-07,1.940383e-07,1.940385e-07,1.940387e-07,1.940389e-07,1.940391e-07,1.940393e-07,1.940395e-07,1.940397e-07,1.940399e-07,1.940401e-07,1.940403e-07,1.940405e-07,1.940407e-07,1.940409e-07,1.940410e-07,1.940412e-07,1.940414e-07,1.940416e-07,1.940418e-07,1.940420e-07,1.940422e-07,1.940424e-07,1.940426e-07,1.940428e-07,1.940430e-07,1.940432e-07,1.940434e-07,1.940436e-07,1.940438e-07,1.940440e-07,1.940442e-07,1.940444e-07,1.940445e-07,1.940447e-07,1.940449e-07,1.940451e-07,1.940453e-07,1.940455e-07,1.940457e-07,1.940459e-07,1.940461e-07,1.940463e-07,1.940465e-07,1.940467e-07,1.940469e-07,1.940471e-07,1.940473e-07,1.940475e-07,1.940477e-07,1.940478e-07,1.940480e-07,1.940482e-07,1.940484e-07,1.940486e-07,1.940488e-07,1.940490e-07,1.940492e-07,1.940494e-07,1.940496e-07,1.940498e-07,1.940500e-07,1.940502e-07,1.940504e-07,1.940506e-07,1.940508e-07,1.940510e-07,1.940511e-07,1.940513e-07,1.940515e-07,1.940517e-07,1.940519e-07,1.940521e-07,1.940523e-07,1.940525e-07,1.940527e-07,1.940529e-07,1.940531e-07,1.940533e-07,1.940535e-07,1.940537e-07,1.940539e-07,1.940541e-07,1.940543e-07,1.940544e-07,1.940546e-07,1.940548e-07,1.940550e-07,1.940552e-07,1.940554e-07,1.940556e-07,1.940558e-07,1.940560e-07,1.940562e-07,1.940564e-07,1.940566e-07,1.940568e-07,1.940570e-07,1.940572e-07,1.940574e-07,1.940576e-07,1.940577e-07,1.940579e-07,1.940581e-07,1.940583e-07,1.940585e-07,1.940587e-07,1.940589e-07,1.940591e-07,1.940593e-07,1.940595e-07,1.940597e-07,1.940599e-07,1.940601e-07,1.940603e-07,1.940605e-07,1.940607e-07,1.940609e-07,1.940610e-07,1.940612e-07,1.940614e-07,1.940616e-07,1.940618e-07,1.940620e-07,1.940622e-07,1.940624e-07,1.940626e-07,1.940628e-07,1.940630e-07,1.940632e-07,1.940634e-07,1.940636e-07,1.940638e-07,1.940640e-07,1.940641e-07,1.940643e-07,1.940645e-07,1.940647e-07,1.940649e-07,1.940651e-07,1.940653e-07,1.940655e-07,1.940657e-07,1.940659e-07,1.940661e-07,1.940663e-07,1.940665e-07,1.940667e-07,1.940669e-07,1.940671e-07,1.940673e-07,1.940674e-07,1.940676e-07,1.940678e-07,1.940680e-07,1.940682e-07,1.940684e-07,1.940686e-07,1.940688e-07,1.940690e-07,1.940692e-07,1.940694e-07,1.940696e-07,1.940698e-07,1.940700e-07,1.940702e-07,1.940704e-07,1.940705e-07,1.940707e-07,1.940709e-07,1.940711e-07,1.940713e-07,1.940715e-07,1.940717e-07,1.940719e-07,1.940721e-07,1.940723e-07,1.940725e-07,1.940727e-07,1.940729e-07,1.940731e-07,1.940733e-07,1.940735e-07,1.940736e-07,1.940738e-07,1.940740e-07,1.940742e-07,1.940744e-07,1.940746e-07,1.940748e-07,1.940750e-07,1.940752e-07,1.940754e-07,1.940756e-07,1.940758e-07,1.940760e-07,1.940762e-07,1.940764e-07,1.940766e-07,1.940767e-07,1.940769e-07,1.940771e-07,1.940773e-07,1.940775e-07,1.940777e-07,1.940779e-07,1.940781e-07,1.940783e-07,1.940785e-07,1.940787e-07,1.940789e-07,1.940791e-07,1.940793e-07,1.940795e-07,1.940797e-07,1.940798e-07,1.940800e-07,1.940802e-07,1.940804e-07,1.940806e-07,1.940808e-07,1.940810e-07,1.940812e-07,1.940814e-07,1.940816e-07,1.940818e-07,1.940820e-07,1.940822e-07,1.940824e-07,1.940826e-07,1.940828e-07,1.940829e-07,1.940831e-07,1.940833e-07,1.940835e-07,1.940837e-07,1.940839e-07,1.940841e-07,1.940843e-07,1.940845e-07,1.940847e-07,1.940849e-07,1.940851e-07,1.940853e-07,1.940855e-07,1.940857e-07,1.940858e-07,1.940860e-07,1.940862e-07,1.940864e-07,1.940866e-07,1.940868e-07,1.940870e-07,1.940872e-07,1.940874e-07,1.940876e-07,1.940878e-07,1.940880e-07,1.940882e-07,1.940884e-07,1.940886e-07,1.940888e-07,1.940889e-07,1.940891e-07,1.940893e-07,1.940895e-07,1.940897e-07,1.940899e-07,1.940901e-07,1.940903e-07,1.940905e-07,1.940907e-07,1.940909e-07,1.940911e-07,1.940913e-07,1.940915e-07,1.940917e-07,1.940918e-07,1.940920e-07,1.940922e-07,1.940924e-07,1.940926e-07,1.940928e-07,1.940930e-07,1.940932e-07,1.940934e-07,1.940936e-07,1.940938e-07,1.940940e-07,1.940942e-07,1.940944e-07,1.940946e-07,1.940948e-07,1.940949e-07,1.940951e-07,1.940953e-07,1.940955e-07,1.940957e-07,1.940959e-07,1.940961e-07,1.940963e-07,1.940965e-07,1.940967e-07,1.940969e-07,1.940971e-07,1.940973e-07,1.940975e-07,1.940977e-07,1.940978e-07,1.940980e-07,1.940982e-07,1.940984e-07,1.940986e-07,1.940988e-07,1.940990e-07,1.940992e-07,1.940994e-07,1.940996e-07,1.940998e-07,1.941000e-07,1.941002e-07,1.941004e-07,1.941006e-07,1.941007e-07,1.941009e-07,1.941011e-07,1.941013e-07,1.941015e-07,1.941017e-07,1.941019e-07,1.941021e-07,1.941023e-07,1.941025e-07,1.941027e-07,1.941029e-07,1.941031e-07,1.941033e-07,1.941035e-07,1.941036e-07,1.941038e-07,1.941040e-07,1.941042e-07,1.941044e-07,1.941046e-07,1.941048e-07,1.941050e-07,1.941052e-07,1.941054e-07,1.941056e-07,1.941058e-07,1.941060e-07,1.941062e-07,1.941063e-07,1.941065e-07,1.941067e-07,1.941069e-07,1.941071e-07,1.941073e-07,1.941075e-07,1.941077e-07,1.941079e-07,1.941081e-07,1.941083e-07,1.941085e-07,1.941087e-07,1.941089e-07,1.941091e-07,1.941092e-07,1.941094e-07,1.941096e-07,1.941098e-07,1.941100e-07,1.941102e-07,1.941104e-07,1.941106e-07,1.941108e-07,1.941110e-07,1.941112e-07,1.941114e-07,1.941116e-07,1.941118e-07,1.941120e-07,1.941121e-07,1.941123e-07,1.941125e-07,1.941127e-07,1.941129e-07,1.941131e-07,1.941133e-07,1.941135e-07,1.941137e-07,1.941139e-07,1.941141e-07,1.941143e-07,1.941145e-07,1.941147e-07,1.941148e-07,1.941150e-07,1.941152e-07,1.941154e-07,1.941156e-07,1.941158e-07,1.941160e-07,1.941162e-07,1.941164e-07,1.941166e-07,1.941168e-07,1.941170e-07,1.941172e-07,1.941174e-07,1.941176e-07,1.941177e-07,1.941179e-07,1.941181e-07,1.941183e-07,1.941185e-07,1.941187e-07,1.941189e-07,1.941191e-07,1.941193e-07,1.941195e-07,1.941197e-07,1.941199e-07,1.941201e-07,1.941203e-07,1.941204e-07,1.941206e-07,1.941208e-07,1.941210e-07,1.941212e-07,1.941214e-07,1.941216e-07,1.941218e-07,1.941220e-07,1.941222e-07,1.941224e-07,1.941226e-07,1.941228e-07,1.941230e-07,1.941231e-07,1.941233e-07,1.941235e-07,1.941237e-07,1.941239e-07,1.941241e-07,1.941243e-07,1.941245e-07,1.941247e-07,1.941249e-07,1.941251e-07,1.941253e-07,1.941255e-07,1.941257e-07,1.941258e-07,1.941260e-07,1.941262e-07,1.941264e-07,1.941266e-07,1.941268e-07,1.941270e-07,1.941272e-07,1.941274e-07,1.941276e-07,1.941278e-07,1.941280e-07,1.941282e-07,1.941284e-07,1.941286e-07,1.941287e-07,1.941289e-07,1.941291e-07,1.941293e-07,1.941295e-07,1.941297e-07,1.941299e-07,1.941301e-07,1.941303e-07,1.941305e-07,1.941307e-07,1.941309e-07,1.941311e-07,1.941313e-07,1.941314e-07,1.941316e-07,1.941318e-07,1.941320e-07,1.941322e-07,1.941324e-07,1.941326e-07,1.941328e-07,1.941330e-07,1.941332e-07,1.941334e-07,1.941336e-07,1.941338e-07,1.941339e-07,1.941341e-07,1.941343e-07,1.941345e-07,1.941347e-07,1.941349e-07,1.941351e-07,1.941353e-07,1.941355e-07,1.941357e-07,1.941359e-07,1.941361e-07,1.941363e-07,1.941365e-07,1.941366e-07,1.941368e-07,1.941370e-07,1.941372e-07,1.941374e-07,1.941376e-07,1.941378e-07,1.941380e-07,1.941382e-07,1.941384e-07,1.941386e-07,1.941388e-07,1.941390e-07,1.941392e-07,1.941393e-07,1.941395e-07,1.941397e-07,1.941399e-07,1.941401e-07,1.941403e-07,1.941405e-07,1.941407e-07,1.941409e-07,1.941411e-07,1.941413e-07,1.941415e-07,1.941417e-07,1.941419e-07,1.941420e-07,1.941422e-07,1.941424e-07,1.941426e-07,1.941428e-07,1.941430e-07,1.941432e-07,1.941434e-07,1.941436e-07,1.941438e-07,1.941440e-07,1.941442e-07,1.941444e-07,1.941445e-07,1.941447e-07,1.941449e-07,1.941451e-07,1.941453e-07,1.941455e-07,1.941457e-07,1.941459e-07,1.941461e-07,1.941463e-07,1.941465e-07,1.941467e-07,1.941469e-07,1.941471e-07,1.941472e-07,1.941474e-07,1.941476e-07,1.941478e-07,1.941480e-07,1.941482e-07,1.941484e-07,1.941486e-07,1.941488e-07,1.941490e-07,1.941492e-07,1.941494e-07,1.941496e-07,1.941497e-07,1.941499e-07,1.941501e-07,1.941503e-07,1.941505e-07,1.941507e-07,1.941509e-07,1.941511e-07,1.941513e-07,1.941515e-07,1.941517e-07,1.941519e-07,1.941521e-07,1.941522e-07,1.941524e-07,1.941526e-07,1.941528e-07,1.941530e-07,1.941532e-07,1.941534e-07,1.941536e-07,1.941538e-07,1.941540e-07,1.941542e-07,1.941544e-07,1.941546e-07,1.941548e-07,1.941549e-07,1.941551e-07,1.941553e-07,1.941555e-07,1.941557e-07,1.941559e-07,1.941561e-07,1.941563e-07,1.941565e-07,1.941567e-07,1.941569e-07,1.941571e-07,1.941573e-07,1.941574e-07,1.941576e-07,1.941578e-07,1.941580e-07,1.941582e-07,1.941584e-07,1.941586e-07,1.941588e-07,1.941590e-07,1.941592e-07,1.941594e-07,1.941596e-07,1.941598e-07,1.941599e-07,1.941601e-07,1.941603e-07,1.941605e-07,1.941607e-07,1.941609e-07,1.941611e-07,1.941613e-07,1.941615e-07,1.941617e-07,1.941619e-07,1.941621e-07,1.941623e-07,1.941624e-07,1.941626e-07,1.941628e-07,1.941630e-07,1.941632e-07,1.941634e-07,1.941636e-07,1.941638e-07,1.941640e-07,1.941642e-07,1.941644e-07,1.941646e-07,1.941648e-07,1.941649e-07,1.941651e-07,1.941653e-07,1.941655e-07,1.941657e-07,1.941659e-07,1.941661e-07,1.941663e-07,1.941665e-07,1.941667e-07,1.941669e-07,1.941671e-07,1.941673e-07,1.941674e-07,1.941676e-07,1.941678e-07,1.941680e-07,1.941682e-07,1.941684e-07,1.941686e-07,1.941688e-07,1.941690e-07,1.941692e-07,1.941694e-07,1.941696e-07,1.941698e-07,1.941699e-07,1.941701e-07,1.941703e-07,1.941705e-07,1.941707e-07,1.941709e-07,1.941711e-07,1.941713e-07,1.941715e-07,1.941717e-07,1.941719e-07,1.941721e-07,1.941722e-07,1.941724e-07,1.941726e-07,1.941728e-07,1.941730e-07,1.941732e-07,1.941734e-07,1.941736e-07,1.941738e-07,1.941740e-07,1.941742e-07,1.941744e-07,1.941746e-07,1.941747e-07,1.941749e-07,1.941751e-07,1.941753e-07,1.941755e-07,1.941757e-07,1.941759e-07,1.941761e-07,1.941763e-07,1.941765e-07,1.941767e-07,1.941769e-07,1.941771e-07,1.941772e-07,1.941774e-07,1.941776e-07,1.941778e-07,1.941780e-07,1.941782e-07,1.941784e-07,1.941786e-07,1.941788e-07,1.941790e-07,1.941792e-07,1.941794e-07,1.941795e-07,1.941797e-07,1.941799e-07,1.941801e-07,1.941803e-07,1.941805e-07,1.941807e-07,1.941809e-07,1.941811e-07,1.941813e-07,1.941815e-07,1.941817e-07,1.941819e-07,1.941820e-07,1.941822e-07,1.941824e-07,1.941826e-07,1.941828e-07,1.941830e-07,1.941832e-07,1.941834e-07,1.941836e-07,1.941838e-07,1.941840e-07,1.941842e-07,1.941843e-07,1.941845e-07,1.941847e-07,1.941849e-07,1.941851e-07,1.941853e-07,1.941855e-07,1.941857e-07,1.941859e-07,1.941861e-07,1.941863e-07,1.941865e-07,1.941867e-07,1.941868e-07,1.941870e-07,1.941872e-07,1.941874e-07,1.941876e-07,1.941878e-07,1.941880e-07,1.941882e-07,1.941884e-07,1.941886e-07,1.941888e-07,1.941890e-07,1.941891e-07,1.941893e-07,1.941895e-07,1.941897e-07,1.941899e-07,1.941901e-07,1.941903e-07,1.941905e-07,1.941907e-07,1.941909e-07,1.941911e-07,1.941913e-07,1.941914e-07,1.941916e-07,1.941918e-07,1.941920e-07,1.941922e-07,1.941924e-07,1.941926e-07,1.941928e-07,1.941930e-07,1.941932e-07,1.941934e-07,1.941936e-07,1.941937e-07,1.941939e-07,1.941941e-07,1.941943e-07,1.941945e-07,1.941947e-07,1.941949e-07,1.941951e-07,1.941953e-07,1.941955e-07,1.941957e-07,1.941959e-07,1.941961e-07,1.941962e-07,1.941964e-07,1.941966e-07,1.941968e-07,1.941970e-07,1.941972e-07,1.941974e-07,1.941976e-07,1.941978e-07,1.941980e-07,1.941982e-07,1.941984e-07,1.941985e-07,1.941987e-07,1.941989e-07,1.941991e-07,1.941993e-07,1.941995e-07,1.941997e-07,1.941999e-07,1.942001e-07,1.942003e-07,1.942005e-07,1.942007e-07,1.942008e-07,1.942010e-07,1.942012e-07,1.942014e-07,1.942016e-07,1.942018e-07,1.942020e-07,1.942022e-07,1.942024e-07,1.942026e-07,1.942028e-07,1.942030e-07,1.942031e-07,1.942033e-07,1.942035e-07,1.942037e-07,1.942039e-07,1.942041e-07,1.942043e-07,1.942045e-07,1.942047e-07,1.942049e-07,1.942051e-07,1.942053e-07,1.942054e-07,1.942056e-07,1.942058e-07,1.942060e-07,1.942062e-07,1.942064e-07,1.942066e-07,1.942068e-07,1.942070e-07,1.942072e-07,1.942074e-07,1.942076e-07,1.942077e-07,1.942079e-07,1.942081e-07,1.942083e-07,1.942085e-07,1.942087e-07,1.942089e-07,1.942091e-07,1.942093e-07,1.942095e-07,1.942097e-07,1.942098e-07,1.942100e-07,1.942102e-07,1.942104e-07,1.942106e-07,1.942108e-07,1.942110e-07,1.942112e-07,1.942114e-07,1.942116e-07,1.942118e-07,1.942120e-07,1.942121e-07,1.942123e-07,1.942125e-07,1.942127e-07,1.942129e-07,1.942131e-07,1.942133e-07,1.942135e-07,1.942137e-07,1.942139e-07,1.942141e-07,1.942143e-07,1.942144e-07,1.942146e-07,1.942148e-07,1.942150e-07,1.942152e-07,1.942154e-07,1.942156e-07,1.942158e-07,1.942160e-07,1.942162e-07,1.942164e-07,1.942166e-07,1.942167e-07,1.942169e-07,1.942171e-07,1.942173e-07,1.942175e-07,1.942177e-07,1.942179e-07,1.942181e-07,1.942183e-07,1.942185e-07,1.942187e-07,1.942188e-07,1.942190e-07,1.942192e-07,1.942194e-07,1.942196e-07,1.942198e-07,1.942200e-07,1.942202e-07,1.942204e-07,1.942206e-07,1.942208e-07,1.942210e-07,1.942211e-07,1.942213e-07,1.942215e-07,1.942217e-07,1.942219e-07,1.942221e-07,1.942223e-07,1.942225e-07,1.942227e-07,1.942229e-07,1.942231e-07,1.942232e-07,1.942234e-07,1.942236e-07,1.942238e-07,1.942240e-07,1.942242e-07,1.942244e-07,1.942246e-07,1.942248e-07,1.942250e-07,1.942252e-07,1.942254e-07,1.942255e-07,1.942257e-07,1.942259e-07,1.942261e-07,1.942263e-07,1.942265e-07,1.942267e-07,1.942269e-07,1.942271e-07,1.942273e-07,1.942275e-07,1.942276e-07,1.942278e-07,1.942280e-07,1.942282e-07,1.942284e-07,1.942286e-07,1.942288e-07,1.942290e-07,1.942292e-07,1.942294e-07,1.942296e-07,1.942298e-07,1.942299e-07,1.942301e-07,1.942303e-07,1.942305e-07,1.942307e-07,1.942309e-07,1.942311e-07,1.942313e-07,1.942315e-07,1.942317e-07,1.942319e-07,1.942320e-07,1.942322e-07,1.942324e-07,1.942326e-07,1.942328e-07,1.942330e-07,1.942332e-07,1.942334e-07,1.942336e-07,1.942338e-07,1.942340e-07,1.942341e-07,1.942343e-07,1.942345e-07,1.942347e-07,1.942349e-07,1.942351e-07,1.942353e-07,1.942355e-07,1.942357e-07,1.942359e-07,1.942361e-07,1.942363e-07,1.942364e-07,1.942366e-07,1.942368e-07,1.942370e-07,1.942372e-07,1.942374e-07,1.942376e-07,1.942378e-07,1.942380e-07,1.942382e-07,1.942384e-07,1.942385e-07,1.942387e-07,1.942389e-07,1.942391e-07,1.942393e-07,1.942395e-07,1.942397e-07,1.942399e-07,1.942401e-07,1.942403e-07,1.942405e-07,1.942406e-07,1.942408e-07,1.942410e-07,1.942412e-07,1.942414e-07,1.942416e-07,1.942418e-07,1.942420e-07,1.942422e-07,1.942424e-07,1.942426e-07,1.942427e-07,1.942429e-07,1.942431e-07,1.942433e-07,1.942435e-07,1.942437e-07,1.942439e-07,1.942441e-07,1.942443e-07,1.942445e-07,1.942447e-07,1.942448e-07,1.942450e-07,1.942452e-07,1.942454e-07,1.942456e-07,1.942458e-07,1.942460e-07,1.942462e-07,1.942464e-07,1.942466e-07,1.942468e-07,1.942469e-07,1.942471e-07,1.942473e-07,1.942475e-07,1.942477e-07,1.942479e-07,1.942481e-07,1.942483e-07,1.942485e-07,1.942487e-07,1.942489e-07,1.942490e-07,1.942492e-07,1.942494e-07,1.942496e-07,1.942498e-07,1.942500e-07,1.942502e-07,1.942504e-07,1.942506e-07,1.942508e-07,1.942510e-07,1.942511e-07,1.942513e-07,1.942515e-07,1.942517e-07,1.942519e-07,1.942521e-07,1.942523e-07,1.942525e-07,1.942527e-07,1.942529e-07,1.942531e-07,1.942532e-07,1.942534e-07,1.942536e-07,1.942538e-07,1.942540e-07,1.942542e-07,1.942544e-07,1.942546e-07,1.942548e-07,1.942550e-07,1.942552e-07,1.942553e-07,1.942555e-07,1.942557e-07,1.942559e-07,1.942561e-07,1.942563e-07,1.942565e-07,1.942567e-07,1.942569e-07,1.942571e-07,1.942573e-07,1.942574e-07,1.942576e-07,1.942578e-07,1.942580e-07,1.942582e-07,1.942584e-07,1.942586e-07,1.942588e-07,1.942590e-07,1.942592e-07,1.942594e-07,1.942595e-07,1.942597e-07,1.942599e-07,1.942601e-07,1.942603e-07,1.942605e-07,1.942607e-07,1.942609e-07,1.942611e-07,1.942613e-07,1.942614e-07,1.942616e-07,1.942618e-07,1.942620e-07,1.942622e-07,1.942624e-07,1.942626e-07,1.942628e-07,1.942630e-07,1.942632e-07,1.942634e-07,1.942635e-07,1.942637e-07,1.942639e-07,1.942641e-07,1.942643e-07,1.942645e-07,1.942647e-07,1.942649e-07,1.942651e-07,1.942653e-07,1.942655e-07,1.942656e-07,1.942658e-07,1.942660e-07,1.942662e-07,1.942664e-07,1.942666e-07,1.942668e-07,1.942670e-07,1.942672e-07,1.942674e-07,1.942675e-07,1.942677e-07,1.942679e-07,1.942681e-07,1.942683e-07,1.942685e-07,1.942687e-07,1.942689e-07,1.942691e-07,1.942693e-07,1.942695e-07,1.942696e-07,1.942698e-07,1.942700e-07,1.942702e-07,1.942704e-07,1.942706e-07,1.942708e-07,1.942710e-07,1.942712e-07,1.942714e-07,1.942716e-07,1.942717e-07,1.942719e-07,1.942721e-07,1.942723e-07,1.942725e-07,1.942727e-07,1.942729e-07,1.942731e-07,1.942733e-07,1.942735e-07,1.942736e-07,1.942738e-07,1.942740e-07,1.942742e-07,1.942744e-07,1.942746e-07,1.942748e-07,1.942750e-07,1.942752e-07,1.942754e-07,1.942756e-07,1.942757e-07,1.942759e-07,1.942761e-07,1.942763e-07,1.942765e-07,1.942767e-07,1.942769e-07,1.942771e-07,1.942773e-07,1.942775e-07,1.942776e-07,1.942778e-07,1.942780e-07,1.942782e-07,1.942784e-07,1.942786e-07,1.942788e-07,1.942790e-07,1.942792e-07,1.942794e-07,1.942795e-07,1.942797e-07,1.942799e-07,1.942801e-07,1.942803e-07,1.942805e-07,1.942807e-07,1.942809e-07,1.942811e-07,1.942813e-07,1.942815e-07,1.942816e-07,1.942818e-07,1.942820e-07,1.942822e-07,1.942824e-07,1.942826e-07,1.942828e-07,1.942830e-07,1.942832e-07,1.942834e-07,1.942835e-07,1.942837e-07,1.942839e-07,1.942841e-07,1.942843e-07,1.942845e-07,1.942847e-07,1.942849e-07,1.942851e-07,1.942853e-07,1.942855e-07,1.942856e-07,1.942858e-07,1.942860e-07,1.942862e-07,1.942864e-07,1.942866e-07,1.942868e-07,1.942870e-07,1.942872e-07,1.942874e-07,1.942875e-07,1.942877e-07,1.942879e-07,1.942881e-07,1.942883e-07,1.942885e-07,1.942887e-07,1.942889e-07,1.942891e-07,1.942893e-07,1.942894e-07,1.942896e-07,1.942898e-07,1.942900e-07,1.942902e-07,1.942904e-07,1.942906e-07,1.942908e-07,1.942910e-07,1.942912e-07,1.942913e-07,1.942915e-07,1.942917e-07,1.942919e-07,1.942921e-07,1.942923e-07,1.942925e-07,1.942927e-07,1.942929e-07,1.942931e-07,1.942933e-07,1.942934e-07,1.942936e-07,1.942938e-07,1.942940e-07,1.942942e-07,1.942944e-07,1.942946e-07,1.942948e-07,1.942950e-07,1.942952e-07,1.942953e-07,1.942955e-07,1.942957e-07,1.942959e-07,1.942961e-07,1.942963e-07,1.942965e-07,1.942967e-07,1.942969e-07,1.942971e-07,1.942972e-07,1.942974e-07,1.942976e-07,1.942978e-07,1.942980e-07,1.942982e-07,1.942984e-07,1.942986e-07,1.942988e-07,1.942990e-07,1.942991e-07,1.942993e-07,1.942995e-07,1.942997e-07,1.942999e-07,1.943001e-07,1.943003e-07,1.943005e-07,1.943007e-07,1.943009e-07,1.943010e-07,1.943012e-07,1.943014e-07,1.943016e-07,1.943018e-07,1.943020e-07,1.943022e-07,1.943024e-07,1.943026e-07,1.943028e-07,1.943029e-07,1.943031e-07,1.943033e-07,1.943035e-07,1.943037e-07,1.943039e-07,1.943041e-07,1.943043e-07,1.943045e-07,1.943047e-07,1.943048e-07,1.943050e-07,1.943052e-07,1.943054e-07,1.943056e-07,1.943058e-07,1.943060e-07,1.943062e-07,1.943064e-07,1.943066e-07,1.943067e-07,1.943069e-07,1.943071e-07,1.943073e-07,1.943075e-07,1.943077e-07,1.943079e-07,1.943081e-07,1.943083e-07,1.943085e-07,1.943086e-07,1.943088e-07,1.943090e-07,1.943092e-07,1.943094e-07,1.943096e-07,1.943098e-07,1.943100e-07,1.943102e-07,1.943104e-07,1.943105e-07,1.943107e-07,1.943109e-07,1.943111e-07,1.943113e-07,1.943115e-07,1.943117e-07,1.943119e-07,1.943121e-07,1.943123e-07,1.943124e-07,1.943126e-07,1.943128e-07,1.943130e-07,1.943132e-07,1.943134e-07,1.943136e-07,1.943138e-07,1.943140e-07,1.943142e-07,1.943143e-07,1.943145e-07,1.943147e-07,1.943149e-07,1.943151e-07,1.943153e-07,1.943155e-07,1.943157e-07,1.943159e-07,1.943160e-07,1.943162e-07,1.943164e-07,1.943166e-07,1.943168e-07,1.943170e-07,1.943172e-07,1.943174e-07,1.943176e-07,1.943178e-07,1.943179e-07,1.943181e-07,1.943183e-07,1.943185e-07,1.943187e-07,1.943189e-07,1.943191e-07,1.943193e-07,1.943195e-07,1.943197e-07,1.943198e-07,1.943200e-07,1.943202e-07,1.943204e-07,1.943206e-07,1.943208e-07,1.943210e-07,1.943212e-07,1.943214e-07,1.943216e-07,1.943217e-07,1.943219e-07,1.943221e-07,1.943223e-07,1.943225e-07,1.943227e-07,1.943229e-07,1.943231e-07,1.943233e-07,1.943234e-07,1.943236e-07,1.943238e-07,1.943240e-07,1.943242e-07,1.943244e-07,1.943246e-07,1.943248e-07,1.943250e-07,1.943252e-07,1.943253e-07,1.943255e-07,1.943257e-07,1.943259e-07,1.943261e-07,1.943263e-07,1.943265e-07,1.943267e-07,1.943269e-07,1.943271e-07,1.943272e-07,1.943274e-07,1.943276e-07,1.943278e-07,1.943280e-07,1.943282e-07,1.943284e-07,1.943286e-07,1.943288e-07,1.943289e-07,1.943291e-07,1.943293e-07,1.943295e-07,1.943297e-07,1.943299e-07,1.943301e-07,1.943303e-07,1.943305e-07,1.943307e-07,1.943308e-07,1.943310e-07,1.943312e-07,1.943314e-07,1.943316e-07,1.943318e-07,1.943320e-07,1.943322e-07,1.943324e-07,1.943325e-07,1.943327e-07,1.943329e-07,1.943331e-07,1.943333e-07,1.943335e-07,1.943337e-07,1.943339e-07,1.943341e-07,1.943343e-07,1.943344e-07,1.943346e-07,1.943348e-07,1.943350e-07,1.943352e-07,1.943354e-07,1.943356e-07,1.943358e-07,1.943360e-07,1.943361e-07,1.943363e-07,1.943365e-07,1.943367e-07,1.943369e-07,1.943371e-07,1.943373e-07,1.943375e-07,1.943377e-07,1.943379e-07,1.943380e-07,1.943382e-07,1.943384e-07,1.943386e-07,1.943388e-07,1.943390e-07,1.943392e-07,1.943394e-07,1.943396e-07,1.943397e-07,1.943399e-07,1.943401e-07,1.943403e-07,1.943405e-07,1.943407e-07,1.943409e-07,1.943411e-07,1.943413e-07,1.943415e-07,1.943416e-07,1.943418e-07,1.943420e-07,1.943422e-07,1.943424e-07,1.943426e-07,1.943428e-07,1.943430e-07,1.943432e-07,1.943433e-07,1.943435e-07,1.943437e-07,1.943439e-07,1.943441e-07,1.943443e-07,1.943445e-07,1.943447e-07,1.943449e-07,1.943451e-07,1.943452e-07,1.943454e-07,1.943456e-07,1.943458e-07,1.943460e-07,1.943462e-07,1.943464e-07,1.943466e-07,1.943468e-07,1.943469e-07,1.943471e-07,1.943473e-07,1.943475e-07,1.943477e-07,1.943479e-07,1.943481e-07,1.943483e-07,1.943485e-07,1.943486e-07,1.943488e-07,1.943490e-07,1.943492e-07,1.943494e-07,1.943496e-07,1.943498e-07,1.943500e-07,1.943502e-07,1.943504e-07,1.943505e-07,1.943507e-07,1.943509e-07,1.943511e-07,1.943513e-07,1.943515e-07,1.943517e-07,1.943519e-07,1.943521e-07,1.943522e-07,1.943524e-07,1.943526e-07,1.943528e-07,1.943530e-07,1.943532e-07,1.943534e-07,1.943536e-07,1.943538e-07,1.943539e-07,1.943541e-07,1.943543e-07,1.943545e-07,1.943547e-07,1.943549e-07,1.943551e-07,1.943553e-07,1.943555e-07,1.943556e-07,1.943558e-07,1.943560e-07,1.943562e-07,1.943564e-07,1.943566e-07,1.943568e-07,1.943570e-07,1.943572e-07,1.943574e-07,1.943575e-07,1.943577e-07,1.943579e-07,1.943581e-07,1.943583e-07,1.943585e-07,1.943587e-07,1.943589e-07,1.943591e-07,1.943592e-07,1.943594e-07,1.943596e-07,1.943598e-07,1.943600e-07,1.943602e-07,1.943604e-07,1.943606e-07,1.943608e-07,1.943609e-07,1.943611e-07,1.943613e-07,1.943615e-07,1.943617e-07,1.943619e-07,1.943621e-07,1.943623e-07,1.943625e-07,1.943626e-07,1.943628e-07,1.943630e-07,1.943632e-07,1.943634e-07,1.943636e-07,1.943638e-07,1.943640e-07,1.943642e-07,1.943643e-07,1.943645e-07,1.943647e-07,1.943649e-07,1.943651e-07,1.943653e-07,1.943655e-07,1.943657e-07,1.943659e-07,1.943660e-07,1.943662e-07,1.943664e-07,1.943666e-07,1.943668e-07,1.943670e-07,1.943672e-07,1.943674e-07,1.943676e-07,1.943677e-07,1.943679e-07,1.943681e-07,1.943683e-07,1.943685e-07,1.943687e-07,1.943689e-07,1.943691e-07,1.943693e-07,1.943695e-07,1.943696e-07,1.943698e-07,1.943700e-07,1.943702e-07,1.943704e-07,1.943706e-07,1.943708e-07,1.943710e-07,1.943712e-07,1.943713e-07,1.943715e-07,1.943717e-07,1.943719e-07,1.943721e-07,1.943723e-07,1.943725e-07,1.943727e-07,1.943729e-07,1.943730e-07,1.943732e-07,1.943734e-07,1.943736e-07,1.943738e-07,1.943740e-07,1.943742e-07,1.943744e-07,1.943746e-07,1.943747e-07,1.943749e-07,1.943751e-07,1.943753e-07,1.943755e-07,1.943757e-07,1.943759e-07,1.943761e-07,1.943762e-07,1.943764e-07,1.943766e-07,1.943768e-07,1.943770e-07,1.943772e-07,1.943774e-07,1.943776e-07,1.943778e-07,1.943779e-07,1.943781e-07,1.943783e-07,1.943785e-07,1.943787e-07,1.943789e-07,1.943791e-07,1.943793e-07,1.943795e-07,1.943796e-07,1.943798e-07,1.943800e-07,1.943802e-07,1.943804e-07,1.943806e-07,1.943808e-07,1.943810e-07,1.943812e-07,1.943813e-07,1.943815e-07,1.943817e-07,1.943819e-07,1.943821e-07,1.943823e-07,1.943825e-07,1.943827e-07,1.943829e-07,1.943830e-07,1.943832e-07,1.943834e-07,1.943836e-07,1.943838e-07,1.943840e-07,1.943842e-07,1.943844e-07,1.943846e-07,1.943847e-07,1.943849e-07,1.943851e-07,1.943853e-07,1.943855e-07,1.943857e-07,1.943859e-07,1.943861e-07,1.943863e-07,1.943864e-07,1.943866e-07,1.943868e-07,1.943870e-07,1.943872e-07,1.943874e-07,1.943876e-07,1.943878e-07,1.943880e-07,1.943881e-07,1.943883e-07,1.943885e-07,1.943887e-07,1.943889e-07,1.943891e-07,1.943893e-07,1.943895e-07,1.943896e-07,1.943898e-07,1.943900e-07,1.943902e-07,1.943904e-07,1.943906e-07,1.943908e-07,1.943910e-07,1.943912e-07,1.943913e-07,1.943915e-07,1.943917e-07,1.943919e-07,1.943921e-07,1.943923e-07,1.943925e-07,1.943927e-07,1.943929e-07,1.943930e-07,1.943932e-07,1.943934e-07,1.943936e-07,1.943938e-07,1.943940e-07,1.943942e-07,1.943944e-07,1.943946e-07,1.943947e-07,1.943949e-07,1.943951e-07,1.943953e-07,1.943955e-07,1.943957e-07,1.943959e-07,1.943961e-07,1.943962e-07,1.943964e-07,1.943966e-07,1.943968e-07,1.943970e-07,1.943972e-07,1.943974e-07,1.943976e-07,1.943978e-07,1.943979e-07,1.943981e-07,1.943983e-07,1.943985e-07,1.943987e-07,1.943989e-07,1.943991e-07,1.943993e-07,1.943995e-07,1.943996e-07,1.943998e-07,1.944000e-07,1.944002e-07,1.944004e-07,1.944006e-07,1.944008e-07,1.944010e-07,1.944011e-07,1.944013e-07,1.944015e-07,1.944017e-07,1.944019e-07,1.944021e-07,1.944023e-07,1.944025e-07,1.944027e-07,1.944028e-07,1.944030e-07,1.944032e-07,1.944034e-07,1.944036e-07,1.944038e-07,1.944040e-07,1.944042e-07,1.944044e-07,1.944045e-07,1.944047e-07,1.944049e-07,1.944051e-07,1.944053e-07,1.944055e-07,1.944057e-07,1.944059e-07,1.944060e-07,1.944062e-07,1.944064e-07,1.944066e-07,1.944068e-07,1.944070e-07,1.944072e-07,1.944074e-07,1.944076e-07,1.944077e-07,1.944079e-07,1.944081e-07,1.944083e-07,1.944085e-07,1.944087e-07,1.944089e-07,1.944091e-07,1.944092e-07,1.944094e-07,1.944096e-07,1.944098e-07,1.944100e-07,1.944102e-07,1.944104e-07,1.944106e-07,1.944108e-07,1.944109e-07,1.944111e-07,1.944113e-07,1.944115e-07,1.944117e-07,1.944119e-07,1.944121e-07,1.944123e-07,1.944124e-07,1.944126e-07,1.944128e-07,1.944130e-07,1.944132e-07,1.944134e-07,1.944136e-07,1.944138e-07,1.944140e-07,1.944141e-07,1.944143e-07,1.944145e-07,1.944147e-07,1.944149e-07,1.944151e-07,1.944153e-07,1.944155e-07,1.944156e-07,1.944158e-07,1.944160e-07,1.944162e-07,1.944164e-07,1.944166e-07,1.944168e-07,1.944170e-07,1.944172e-07,1.944173e-07,1.944175e-07,1.944177e-07,1.944179e-07,1.944181e-07,1.944183e-07,1.944185e-07,1.944187e-07,1.944188e-07,1.944190e-07,1.944192e-07,1.944194e-07,1.944196e-07,1.944198e-07,1.944200e-07,1.944202e-07,1.944204e-07,1.944205e-07,1.944207e-07,1.944209e-07,1.944211e-07,1.944213e-07,1.944215e-07,1.944217e-07,1.944219e-07,1.944220e-07,1.944222e-07,1.944224e-07,1.944226e-07,1.944228e-07,1.944230e-07,1.944232e-07,1.944234e-07,1.944235e-07,1.944237e-07,1.944239e-07,1.944241e-07,1.944243e-07,1.944245e-07,1.944247e-07,1.944249e-07,1.944251e-07,1.944252e-07,1.944254e-07,1.944256e-07,1.944258e-07,1.944260e-07,1.944262e-07,1.944264e-07,1.944266e-07,1.944267e-07,1.944269e-07,1.944271e-07,1.944273e-07,1.944275e-07,1.944277e-07,1.944279e-07,1.944281e-07,1.944283e-07,1.944284e-07,1.944286e-07,1.944288e-07,1.944290e-07,1.944292e-07,1.944294e-07,1.944296e-07,1.944298e-07,1.944299e-07,1.944301e-07,1.944303e-07,1.944305e-07,1.944307e-07,1.944309e-07,1.944311e-07,1.944313e-07,1.944314e-07,1.944316e-07,1.944318e-07,1.944320e-07,1.944322e-07,1.944324e-07,1.944326e-07,1.944328e-07,1.944329e-07,1.944331e-07,1.944333e-07,1.944335e-07,1.944337e-07,1.944339e-07,1.944341e-07,1.944343e-07,1.944345e-07,1.944346e-07,1.944348e-07,1.944350e-07,1.944352e-07,1.944354e-07,1.944356e-07,1.944358e-07,1.944360e-07,1.944361e-07,1.944363e-07,1.944365e-07,1.944367e-07,1.944369e-07,1.944371e-07,1.944373e-07,1.944375e-07,1.944376e-07,1.944378e-07,1.944380e-07,1.944382e-07,1.944384e-07,1.944386e-07,1.944388e-07,1.944390e-07,1.944391e-07,1.944393e-07,1.944395e-07,1.944397e-07,1.944399e-07,1.944401e-07,1.944403e-07,1.944405e-07,1.944407e-07,1.944408e-07,1.944410e-07,1.944412e-07,1.944414e-07,1.944416e-07,1.944418e-07,1.944420e-07,1.944422e-07,1.944423e-07,1.944425e-07,1.944427e-07,1.944429e-07,1.944431e-07,1.944433e-07,1.944435e-07,1.944437e-07,1.944438e-07,1.944440e-07,1.944442e-07,1.944444e-07,1.944446e-07,1.944448e-07,1.944450e-07,1.944452e-07,1.944453e-07,1.944455e-07,1.944457e-07,1.944459e-07,1.944461e-07,1.944463e-07,1.944465e-07,1.944467e-07,1.944468e-07,1.944470e-07,1.944472e-07,1.944474e-07,1.944476e-07,1.944478e-07,1.944480e-07,1.944482e-07,1.944483e-07,1.944485e-07,1.944487e-07,1.944489e-07,1.944491e-07,1.944493e-07,1.944495e-07,1.944497e-07,1.944498e-07,1.944500e-07,1.944502e-07,1.944504e-07,1.944506e-07,1.944508e-07,1.944510e-07,1.944512e-07,1.944514e-07,1.944515e-07,1.944517e-07,1.944519e-07,1.944521e-07,1.944523e-07,1.944525e-07,1.944527e-07,1.944529e-07,1.944530e-07,1.944532e-07,1.944534e-07,1.944536e-07,1.944538e-07,1.944540e-07,1.944542e-07,1.944544e-07,1.944545e-07,1.944547e-07,1.944549e-07,1.944551e-07,1.944553e-07,1.944555e-07,1.944557e-07,1.944559e-07,1.944560e-07,1.944562e-07,1.944564e-07,1.944566e-07,1.944568e-07,1.944570e-07,1.944572e-07,1.944574e-07,1.944575e-07,1.944577e-07,1.944579e-07,1.944581e-07,1.944583e-07,1.944585e-07,1.944587e-07,1.944589e-07,1.944590e-07,1.944592e-07,1.944594e-07,1.944596e-07,1.944598e-07,1.944600e-07,1.944602e-07,1.944604e-07,1.944605e-07,1.944607e-07,1.944609e-07,1.944611e-07,1.944613e-07,1.944615e-07,1.944617e-07,1.944619e-07,1.944620e-07,1.944622e-07,1.944624e-07,1.944626e-07,1.944628e-07,1.944630e-07,1.944632e-07,1.944634e-07,1.944635e-07,1.944637e-07,1.944639e-07,1.944641e-07,1.944643e-07,1.944645e-07,1.944647e-07,1.944649e-07,1.944650e-07,1.944652e-07,1.944654e-07,1.944656e-07,1.944658e-07,1.944660e-07,1.944662e-07,1.944664e-07,1.944665e-07,1.944667e-07,1.944669e-07,1.944671e-07,1.944673e-07,1.944675e-07,1.944677e-07,1.944678e-07,1.944680e-07,1.944682e-07,1.944684e-07,1.944686e-07,1.944688e-07,1.944690e-07,1.944692e-07,1.944693e-07,1.944695e-07,1.944697e-07,1.944699e-07,1.944701e-07,1.944703e-07,1.944705e-07,1.944707e-07,1.944708e-07,1.944710e-07,1.944712e-07,1.944714e-07,1.944716e-07,1.944718e-07,1.944720e-07,1.944722e-07,1.944723e-07,1.944725e-07,1.944727e-07,1.944729e-07,1.944731e-07,1.944733e-07,1.944735e-07,1.944737e-07,1.944738e-07,1.944740e-07,1.944742e-07,1.944744e-07,1.944746e-07,1.944748e-07,1.944750e-07,1.944752e-07,1.944753e-07,1.944755e-07,1.944757e-07,1.944759e-07,1.944761e-07,1.944763e-07,1.944765e-07,1.944767e-07,1.944768e-07,1.944770e-07,1.944772e-07,1.944774e-07,1.944776e-07,1.944778e-07,1.944780e-07,1.944781e-07,1.944783e-07,1.944785e-07,1.944787e-07,1.944789e-07,1.944791e-07,1.944793e-07,1.944795e-07,1.944796e-07,1.944798e-07,1.944800e-07,1.944802e-07,1.944804e-07,1.944806e-07,1.944808e-07,1.944810e-07,1.944811e-07,1.944813e-07,1.944815e-07,1.944817e-07,1.944819e-07,1.944821e-07,1.944823e-07,1.944825e-07,1.944826e-07,1.944828e-07,1.944830e-07,1.944832e-07,1.944834e-07,1.944836e-07,1.944838e-07,1.944840e-07,1.944841e-07,1.944843e-07,1.944845e-07,1.944847e-07,1.944849e-07,1.944851e-07,1.944853e-07,1.944854e-07,1.944856e-07,1.944858e-07,1.944860e-07,1.944862e-07,1.944864e-07,1.944866e-07,1.944868e-07,1.944869e-07,1.944871e-07,1.944873e-07,1.944875e-07,1.944877e-07,1.944879e-07,1.944881e-07,1.944883e-07,1.944884e-07,1.944886e-07,1.944888e-07,1.944890e-07,1.944892e-07,1.944894e-07,1.944896e-07,1.944897e-07,1.944899e-07,1.944901e-07,1.944903e-07,1.944905e-07,1.944907e-07,1.944909e-07,1.944911e-07,1.944912e-07,1.944914e-07,1.944916e-07,1.944918e-07,1.944920e-07,1.944922e-07,1.944924e-07,1.944926e-07,1.944927e-07,1.944929e-07,1.944931e-07,1.944933e-07,1.944935e-07,1.944937e-07,1.944939e-07,1.944940e-07,1.944942e-07,1.944944e-07,1.944946e-07,1.944948e-07,1.944950e-07,1.944952e-07,1.944954e-07,1.944955e-07,1.944957e-07,1.944959e-07,1.944961e-07,1.944963e-07,1.944965e-07,1.944967e-07,1.944969e-07,1.944970e-07,1.944972e-07,1.944974e-07,1.944976e-07,1.944978e-07,1.944980e-07,1.944982e-07,1.944983e-07,1.944985e-07,1.944987e-07,1.944989e-07,1.944991e-07,1.944993e-07,1.944995e-07,1.944997e-07,1.944998e-07,1.945000e-07,1.945002e-07,1.945004e-07,1.945006e-07,1.945008e-07,1.945010e-07,1.945012e-07,1.945013e-07,1.945015e-07,1.945017e-07,1.945019e-07,1.945021e-07,1.945023e-07,1.945025e-07,1.945026e-07,1.945028e-07,1.945030e-07,1.945032e-07,1.945034e-07,1.945036e-07,1.945038e-07,1.945040e-07,1.945041e-07,1.945043e-07,1.945045e-07,1.945047e-07,1.945049e-07,1.945051e-07,1.945053e-07,1.945054e-07,1.945056e-07,1.945058e-07,1.945060e-07,1.945062e-07,1.945064e-07,1.945066e-07,1.945068e-07,1.945069e-07,1.945071e-07,1.945073e-07,1.945075e-07,1.945077e-07,1.945079e-07,1.945081e-07,1.945082e-07,1.945084e-07,1.945086e-07,1.945088e-07,1.945090e-07,1.945092e-07,1.945094e-07,1.945096e-07,1.945097e-07,1.945099e-07,1.945101e-07,1.945103e-07,1.945105e-07,1.945107e-07,1.945109e-07,1.945110e-07,1.945112e-07,1.945114e-07,1.945116e-07,1.945118e-07,1.945120e-07,1.945122e-07,1.945124e-07,1.945125e-07,1.945127e-07,1.945129e-07,1.945131e-07,1.945133e-07,1.945135e-07,1.945137e-07,1.945138e-07,1.945140e-07,1.945142e-07,1.945144e-07,1.945146e-07,1.945148e-07,1.945150e-07,1.945152e-07,1.945153e-07,1.945155e-07,1.945157e-07,1.945159e-07,1.945161e-07,1.945163e-07,1.945165e-07,1.945166e-07,1.945168e-07,1.945170e-07,1.945172e-07,1.945174e-07,1.945176e-07,1.945178e-07,1.945180e-07,1.945181e-07,1.945183e-07,1.945185e-07,1.945187e-07,1.945189e-07,1.945191e-07,1.945193e-07,1.945194e-07,1.945196e-07,1.945198e-07,1.945200e-07,1.945202e-07,1.945204e-07,1.945206e-07,1.945208e-07,1.945209e-07,1.945211e-07,1.945213e-07,1.945215e-07,1.945217e-07,1.945219e-07,1.945221e-07,1.945222e-07,1.945224e-07,1.945226e-07,1.945228e-07,1.945230e-07,1.945232e-07,1.945234e-07,1.945235e-07,1.945237e-07,1.945239e-07,1.945241e-07,1.945243e-07,1.945245e-07,1.945247e-07,1.945249e-07,1.945250e-07,1.945252e-07,1.945254e-07,1.945256e-07,1.945258e-07,1.945260e-07,1.945262e-07,1.945263e-07,1.945265e-07,1.945267e-07,1.945269e-07,1.945271e-07,1.945273e-07,1.945275e-07,1.945276e-07,1.945278e-07,1.945280e-07,1.945282e-07,1.945284e-07,1.945286e-07,1.945288e-07,1.945290e-07,1.945291e-07,1.945293e-07,1.945295e-07,1.945297e-07,1.945299e-07,1.945301e-07,1.945303e-07,1.945304e-07,1.945306e-07,1.945308e-07,1.945310e-07,1.945312e-07,1.945314e-07,1.945316e-07,1.945317e-07,1.945319e-07,1.945321e-07,1.945323e-07,1.945325e-07,1.945327e-07,1.945329e-07,1.945331e-07,1.945332e-07,1.945334e-07,1.945336e-07,1.945338e-07,1.945340e-07,1.945342e-07,1.945344e-07,1.945345e-07,1.945347e-07,1.945349e-07,1.945351e-07,1.945353e-07,1.945355e-07,1.945357e-07,1.945358e-07,1.945360e-07,1.945362e-07,1.945364e-07,1.945366e-07,1.945368e-07,1.945370e-07,1.945372e-07,1.945373e-07,1.945375e-07,1.945377e-07,1.945379e-07,1.945381e-07,1.945383e-07,1.945385e-07,1.945386e-07,1.945388e-07,1.945390e-07,1.945392e-07,1.945394e-07,1.945396e-07,1.945398e-07,1.945399e-07,1.945401e-07,1.945403e-07,1.945405e-07,1.945407e-07,1.945409e-07,1.945411e-07,1.945412e-07,1.945414e-07,1.945416e-07,1.945418e-07,1.945420e-07,1.945422e-07,1.945424e-07,1.945426e-07,1.945427e-07,1.945429e-07,1.945431e-07,1.945433e-07,1.945435e-07,1.945437e-07,1.945439e-07,1.945440e-07,1.945442e-07,1.945444e-07,1.945446e-07,1.945448e-07,1.945450e-07,1.945452e-07,1.945453e-07,1.945455e-07,1.945457e-07,1.945459e-07,1.945461e-07,1.945463e-07,1.945465e-07,1.945466e-07,1.945468e-07,1.945470e-07,1.945472e-07,1.945474e-07,1.945476e-07,1.945478e-07,1.945479e-07,1.945481e-07,1.945483e-07,1.945485e-07,1.945487e-07,1.945489e-07,1.945491e-07,1.945493e-07,1.945494e-07,1.945496e-07,1.945498e-07,1.945500e-07,1.945502e-07,1.945504e-07,1.945506e-07,1.945507e-07,1.945509e-07,1.945511e-07,1.945513e-07,1.945515e-07,1.945517e-07,1.945519e-07,1.945520e-07,1.945522e-07,1.945524e-07,1.945526e-07,1.945528e-07,1.945530e-07,1.945532e-07,1.945533e-07,1.945535e-07,1.945537e-07,1.945539e-07,1.945541e-07,1.945543e-07,1.945545e-07,1.945546e-07,1.945548e-07,1.945550e-07,1.945552e-07,1.945554e-07,1.945556e-07,1.945558e-07,1.945559e-07,1.945561e-07,1.945563e-07,1.945565e-07,1.945567e-07,1.945569e-07,1.945571e-07,1.945572e-07,1.945574e-07,1.945576e-07,1.945578e-07,1.945580e-07,1.945582e-07,1.945584e-07,1.945586e-07,1.945587e-07,1.945589e-07,1.945591e-07,1.945593e-07,1.945595e-07,1.945597e-07,1.945599e-07,1.945600e-07,1.945602e-07,1.945604e-07,1.945606e-07,1.945608e-07,1.945610e-07,1.945612e-07,1.945613e-07,1.945615e-07,1.945617e-07,1.945619e-07,1.945621e-07,1.945623e-07,1.945625e-07,1.945626e-07,1.945628e-07,1.945630e-07,1.945632e-07,1.945634e-07,1.945636e-07,1.945638e-07,1.945639e-07,1.945641e-07,1.945643e-07,1.945645e-07,1.945647e-07,1.945649e-07,1.945651e-07,1.945652e-07,1.945654e-07,1.945656e-07,1.945658e-07,1.945660e-07,1.945662e-07,1.945664e-07,1.945665e-07,1.945667e-07,1.945669e-07,1.945671e-07,1.945673e-07,1.945675e-07,1.945677e-07,1.945678e-07,1.945680e-07,1.945682e-07,1.945684e-07,1.945686e-07,1.945688e-07,1.945690e-07,1.945691e-07,1.945693e-07,1.945695e-07,1.945697e-07,1.945699e-07,1.945701e-07,1.945703e-07,1.945704e-07,1.945706e-07,1.945708e-07,1.945710e-07,1.945712e-07,1.945714e-07,1.945716e-07,1.945717e-07,1.945719e-07,1.945721e-07,1.945723e-07,1.945725e-07,1.945727e-07,1.945729e-07,1.945730e-07,1.945732e-07,1.945734e-07,1.945736e-07,1.945738e-07,1.945740e-07,1.945742e-07,1.945743e-07,1.945745e-07,1.945747e-07,1.945749e-07,1.945751e-07,1.945753e-07,1.945755e-07,1.945756e-07,1.945758e-07,1.945760e-07,1.945762e-07,1.945764e-07,1.945766e-07,1.945768e-07,1.945769e-07,1.945771e-07,1.945773e-07,1.945775e-07,1.945777e-07,1.945779e-07,1.945781e-07,1.945782e-07,1.945784e-07,1.945786e-07,1.945788e-07,1.945790e-07,1.945792e-07,1.945794e-07,1.945795e-07,1.945797e-07,1.945799e-07,1.945801e-07,1.945803e-07,1.945805e-07,1.945807e-07,1.945808e-07,1.945810e-07,1.945812e-07,1.945814e-07,1.945816e-07,1.945818e-07,1.945820e-07,1.945821e-07,1.945823e-07,1.945825e-07,1.945827e-07,1.945829e-07,1.945831e-07,1.945833e-07,1.945834e-07,1.945836e-07,1.945838e-07,1.945840e-07,1.945842e-07,1.945844e-07,1.945845e-07,1.945847e-07,1.945849e-07,1.945851e-07,1.945853e-07,1.945855e-07,1.945857e-07,1.945858e-07,1.945860e-07,1.945862e-07,1.945864e-07,1.945866e-07,1.945868e-07,1.945870e-07,1.945871e-07,1.945873e-07,1.945875e-07,1.945877e-07,1.945879e-07,1.945881e-07,1.945883e-07,1.945884e-07,1.945886e-07,1.945888e-07,1.945890e-07,1.945892e-07,1.945894e-07,1.945896e-07,1.945897e-07,1.945899e-07,1.945901e-07,1.945903e-07,1.945905e-07,1.945907e-07,1.945909e-07,1.945910e-07,1.945912e-07,1.945914e-07,1.945916e-07,1.945918e-07,1.945920e-07,1.945922e-07,1.945923e-07,1.945925e-07,1.945927e-07,1.945929e-07,1.945931e-07,1.945933e-07,1.945935e-07,1.945936e-07,1.945938e-07,1.945940e-07,1.945942e-07,1.945944e-07,1.945946e-07,1.945947e-07,1.945949e-07,1.945951e-07,1.945953e-07,1.945955e-07,1.945957e-07,1.945959e-07,1.945960e-07,1.945962e-07,1.945964e-07,1.945966e-07,1.945968e-07,1.945970e-07,1.945972e-07,1.945973e-07,1.945975e-07,1.945977e-07,1.945979e-07,1.945981e-07,1.945983e-07,1.945985e-07,1.945986e-07,1.945988e-07,1.945990e-07,1.945992e-07,1.945994e-07,1.945996e-07,1.945998e-07,1.945999e-07,1.946001e-07,1.946003e-07,1.946005e-07,1.946007e-07,1.946009e-07,1.946010e-07,1.946012e-07,1.946014e-07,1.946016e-07,1.946018e-07,1.946020e-07,1.946022e-07,1.946023e-07,1.946025e-07,1.946027e-07,1.946029e-07,1.946031e-07,1.946033e-07,1.946035e-07,1.946036e-07,1.946038e-07,1.946040e-07,1.946042e-07,1.946044e-07,1.946046e-07,1.946048e-07,1.946049e-07,1.946051e-07,1.946053e-07,1.946055e-07,1.946057e-07,1.946059e-07,1.946060e-07,1.946062e-07,1.946064e-07,1.946066e-07,1.946068e-07,1.946070e-07,1.946072e-07,1.946073e-07,1.946075e-07,1.946077e-07,1.946079e-07,1.946081e-07,1.946083e-07,1.946085e-07,1.946086e-07,1.946088e-07,1.946090e-07,1.946092e-07,1.946094e-07,1.946096e-07,1.946098e-07,1.946099e-07,1.946101e-07,1.946103e-07,1.946105e-07,1.946107e-07,1.946109e-07,1.946110e-07,1.946112e-07,1.946114e-07,1.946116e-07,1.946118e-07,1.946120e-07,1.946122e-07,1.946123e-07,1.946125e-07,1.946127e-07,1.946129e-07,1.946131e-07,1.946133e-07,1.946135e-07,1.946136e-07,1.946138e-07,1.946140e-07,1.946142e-07,1.946144e-07,1.946146e-07,1.946147e-07,1.946149e-07,1.946151e-07,1.946153e-07,1.946155e-07,1.946157e-07,1.946159e-07,1.946160e-07,1.946162e-07,1.946164e-07,1.946166e-07,1.946168e-07,1.946170e-07,1.946172e-07,1.946173e-07,1.946175e-07,1.946177e-07,1.946179e-07,1.946181e-07,1.946183e-07,1.946184e-07,1.946186e-07,1.946188e-07,1.946190e-07,1.946192e-07,1.946194e-07,1.946196e-07,1.946197e-07,1.946199e-07,1.946201e-07,1.946203e-07,1.946205e-07,1.946207e-07,1.946209e-07,1.946210e-07,1.946212e-07,1.946214e-07,1.946216e-07,1.946218e-07,1.946220e-07,1.946221e-07,1.946223e-07,1.946225e-07,1.946227e-07,1.946229e-07,1.946231e-07,1.946233e-07,1.946234e-07,1.946236e-07,1.946238e-07,1.946240e-07,1.946242e-07,1.946244e-07,1.946245e-07,1.946247e-07,1.946249e-07,1.946251e-07,1.946253e-07,1.946255e-07,1.946257e-07,1.946258e-07,1.946260e-07,1.946262e-07,1.946264e-07,1.946266e-07,1.946268e-07,1.946270e-07,1.946271e-07,1.946273e-07,1.946275e-07,1.946277e-07,1.946279e-07,1.946281e-07,1.946282e-07,1.946284e-07,1.946286e-07,1.946288e-07,1.946290e-07,1.946292e-07,1.946294e-07,1.946295e-07,1.946297e-07,1.946299e-07,1.946301e-07,1.946303e-07,1.946305e-07,1.946306e-07,1.946308e-07,1.946310e-07,1.946312e-07,1.946314e-07,1.946316e-07,1.946318e-07,1.946319e-07,1.946321e-07,1.946323e-07,1.946325e-07,1.946327e-07,1.946329e-07,1.946330e-07,1.946332e-07,1.946334e-07,1.946336e-07,1.946338e-07,1.946340e-07,1.946342e-07,1.946343e-07,1.946345e-07,1.946347e-07,1.946349e-07,1.946351e-07,1.946353e-07,1.946355e-07,1.946356e-07,1.946358e-07,1.946360e-07,1.946362e-07,1.946364e-07,1.946366e-07,1.946367e-07,1.946369e-07,1.946371e-07,1.946373e-07,1.946375e-07,1.946377e-07,1.946379e-07,1.946380e-07,1.946382e-07,1.946384e-07,1.946386e-07,1.946388e-07,1.946390e-07,1.946391e-07,1.946393e-07,1.946395e-07,1.946397e-07,1.946399e-07,1.946401e-07,1.946403e-07,1.946404e-07,1.946406e-07,1.946408e-07,1.946410e-07,1.946412e-07,1.946414e-07,1.946415e-07,1.946417e-07,1.946419e-07,1.946421e-07,1.946423e-07,1.946425e-07,1.946427e-07,1.946428e-07,1.946430e-07,1.946432e-07,1.946434e-07,1.946436e-07,1.946438e-07,1.946439e-07,1.946441e-07,1.946443e-07,1.946445e-07,1.946447e-07,1.946449e-07,1.946451e-07,1.946452e-07,1.946454e-07,1.946456e-07,1.946458e-07,1.946460e-07,1.946462e-07,1.946463e-07,1.946465e-07,1.946467e-07,1.946469e-07,1.946471e-07,1.946473e-07,1.946474e-07,1.946476e-07,1.946478e-07,1.946480e-07,1.946482e-07,1.946484e-07,1.946486e-07,1.946487e-07,1.946489e-07,1.946491e-07,1.946493e-07,1.946495e-07,1.946497e-07,1.946498e-07,1.946500e-07,1.946502e-07,1.946504e-07,1.946506e-07,1.946508e-07,1.946510e-07,1.946511e-07,1.946513e-07,1.946515e-07,1.946517e-07,1.946519e-07,1.946521e-07,1.946522e-07,1.946524e-07,1.946526e-07,1.946528e-07,1.946530e-07,1.946532e-07,1.946534e-07,1.946535e-07,1.946537e-07,1.946539e-07,1.946541e-07,1.946543e-07,1.946545e-07,1.946546e-07,1.946548e-07,1.946550e-07,1.946552e-07,1.946554e-07,1.946556e-07,1.946557e-07,1.946559e-07,1.946561e-07,1.946563e-07,1.946565e-07,1.946567e-07,1.946569e-07,1.946570e-07,1.946572e-07,1.946574e-07,1.946576e-07,1.946578e-07,1.946580e-07,1.946581e-07,1.946583e-07,1.946585e-07,1.946587e-07,1.946589e-07,1.946591e-07,1.946593e-07,1.946594e-07,1.946596e-07,1.946598e-07,1.946600e-07,1.946602e-07,1.946604e-07,1.946605e-07,1.946607e-07,1.946609e-07,1.946611e-07,1.946613e-07,1.946615e-07,1.946616e-07,1.946618e-07,1.946620e-07,1.946622e-07,1.946624e-07,1.946626e-07,1.946628e-07,1.946629e-07,1.946631e-07,1.946633e-07,1.946635e-07,1.946637e-07,1.946639e-07,1.946640e-07,1.946642e-07,1.946644e-07,1.946646e-07,1.946648e-07,1.946650e-07,1.946651e-07,1.946653e-07,1.946655e-07,1.946657e-07,1.946659e-07,1.946661e-07,1.946663e-07,1.946664e-07,1.946666e-07,1.946668e-07,1.946670e-07,1.946672e-07,1.946674e-07,1.946675e-07,1.946677e-07,1.946679e-07,1.946681e-07,1.946683e-07,1.946685e-07,1.946686e-07,1.946688e-07,1.946690e-07,1.946692e-07,1.946694e-07,1.946696e-07,1.946698e-07,1.946699e-07,1.946701e-07,1.946703e-07,1.946705e-07,1.946707e-07,1.946709e-07,1.946710e-07,1.946712e-07,1.946714e-07,1.946716e-07,1.946718e-07,1.946720e-07,1.946721e-07,1.946723e-07,1.946725e-07,1.946727e-07,1.946729e-07,1.946731e-07,1.946733e-07,1.946734e-07,1.946736e-07,1.946738e-07,1.946740e-07,1.946742e-07,1.946744e-07,1.946745e-07,1.946747e-07,1.946749e-07,1.946751e-07,1.946753e-07,1.946755e-07,1.946756e-07,1.946758e-07,1.946760e-07,1.946762e-07,1.946764e-07,1.946766e-07,1.946767e-07,1.946769e-07,1.946771e-07,1.946773e-07,1.946775e-07,1.946777e-07,1.946779e-07,1.946780e-07,1.946782e-07,1.946784e-07,1.946786e-07,1.946788e-07,1.946790e-07,1.946791e-07,1.946793e-07,1.946795e-07,1.946797e-07,1.946799e-07,1.946801e-07,1.946802e-07,1.946804e-07,1.946806e-07,1.946808e-07,1.946810e-07,1.946812e-07,1.946813e-07,1.946815e-07,1.946817e-07,1.946819e-07,1.946821e-07,1.946823e-07,1.946825e-07,1.946826e-07,1.946828e-07,1.946830e-07,1.946832e-07,1.946834e-07,1.946836e-07,1.946837e-07,1.946839e-07,1.946841e-07,1.946843e-07,1.946845e-07,1.946847e-07,1.946848e-07,1.946850e-07,1.946852e-07,1.946854e-07,1.946856e-07,1.946858e-07,1.946859e-07,1.946861e-07,1.946863e-07,1.946865e-07,1.946867e-07,1.946869e-07,1.946871e-07,1.946872e-07,1.946874e-07,1.946876e-07,1.946878e-07,1.946880e-07,1.946882e-07,1.946883e-07,1.946885e-07,1.946887e-07,1.946889e-07,1.946891e-07,1.946893e-07,1.946894e-07,1.946896e-07,1.946898e-07,1.946900e-07,1.946902e-07,1.946904e-07,1.946905e-07,1.946907e-07,1.946909e-07,1.946911e-07,1.946913e-07,1.946915e-07,1.946916e-07,1.946918e-07,1.946920e-07,1.946922e-07,1.946924e-07,1.946926e-07,1.946927e-07,1.946929e-07,1.946931e-07,1.946933e-07,1.946935e-07,1.946937e-07,1.946939e-07,1.946940e-07,1.946942e-07,1.946944e-07,1.946946e-07,1.946948e-07,1.946950e-07,1.946951e-07,1.946953e-07,1.946955e-07,1.946957e-07,1.946959e-07,1.946961e-07,1.946962e-07,1.946964e-07,1.946966e-07,1.946968e-07,1.946970e-07,1.946972e-07,1.946973e-07,1.946975e-07,1.946977e-07,1.946979e-07,1.946981e-07,1.946983e-07,1.946984e-07,1.946986e-07,1.946988e-07,1.946990e-07,1.946992e-07,1.946994e-07,1.946995e-07,1.946997e-07,1.946999e-07,1.947001e-07,1.947003e-07,1.947005e-07,1.947006e-07,1.947008e-07,1.947010e-07,1.947012e-07,1.947014e-07,1.947016e-07,1.947018e-07,1.947019e-07,1.947021e-07,1.947023e-07,1.947025e-07,1.947027e-07,1.947029e-07,1.947030e-07,1.947032e-07,1.947034e-07,1.947036e-07,1.947038e-07,1.947040e-07,1.947041e-07,1.947043e-07,1.947045e-07,1.947047e-07,1.947049e-07,1.947051e-07,1.947052e-07,1.947054e-07,1.947056e-07,1.947058e-07,1.947060e-07,1.947062e-07,1.947063e-07,1.947065e-07,1.947067e-07,1.947069e-07,1.947071e-07,1.947073e-07,1.947074e-07,1.947076e-07,1.947078e-07,1.947080e-07,1.947082e-07,1.947084e-07,1.947085e-07,1.947087e-07,1.947089e-07,1.947091e-07,1.947093e-07,1.947095e-07,1.947096e-07,1.947098e-07,1.947100e-07,1.947102e-07,1.947104e-07,1.947106e-07,1.947107e-07,1.947109e-07,1.947111e-07,1.947113e-07,1.947115e-07,1.947117e-07,1.947118e-07,1.947120e-07,1.947122e-07,1.947124e-07,1.947126e-07,1.947128e-07,1.947129e-07,1.947131e-07,1.947133e-07,1.947135e-07,1.947137e-07,1.947139e-07,1.947140e-07,1.947142e-07,1.947144e-07,1.947146e-07,1.947148e-07,1.947150e-07,1.947151e-07,1.947153e-07,1.947155e-07,1.947157e-07,1.947159e-07,1.947161e-07,1.947163e-07,1.947164e-07,1.947166e-07,1.947168e-07,1.947170e-07,1.947172e-07,1.947174e-07,1.947175e-07,1.947177e-07,1.947179e-07,1.947181e-07,1.947183e-07,1.947185e-07,1.947186e-07,1.947188e-07,1.947190e-07,1.947192e-07,1.947194e-07,1.947196e-07,1.947197e-07,1.947199e-07,1.947201e-07,1.947203e-07,1.947205e-07,1.947207e-07,1.947208e-07,1.947210e-07,1.947212e-07,1.947214e-07,1.947216e-07,1.947218e-07,1.947219e-07,1.947221e-07,1.947223e-07,1.947225e-07,1.947227e-07,1.947229e-07,1.947230e-07,1.947232e-07,1.947234e-07,1.947236e-07,1.947238e-07,1.947240e-07,1.947241e-07,1.947243e-07,1.947245e-07,1.947247e-07,1.947249e-07,1.947251e-07,1.947252e-07,1.947254e-07,1.947256e-07,1.947258e-07,1.947260e-07,1.947262e-07,1.947263e-07,1.947265e-07,1.947267e-07,1.947269e-07,1.947271e-07,1.947273e-07,1.947274e-07,1.947276e-07,1.947278e-07,1.947280e-07,1.947282e-07,1.947284e-07,1.947285e-07,1.947287e-07,1.947289e-07,1.947291e-07,1.947293e-07,1.947294e-07,1.947296e-07,1.947298e-07,1.947300e-07,1.947302e-07,1.947304e-07,1.947305e-07,1.947307e-07,1.947309e-07,1.947311e-07,1.947313e-07,1.947315e-07,1.947316e-07,1.947318e-07,1.947320e-07,1.947322e-07,1.947324e-07,1.947326e-07,1.947327e-07,1.947329e-07,1.947331e-07,1.947333e-07,1.947335e-07,1.947337e-07,1.947338e-07,1.947340e-07,1.947342e-07,1.947344e-07,1.947346e-07,1.947348e-07,1.947349e-07,1.947351e-07,1.947353e-07,1.947355e-07,1.947357e-07,1.947359e-07,1.947360e-07,1.947362e-07,1.947364e-07,1.947366e-07,1.947368e-07,1.947370e-07,1.947371e-07,1.947373e-07,1.947375e-07,1.947377e-07,1.947379e-07,1.947381e-07,1.947382e-07,1.947384e-07,1.947386e-07,1.947388e-07,1.947390e-07,1.947392e-07,1.947393e-07,1.947395e-07,1.947397e-07,1.947399e-07,1.947401e-07,1.947403e-07,1.947404e-07,1.947406e-07,1.947408e-07,1.947410e-07,1.947412e-07,1.947414e-07,1.947415e-07,1.947417e-07,1.947419e-07,1.947421e-07,1.947423e-07,1.947425e-07,1.947426e-07,1.947428e-07,1.947430e-07,1.947432e-07,1.947434e-07,1.947435e-07,1.947437e-07,1.947439e-07,1.947441e-07,1.947443e-07,1.947445e-07,1.947446e-07,1.947448e-07,1.947450e-07,1.947452e-07,1.947454e-07,1.947456e-07,1.947457e-07,1.947459e-07,1.947461e-07,1.947463e-07,1.947465e-07,1.947467e-07,1.947468e-07,1.947470e-07,1.947472e-07,1.947474e-07,1.947476e-07,1.947478e-07,1.947479e-07,1.947481e-07,1.947483e-07,1.947485e-07,1.947487e-07,1.947489e-07,1.947490e-07,1.947492e-07,1.947494e-07,1.947496e-07,1.947498e-07,1.947500e-07,1.947501e-07,1.947503e-07,1.947505e-07,1.947507e-07,1.947509e-07,1.947510e-07,1.947512e-07,1.947514e-07,1.947516e-07,1.947518e-07,1.947520e-07,1.947521e-07,1.947523e-07,1.947525e-07,1.947527e-07,1.947529e-07,1.947531e-07,1.947532e-07,1.947534e-07,1.947536e-07,1.947538e-07,1.947540e-07,1.947542e-07,1.947543e-07,1.947545e-07,1.947547e-07,1.947549e-07,1.947551e-07,1.947553e-07,1.947554e-07,1.947556e-07,1.947558e-07,1.947560e-07,1.947562e-07,1.947564e-07,1.947565e-07,1.947567e-07,1.947569e-07,1.947571e-07,1.947573e-07,1.947574e-07,1.947576e-07,1.947578e-07,1.947580e-07,1.947582e-07,1.947584e-07,1.947585e-07,1.947587e-07,1.947589e-07,1.947591e-07,1.947593e-07,1.947595e-07,1.947596e-07,1.947598e-07,1.947600e-07,1.947602e-07,1.947604e-07,1.947606e-07,1.947607e-07,1.947609e-07,1.947611e-07,1.947613e-07,1.947615e-07,1.947617e-07,1.947618e-07,1.947620e-07,1.947622e-07,1.947624e-07,1.947626e-07,1.947627e-07,1.947629e-07,1.947631e-07,1.947633e-07,1.947635e-07,1.947637e-07,1.947638e-07,1.947640e-07,1.947642e-07,1.947644e-07,1.947646e-07,1.947648e-07,1.947649e-07,1.947651e-07,1.947653e-07,1.947655e-07,1.947657e-07,1.947659e-07,1.947660e-07,1.947662e-07,1.947664e-07,1.947666e-07,1.947668e-07,1.947669e-07,1.947671e-07,1.947673e-07,1.947675e-07,1.947677e-07,1.947679e-07,1.947680e-07,1.947682e-07,1.947684e-07,1.947686e-07,1.947688e-07,1.947690e-07,1.947691e-07,1.947693e-07,1.947695e-07,1.947697e-07,1.947699e-07,1.947701e-07,1.947702e-07,1.947704e-07,1.947706e-07,1.947708e-07,1.947710e-07,1.947711e-07,1.947713e-07,1.947715e-07,1.947717e-07,1.947719e-07,1.947721e-07,1.947722e-07,1.947724e-07,1.947726e-07,1.947728e-07,1.947730e-07,1.947732e-07,1.947733e-07,1.947735e-07,1.947737e-07,1.947739e-07,1.947741e-07,1.947743e-07,1.947744e-07,1.947746e-07,1.947748e-07,1.947750e-07,1.947752e-07,1.947753e-07,1.947755e-07,1.947757e-07,1.947759e-07,1.947761e-07,1.947763e-07,1.947764e-07,1.947766e-07,1.947768e-07,1.947770e-07,1.947772e-07,1.947774e-07,1.947775e-07,1.947777e-07,1.947779e-07,1.947781e-07,1.947783e-07,1.947784e-07,1.947786e-07,1.947788e-07,1.947790e-07,1.947792e-07,1.947794e-07,1.947795e-07,1.947797e-07,1.947799e-07,1.947801e-07,1.947803e-07,1.947805e-07,1.947806e-07,1.947808e-07,1.947810e-07,1.947812e-07,1.947814e-07,1.947815e-07,1.947817e-07,1.947819e-07,1.947821e-07,1.947823e-07,1.947825e-07,1.947826e-07,1.947828e-07,1.947830e-07,1.947832e-07,1.947834e-07,1.947836e-07,1.947837e-07,1.947839e-07,1.947841e-07,1.947843e-07,1.947845e-07,1.947846e-07,1.947848e-07,1.947850e-07,1.947852e-07,1.947854e-07,1.947856e-07,1.947857e-07,1.947859e-07,1.947861e-07,1.947863e-07,1.947865e-07,1.947867e-07,1.947868e-07,1.947870e-07,1.947872e-07,1.947874e-07,1.947876e-07,1.947877e-07,1.947879e-07,1.947881e-07,1.947883e-07,1.947885e-07,1.947887e-07,1.947888e-07,1.947890e-07,1.947892e-07,1.947894e-07,1.947896e-07,1.947898e-07,1.947899e-07,1.947901e-07,1.947903e-07,1.947905e-07,1.947907e-07,1.947908e-07,1.947910e-07,1.947912e-07,1.947914e-07,1.947916e-07,1.947918e-07,1.947919e-07,1.947921e-07,1.947923e-07,1.947925e-07,1.947927e-07,1.947929e-07,1.947930e-07,1.947932e-07,1.947934e-07,1.947936e-07,1.947938e-07,1.947939e-07,1.947941e-07,1.947943e-07,1.947945e-07,1.947947e-07,1.947949e-07,1.947950e-07,1.947952e-07,1.947954e-07,1.947956e-07,1.947958e-07,1.947960e-07,1.947961e-07,1.947963e-07,1.947965e-07,1.947967e-07,1.947969e-07,1.947970e-07,1.947972e-07,1.947974e-07,1.947976e-07,1.947978e-07,1.947980e-07,1.947981e-07,1.947983e-07,1.947985e-07,1.947987e-07,1.947989e-07,1.947990e-07,1.947992e-07,1.947994e-07,1.947996e-07,1.947998e-07,1.948000e-07,1.948001e-07,1.948003e-07,1.948005e-07,1.948007e-07,1.948009e-07,1.948011e-07,1.948012e-07,1.948014e-07,1.948016e-07,1.948018e-07,1.948020e-07,1.948021e-07,1.948023e-07,1.948025e-07,1.948027e-07,1.948029e-07,1.948031e-07,1.948032e-07,1.948034e-07,1.948036e-07,1.948038e-07,1.948040e-07,1.948041e-07,1.948043e-07,1.948045e-07,1.948047e-07,1.948049e-07,1.948051e-07,1.948052e-07,1.948054e-07,1.948056e-07,1.948058e-07,1.948060e-07,1.948061e-07,1.948063e-07,1.948065e-07,1.948067e-07,1.948069e-07,1.948071e-07,1.948072e-07,1.948074e-07,1.948076e-07,1.948078e-07,1.948080e-07,1.948081e-07,1.948083e-07,1.948085e-07,1.948087e-07,1.948089e-07,1.948091e-07,1.948092e-07,1.948094e-07,1.948096e-07,1.948098e-07,1.948100e-07,1.948102e-07,1.948103e-07,1.948105e-07,1.948107e-07,1.948109e-07,1.948111e-07,1.948112e-07,1.948114e-07,1.948116e-07,1.948118e-07,1.948120e-07,1.948122e-07,1.948123e-07,1.948125e-07,1.948127e-07,1.948129e-07,1.948131e-07,1.948132e-07,1.948134e-07,1.948136e-07,1.948138e-07,1.948140e-07,1.948142e-07,1.948143e-07,1.948145e-07,1.948147e-07,1.948149e-07,1.948151e-07,1.948152e-07,1.948154e-07,1.948156e-07,1.948158e-07,1.948160e-07,1.948162e-07,1.948163e-07,1.948165e-07,1.948167e-07,1.948169e-07,1.948171e-07,1.948172e-07,1.948174e-07,1.948176e-07,1.948178e-07,1.948180e-07,1.948182e-07,1.948183e-07,1.948185e-07,1.948187e-07,1.948189e-07,1.948191e-07,1.948192e-07,1.948194e-07,1.948196e-07,1.948198e-07,1.948200e-07,1.948202e-07,1.948203e-07,1.948205e-07,1.948207e-07,1.948209e-07,1.948211e-07,1.948212e-07,1.948214e-07,1.948216e-07,1.948218e-07,1.948220e-07,1.948222e-07,1.948223e-07,1.948225e-07,1.948227e-07,1.948229e-07,1.948231e-07,1.948232e-07,1.948234e-07,1.948236e-07,1.948238e-07,1.948240e-07,1.948242e-07,1.948243e-07,1.948245e-07,1.948247e-07,1.948249e-07,1.948251e-07,1.948252e-07,1.948254e-07,1.948256e-07,1.948258e-07,1.948260e-07,1.948262e-07,1.948263e-07,1.948265e-07,1.948267e-07,1.948269e-07,1.948271e-07,1.948272e-07,1.948274e-07,1.948276e-07,1.948278e-07,1.948280e-07,1.948282e-07,1.948283e-07,1.948285e-07,1.948287e-07,1.948289e-07,1.948291e-07,1.948292e-07,1.948294e-07,1.948296e-07,1.948298e-07,1.948300e-07,1.948301e-07,1.948303e-07,1.948305e-07,1.948307e-07,1.948309e-07,1.948311e-07,1.948312e-07,1.948314e-07,1.948316e-07,1.948318e-07,1.948320e-07,1.948321e-07,1.948323e-07,1.948325e-07,1.948327e-07,1.948329e-07,1.948331e-07,1.948332e-07,1.948334e-07,1.948336e-07,1.948338e-07,1.948340e-07,1.948341e-07,1.948343e-07,1.948345e-07,1.948347e-07,1.948349e-07,1.948351e-07,1.948352e-07,1.948354e-07,1.948356e-07,1.948358e-07,1.948360e-07,1.948361e-07,1.948363e-07,1.948365e-07,1.948367e-07,1.948369e-07,1.948371e-07,1.948372e-07,1.948374e-07,1.948376e-07,1.948378e-07,1.948380e-07,1.948381e-07,1.948383e-07,1.948385e-07,1.948387e-07,1.948389e-07,1.948390e-07,1.948392e-07,1.948394e-07,1.948396e-07,1.948398e-07,1.948400e-07,1.948401e-07,1.948403e-07,1.948405e-07,1.948407e-07,1.948409e-07,1.948410e-07,1.948412e-07,1.948414e-07,1.948416e-07,1.948418e-07,1.948420e-07,1.948421e-07,1.948423e-07,1.948425e-07,1.948427e-07,1.948429e-07,1.948430e-07,1.948432e-07,1.948434e-07,1.948436e-07,1.948438e-07,1.948439e-07,1.948441e-07,1.948443e-07,1.948445e-07,1.948447e-07,1.948449e-07,1.948450e-07,1.948452e-07,1.948454e-07,1.948456e-07,1.948458e-07,1.948459e-07,1.948461e-07,1.948463e-07,1.948465e-07,1.948467e-07,1.948468e-07,1.948470e-07,1.948472e-07,1.948474e-07,1.948476e-07,1.948478e-07,1.948479e-07,1.948481e-07,1.948483e-07,1.948485e-07,1.948487e-07,1.948488e-07,1.948490e-07,1.948492e-07,1.948494e-07,1.948496e-07,1.948498e-07,1.948499e-07,1.948501e-07,1.948503e-07,1.948505e-07,1.948507e-07,1.948508e-07,1.948510e-07,1.948512e-07,1.948514e-07,1.948516e-07,1.948517e-07,1.948519e-07,1.948521e-07,1.948523e-07,1.948525e-07,1.948527e-07,1.948528e-07,1.948530e-07,1.948532e-07,1.948534e-07,1.948536e-07,1.948537e-07,1.948539e-07,1.948541e-07,1.948543e-07,1.948545e-07,1.948546e-07,1.948548e-07,1.948550e-07,1.948552e-07,1.948554e-07,1.948556e-07,1.948557e-07,1.948559e-07,1.948561e-07,1.948563e-07,1.948565e-07,1.948566e-07,1.948568e-07,1.948570e-07,1.948572e-07,1.948574e-07,1.948575e-07,1.948577e-07,1.948579e-07,1.948581e-07,1.948583e-07,1.948585e-07,1.948586e-07,1.948588e-07,1.948590e-07,1.948592e-07,1.948594e-07,1.948595e-07,1.948597e-07,1.948599e-07,1.948601e-07,1.948603e-07,1.948604e-07,1.948606e-07,1.948608e-07,1.948610e-07,1.948612e-07,1.948614e-07,1.948615e-07,1.948617e-07,1.948619e-07,1.948621e-07,1.948623e-07,1.948624e-07,1.948626e-07,1.948628e-07,1.948630e-07,1.948632e-07,1.948633e-07,1.948635e-07,1.948637e-07,1.948639e-07,1.948641e-07,1.948642e-07,1.948644e-07,1.948646e-07,1.948648e-07,1.948650e-07,1.948652e-07,1.948653e-07,1.948655e-07,1.948657e-07,1.948659e-07,1.948661e-07,1.948662e-07,1.948664e-07,1.948666e-07,1.948668e-07,1.948670e-07,1.948671e-07,1.948673e-07,1.948675e-07,1.948677e-07,1.948679e-07,1.948681e-07,1.948682e-07,1.948684e-07,1.948686e-07,1.948688e-07,1.948690e-07,1.948691e-07,1.948693e-07,1.948695e-07,1.948697e-07,1.948699e-07,1.948700e-07,1.948702e-07,1.948704e-07,1.948706e-07,1.948708e-07,1.948709e-07,1.948711e-07,1.948713e-07,1.948715e-07,1.948717e-07,1.948719e-07,1.948720e-07,1.948722e-07,1.948724e-07,1.948726e-07,1.948728e-07,1.948729e-07,1.948731e-07,1.948733e-07,1.948735e-07,1.948737e-07,1.948738e-07,1.948740e-07,1.948742e-07,1.948744e-07,1.948746e-07,1.948747e-07,1.948749e-07,1.948751e-07,1.948753e-07,1.948755e-07,1.948757e-07,1.948758e-07,1.948760e-07,1.948762e-07,1.948764e-07,1.948766e-07,1.948767e-07,1.948769e-07,1.948771e-07,1.948773e-07,1.948775e-07,1.948776e-07,1.948778e-07,1.948780e-07,1.948782e-07,1.948784e-07,1.948785e-07,1.948787e-07,1.948789e-07,1.948791e-07,1.948793e-07,1.948795e-07,1.948796e-07,1.948798e-07,1.948800e-07,1.948802e-07,1.948804e-07,1.948805e-07,1.948807e-07,1.948809e-07,1.948811e-07,1.948813e-07,1.948814e-07,1.948816e-07,1.948818e-07,1.948820e-07,1.948822e-07,1.948823e-07,1.948825e-07,1.948827e-07,1.948829e-07,1.948831e-07,1.948833e-07,1.948834e-07,1.948836e-07,1.948838e-07,1.948840e-07,1.948842e-07,1.948843e-07,1.948845e-07,1.948847e-07,1.948849e-07,1.948851e-07,1.948852e-07,1.948854e-07,1.948856e-07,1.948858e-07,1.948860e-07,1.948861e-07,1.948863e-07,1.948865e-07,1.948867e-07,1.948869e-07,1.948870e-07,1.948872e-07,1.948874e-07,1.948876e-07,1.948878e-07,1.948880e-07,1.948881e-07,1.948883e-07,1.948885e-07,1.948887e-07,1.948889e-07,1.948890e-07,1.948892e-07,1.948894e-07,1.948896e-07,1.948898e-07,1.948899e-07,1.948901e-07,1.948903e-07,1.948905e-07,1.948907e-07,1.948908e-07,1.948910e-07,1.948912e-07,1.948914e-07,1.948916e-07,1.948917e-07,1.948919e-07,1.948921e-07,1.948923e-07,1.948925e-07,1.948927e-07,1.948928e-07,1.948930e-07,1.948932e-07,1.948934e-07,1.948936e-07,1.948937e-07,1.948939e-07,1.948941e-07,1.948943e-07,1.948945e-07,1.948946e-07,1.948948e-07,1.948950e-07,1.948952e-07,1.948954e-07,1.948955e-07,1.948957e-07,1.948959e-07,1.948961e-07,1.948963e-07,1.948964e-07,1.948966e-07,1.948968e-07,1.948970e-07,1.948972e-07,1.948973e-07,1.948975e-07,1.948977e-07,1.948979e-07,1.948981e-07,1.948982e-07,1.948984e-07,1.948986e-07,1.948988e-07,1.948990e-07,1.948992e-07,1.948993e-07,1.948995e-07,1.948997e-07,1.948999e-07,1.949001e-07,1.949002e-07,1.949004e-07,1.949006e-07,1.949008e-07,1.949010e-07,1.949011e-07,1.949013e-07,1.949015e-07,1.949017e-07,1.949019e-07,1.949020e-07,1.949022e-07,1.949024e-07,1.949026e-07,1.949028e-07,1.949029e-07,1.949031e-07,1.949033e-07,1.949035e-07,1.949037e-07,1.949038e-07,1.949040e-07,1.949042e-07,1.949044e-07,1.949046e-07,1.949047e-07,1.949049e-07,1.949051e-07,1.949053e-07,1.949055e-07,1.949057e-07,1.949058e-07,1.949060e-07,1.949062e-07,1.949064e-07,1.949066e-07,1.949067e-07,1.949069e-07,1.949071e-07,1.949073e-07,1.949075e-07,1.949076e-07,1.949078e-07,1.949080e-07,1.949082e-07,1.949084e-07,1.949085e-07,1.949087e-07,1.949089e-07,1.949091e-07,1.949093e-07,1.949094e-07,1.949096e-07,1.949098e-07,1.949100e-07,1.949102e-07,1.949103e-07,1.949105e-07,1.949107e-07,1.949109e-07,1.949111e-07,1.949112e-07,1.949114e-07,1.949116e-07,1.949118e-07,1.949120e-07,1.949121e-07,1.949123e-07,1.949125e-07,1.949127e-07,1.949129e-07,1.949130e-07,1.949132e-07,1.949134e-07,1.949136e-07,1.949138e-07,1.949140e-07,1.949141e-07,1.949143e-07,1.949145e-07,1.949147e-07,1.949149e-07,1.949150e-07,1.949152e-07,1.949154e-07,1.949156e-07,1.949158e-07,1.949159e-07,1.949161e-07,1.949163e-07,1.949165e-07,1.949167e-07,1.949168e-07,1.949170e-07,1.949172e-07,1.949174e-07,1.949176e-07,1.949177e-07,1.949179e-07,1.949181e-07,1.949183e-07,1.949185e-07,1.949186e-07,1.949188e-07,1.949190e-07,1.949192e-07,1.949194e-07,1.949195e-07,1.949197e-07,1.949199e-07,1.949201e-07,1.949203e-07,1.949204e-07,1.949206e-07,1.949208e-07,1.949210e-07,1.949212e-07,1.949213e-07,1.949215e-07,1.949217e-07,1.949219e-07,1.949221e-07,1.949222e-07,1.949224e-07,1.949226e-07,1.949228e-07,1.949230e-07,1.949231e-07,1.949233e-07,1.949235e-07,1.949237e-07,1.949239e-07,1.949240e-07,1.949242e-07,1.949244e-07,1.949246e-07,1.949248e-07,1.949249e-07,1.949251e-07,1.949253e-07,1.949255e-07,1.949257e-07,1.949258e-07,1.949260e-07,1.949262e-07,1.949264e-07,1.949266e-07,1.949267e-07,1.949269e-07,1.949271e-07,1.949273e-07,1.949275e-07,1.949276e-07,1.949278e-07,1.949280e-07,1.949282e-07,1.949284e-07,1.949286e-07,1.949287e-07,1.949289e-07,1.949291e-07,1.949293e-07,1.949295e-07,1.949296e-07,1.949298e-07,1.949300e-07,1.949302e-07,1.949304e-07,1.949305e-07,1.949307e-07,1.949309e-07,1.949311e-07,1.949313e-07,1.949314e-07,1.949316e-07,1.949318e-07,1.949320e-07,1.949322e-07,1.949323e-07,1.949325e-07,1.949327e-07,1.949329e-07,1.949331e-07,1.949332e-07,1.949334e-07,1.949336e-07,1.949338e-07,1.949340e-07,1.949341e-07,1.949343e-07,1.949345e-07,1.949347e-07,1.949349e-07,1.949350e-07,1.949352e-07,1.949354e-07,1.949356e-07,1.949358e-07,1.949359e-07,1.949361e-07,1.949363e-07,1.949365e-07,1.949367e-07,1.949368e-07,1.949370e-07,1.949372e-07,1.949374e-07,1.949376e-07,1.949377e-07,1.949379e-07,1.949381e-07,1.949383e-07,1.949385e-07,1.949386e-07,1.949388e-07,1.949390e-07,1.949392e-07,1.949394e-07,1.949395e-07,1.949397e-07,1.949399e-07,1.949401e-07,1.949403e-07,1.949404e-07,1.949406e-07,1.949408e-07,1.949410e-07,1.949412e-07,1.949413e-07,1.949415e-07,1.949417e-07,1.949419e-07,1.949421e-07,1.949422e-07,1.949424e-07,1.949426e-07,1.949428e-07,1.949430e-07,1.949431e-07,1.949433e-07,1.949435e-07,1.949437e-07,1.949439e-07,1.949440e-07,1.949442e-07,1.949444e-07,1.949446e-07,1.949448e-07,1.949449e-07,1.949451e-07,1.949453e-07,1.949455e-07,1.949456e-07,1.949458e-07,1.949460e-07,1.949462e-07,1.949464e-07,1.949465e-07,1.949467e-07,1.949469e-07,1.949471e-07,1.949473e-07,1.949474e-07,1.949476e-07,1.949478e-07,1.949480e-07,1.949482e-07,1.949483e-07,1.949485e-07,1.949487e-07,1.949489e-07,1.949491e-07,1.949492e-07,1.949494e-07,1.949496e-07,1.949498e-07,1.949500e-07,1.949501e-07,1.949503e-07,1.949505e-07,1.949507e-07,1.949509e-07,1.949510e-07,1.949512e-07,1.949514e-07,1.949516e-07,1.949518e-07,1.949519e-07,1.949521e-07,1.949523e-07,1.949525e-07,1.949527e-07,1.949528e-07,1.949530e-07,1.949532e-07,1.949534e-07,1.949536e-07,1.949537e-07,1.949539e-07,1.949541e-07,1.949543e-07,1.949545e-07,1.949546e-07,1.949548e-07,1.949550e-07,1.949552e-07,1.949554e-07,1.949555e-07,1.949557e-07,1.949559e-07,1.949561e-07,1.949563e-07,1.949564e-07,1.949566e-07,1.949568e-07,1.949570e-07,1.949572e-07,1.949573e-07,1.949575e-07,1.949577e-07,1.949579e-07,1.949581e-07,1.949582e-07,1.949584e-07,1.949586e-07,1.949588e-07,1.949590e-07,1.949591e-07,1.949593e-07,1.949595e-07,1.949597e-07,1.949599e-07,1.949600e-07,1.949602e-07,1.949604e-07,1.949606e-07,1.949607e-07,1.949609e-07,1.949611e-07,1.949613e-07,1.949615e-07,1.949616e-07,1.949618e-07,1.949620e-07,1.949622e-07,1.949624e-07,1.949625e-07,1.949627e-07,1.949629e-07,1.949631e-07,1.949633e-07,1.949634e-07,1.949636e-07,1.949638e-07,1.949640e-07,1.949642e-07,1.949643e-07,1.949645e-07,1.949647e-07,1.949649e-07,1.949651e-07,1.949652e-07,1.949654e-07,1.949656e-07,1.949658e-07,1.949660e-07,1.949661e-07,1.949663e-07,1.949665e-07,1.949667e-07,1.949669e-07,1.949670e-07,1.949672e-07,1.949674e-07,1.949676e-07,1.949678e-07,1.949679e-07,1.949681e-07,1.949683e-07,1.949685e-07,1.949686e-07,1.949688e-07,1.949690e-07,1.949692e-07,1.949694e-07,1.949695e-07,1.949697e-07,1.949699e-07,1.949701e-07,1.949703e-07,1.949704e-07,1.949706e-07,1.949708e-07,1.949710e-07,1.949712e-07,1.949713e-07,1.949715e-07,1.949717e-07,1.949719e-07,1.949721e-07,1.949722e-07,1.949724e-07,1.949726e-07,1.949728e-07,1.949730e-07,1.949731e-07,1.949733e-07,1.949735e-07,1.949737e-07,1.949739e-07,1.949740e-07,1.949742e-07,1.949744e-07,1.949746e-07,1.949748e-07,1.949749e-07,1.949751e-07,1.949753e-07,1.949755e-07,1.949756e-07,1.949758e-07,1.949760e-07,1.949762e-07,1.949764e-07,1.949765e-07,1.949767e-07,1.949769e-07,1.949771e-07,1.949773e-07,1.949774e-07,1.949776e-07,1.949778e-07,1.949780e-07,1.949782e-07,1.949783e-07,1.949785e-07,1.949787e-07,1.949789e-07,1.949791e-07,1.949792e-07,1.949794e-07,1.949796e-07,1.949798e-07,1.949800e-07,1.949801e-07,1.949803e-07,1.949805e-07,1.949807e-07,1.949808e-07,1.949810e-07,1.949812e-07,1.949814e-07,1.949816e-07,1.949817e-07,1.949819e-07,1.949821e-07,1.949823e-07,1.949825e-07,1.949826e-07,1.949828e-07,1.949830e-07,1.949832e-07,1.949834e-07,1.949835e-07,1.949837e-07,1.949839e-07,1.949841e-07,1.949843e-07,1.949844e-07,1.949846e-07,1.949848e-07,1.949850e-07,1.949852e-07,1.949853e-07,1.949855e-07,1.949857e-07,1.949859e-07,1.949860e-07,1.949862e-07,1.949864e-07,1.949866e-07,1.949868e-07,1.949869e-07,1.949871e-07,1.949873e-07,1.949875e-07,1.949877e-07,1.949878e-07,1.949880e-07,1.949882e-07,1.949884e-07,1.949886e-07,1.949887e-07,1.949889e-07,1.949891e-07,1.949893e-07,1.949895e-07,1.949896e-07,1.949898e-07,1.949900e-07,1.949902e-07,1.949903e-07,1.949905e-07,1.949907e-07,1.949909e-07,1.949911e-07,1.949912e-07,1.949914e-07,1.949916e-07,1.949918e-07,1.949920e-07,1.949921e-07,1.949923e-07,1.949925e-07,1.949927e-07,1.949929e-07,1.949930e-07,1.949932e-07,1.949934e-07,1.949936e-07,1.949938e-07,1.949939e-07,1.949941e-07,1.949943e-07,1.949945e-07,1.949946e-07,1.949948e-07,1.949950e-07,1.949952e-07,1.949954e-07,1.949955e-07,1.949957e-07,1.949959e-07,1.949961e-07,1.949963e-07,1.949964e-07,1.949966e-07,1.949968e-07,1.949970e-07,1.949972e-07,1.949973e-07,1.949975e-07,1.949977e-07,1.949979e-07,1.949981e-07,1.949982e-07,1.949984e-07,1.949986e-07,1.949988e-07,1.949989e-07,1.949991e-07,1.949993e-07,1.949995e-07,1.949997e-07,1.949998e-07,1.950000e-07,1.950002e-07,1.950004e-07,1.950006e-07,1.950007e-07,1.950009e-07,1.950011e-07,1.950013e-07,1.950015e-07,1.950016e-07,1.950018e-07,1.950020e-07,1.950022e-07,1.950023e-07,1.950025e-07,1.950027e-07,1.950029e-07,1.950031e-07,1.950032e-07,1.950034e-07,1.950036e-07,1.950038e-07,1.950040e-07,1.950041e-07,1.950043e-07,1.950045e-07,1.950047e-07,1.950049e-07,1.950050e-07,1.950052e-07,1.950054e-07,1.950056e-07,1.950057e-07,1.950059e-07,1.950061e-07,1.950063e-07,1.950065e-07,1.950066e-07,1.950068e-07,1.950070e-07,1.950072e-07,1.950074e-07,1.950075e-07,1.950077e-07,1.950079e-07,1.950081e-07,1.950083e-07,1.950084e-07,1.950086e-07,1.950088e-07,1.950090e-07,1.950091e-07,1.950093e-07,1.950095e-07,1.950097e-07,1.950099e-07,1.950100e-07,1.950102e-07,1.950104e-07,1.950106e-07,1.950108e-07,1.950109e-07,1.950111e-07,1.950113e-07,1.950115e-07,1.950117e-07,1.950118e-07,1.950120e-07,1.950122e-07,1.950124e-07,1.950125e-07,1.950127e-07,1.950129e-07,1.950131e-07,1.950133e-07,1.950134e-07,1.950136e-07,1.950138e-07,1.950140e-07,1.950142e-07,1.950143e-07,1.950145e-07,1.950147e-07,1.950149e-07,1.950151e-07,1.950152e-07,1.950154e-07,1.950156e-07,1.950158e-07,1.950159e-07,1.950161e-07,1.950163e-07,1.950165e-07,1.950167e-07,1.950168e-07,1.950170e-07,1.950172e-07,1.950174e-07,1.950176e-07,1.950177e-07,1.950179e-07,1.950181e-07,1.950183e-07,1.950184e-07,1.950186e-07,1.950188e-07,1.950190e-07,1.950192e-07,1.950193e-07,1.950195e-07,1.950197e-07,1.950199e-07,1.950201e-07,1.950202e-07,1.950204e-07,1.950206e-07,1.950208e-07,1.950209e-07,1.950211e-07,1.950213e-07,1.950215e-07,1.950217e-07,1.950218e-07,1.950220e-07,1.950222e-07,1.950224e-07,1.950226e-07,1.950227e-07,1.950229e-07,1.950231e-07,1.950233e-07,1.950235e-07,1.950236e-07,1.950238e-07,1.950240e-07,1.950242e-07,1.950243e-07,1.950245e-07,1.950247e-07,1.950249e-07,1.950251e-07,1.950252e-07,1.950254e-07,1.950256e-07,1.950258e-07,1.950260e-07,1.950261e-07,1.950263e-07,1.950265e-07,1.950267e-07,1.950268e-07,1.950270e-07,1.950272e-07,1.950274e-07,1.950276e-07,1.950277e-07,1.950279e-07,1.950281e-07,1.950283e-07,1.950285e-07,1.950286e-07,1.950288e-07,1.950290e-07,1.950292e-07,1.950293e-07,1.950295e-07,1.950297e-07,1.950299e-07,1.950301e-07,1.950302e-07,1.950304e-07,1.950306e-07,1.950308e-07,1.950310e-07,1.950311e-07,1.950313e-07,1.950315e-07,1.950317e-07,1.950318e-07,1.950320e-07,1.950322e-07,1.950324e-07,1.950326e-07,1.950327e-07,1.950329e-07,1.950331e-07,1.950333e-07,1.950335e-07,1.950336e-07,1.950338e-07,1.950340e-07,1.950342e-07,1.950343e-07,1.950345e-07,1.950347e-07,1.950349e-07,1.950351e-07,1.950352e-07,1.950354e-07,1.950356e-07,1.950358e-07,1.950360e-07,1.950361e-07,1.950363e-07,1.950365e-07,1.950367e-07,1.950368e-07,1.950370e-07,1.950372e-07,1.950374e-07,1.950376e-07,1.950377e-07,1.950379e-07,1.950381e-07,1.950383e-07,1.950384e-07,1.950386e-07,1.950388e-07,1.950390e-07,1.950392e-07,1.950393e-07,1.950395e-07,1.950397e-07,1.950399e-07,1.950401e-07,1.950402e-07,1.950404e-07,1.950406e-07,1.950408e-07,1.950409e-07,1.950411e-07,1.950413e-07,1.950415e-07,1.950417e-07,1.950418e-07,1.950420e-07,1.950422e-07,1.950424e-07,1.950426e-07,1.950427e-07,1.950429e-07,1.950431e-07,1.950433e-07,1.950434e-07,1.950436e-07,1.950438e-07,1.950440e-07,1.950442e-07,1.950443e-07,1.950445e-07,1.950447e-07,1.950449e-07,1.950451e-07,1.950452e-07,1.950454e-07,1.950456e-07,1.950458e-07,1.950459e-07,1.950461e-07,1.950463e-07,1.950465e-07,1.950467e-07,1.950468e-07,1.950470e-07,1.950472e-07,1.950474e-07,1.950475e-07,1.950477e-07,1.950479e-07,1.950481e-07,1.950483e-07,1.950484e-07,1.950486e-07,1.950488e-07,1.950490e-07,1.950492e-07,1.950493e-07,1.950495e-07,1.950497e-07,1.950499e-07,1.950500e-07,1.950502e-07,1.950504e-07,1.950506e-07,1.950508e-07,1.950509e-07,1.950511e-07,1.950513e-07,1.950515e-07,1.950516e-07,1.950518e-07,1.950520e-07,1.950522e-07,1.950524e-07,1.950525e-07,1.950527e-07,1.950529e-07,1.950531e-07,1.950533e-07,1.950534e-07,1.950536e-07,1.950538e-07,1.950540e-07,1.950541e-07,1.950543e-07,1.950545e-07,1.950547e-07,1.950549e-07,1.950550e-07,1.950552e-07,1.950554e-07,1.950556e-07,1.950557e-07,1.950559e-07,1.950561e-07,1.950563e-07,1.950565e-07,1.950566e-07,1.950568e-07,1.950570e-07,1.950572e-07,1.950573e-07,1.950575e-07,1.950577e-07,1.950579e-07,1.950581e-07,1.950582e-07,1.950584e-07,1.950586e-07,1.950588e-07,1.950590e-07,1.950591e-07,1.950593e-07,1.950595e-07,1.950597e-07,1.950598e-07,1.950600e-07,1.950602e-07,1.950604e-07,1.950606e-07,1.950607e-07,1.950609e-07,1.950611e-07,1.950613e-07,1.950614e-07,1.950616e-07,1.950618e-07,1.950620e-07,1.950622e-07,1.950623e-07,1.950625e-07,1.950627e-07,1.950629e-07,1.950630e-07,1.950632e-07,1.950634e-07,1.950636e-07,1.950638e-07,1.950639e-07,1.950641e-07,1.950643e-07,1.950645e-07,1.950647e-07,1.950648e-07,1.950650e-07,1.950652e-07,1.950654e-07,1.950655e-07,1.950657e-07,1.950659e-07,1.950661e-07,1.950663e-07,1.950664e-07,1.950666e-07,1.950668e-07,1.950670e-07,1.950671e-07,1.950673e-07,1.950675e-07,1.950677e-07,1.950679e-07,1.950680e-07,1.950682e-07,1.950684e-07,1.950686e-07,1.950687e-07,1.950689e-07,1.950691e-07,1.950693e-07,1.950695e-07,1.950696e-07,1.950698e-07,1.950700e-07,1.950702e-07,1.950703e-07,1.950705e-07,1.950707e-07,1.950709e-07,1.950711e-07,1.950712e-07,1.950714e-07,1.950716e-07,1.950718e-07,1.950719e-07,1.950721e-07,1.950723e-07,1.950725e-07,1.950727e-07,1.950728e-07,1.950730e-07,1.950732e-07,1.950734e-07,1.950736e-07,1.950737e-07,1.950739e-07,1.950741e-07,1.950743e-07,1.950744e-07,1.950746e-07,1.950748e-07,1.950750e-07,1.950752e-07,1.950753e-07,1.950755e-07,1.950757e-07,1.950759e-07,1.950760e-07,1.950762e-07,1.950764e-07,1.950766e-07,1.950768e-07,1.950769e-07,1.950771e-07,1.950773e-07,1.950775e-07,1.950776e-07,1.950778e-07,1.950780e-07,1.950782e-07,1.950784e-07,1.950785e-07,1.950787e-07,1.950789e-07,1.950791e-07,1.950792e-07,1.950794e-07,1.950796e-07,1.950798e-07,1.950800e-07,1.950801e-07,1.950803e-07,1.950805e-07,1.950807e-07,1.950808e-07,1.950810e-07,1.950812e-07,1.950814e-07,1.950816e-07,1.950817e-07,1.950819e-07,1.950821e-07,1.950823e-07,1.950824e-07,1.950826e-07,1.950828e-07,1.950830e-07,1.950832e-07,1.950833e-07,1.950835e-07,1.950837e-07,1.950839e-07,1.950840e-07,1.950842e-07,1.950844e-07,1.950846e-07,1.950848e-07,1.950849e-07,1.950851e-07,1.950853e-07,1.950855e-07,1.950856e-07,1.950858e-07,1.950860e-07,1.950862e-07,1.950864e-07,1.950865e-07,1.950867e-07,1.950869e-07,1.950871e-07,1.950872e-07,1.950874e-07,1.950876e-07,1.950878e-07,1.950880e-07,1.950881e-07,1.950883e-07,1.950885e-07,1.950887e-07,1.950888e-07,1.950890e-07,1.950892e-07,1.950894e-07,1.950896e-07,1.950897e-07,1.950899e-07,1.950901e-07,1.950903e-07,1.950904e-07,1.950906e-07,1.950908e-07,1.950910e-07,1.950911e-07,1.950913e-07,1.950915e-07,1.950917e-07,1.950919e-07,1.950920e-07,1.950922e-07,1.950924e-07,1.950926e-07,1.950927e-07,1.950929e-07,1.950931e-07,1.950933e-07,1.950935e-07,1.950936e-07,1.950938e-07,1.950940e-07,1.950942e-07,1.950943e-07,1.950945e-07,1.950947e-07,1.950949e-07,1.950951e-07,1.950952e-07,1.950954e-07,1.950956e-07,1.950958e-07,1.950959e-07,1.950961e-07,1.950963e-07,1.950965e-07,1.950967e-07,1.950968e-07,1.950970e-07,1.950972e-07,1.950974e-07,1.950975e-07,1.950977e-07,1.950979e-07,1.950981e-07,1.950983e-07,1.950984e-07,1.950986e-07,1.950988e-07,1.950990e-07,1.950991e-07,1.950993e-07,1.950995e-07,1.950997e-07,1.950999e-07,1.951000e-07,1.951002e-07,1.951004e-07,1.951006e-07,1.951007e-07,1.951009e-07,1.951011e-07,1.951013e-07,1.951014e-07,1.951016e-07,1.951018e-07,1.951020e-07,1.951022e-07,1.951023e-07,1.951025e-07,1.951027e-07,1.951029e-07,1.951030e-07,1.951032e-07,1.951034e-07,1.951036e-07,1.951038e-07,1.951039e-07,1.951041e-07,1.951043e-07,1.951045e-07,1.951046e-07,1.951048e-07,1.951050e-07,1.951052e-07,1.951054e-07,1.951055e-07,1.951057e-07,1.951059e-07,1.951061e-07,1.951062e-07,1.951064e-07,1.951066e-07,1.951068e-07,1.951069e-07,1.951071e-07,1.951073e-07,1.951075e-07,1.951077e-07,1.951078e-07,1.951080e-07,1.951082e-07,1.951084e-07,1.951085e-07,1.951087e-07,1.951089e-07,1.951091e-07,1.951093e-07,1.951094e-07,1.951096e-07,1.951098e-07,1.951100e-07,1.951101e-07,1.951103e-07,1.951105e-07,1.951107e-07,1.951109e-07,1.951110e-07,1.951112e-07,1.951114e-07,1.951116e-07,1.951117e-07,1.951119e-07,1.951121e-07,1.951123e-07,1.951124e-07,1.951126e-07,1.951128e-07,1.951130e-07,1.951132e-07,1.951133e-07,1.951135e-07,1.951137e-07,1.951139e-07,1.951140e-07,1.951142e-07,1.951144e-07,1.951146e-07,1.951148e-07,1.951149e-07,1.951151e-07,1.951153e-07,1.951155e-07,1.951156e-07,1.951158e-07,1.951160e-07,1.951162e-07,1.951163e-07,1.951165e-07,1.951167e-07,1.951169e-07,1.951171e-07,1.951172e-07,1.951174e-07,1.951176e-07,1.951178e-07,1.951179e-07,1.951181e-07,1.951183e-07,1.951185e-07,1.951187e-07,1.951188e-07,1.951190e-07,1.951192e-07,1.951194e-07,1.951195e-07,1.951197e-07,1.951199e-07,1.951201e-07,1.951202e-07,1.951204e-07,1.951206e-07,1.951208e-07,1.951210e-07,1.951211e-07,1.951213e-07,1.951215e-07,1.951217e-07,1.951218e-07,1.951220e-07,1.951222e-07,1.951224e-07,1.951226e-07,1.951227e-07,1.951229e-07,1.951231e-07,1.951233e-07,1.951234e-07,1.951236e-07,1.951238e-07,1.951240e-07,1.951241e-07,1.951243e-07,1.951245e-07,1.951247e-07,1.951249e-07,1.951250e-07,1.951252e-07,1.951254e-07,1.951256e-07,1.951257e-07,1.951259e-07,1.951261e-07,1.951263e-07,1.951264e-07,1.951266e-07,1.951268e-07,1.951270e-07,1.951272e-07,1.951273e-07,1.951275e-07,1.951277e-07,1.951279e-07,1.951280e-07,1.951282e-07,1.951284e-07,1.951286e-07,1.951287e-07,1.951289e-07,1.951291e-07,1.951293e-07,1.951295e-07,1.951296e-07,1.951298e-07,1.951300e-07,1.951302e-07,1.951303e-07,1.951305e-07,1.951307e-07,1.951309e-07,1.951311e-07,1.951312e-07,1.951314e-07,1.951316e-07,1.951318e-07,1.951319e-07,1.951321e-07,1.951323e-07,1.951325e-07,1.951326e-07,1.951328e-07,1.951330e-07,1.951332e-07,1.951334e-07,1.951335e-07,1.951337e-07,1.951339e-07,1.951341e-07,1.951342e-07,1.951344e-07,1.951346e-07,1.951348e-07,1.951349e-07,1.951351e-07,1.951353e-07,1.951355e-07,1.951357e-07,1.951358e-07,1.951360e-07,1.951362e-07,1.951364e-07,1.951365e-07,1.951367e-07,1.951369e-07,1.951371e-07,1.951372e-07,1.951374e-07,1.951376e-07,1.951378e-07,1.951380e-07,1.951381e-07,1.951383e-07,1.951385e-07,1.951387e-07,1.951388e-07,1.951390e-07,1.951392e-07,1.951394e-07,1.951395e-07,1.951397e-07,1.951399e-07,1.951401e-07,1.951403e-07,1.951404e-07,1.951406e-07,1.951408e-07,1.951410e-07,1.951411e-07,1.951413e-07,1.951415e-07,1.951417e-07,1.951418e-07,1.951420e-07,1.951422e-07,1.951424e-07,1.951426e-07,1.951427e-07,1.951429e-07,1.951431e-07,1.951433e-07,1.951434e-07,1.951436e-07,1.951438e-07,1.951440e-07,1.951441e-07,1.951443e-07,1.951445e-07,1.951447e-07,1.951449e-07,1.951450e-07,1.951452e-07,1.951454e-07,1.951456e-07,1.951457e-07,1.951459e-07,1.951461e-07,1.951463e-07,1.951464e-07,1.951466e-07,1.951468e-07,1.951470e-07,1.951472e-07,1.951473e-07,1.951475e-07,1.951477e-07,1.951479e-07,1.951480e-07,1.951482e-07,1.951484e-07,1.951486e-07,1.951487e-07,1.951489e-07,1.951491e-07,1.951493e-07,1.951494e-07,1.951496e-07,1.951498e-07,1.951500e-07,1.951502e-07,1.951503e-07,1.951505e-07,1.951507e-07,1.951509e-07,1.951510e-07,1.951512e-07,1.951514e-07,1.951516e-07,1.951517e-07,1.951519e-07,1.951521e-07,1.951523e-07,1.951525e-07,1.951526e-07,1.951528e-07,1.951530e-07,1.951532e-07,1.951533e-07,1.951535e-07,1.951537e-07,1.951539e-07,1.951540e-07,1.951542e-07,1.951544e-07,1.951546e-07,1.951547e-07,1.951549e-07,1.951551e-07,1.951553e-07,1.951555e-07,1.951556e-07,1.951558e-07,1.951560e-07,1.951562e-07,1.951563e-07,1.951565e-07,1.951567e-07,1.951569e-07,1.951570e-07,1.951572e-07,1.951574e-07,1.951576e-07,1.951578e-07,1.951579e-07,1.951581e-07,1.951583e-07,1.951585e-07,1.951586e-07,1.951588e-07,1.951590e-07,1.951592e-07,1.951593e-07,1.951595e-07,1.951597e-07,1.951599e-07,1.951600e-07,1.951602e-07,1.951604e-07,1.951606e-07,1.951608e-07,1.951609e-07,1.951611e-07,1.951613e-07,1.951615e-07,1.951616e-07,1.951618e-07,1.951620e-07,1.951622e-07,1.951623e-07,1.951625e-07,1.951627e-07,1.951629e-07,1.951631e-07,1.951632e-07,1.951634e-07,1.951636e-07,1.951638e-07,1.951639e-07,1.951641e-07,1.951643e-07,1.951645e-07,1.951646e-07,1.951648e-07,1.951650e-07,1.951652e-07,1.951653e-07,1.951655e-07,1.951657e-07,1.951659e-07,1.951661e-07,1.951662e-07,1.951664e-07,1.951666e-07,1.951668e-07,1.951669e-07,1.951671e-07,1.951673e-07,1.951675e-07,1.951676e-07,1.951678e-07,1.951680e-07,1.951682e-07,1.951683e-07,1.951685e-07,1.951687e-07,1.951689e-07,1.951691e-07,1.951692e-07,1.951694e-07,1.951696e-07,1.951698e-07,1.951699e-07,1.951701e-07,1.951703e-07,1.951705e-07,1.951706e-07,1.951708e-07,1.951710e-07,1.951712e-07,1.951713e-07,1.951715e-07,1.951717e-07,1.951719e-07,1.951721e-07,1.951722e-07,1.951724e-07,1.951726e-07,1.951728e-07,1.951729e-07,1.951731e-07,1.951733e-07,1.951735e-07,1.951736e-07,1.951738e-07,1.951740e-07,1.951742e-07,1.951743e-07,1.951745e-07,1.951747e-07,1.951749e-07,1.951751e-07,1.951752e-07,1.951754e-07,1.951756e-07,1.951758e-07,1.951759e-07,1.951761e-07,1.951763e-07,1.951765e-07,1.951766e-07,1.951768e-07,1.951770e-07,1.951772e-07,1.951773e-07,1.951775e-07,1.951777e-07,1.951779e-07,1.951780e-07,1.951782e-07,1.951784e-07,1.951786e-07,1.951788e-07,1.951789e-07,1.951791e-07,1.951793e-07,1.951795e-07,1.951796e-07,1.951798e-07,1.951800e-07,1.951802e-07,1.951803e-07,1.951805e-07,1.951807e-07,1.951809e-07,1.951810e-07,1.951812e-07,1.951814e-07,1.951816e-07,1.951818e-07,1.951819e-07,1.951821e-07,1.951823e-07,1.951825e-07,1.951826e-07,1.951828e-07,1.951830e-07,1.951832e-07,1.951833e-07,1.951835e-07,1.951837e-07,1.951839e-07,1.951840e-07,1.951842e-07,1.951844e-07,1.951846e-07,1.951847e-07,1.951849e-07,1.951851e-07,1.951853e-07,1.951855e-07,1.951856e-07,1.951858e-07,1.951860e-07,1.951862e-07,1.951863e-07,1.951865e-07,1.951867e-07,1.951869e-07,1.951870e-07,1.951872e-07,1.951874e-07,1.951876e-07,1.951877e-07,1.951879e-07,1.951881e-07,1.951883e-07,1.951884e-07,1.951886e-07,1.951888e-07,1.951890e-07,1.951892e-07,1.951893e-07,1.951895e-07,1.951897e-07,1.951899e-07,1.951900e-07,1.951902e-07,1.951904e-07,1.951906e-07,1.951907e-07,1.951909e-07,1.951911e-07,1.951913e-07,1.951914e-07,1.951916e-07,1.951918e-07,1.951920e-07,1.951921e-07,1.951923e-07,1.951925e-07,1.951927e-07,1.951929e-07,1.951930e-07,1.951932e-07,1.951934e-07,1.951936e-07,1.951937e-07,1.951939e-07,1.951941e-07,1.951943e-07,1.951944e-07,1.951946e-07,1.951948e-07,1.951950e-07,1.951951e-07,1.951953e-07,1.951955e-07,1.951957e-07,1.951958e-07,1.951960e-07,1.951962e-07,1.951964e-07,1.951965e-07,1.951967e-07,1.951969e-07,1.951971e-07,1.951973e-07,1.951974e-07,1.951976e-07,1.951978e-07,1.951980e-07,1.951981e-07,1.951983e-07,1.951985e-07,1.951987e-07,1.951988e-07,1.951990e-07,1.951992e-07,1.951994e-07,1.951995e-07,1.951997e-07,1.951999e-07,1.952001e-07,1.952002e-07,1.952004e-07,1.952006e-07,1.952008e-07,1.952009e-07,1.952011e-07,1.952013e-07,1.952015e-07,1.952017e-07,1.952018e-07,1.952020e-07,1.952022e-07,1.952024e-07,1.952025e-07,1.952027e-07,1.952029e-07,1.952031e-07,1.952032e-07,1.952034e-07,1.952036e-07,1.952038e-07,1.952039e-07,1.952041e-07,1.952043e-07,1.952045e-07,1.952046e-07,1.952048e-07,1.952050e-07,1.952052e-07,1.952053e-07,1.952055e-07,1.952057e-07,1.952059e-07,1.952061e-07,1.952062e-07,1.952064e-07,1.952066e-07,1.952068e-07,1.952069e-07,1.952071e-07,1.952073e-07,1.952075e-07,1.952076e-07,1.952078e-07,1.952080e-07,1.952082e-07,1.952083e-07,1.952085e-07,1.952087e-07,1.952089e-07,1.952090e-07,1.952092e-07,1.952094e-07,1.952096e-07,1.952097e-07,1.952099e-07,1.952101e-07,1.952103e-07,1.952104e-07,1.952106e-07,1.952108e-07,1.952110e-07,1.952112e-07,1.952113e-07,1.952115e-07,1.952117e-07,1.952119e-07,1.952120e-07,1.952122e-07,1.952124e-07,1.952126e-07,1.952127e-07,1.952129e-07,1.952131e-07,1.952133e-07,1.952134e-07,1.952136e-07,1.952138e-07,1.952140e-07,1.952141e-07,1.952143e-07,1.952145e-07,1.952147e-07,1.952148e-07,1.952150e-07,1.952152e-07,1.952154e-07,1.952155e-07,1.952157e-07,1.952159e-07,1.952161e-07,1.952162e-07,1.952164e-07,1.952166e-07,1.952168e-07,1.952170e-07,1.952171e-07,1.952173e-07,1.952175e-07,1.952177e-07,1.952178e-07,1.952180e-07,1.952182e-07,1.952184e-07,1.952185e-07,1.952187e-07,1.952189e-07,1.952191e-07,1.952192e-07,1.952194e-07,1.952196e-07,1.952198e-07,1.952199e-07,1.952201e-07,1.952203e-07,1.952205e-07,1.952206e-07,1.952208e-07,1.952210e-07,1.952212e-07,1.952213e-07,1.952215e-07,1.952217e-07,1.952219e-07,1.952220e-07,1.952222e-07,1.952224e-07,1.952226e-07,1.952227e-07,1.952229e-07,1.952231e-07,1.952233e-07,1.952235e-07,1.952236e-07,1.952238e-07,1.952240e-07,1.952242e-07,1.952243e-07,1.952245e-07,1.952247e-07,1.952249e-07,1.952250e-07,1.952252e-07,1.952254e-07,1.952256e-07,1.952257e-07,1.952259e-07,1.952261e-07,1.952263e-07,1.952264e-07,1.952266e-07,1.952268e-07,1.952270e-07,1.952271e-07,1.952273e-07,1.952275e-07,1.952277e-07,1.952278e-07,1.952280e-07,1.952282e-07,1.952284e-07,1.952285e-07,1.952287e-07,1.952289e-07,1.952291e-07,1.952292e-07,1.952294e-07,1.952296e-07,1.952298e-07,1.952299e-07,1.952301e-07,1.952303e-07,1.952305e-07,1.952307e-07,1.952308e-07,1.952310e-07,1.952312e-07,1.952314e-07,1.952315e-07,1.952317e-07,1.952319e-07,1.952321e-07,1.952322e-07,1.952324e-07,1.952326e-07,1.952328e-07,1.952329e-07,1.952331e-07,1.952333e-07,1.952335e-07,1.952336e-07,1.952338e-07,1.952340e-07,1.952342e-07,1.952343e-07,1.952345e-07,1.952347e-07,1.952349e-07,1.952350e-07,1.952352e-07,1.952354e-07,1.952356e-07,1.952357e-07,1.952359e-07,1.952361e-07,1.952363e-07,1.952364e-07,1.952366e-07,1.952368e-07,1.952370e-07,1.952371e-07,1.952373e-07,1.952375e-07,1.952377e-07,1.952378e-07,1.952380e-07,1.952382e-07,1.952384e-07,1.952385e-07,1.952387e-07,1.952389e-07,1.952391e-07,1.952392e-07,1.952394e-07,1.952396e-07,1.952398e-07,1.952400e-07,1.952401e-07,1.952403e-07,1.952405e-07,1.952407e-07,1.952408e-07,1.952410e-07,1.952412e-07,1.952414e-07,1.952415e-07,1.952417e-07,1.952419e-07,1.952421e-07,1.952422e-07,1.952424e-07,1.952426e-07,1.952428e-07,1.952429e-07,1.952431e-07,1.952433e-07,1.952435e-07,1.952436e-07,1.952438e-07,1.952440e-07,1.952442e-07,1.952443e-07,1.952445e-07,1.952447e-07,1.952449e-07,1.952450e-07,1.952452e-07,1.952454e-07,1.952456e-07,1.952457e-07,1.952459e-07,1.952461e-07,1.952463e-07,1.952464e-07,1.952466e-07,1.952468e-07,1.952470e-07,1.952471e-07,1.952473e-07,1.952475e-07,1.952477e-07,1.952478e-07,1.952480e-07,1.952482e-07,1.952484e-07,1.952485e-07,1.952487e-07,1.952489e-07,1.952491e-07,1.952492e-07,1.952494e-07,1.952496e-07,1.952498e-07,1.952499e-07,1.952501e-07,1.952503e-07,1.952505e-07,1.952506e-07,1.952508e-07,1.952510e-07,1.952512e-07,1.952513e-07,1.952515e-07,1.952517e-07,1.952519e-07,1.952520e-07,1.952522e-07,1.952524e-07,1.952526e-07,1.952527e-07,1.952529e-07,1.952531e-07,1.952533e-07,1.952534e-07,1.952536e-07,1.952538e-07,1.952540e-07,1.952542e-07,1.952543e-07,1.952545e-07,1.952547e-07,1.952549e-07,1.952550e-07,1.952552e-07,1.952554e-07,1.952556e-07,1.952557e-07,1.952559e-07,1.952561e-07,1.952563e-07,1.952564e-07,1.952566e-07,1.952568e-07,1.952570e-07,1.952571e-07,1.952573e-07,1.952575e-07,1.952577e-07,1.952578e-07,1.952580e-07,1.952582e-07,1.952584e-07,1.952585e-07,1.952587e-07,1.952589e-07,1.952591e-07,1.952592e-07,1.952594e-07,1.952596e-07,1.952598e-07,1.952599e-07,1.952601e-07,1.952603e-07,1.952605e-07,1.952606e-07,1.952608e-07,1.952610e-07,1.952612e-07,1.952613e-07,1.952615e-07,1.952617e-07,1.952619e-07,1.952620e-07,1.952622e-07,1.952624e-07,1.952626e-07,1.952627e-07,1.952629e-07,1.952631e-07,1.952633e-07,1.952634e-07,1.952636e-07,1.952638e-07,1.952640e-07,1.952641e-07,1.952643e-07,1.952645e-07,1.952647e-07,1.952648e-07,1.952650e-07,1.952652e-07,1.952654e-07,1.952655e-07,1.952657e-07,1.952659e-07,1.952661e-07,1.952662e-07,1.952664e-07,1.952666e-07,1.952668e-07,1.952669e-07,1.952671e-07,1.952673e-07,1.952675e-07,1.952676e-07,1.952678e-07,1.952680e-07,1.952682e-07,1.952683e-07,1.952685e-07,1.952687e-07,1.952689e-07,1.952690e-07,1.952692e-07,1.952694e-07,1.952696e-07,1.952697e-07,1.952699e-07,1.952701e-07,1.952703e-07,1.952704e-07,1.952706e-07,1.952708e-07,1.952710e-07,1.952711e-07,1.952713e-07,1.952715e-07,1.952717e-07,1.952718e-07,1.952720e-07,1.952722e-07,1.952724e-07,1.952725e-07,1.952727e-07,1.952729e-07,1.952731e-07,1.952732e-07,1.952734e-07,1.952736e-07,1.952738e-07,1.952739e-07,1.952741e-07,1.952743e-07,1.952745e-07,1.952746e-07,1.952748e-07,1.952750e-07,1.952752e-07,1.952753e-07,1.952755e-07,1.952757e-07,1.952759e-07,1.952760e-07,1.952762e-07,1.952764e-07,1.952766e-07,1.952767e-07,1.952769e-07,1.952771e-07,1.952773e-07,1.952774e-07,1.952776e-07,1.952778e-07,1.952780e-07,1.952781e-07,1.952783e-07,1.952785e-07,1.952787e-07,1.952788e-07,1.952790e-07,1.952792e-07,1.952793e-07,1.952795e-07,1.952797e-07,1.952799e-07,1.952800e-07,1.952802e-07,1.952804e-07,1.952806e-07,1.952807e-07,1.952809e-07,1.952811e-07,1.952813e-07,1.952814e-07,1.952816e-07,1.952818e-07,1.952820e-07,1.952821e-07,1.952823e-07,1.952825e-07,1.952827e-07,1.952828e-07,1.952830e-07,1.952832e-07,1.952834e-07,1.952835e-07,1.952837e-07,1.952839e-07,1.952841e-07,1.952842e-07,1.952844e-07,1.952846e-07,1.952848e-07,1.952849e-07,1.952851e-07,1.952853e-07,1.952855e-07,1.952856e-07,1.952858e-07,1.952860e-07,1.952862e-07,1.952863e-07,1.952865e-07,1.952867e-07,1.952869e-07,1.952870e-07,1.952872e-07,1.952874e-07,1.952876e-07,1.952877e-07,1.952879e-07,1.952881e-07,1.952883e-07,1.952884e-07,1.952886e-07,1.952888e-07,1.952890e-07,1.952891e-07,1.952893e-07,1.952895e-07,1.952897e-07,1.952898e-07,1.952900e-07,1.952902e-07,1.952904e-07,1.952905e-07,1.952907e-07,1.952909e-07,1.952911e-07,1.952912e-07,1.952914e-07,1.952916e-07,1.952918e-07,1.952919e-07,1.952921e-07,1.952923e-07,1.952925e-07,1.952926e-07,1.952928e-07,1.952930e-07,1.952932e-07,1.952933e-07,1.952935e-07,1.952937e-07,1.952938e-07,1.952940e-07,1.952942e-07,1.952944e-07,1.952945e-07,1.952947e-07,1.952949e-07,1.952951e-07,1.952952e-07,1.952954e-07,1.952956e-07,1.952958e-07,1.952959e-07,1.952961e-07,1.952963e-07,1.952965e-07,1.952966e-07,1.952968e-07,1.952970e-07,1.952972e-07,1.952973e-07,1.952975e-07,1.952977e-07,1.952979e-07,1.952980e-07,1.952982e-07,1.952984e-07,1.952986e-07,1.952987e-07,1.952989e-07,1.952991e-07,1.952993e-07,1.952994e-07,1.952996e-07,1.952998e-07,1.953000e-07,1.953001e-07,1.953003e-07,1.953005e-07,1.953007e-07,1.953008e-07,1.953010e-07,1.953012e-07,1.953014e-07,1.953015e-07,1.953017e-07,1.953019e-07,1.953021e-07,1.953022e-07,1.953024e-07,1.953026e-07,1.953028e-07,1.953029e-07,1.953031e-07,1.953033e-07,1.953034e-07,1.953036e-07,1.953038e-07,1.953040e-07,1.953041e-07,1.953043e-07,1.953045e-07,1.953047e-07,1.953048e-07,1.953050e-07,1.953052e-07,1.953054e-07,1.953055e-07,1.953057e-07,1.953059e-07,1.953061e-07,1.953062e-07,1.953064e-07,1.953066e-07,1.953068e-07,1.953069e-07,1.953071e-07,1.953073e-07,1.953075e-07,1.953076e-07,1.953078e-07,1.953080e-07,1.953082e-07,1.953083e-07,1.953085e-07,1.953087e-07,1.953089e-07,1.953090e-07,1.953092e-07,1.953094e-07,1.953096e-07,1.953097e-07,1.953099e-07,1.953101e-07,1.953102e-07,1.953104e-07,1.953106e-07,1.953108e-07,1.953109e-07,1.953111e-07,1.953113e-07,1.953115e-07,1.953116e-07,1.953118e-07,1.953120e-07,1.953122e-07,1.953123e-07,1.953125e-07,1.953127e-07,1.953129e-07,1.953130e-07,1.953132e-07,1.953134e-07,1.953136e-07,1.953137e-07,1.953139e-07,1.953141e-07,1.953143e-07,1.953144e-07,1.953146e-07,1.953148e-07,1.953150e-07,1.953151e-07,1.953153e-07,1.953155e-07,1.953157e-07,1.953158e-07,1.953160e-07,1.953162e-07,1.953164e-07,1.953165e-07,1.953167e-07,1.953169e-07,1.953170e-07,1.953172e-07,1.953174e-07,1.953176e-07,1.953177e-07,1.953179e-07,1.953181e-07,1.953183e-07,1.953184e-07,1.953186e-07,1.953188e-07,1.953190e-07,1.953191e-07,1.953193e-07,1.953195e-07,1.953197e-07,1.953198e-07,1.953200e-07,1.953202e-07,1.953204e-07,1.953205e-07,1.953207e-07,1.953209e-07,1.953211e-07,1.953212e-07,1.953214e-07,1.953216e-07,1.953218e-07,1.953219e-07,1.953221e-07,1.953223e-07,1.953224e-07,1.953226e-07,1.953228e-07,1.953230e-07,1.953231e-07,1.953233e-07,1.953235e-07,1.953237e-07,1.953238e-07,1.953240e-07,1.953242e-07,1.953244e-07,1.953245e-07,1.953247e-07,1.953249e-07,1.953251e-07,1.953252e-07,1.953254e-07,1.953256e-07,1.953258e-07,1.953259e-07,1.953261e-07,1.953263e-07,1.953265e-07,1.953266e-07,1.953268e-07,1.953270e-07,1.953271e-07,1.953273e-07,1.953275e-07,1.953277e-07,1.953278e-07,1.953280e-07,1.953282e-07,1.953284e-07,1.953285e-07,1.953287e-07,1.953289e-07,1.953291e-07,1.953292e-07,1.953294e-07,1.953296e-07,1.953298e-07,1.953299e-07,1.953301e-07,1.953303e-07,1.953305e-07,1.953306e-07,1.953308e-07,1.953310e-07,1.953312e-07,1.953313e-07,1.953315e-07,1.953317e-07,1.953318e-07,1.953320e-07,1.953322e-07,1.953324e-07,1.953325e-07,1.953327e-07,1.953329e-07,1.953331e-07,1.953332e-07,1.953334e-07,1.953336e-07,1.953338e-07,1.953339e-07,1.953341e-07,1.953343e-07,1.953345e-07,1.953346e-07,1.953348e-07,1.953350e-07,1.953352e-07,1.953353e-07,1.953355e-07,1.953357e-07,1.953359e-07,1.953360e-07,1.953362e-07,1.953364e-07,1.953365e-07,1.953367e-07,1.953369e-07,1.953371e-07,1.953372e-07,1.953374e-07,1.953376e-07,1.953378e-07,1.953379e-07,1.953381e-07,1.953383e-07,1.953385e-07,1.953386e-07,1.953388e-07,1.953390e-07,1.953392e-07,1.953393e-07,1.953395e-07,1.953397e-07,1.953399e-07,1.953400e-07,1.953402e-07,1.953404e-07,1.953405e-07,1.953407e-07,1.953409e-07,1.953411e-07,1.953412e-07,1.953414e-07,1.953416e-07,1.953418e-07,1.953419e-07,1.953421e-07,1.953423e-07,1.953425e-07,1.953426e-07,1.953428e-07,1.953430e-07,1.953432e-07,1.953433e-07,1.953435e-07,1.953437e-07,1.953439e-07,1.953440e-07,1.953442e-07,1.953444e-07,1.953445e-07,1.953447e-07,1.953449e-07,1.953451e-07,1.953452e-07,1.953454e-07,1.953456e-07,1.953458e-07,1.953459e-07,1.953461e-07,1.953463e-07,1.953465e-07,1.953466e-07,1.953468e-07,1.953470e-07,1.953472e-07,1.953473e-07,1.953475e-07,1.953477e-07,1.953478e-07,1.953480e-07,1.953482e-07,1.953484e-07,1.953485e-07,1.953487e-07,1.953489e-07,1.953491e-07,1.953492e-07,1.953494e-07,1.953496e-07,1.953498e-07,1.953499e-07,1.953501e-07,1.953503e-07,1.953505e-07,1.953506e-07,1.953508e-07,1.953510e-07,1.953512e-07,1.953513e-07,1.953515e-07,1.953517e-07,1.953518e-07,1.953520e-07,1.953522e-07,1.953524e-07,1.953525e-07,1.953527e-07,1.953529e-07,1.953531e-07,1.953532e-07,1.953534e-07,1.953536e-07,1.953538e-07,1.953539e-07,1.953541e-07,1.953543e-07,1.953545e-07,1.953546e-07,1.953548e-07,1.953550e-07,1.953551e-07,1.953553e-07,1.953555e-07,1.953557e-07,1.953558e-07,1.953560e-07,1.953562e-07,1.953564e-07,1.953565e-07,1.953567e-07,1.953569e-07,1.953571e-07,1.953572e-07,1.953574e-07,1.953576e-07,1.953578e-07,1.953579e-07,1.953581e-07,1.953583e-07,1.953584e-07,1.953586e-07,1.953588e-07,1.953590e-07,1.953591e-07,1.953593e-07,1.953595e-07,1.953597e-07,1.953598e-07,1.953600e-07,1.953602e-07,1.953604e-07,1.953605e-07,1.953607e-07,1.953609e-07,1.953610e-07,1.953612e-07,1.953614e-07,1.953616e-07,1.953617e-07,1.953619e-07,1.953621e-07,1.953623e-07,1.953624e-07,1.953626e-07,1.953628e-07,1.953630e-07,1.953631e-07,1.953633e-07,1.953635e-07,1.953637e-07,1.953638e-07,1.953640e-07,1.953642e-07,1.953643e-07,1.953645e-07,1.953647e-07,1.953649e-07,1.953650e-07,1.953652e-07,1.953654e-07,1.953656e-07,1.953657e-07,1.953659e-07,1.953661e-07,1.953663e-07,1.953664e-07,1.953666e-07,1.953668e-07,1.953669e-07,1.953671e-07,1.953673e-07,1.953675e-07,1.953676e-07,1.953678e-07,1.953680e-07,1.953682e-07,1.953683e-07,1.953685e-07,1.953687e-07,1.953689e-07,1.953690e-07,1.953692e-07,1.953694e-07,1.953696e-07,1.953697e-07,1.953699e-07,1.953701e-07,1.953702e-07,1.953704e-07,1.953706e-07,1.953708e-07,1.953709e-07,1.953711e-07,1.953713e-07,1.953715e-07,1.953716e-07,1.953718e-07,1.953720e-07,1.953722e-07,1.953723e-07,1.953725e-07,1.953727e-07,1.953728e-07,1.953730e-07,1.953732e-07,1.953734e-07,1.953735e-07,1.953737e-07,1.953739e-07,1.953741e-07,1.953742e-07,1.953744e-07,1.953746e-07,1.953748e-07,1.953749e-07,1.953751e-07,1.953753e-07,1.953754e-07,1.953756e-07,1.953758e-07,1.953760e-07,1.953761e-07,1.953763e-07,1.953765e-07,1.953767e-07,1.953768e-07,1.953770e-07,1.953772e-07,1.953774e-07,1.953775e-07,1.953777e-07,1.953779e-07,1.953780e-07,1.953782e-07,1.953784e-07,1.953786e-07,1.953787e-07,1.953789e-07,1.953791e-07,1.953793e-07,1.953794e-07,1.953796e-07,1.953798e-07,1.953800e-07,1.953801e-07,1.953803e-07,1.953805e-07,1.953806e-07,1.953808e-07,1.953810e-07,1.953812e-07,1.953813e-07,1.953815e-07,1.953817e-07,1.953819e-07,1.953820e-07,1.953822e-07,1.953824e-07,1.953826e-07,1.953827e-07,1.953829e-07,1.953831e-07,1.953832e-07,1.953834e-07,1.953836e-07,1.953838e-07,1.953839e-07,1.953841e-07,1.953843e-07,1.953845e-07,1.953846e-07,1.953848e-07,1.953850e-07,1.953852e-07,1.953853e-07,1.953855e-07,1.953857e-07,1.953858e-07,1.953860e-07,1.953862e-07,1.953864e-07,1.953865e-07,1.953867e-07,1.953869e-07,1.953871e-07,1.953872e-07,1.953874e-07,1.953876e-07,1.953878e-07,1.953879e-07,1.953881e-07,1.953883e-07,1.953884e-07,1.953886e-07,1.953888e-07,1.953890e-07,1.953891e-07,1.953893e-07,1.953895e-07,1.953897e-07,1.953898e-07,1.953900e-07,1.953902e-07,1.953903e-07,1.953905e-07,1.953907e-07,1.953909e-07,1.953910e-07,1.953912e-07,1.953914e-07,1.953916e-07,1.953917e-07,1.953919e-07,1.953921e-07,1.953923e-07,1.953924e-07,1.953926e-07,1.953928e-07,1.953929e-07,1.953931e-07,1.953933e-07,1.953935e-07,1.953936e-07,1.953938e-07,1.953940e-07,1.953942e-07,1.953943e-07,1.953945e-07,1.953947e-07,1.953949e-07,1.953950e-07,1.953952e-07,1.953954e-07,1.953955e-07,1.953957e-07,1.953959e-07,1.953961e-07,1.953962e-07,1.953964e-07,1.953966e-07,1.953968e-07,1.953969e-07,1.953971e-07,1.953973e-07,1.953974e-07,1.953976e-07,1.953978e-07,1.953980e-07,1.953981e-07,1.953983e-07,1.953985e-07,1.953987e-07,1.953988e-07,1.953990e-07,1.953992e-07,1.953994e-07,1.953995e-07,1.953997e-07,1.953999e-07,1.954000e-07,1.954002e-07,1.954004e-07,1.954006e-07,1.954007e-07,1.954009e-07,1.954011e-07,1.954013e-07,1.954014e-07,1.954016e-07,1.954018e-07,1.954019e-07,1.954021e-07,1.954023e-07,1.954025e-07,1.954026e-07,1.954028e-07,1.954030e-07,1.954032e-07,1.954033e-07,1.954035e-07,1.954037e-07,1.954038e-07,1.954040e-07,1.954042e-07,1.954044e-07,1.954045e-07,1.954047e-07,1.954049e-07,1.954051e-07,1.954052e-07,1.954054e-07,1.954056e-07,1.954058e-07,1.954059e-07,1.954061e-07,1.954063e-07,1.954064e-07,1.954066e-07,1.954068e-07,1.954070e-07,1.954071e-07,1.954073e-07,1.954075e-07,1.954077e-07,1.954078e-07,1.954080e-07,1.954082e-07,1.954083e-07,1.954085e-07,1.954087e-07,1.954089e-07,1.954090e-07,1.954092e-07,1.954094e-07,1.954096e-07,1.954097e-07,1.954099e-07,1.954101e-07,1.954102e-07,1.954104e-07,1.954106e-07,1.954108e-07,1.954109e-07,1.954111e-07,1.954113e-07,1.954115e-07,1.954116e-07,1.954118e-07,1.954120e-07,1.954121e-07,1.954123e-07,1.954125e-07,1.954127e-07,1.954128e-07,1.954130e-07,1.954132e-07,1.954134e-07,1.954135e-07,1.954137e-07,1.954139e-07,1.954140e-07,1.954142e-07,1.954144e-07,1.954146e-07,1.954147e-07,1.954149e-07,1.954151e-07,1.954153e-07,1.954154e-07,1.954156e-07,1.954158e-07,1.954159e-07,1.954161e-07,1.954163e-07,1.954165e-07,1.954166e-07,1.954168e-07,1.954170e-07,1.954172e-07,1.954173e-07,1.954175e-07,1.954177e-07,1.954178e-07,1.954180e-07,1.954182e-07,1.954184e-07,1.954185e-07,1.954187e-07,1.954189e-07,1.954191e-07,1.954192e-07,1.954194e-07,1.954196e-07,1.954197e-07,1.954199e-07,1.954201e-07,1.954203e-07,1.954204e-07,1.954206e-07,1.954208e-07,1.954210e-07,1.954211e-07,1.954213e-07,1.954215e-07,1.954216e-07,1.954218e-07,1.954220e-07,1.954222e-07,1.954223e-07,1.954225e-07,1.954227e-07,1.954229e-07,1.954230e-07,1.954232e-07,1.954234e-07,1.954235e-07,1.954237e-07,1.954239e-07,1.954241e-07,1.954242e-07,1.954244e-07,1.954246e-07,1.954248e-07,1.954249e-07,1.954251e-07,1.954253e-07,1.954254e-07,1.954256e-07,1.954258e-07,1.954260e-07,1.954261e-07,1.954263e-07,1.954265e-07,1.954267e-07,1.954268e-07,1.954270e-07,1.954272e-07,1.954273e-07,1.954275e-07,1.954277e-07,1.954279e-07,1.954280e-07,1.954282e-07,1.954284e-07,1.954286e-07,1.954287e-07,1.954289e-07,1.954291e-07,1.954292e-07,1.954294e-07,1.954296e-07,1.954298e-07,1.954299e-07,1.954301e-07,1.954303e-07,1.954305e-07,1.954306e-07,1.954308e-07,1.954310e-07,1.954311e-07,1.954313e-07,1.954315e-07,1.954317e-07,1.954318e-07,1.954320e-07,1.954322e-07,1.954324e-07,1.954325e-07,1.954327e-07,1.954329e-07,1.954330e-07,1.954332e-07,1.954334e-07,1.954336e-07,1.954337e-07,1.954339e-07,1.954341e-07,1.954342e-07,1.954344e-07,1.954346e-07,1.954348e-07,1.954349e-07,1.954351e-07,1.954353e-07,1.954355e-07,1.954356e-07,1.954358e-07,1.954360e-07,1.954361e-07,1.954363e-07,1.954365e-07,1.954367e-07,1.954368e-07,1.954370e-07,1.954372e-07,1.954374e-07,1.954375e-07,1.954377e-07,1.954379e-07,1.954380e-07,1.954382e-07,1.954384e-07,1.954386e-07,1.954387e-07,1.954389e-07,1.954391e-07,1.954393e-07,1.954394e-07,1.954396e-07,1.954398e-07,1.954399e-07,1.954401e-07,1.954403e-07,1.954405e-07,1.954406e-07,1.954408e-07,1.954410e-07,1.954411e-07,1.954413e-07,1.954415e-07,1.954417e-07,1.954418e-07,1.954420e-07,1.954422e-07,1.954424e-07,1.954425e-07,1.954427e-07,1.954429e-07,1.954430e-07,1.954432e-07,1.954434e-07,1.954436e-07,1.954437e-07,1.954439e-07,1.954441e-07,1.954443e-07,1.954444e-07,1.954446e-07,1.954448e-07,1.954449e-07,1.954451e-07,1.954453e-07,1.954455e-07,1.954456e-07,1.954458e-07,1.954460e-07,1.954461e-07,1.954463e-07,1.954465e-07,1.954467e-07,1.954468e-07,1.954470e-07,1.954472e-07,1.954474e-07,1.954475e-07,1.954477e-07,1.954479e-07,1.954480e-07,1.954482e-07,1.954484e-07,1.954486e-07,1.954487e-07,1.954489e-07,1.954491e-07,1.954492e-07,1.954494e-07,1.954496e-07,1.954498e-07,1.954499e-07,1.954501e-07,1.954503e-07,1.954505e-07,1.954506e-07,1.954508e-07,1.954510e-07,1.954511e-07,1.954513e-07,1.954515e-07,1.954517e-07,1.954518e-07,1.954520e-07,1.954522e-07,1.954523e-07,1.954525e-07,1.954527e-07,1.954529e-07,1.954530e-07,1.954532e-07,1.954534e-07,1.954536e-07,1.954537e-07,1.954539e-07,1.954541e-07,1.954542e-07,1.954544e-07,1.954546e-07,1.954548e-07,1.954549e-07,1.954551e-07,1.954553e-07,1.954554e-07,1.954556e-07,1.954558e-07,1.954560e-07,1.954561e-07,1.954563e-07,1.954565e-07,1.954567e-07,1.954568e-07,1.954570e-07,1.954572e-07,1.954573e-07,1.954575e-07,1.954577e-07,1.954579e-07,1.954580e-07,1.954582e-07,1.954584e-07,1.954585e-07,1.954587e-07,1.954589e-07,1.954591e-07,1.954592e-07,1.954594e-07,1.954596e-07,1.954598e-07,1.954599e-07,1.954601e-07,1.954603e-07,1.954604e-07,1.954606e-07,1.954608e-07,1.954610e-07,1.954611e-07,1.954613e-07,1.954615e-07,1.954616e-07,1.954618e-07,1.954620e-07,1.954622e-07,1.954623e-07,1.954625e-07,1.954627e-07,1.954629e-07,1.954630e-07,1.954632e-07,1.954634e-07,1.954635e-07,1.954637e-07,1.954639e-07,1.954641e-07,1.954642e-07,1.954644e-07,1.954646e-07,1.954647e-07,1.954649e-07,1.954651e-07,1.954653e-07,1.954654e-07,1.954656e-07,1.954658e-07,1.954659e-07,1.954661e-07,1.954663e-07,1.954665e-07,1.954666e-07,1.954668e-07,1.954670e-07,1.954672e-07,1.954673e-07,1.954675e-07,1.954677e-07,1.954678e-07,1.954680e-07,1.954682e-07,1.954684e-07,1.954685e-07,1.954687e-07,1.954689e-07,1.954690e-07,1.954692e-07,1.954694e-07,1.954696e-07,1.954697e-07,1.954699e-07,1.954701e-07,1.954702e-07,1.954704e-07,1.954706e-07,1.954708e-07,1.954709e-07,1.954711e-07,1.954713e-07,1.954715e-07,1.954716e-07,1.954718e-07,1.954720e-07,1.954721e-07,1.954723e-07,1.954725e-07,1.954727e-07,1.954728e-07,1.954730e-07,1.954732e-07,1.954733e-07,1.954735e-07,1.954737e-07,1.954739e-07,1.954740e-07,1.954742e-07,1.954744e-07,1.954745e-07,1.954747e-07,1.954749e-07,1.954751e-07,1.954752e-07,1.954754e-07,1.954756e-07,1.954758e-07,1.954759e-07,1.954761e-07,1.954763e-07,1.954764e-07,1.954766e-07,1.954768e-07,1.954770e-07,1.954771e-07,1.954773e-07,1.954775e-07,1.954776e-07,1.954778e-07,1.954780e-07,1.954782e-07,1.954783e-07,1.954785e-07,1.954787e-07,1.954788e-07,1.954790e-07,1.954792e-07,1.954794e-07,1.954795e-07,1.954797e-07,1.954799e-07,1.954800e-07,1.954802e-07,1.954804e-07,1.954806e-07,1.954807e-07,1.954809e-07,1.954811e-07,1.954813e-07,1.954814e-07,1.954816e-07,1.954818e-07,1.954819e-07,1.954821e-07,1.954823e-07,1.954825e-07,1.954826e-07,1.954828e-07,1.954830e-07,1.954831e-07,1.954833e-07,1.954835e-07,1.954837e-07,1.954838e-07,1.954840e-07,1.954842e-07,1.954843e-07,1.954845e-07,1.954847e-07,1.954849e-07,1.954850e-07,1.954852e-07,1.954854e-07,1.954855e-07,1.954857e-07,1.954859e-07,1.954861e-07,1.954862e-07,1.954864e-07,1.954866e-07,1.954867e-07,1.954869e-07,1.954871e-07,1.954873e-07,1.954874e-07,1.954876e-07,1.954878e-07,1.954879e-07,1.954881e-07,1.954883e-07,1.954885e-07,1.954886e-07,1.954888e-07,1.954890e-07,1.954892e-07,1.954893e-07,1.954895e-07,1.954897e-07,1.954898e-07,1.954900e-07,1.954902e-07,1.954904e-07,1.954905e-07,1.954907e-07,1.954909e-07,1.954910e-07,1.954912e-07,1.954914e-07,1.954916e-07,1.954917e-07,1.954919e-07,1.954921e-07,1.954922e-07,1.954924e-07,1.954926e-07,1.954928e-07,1.954929e-07,1.954931e-07,1.954933e-07,1.954934e-07,1.954936e-07,1.954938e-07,1.954940e-07,1.954941e-07,1.954943e-07,1.954945e-07,1.954946e-07,1.954948e-07,1.954950e-07,1.954952e-07,1.954953e-07,1.954955e-07,1.954957e-07,1.954958e-07,1.954960e-07,1.954962e-07,1.954964e-07,1.954965e-07,1.954967e-07,1.954969e-07,1.954970e-07,1.954972e-07,1.954974e-07,1.954976e-07,1.954977e-07,1.954979e-07,1.954981e-07,1.954982e-07,1.954984e-07,1.954986e-07,1.954988e-07,1.954989e-07,1.954991e-07,1.954993e-07,1.954994e-07,1.954996e-07,1.954998e-07,1.955000e-07,1.955001e-07,1.955003e-07,1.955005e-07,1.955007e-07,1.955008e-07,1.955010e-07,1.955012e-07,1.955013e-07,1.955015e-07,1.955017e-07,1.955019e-07,1.955020e-07,1.955022e-07,1.955024e-07,1.955025e-07,1.955027e-07,1.955029e-07,1.955031e-07,1.955032e-07,1.955034e-07,1.955036e-07,1.955037e-07,1.955039e-07,1.955041e-07,1.955043e-07,1.955044e-07,1.955046e-07,1.955048e-07,1.955049e-07,1.955051e-07,1.955053e-07,1.955055e-07,1.955056e-07,1.955058e-07,1.955060e-07,1.955061e-07,1.955063e-07,1.955065e-07,1.955067e-07,1.955068e-07,1.955070e-07,1.955072e-07,1.955073e-07,1.955075e-07,1.955077e-07,1.955079e-07,1.955080e-07,1.955082e-07,1.955084e-07,1.955085e-07,1.955087e-07,1.955089e-07,1.955091e-07,1.955092e-07,1.955094e-07,1.955096e-07,1.955097e-07,1.955099e-07,1.955101e-07,1.955103e-07,1.955104e-07,1.955106e-07,1.955108e-07,1.955109e-07,1.955111e-07,1.955113e-07,1.955115e-07,1.955116e-07,1.955118e-07,1.955120e-07,1.955121e-07,1.955123e-07,1.955125e-07,1.955127e-07,1.955128e-07,1.955130e-07,1.955132e-07,1.955133e-07,1.955135e-07,1.955137e-07,1.955139e-07,1.955140e-07,1.955142e-07,1.955144e-07,1.955145e-07,1.955147e-07,1.955149e-07,1.955151e-07,1.955152e-07,1.955154e-07,1.955156e-07,1.955157e-07,1.955159e-07,1.955161e-07,1.955162e-07,1.955164e-07,1.955166e-07,1.955168e-07,1.955169e-07,1.955171e-07,1.955173e-07,1.955174e-07,1.955176e-07,1.955178e-07,1.955180e-07,1.955181e-07,1.955183e-07,1.955185e-07,1.955186e-07,1.955188e-07,1.955190e-07,1.955192e-07,1.955193e-07,1.955195e-07,1.955197e-07,1.955198e-07,1.955200e-07,1.955202e-07,1.955204e-07,1.955205e-07,1.955207e-07,1.955209e-07,1.955210e-07,1.955212e-07,1.955214e-07,1.955216e-07,1.955217e-07,1.955219e-07,1.955221e-07,1.955222e-07,1.955224e-07,1.955226e-07,1.955228e-07,1.955229e-07,1.955231e-07,1.955233e-07,1.955234e-07,1.955236e-07,1.955238e-07,1.955240e-07,1.955241e-07,1.955243e-07,1.955245e-07,1.955246e-07,1.955248e-07,1.955250e-07,1.955252e-07,1.955253e-07,1.955255e-07,1.955257e-07,1.955258e-07,1.955260e-07,1.955262e-07,1.955264e-07,1.955265e-07,1.955267e-07,1.955269e-07,1.955270e-07,1.955272e-07,1.955274e-07,1.955276e-07,1.955277e-07,1.955279e-07,1.955281e-07,1.955282e-07,1.955284e-07,1.955286e-07,1.955287e-07,1.955289e-07,1.955291e-07,1.955293e-07,1.955294e-07,1.955296e-07,1.955298e-07,1.955299e-07,1.955301e-07,1.955303e-07,1.955305e-07,1.955306e-07,1.955308e-07,1.955310e-07,1.955311e-07,1.955313e-07,1.955315e-07,1.955317e-07,1.955318e-07,1.955320e-07,1.955322e-07,1.955323e-07,1.955325e-07,1.955327e-07,1.955329e-07,1.955330e-07,1.955332e-07,1.955334e-07,1.955335e-07,1.955337e-07,1.955339e-07,1.955341e-07,1.955342e-07,1.955344e-07,1.955346e-07,1.955347e-07,1.955349e-07,1.955351e-07,1.955352e-07,1.955354e-07,1.955356e-07,1.955358e-07,1.955359e-07,1.955361e-07,1.955363e-07,1.955364e-07,1.955366e-07,1.955368e-07,1.955370e-07,1.955371e-07,1.955373e-07,1.955375e-07,1.955376e-07,1.955378e-07,1.955380e-07,1.955382e-07,1.955383e-07,1.955385e-07,1.955387e-07,1.955388e-07,1.955390e-07,1.955392e-07,1.955394e-07,1.955395e-07,1.955397e-07,1.955399e-07,1.955400e-07,1.955402e-07,1.955404e-07,1.955406e-07,1.955407e-07,1.955409e-07,1.955411e-07,1.955412e-07,1.955414e-07,1.955416e-07,1.955417e-07,1.955419e-07,1.955421e-07,1.955423e-07,1.955424e-07,1.955426e-07,1.955428e-07,1.955429e-07,1.955431e-07,1.955433e-07,1.955435e-07,1.955436e-07,1.955438e-07,1.955440e-07,1.955441e-07,1.955443e-07,1.955445e-07,1.955447e-07,1.955448e-07,1.955450e-07,1.955452e-07,1.955453e-07,1.955455e-07,1.955457e-07,1.955458e-07,1.955460e-07,1.955462e-07,1.955464e-07,1.955465e-07,1.955467e-07,1.955469e-07,1.955470e-07,1.955472e-07,1.955474e-07,1.955476e-07,1.955477e-07,1.955479e-07,1.955481e-07,1.955482e-07,1.955484e-07,1.955486e-07,1.955488e-07,1.955489e-07,1.955491e-07,1.955493e-07,1.955494e-07,1.955496e-07,1.955498e-07,1.955499e-07,1.955501e-07,1.955503e-07,1.955505e-07,1.955506e-07,1.955508e-07,1.955510e-07,1.955511e-07,1.955513e-07,1.955515e-07,1.955517e-07,1.955518e-07,1.955520e-07,1.955522e-07,1.955523e-07,1.955525e-07,1.955527e-07,1.955529e-07,1.955530e-07,1.955532e-07,1.955534e-07,1.955535e-07,1.955537e-07,1.955539e-07,1.955540e-07,1.955542e-07,1.955544e-07,1.955546e-07,1.955547e-07,1.955549e-07,1.955551e-07,1.955552e-07,1.955554e-07,1.955556e-07,1.955558e-07,1.955559e-07,1.955561e-07,1.955563e-07,1.955564e-07,1.955566e-07,1.955568e-07,1.955569e-07,1.955571e-07,1.955573e-07,1.955575e-07,1.955576e-07,1.955578e-07,1.955580e-07,1.955581e-07,1.955583e-07,1.955585e-07,1.955587e-07,1.955588e-07,1.955590e-07,1.955592e-07,1.955593e-07,1.955595e-07,1.955597e-07,1.955599e-07,1.955600e-07,1.955602e-07,1.955604e-07,1.955605e-07,1.955607e-07,1.955609e-07,1.955610e-07,1.955612e-07,1.955614e-07,1.955616e-07,1.955617e-07,1.955619e-07,1.955621e-07,1.955622e-07,1.955624e-07,1.955626e-07,1.955628e-07,1.955629e-07,1.955631e-07,1.955633e-07,1.955634e-07,1.955636e-07,1.955638e-07,1.955639e-07,1.955641e-07,1.955643e-07,1.955645e-07,1.955646e-07,1.955648e-07,1.955650e-07,1.955651e-07,1.955653e-07,1.955655e-07,1.955657e-07,1.955658e-07,1.955660e-07,1.955662e-07,1.955663e-07,1.955665e-07,1.955667e-07,1.955668e-07,1.955670e-07,1.955672e-07,1.955674e-07,1.955675e-07,1.955677e-07,1.955679e-07,1.955680e-07,1.955682e-07,1.955684e-07,1.955686e-07,1.955687e-07,1.955689e-07,1.955691e-07,1.955692e-07,1.955694e-07,1.955696e-07,1.955697e-07,1.955699e-07,1.955701e-07,1.955703e-07,1.955704e-07,1.955706e-07,1.955708e-07,1.955709e-07,1.955711e-07,1.955713e-07,1.955715e-07,1.955716e-07,1.955718e-07,1.955720e-07,1.955721e-07,1.955723e-07,1.955725e-07,1.955726e-07,1.955728e-07,1.955730e-07,1.955732e-07,1.955733e-07,1.955735e-07,1.955737e-07,1.955738e-07,1.955740e-07,1.955742e-07,1.955743e-07,1.955745e-07,1.955747e-07,1.955749e-07,1.955750e-07,1.955752e-07,1.955754e-07,1.955755e-07,1.955757e-07,1.955759e-07,1.955761e-07,1.955762e-07,1.955764e-07,1.955766e-07,1.955767e-07,1.955769e-07,1.955771e-07,1.955772e-07,1.955774e-07,1.955776e-07,1.955778e-07,1.955779e-07,1.955781e-07,1.955783e-07,1.955784e-07,1.955786e-07,1.955788e-07,1.955790e-07,1.955791e-07,1.955793e-07,1.955795e-07,1.955796e-07,1.955798e-07,1.955800e-07,1.955801e-07,1.955803e-07,1.955805e-07,1.955807e-07,1.955808e-07,1.955810e-07,1.955812e-07,1.955813e-07,1.955815e-07,1.955817e-07,1.955818e-07,1.955820e-07,1.955822e-07,1.955824e-07,1.955825e-07,1.955827e-07,1.955829e-07,1.955830e-07,1.955832e-07,1.955834e-07,1.955836e-07,1.955837e-07,1.955839e-07,1.955841e-07,1.955842e-07,1.955844e-07,1.955846e-07,1.955847e-07,1.955849e-07,1.955851e-07,1.955853e-07,1.955854e-07,1.955856e-07,1.955858e-07,1.955859e-07,1.955861e-07,1.955863e-07,1.955864e-07,1.955866e-07,1.955868e-07,1.955870e-07,1.955871e-07,1.955873e-07,1.955875e-07,1.955876e-07,1.955878e-07,1.955880e-07,1.955881e-07,1.955883e-07,1.955885e-07,1.955887e-07,1.955888e-07,1.955890e-07,1.955892e-07,1.955893e-07,1.955895e-07,1.955897e-07,1.955899e-07,1.955900e-07,1.955902e-07,1.955904e-07,1.955905e-07,1.955907e-07,1.955909e-07,1.955910e-07,1.955912e-07,1.955914e-07,1.955916e-07,1.955917e-07,1.955919e-07,1.955921e-07,1.955922e-07,1.955924e-07,1.955926e-07,1.955927e-07,1.955929e-07,1.955931e-07,1.955933e-07,1.955934e-07,1.955936e-07,1.955938e-07,1.955939e-07,1.955941e-07,1.955943e-07,1.955944e-07,1.955946e-07,1.955948e-07,1.955950e-07,1.955951e-07,1.955953e-07,1.955955e-07,1.955956e-07,1.955958e-07,1.955960e-07,1.955961e-07,1.955963e-07,1.955965e-07,1.955967e-07,1.955968e-07,1.955970e-07,1.955972e-07,1.955973e-07,1.955975e-07,1.955977e-07,1.955978e-07,1.955980e-07,1.955982e-07,1.955984e-07,1.955985e-07,1.955987e-07,1.955989e-07,1.955990e-07,1.955992e-07,1.955994e-07,1.955996e-07,1.955997e-07,1.955999e-07,1.956001e-07,1.956002e-07,1.956004e-07,1.956006e-07,1.956007e-07,1.956009e-07,1.956011e-07,1.956013e-07,1.956014e-07,1.956016e-07,1.956018e-07,1.956019e-07,1.956021e-07,1.956023e-07,1.956024e-07,1.956026e-07,1.956028e-07,1.956030e-07,1.956031e-07,1.956033e-07,1.956035e-07,1.956036e-07,1.956038e-07,1.956040e-07,1.956041e-07,1.956043e-07,1.956045e-07,1.956047e-07,1.956048e-07,1.956050e-07,1.956052e-07,1.956053e-07,1.956055e-07,1.956057e-07,1.956058e-07,1.956060e-07,1.956062e-07,1.956064e-07,1.956065e-07,1.956067e-07,1.956069e-07,1.956070e-07,1.956072e-07,1.956074e-07,1.956075e-07,1.956077e-07,1.956079e-07,1.956081e-07,1.956082e-07,1.956084e-07,1.956086e-07,1.956087e-07,1.956089e-07,1.956091e-07,1.956092e-07,1.956094e-07,1.956096e-07,1.956098e-07,1.956099e-07,1.956101e-07,1.956103e-07,1.956104e-07,1.956106e-07,1.956108e-07,1.956109e-07,1.956111e-07,1.956113e-07,1.956115e-07,1.956116e-07,1.956118e-07,1.956120e-07,1.956121e-07,1.956123e-07,1.956125e-07,1.956126e-07,1.956128e-07,1.956130e-07,1.956132e-07,1.956133e-07,1.956135e-07,1.956137e-07,1.956138e-07,1.956140e-07,1.956142e-07,1.956143e-07,1.956145e-07,1.956147e-07,1.956148e-07,1.956150e-07,1.956152e-07,1.956154e-07,1.956155e-07,1.956157e-07,1.956159e-07,1.956160e-07,1.956162e-07,1.956164e-07,1.956165e-07,1.956167e-07,1.956169e-07,1.956171e-07,1.956172e-07,1.956174e-07,1.956176e-07,1.956177e-07,1.956179e-07,1.956181e-07,1.956182e-07,1.956184e-07,1.956186e-07,1.956188e-07,1.956189e-07,1.956191e-07,1.956193e-07,1.956194e-07,1.956196e-07,1.956198e-07,1.956199e-07,1.956201e-07,1.956203e-07,1.956205e-07,1.956206e-07,1.956208e-07,1.956210e-07,1.956211e-07,1.956213e-07,1.956215e-07,1.956216e-07,1.956218e-07,1.956220e-07,1.956222e-07,1.956223e-07,1.956225e-07,1.956227e-07,1.956228e-07,1.956230e-07,1.956232e-07,1.956233e-07,1.956235e-07,1.956237e-07,1.956238e-07,1.956240e-07,1.956242e-07,1.956244e-07,1.956245e-07,1.956247e-07,1.956249e-07,1.956250e-07,1.956252e-07,1.956254e-07,1.956255e-07,1.956257e-07,1.956259e-07,1.956261e-07,1.956262e-07,1.956264e-07,1.956266e-07,1.956267e-07,1.956269e-07,1.956271e-07,1.956272e-07,1.956274e-07,1.956276e-07,1.956278e-07,1.956279e-07,1.956281e-07,1.956283e-07,1.956284e-07,1.956286e-07,1.956288e-07,1.956289e-07,1.956291e-07,1.956293e-07,1.956294e-07,1.956296e-07,1.956298e-07,1.956300e-07,1.956301e-07,1.956303e-07,1.956305e-07,1.956306e-07,1.956308e-07,1.956310e-07,1.956311e-07,1.956313e-07,1.956315e-07,1.956317e-07,1.956318e-07,1.956320e-07,1.956322e-07,1.956323e-07,1.956325e-07,1.956327e-07,1.956328e-07,1.956330e-07,1.956332e-07,1.956334e-07,1.956335e-07,1.956337e-07,1.956339e-07,1.956340e-07,1.956342e-07,1.956344e-07,1.956345e-07,1.956347e-07,1.956349e-07,1.956350e-07,1.956352e-07,1.956354e-07,1.956356e-07,1.956357e-07,1.956359e-07,1.956361e-07,1.956362e-07,1.956364e-07,1.956366e-07,1.956367e-07,1.956369e-07,1.956371e-07,1.956373e-07,1.956374e-07,1.956376e-07,1.956378e-07,1.956379e-07,1.956381e-07,1.956383e-07,1.956384e-07,1.956386e-07,1.956388e-07,1.956389e-07,1.956391e-07,1.956393e-07,1.956395e-07,1.956396e-07,1.956398e-07,1.956400e-07,1.956401e-07,1.956403e-07,1.956405e-07,1.956406e-07,1.956408e-07,1.956410e-07,1.956411e-07,1.956413e-07,1.956415e-07,1.956417e-07,1.956418e-07,1.956420e-07,1.956422e-07,1.956423e-07,1.956425e-07,1.956427e-07,1.956428e-07,1.956430e-07,1.956432e-07,1.956434e-07,1.956435e-07,1.956437e-07,1.956439e-07,1.956440e-07,1.956442e-07,1.956444e-07,1.956445e-07,1.956447e-07,1.956449e-07,1.956450e-07,1.956452e-07,1.956454e-07,1.956456e-07,1.956457e-07,1.956459e-07,1.956461e-07,1.956462e-07,1.956464e-07,1.956466e-07,1.956467e-07,1.956469e-07,1.956471e-07,1.956472e-07,1.956474e-07,1.956476e-07,1.956478e-07,1.956479e-07,1.956481e-07,1.956483e-07,1.956484e-07,1.956486e-07,1.956488e-07,1.956489e-07,1.956491e-07,1.956493e-07,1.956495e-07,1.956496e-07,1.956498e-07,1.956500e-07,1.956501e-07,1.956503e-07,1.956505e-07,1.956506e-07,1.956508e-07,1.956510e-07,1.956511e-07,1.956513e-07,1.956515e-07,1.956517e-07,1.956518e-07,1.956520e-07,1.956522e-07,1.956523e-07,1.956525e-07,1.956527e-07,1.956528e-07,1.956530e-07,1.956532e-07,1.956533e-07,1.956535e-07,1.956537e-07,1.956539e-07,1.956540e-07,1.956542e-07,1.956544e-07,1.956545e-07,1.956547e-07,1.956549e-07,1.956550e-07,1.956552e-07,1.956554e-07,1.956555e-07,1.956557e-07,1.956559e-07,1.956561e-07,1.956562e-07,1.956564e-07,1.956566e-07,1.956567e-07,1.956569e-07,1.956571e-07,1.956572e-07,1.956574e-07,1.956576e-07,1.956577e-07,1.956579e-07,1.956581e-07,1.956583e-07,1.956584e-07,1.956586e-07,1.956588e-07,1.956589e-07,1.956591e-07,1.956593e-07,1.956594e-07,1.956596e-07,1.956598e-07,1.956599e-07,1.956601e-07,1.956603e-07,1.956605e-07,1.956606e-07,1.956608e-07,1.956610e-07,1.956611e-07,1.956613e-07,1.956615e-07,1.956616e-07,1.956618e-07,1.956620e-07,1.956621e-07,1.956623e-07,1.956625e-07,1.956627e-07,1.956628e-07,1.956630e-07,1.956632e-07,1.956633e-07,1.956635e-07,1.956637e-07,1.956638e-07,1.956640e-07,1.956642e-07,1.956643e-07,1.956645e-07,1.956647e-07,1.956649e-07,1.956650e-07,1.956652e-07,1.956654e-07,1.956655e-07,1.956657e-07,1.956659e-07,1.956660e-07,1.956662e-07,1.956664e-07,1.956665e-07,1.956667e-07,1.956669e-07,1.956671e-07,1.956672e-07,1.956674e-07,1.956676e-07,1.956677e-07,1.956679e-07,1.956681e-07,1.956682e-07,1.956684e-07,1.956686e-07,1.956687e-07,1.956689e-07,1.956691e-07,1.956693e-07,1.956694e-07,1.956696e-07,1.956698e-07,1.956699e-07,1.956701e-07,1.956703e-07,1.956704e-07,1.956706e-07,1.956708e-07,1.956709e-07,1.956711e-07,1.956713e-07,1.956714e-07,1.956716e-07,1.956718e-07,1.956720e-07,1.956721e-07,1.956723e-07,1.956725e-07,1.956726e-07,1.956728e-07,1.956730e-07,1.956731e-07,1.956733e-07,1.956735e-07,1.956736e-07,1.956738e-07,1.956740e-07,1.956742e-07,1.956743e-07,1.956745e-07,1.956747e-07,1.956748e-07,1.956750e-07,1.956752e-07,1.956753e-07,1.956755e-07,1.956757e-07,1.956758e-07,1.956760e-07,1.956762e-07,1.956764e-07,1.956765e-07,1.956767e-07,1.956769e-07,1.956770e-07,1.956772e-07,1.956774e-07,1.956775e-07,1.956777e-07,1.956779e-07,1.956780e-07,1.956782e-07,1.956784e-07,1.956785e-07,1.956787e-07,1.956789e-07,1.956791e-07,1.956792e-07,1.956794e-07,1.956796e-07,1.956797e-07,1.956799e-07,1.956801e-07,1.956802e-07,1.956804e-07,1.956806e-07,1.956807e-07,1.956809e-07,1.956811e-07,1.956812e-07,1.956814e-07,1.956816e-07,1.956818e-07,1.956819e-07,1.956821e-07,1.956823e-07,1.956824e-07,1.956826e-07,1.956828e-07,1.956829e-07,1.956831e-07,1.956833e-07,1.956834e-07,1.956836e-07,1.956838e-07,1.956840e-07,1.956841e-07,1.956843e-07,1.956845e-07,1.956846e-07,1.956848e-07,1.956850e-07,1.956851e-07,1.956853e-07,1.956855e-07,1.956856e-07,1.956858e-07,1.956860e-07,1.956861e-07,1.956863e-07,1.956865e-07,1.956867e-07,1.956868e-07,1.956870e-07,1.956872e-07,1.956873e-07,1.956875e-07,1.956877e-07,1.956878e-07,1.956880e-07,1.956882e-07,1.956883e-07,1.956885e-07,1.956887e-07,1.956888e-07,1.956890e-07,1.956892e-07,1.956894e-07,1.956895e-07,1.956897e-07,1.956899e-07,1.956900e-07,1.956902e-07,1.956904e-07,1.956905e-07,1.956907e-07,1.956909e-07,1.956910e-07,1.956912e-07,1.956914e-07,1.956915e-07,1.956917e-07,1.956919e-07,1.956921e-07,1.956922e-07,1.956924e-07,1.956926e-07,1.956927e-07,1.956929e-07,1.956931e-07,1.956932e-07,1.956934e-07,1.956936e-07,1.956937e-07,1.956939e-07,1.956941e-07,1.956942e-07,1.956944e-07,1.956946e-07,1.956948e-07,1.956949e-07,1.956951e-07,1.956953e-07,1.956954e-07,1.956956e-07,1.956958e-07,1.956959e-07,1.956961e-07,1.956963e-07,1.956964e-07,1.956966e-07,1.956968e-07,1.956969e-07,1.956971e-07,1.956973e-07,1.956975e-07,1.956976e-07,1.956978e-07,1.956980e-07,1.956981e-07,1.956983e-07,1.956985e-07,1.956986e-07,1.956988e-07,1.956990e-07,1.956991e-07,1.956993e-07,1.956995e-07,1.956996e-07,1.956998e-07,1.957000e-07,1.957002e-07,1.957003e-07,1.957005e-07,1.957007e-07,1.957008e-07,1.957010e-07,1.957012e-07,1.957013e-07,1.957015e-07,1.957017e-07,1.957018e-07,1.957020e-07,1.957022e-07,1.957023e-07,1.957025e-07,1.957027e-07,1.957029e-07,1.957030e-07,1.957032e-07,1.957034e-07,1.957035e-07,1.957037e-07,1.957039e-07,1.957040e-07,1.957042e-07,1.957044e-07,1.957045e-07,1.957047e-07,1.957049e-07,1.957050e-07,1.957052e-07,1.957054e-07,1.957055e-07,1.957057e-07,1.957059e-07,1.957061e-07,1.957062e-07,1.957064e-07,1.957066e-07,1.957067e-07,1.957069e-07,1.957071e-07,1.957072e-07,1.957074e-07,1.957076e-07,1.957077e-07,1.957079e-07,1.957081e-07,1.957082e-07,1.957084e-07,1.957086e-07,1.957087e-07,1.957089e-07,1.957091e-07,1.957093e-07,1.957094e-07,1.957096e-07,1.957098e-07,1.957099e-07,1.957101e-07,1.957103e-07,1.957104e-07,1.957106e-07,1.957108e-07,1.957109e-07,1.957111e-07,1.957113e-07,1.957114e-07,1.957116e-07,1.957118e-07,1.957120e-07,1.957121e-07,1.957123e-07,1.957125e-07,1.957126e-07,1.957128e-07,1.957130e-07,1.957131e-07,1.957133e-07,1.957135e-07,1.957136e-07,1.957138e-07,1.957140e-07,1.957141e-07,1.957143e-07,1.957145e-07,1.957146e-07,1.957148e-07,1.957150e-07,1.957152e-07,1.957153e-07,1.957155e-07,1.957157e-07,1.957158e-07,1.957160e-07,1.957162e-07,1.957163e-07,1.957165e-07,1.957167e-07,1.957168e-07,1.957170e-07,1.957172e-07,1.957173e-07,1.957175e-07,1.957177e-07,1.957178e-07,1.957180e-07,1.957182e-07,1.957184e-07,1.957185e-07,1.957187e-07,1.957189e-07,1.957190e-07,1.957192e-07,1.957194e-07,1.957195e-07,1.957197e-07,1.957199e-07,1.957200e-07,1.957202e-07,1.957204e-07,1.957205e-07,1.957207e-07,1.957209e-07,1.957210e-07,1.957212e-07,1.957214e-07,1.957215e-07,1.957217e-07,1.957219e-07,1.957221e-07,1.957222e-07,1.957224e-07,1.957226e-07,1.957227e-07,1.957229e-07,1.957231e-07,1.957232e-07,1.957234e-07,1.957236e-07,1.957237e-07,1.957239e-07,1.957241e-07,1.957242e-07,1.957244e-07,1.957246e-07,1.957247e-07,1.957249e-07,1.957251e-07,1.957253e-07,1.957254e-07,1.957256e-07,1.957258e-07,1.957259e-07,1.957261e-07,1.957263e-07,1.957264e-07,1.957266e-07,1.957268e-07,1.957269e-07,1.957271e-07,1.957273e-07,1.957274e-07,1.957276e-07,1.957278e-07,1.957279e-07,1.957281e-07,1.957283e-07,1.957284e-07,1.957286e-07,1.957288e-07,1.957290e-07,1.957291e-07,1.957293e-07,1.957295e-07,1.957296e-07,1.957298e-07,1.957300e-07,1.957301e-07,1.957303e-07,1.957305e-07,1.957306e-07,1.957308e-07,1.957310e-07,1.957311e-07,1.957313e-07,1.957315e-07,1.957316e-07,1.957318e-07,1.957320e-07,1.957321e-07,1.957323e-07,1.957325e-07,1.957327e-07,1.957328e-07,1.957330e-07,1.957332e-07,1.957333e-07,1.957335e-07,1.957337e-07,1.957338e-07,1.957340e-07,1.957342e-07,1.957343e-07,1.957345e-07,1.957347e-07,1.957348e-07,1.957350e-07,1.957352e-07,1.957353e-07,1.957355e-07,1.957357e-07,1.957358e-07,1.957360e-07,1.957362e-07,1.957364e-07,1.957365e-07,1.957367e-07,1.957369e-07,1.957370e-07,1.957372e-07,1.957374e-07,1.957375e-07,1.957377e-07,1.957379e-07,1.957380e-07,1.957382e-07,1.957384e-07,1.957385e-07,1.957387e-07,1.957389e-07,1.957390e-07,1.957392e-07,1.957394e-07,1.957395e-07,1.957397e-07,1.957399e-07,1.957401e-07,1.957402e-07,1.957404e-07,1.957406e-07,1.957407e-07,1.957409e-07,1.957411e-07,1.957412e-07,1.957414e-07,1.957416e-07,1.957417e-07,1.957419e-07,1.957421e-07,1.957422e-07,1.957424e-07,1.957426e-07,1.957427e-07,1.957429e-07,1.957431e-07,1.957432e-07,1.957434e-07,1.957436e-07,1.957437e-07,1.957439e-07,1.957441e-07,1.957443e-07,1.957444e-07,1.957446e-07,1.957448e-07,1.957449e-07,1.957451e-07,1.957453e-07,1.957454e-07,1.957456e-07,1.957458e-07,1.957459e-07,1.957461e-07,1.957463e-07,1.957464e-07,1.957466e-07,1.957468e-07,1.957469e-07,1.957471e-07,1.957473e-07,1.957474e-07,1.957476e-07,1.957478e-07,1.957479e-07,1.957481e-07,1.957483e-07,1.957485e-07,1.957486e-07,1.957488e-07,1.957490e-07,1.957491e-07,1.957493e-07,1.957495e-07,1.957496e-07,1.957498e-07,1.957500e-07,1.957501e-07,1.957503e-07,1.957505e-07,1.957506e-07,1.957508e-07,1.957510e-07,1.957511e-07,1.957513e-07,1.957515e-07,1.957516e-07,1.957518e-07,1.957520e-07,1.957521e-07,1.957523e-07,1.957525e-07,1.957526e-07,1.957528e-07,1.957530e-07,1.957532e-07,1.957533e-07,1.957535e-07,1.957537e-07,1.957538e-07,1.957540e-07,1.957542e-07,1.957543e-07,1.957545e-07,1.957547e-07,1.957548e-07,1.957550e-07,1.957552e-07,1.957553e-07,1.957555e-07,1.957557e-07,1.957558e-07,1.957560e-07,1.957562e-07,1.957563e-07,1.957565e-07,1.957567e-07,1.957568e-07,1.957570e-07,1.957572e-07,1.957573e-07,1.957575e-07,1.957577e-07,1.957579e-07,1.957580e-07,1.957582e-07,1.957584e-07,1.957585e-07,1.957587e-07,1.957589e-07,1.957590e-07,1.957592e-07,1.957594e-07,1.957595e-07,1.957597e-07,1.957599e-07,1.957600e-07,1.957602e-07,1.957604e-07,1.957605e-07,1.957607e-07,1.957609e-07,1.957610e-07,1.957612e-07,1.957614e-07,1.957615e-07,1.957617e-07,1.957619e-07,1.957620e-07,1.957622e-07,1.957624e-07,1.957626e-07,1.957627e-07,1.957629e-07,1.957631e-07,1.957632e-07,1.957634e-07,1.957636e-07,1.957637e-07,1.957639e-07,1.957641e-07,1.957642e-07,1.957644e-07,1.957646e-07,1.957647e-07,1.957649e-07,1.957651e-07,1.957652e-07,1.957654e-07,1.957656e-07,1.957657e-07,1.957659e-07,1.957661e-07,1.957662e-07,1.957664e-07,1.957666e-07,1.957667e-07,1.957669e-07,1.957671e-07,1.957672e-07,1.957674e-07,1.957676e-07,1.957677e-07,1.957679e-07,1.957681e-07,1.957683e-07,1.957684e-07,1.957686e-07,1.957688e-07,1.957689e-07,1.957691e-07,1.957693e-07,1.957694e-07,1.957696e-07,1.957698e-07,1.957699e-07,1.957701e-07,1.957703e-07,1.957704e-07,1.957706e-07,1.957708e-07,1.957709e-07,1.957711e-07,1.957713e-07,1.957714e-07,1.957716e-07,1.957718e-07,1.957719e-07,1.957721e-07,1.957723e-07,1.957724e-07,1.957726e-07,1.957728e-07,1.957729e-07,1.957731e-07,1.957733e-07,1.957734e-07,1.957736e-07,1.957738e-07,1.957740e-07,1.957741e-07,1.957743e-07,1.957745e-07,1.957746e-07,1.957748e-07,1.957750e-07,1.957751e-07,1.957753e-07,1.957755e-07,1.957756e-07,1.957758e-07,1.957760e-07,1.957761e-07,1.957763e-07,1.957765e-07,1.957766e-07,1.957768e-07,1.957770e-07,1.957771e-07,1.957773e-07,1.957775e-07,1.957776e-07,1.957778e-07,1.957780e-07,1.957781e-07,1.957783e-07,1.957785e-07,1.957786e-07,1.957788e-07,1.957790e-07,1.957791e-07,1.957793e-07,1.957795e-07,1.957796e-07,1.957798e-07,1.957800e-07,1.957802e-07,1.957803e-07,1.957805e-07,1.957807e-07,1.957808e-07,1.957810e-07,1.957812e-07,1.957813e-07,1.957815e-07,1.957817e-07,1.957818e-07,1.957820e-07,1.957822e-07,1.957823e-07,1.957825e-07,1.957827e-07,1.957828e-07,1.957830e-07,1.957832e-07,1.957833e-07,1.957835e-07,1.957837e-07,1.957838e-07,1.957840e-07,1.957842e-07,1.957843e-07,1.957845e-07,1.957847e-07,1.957848e-07,1.957850e-07,1.957852e-07,1.957853e-07,1.957855e-07,1.957857e-07,1.957858e-07,1.957860e-07,1.957862e-07,1.957863e-07,1.957865e-07,1.957867e-07,1.957868e-07,1.957870e-07,1.957872e-07,1.957874e-07,1.957875e-07,1.957877e-07,1.957879e-07,1.957880e-07,1.957882e-07,1.957884e-07,1.957885e-07,1.957887e-07,1.957889e-07,1.957890e-07,1.957892e-07,1.957894e-07,1.957895e-07,1.957897e-07,1.957899e-07,1.957900e-07,1.957902e-07,1.957904e-07,1.957905e-07,1.957907e-07,1.957909e-07,1.957910e-07,1.957912e-07,1.957914e-07,1.957915e-07,1.957917e-07,1.957919e-07,1.957920e-07,1.957922e-07,1.957924e-07,1.957925e-07,1.957927e-07,1.957929e-07,1.957930e-07,1.957932e-07,1.957934e-07,1.957935e-07,1.957937e-07,1.957939e-07,1.957940e-07,1.957942e-07,1.957944e-07,1.957945e-07,1.957947e-07,1.957949e-07,1.957950e-07,1.957952e-07,1.957954e-07,1.957955e-07,1.957957e-07,1.957959e-07,1.957961e-07,1.957962e-07,1.957964e-07,1.957966e-07,1.957967e-07,1.957969e-07,1.957971e-07,1.957972e-07,1.957974e-07,1.957976e-07,1.957977e-07,1.957979e-07,1.957981e-07,1.957982e-07,1.957984e-07,1.957986e-07,1.957987e-07,1.957989e-07,1.957991e-07,1.957992e-07,1.957994e-07,1.957996e-07,1.957997e-07,1.957999e-07,1.958001e-07,1.958002e-07,1.958004e-07,1.958006e-07,1.958007e-07,1.958009e-07,1.958011e-07,1.958012e-07,1.958014e-07,1.958016e-07,1.958017e-07,1.958019e-07,1.958021e-07,1.958022e-07,1.958024e-07,1.958026e-07,1.958027e-07,1.958029e-07,1.958031e-07,1.958032e-07,1.958034e-07,1.958036e-07,1.958037e-07,1.958039e-07,1.958041e-07,1.958042e-07,1.958044e-07,1.958046e-07,1.958047e-07,1.958049e-07,1.958051e-07,1.958052e-07,1.958054e-07,1.958056e-07,1.958057e-07,1.958059e-07,1.958061e-07,1.958062e-07,1.958064e-07,1.958066e-07,1.958068e-07,1.958069e-07,1.958071e-07,1.958073e-07,1.958074e-07,1.958076e-07,1.958078e-07,1.958079e-07,1.958081e-07,1.958083e-07,1.958084e-07,1.958086e-07,1.958088e-07,1.958089e-07,1.958091e-07,1.958093e-07,1.958094e-07,1.958096e-07,1.958098e-07,1.958099e-07,1.958101e-07,1.958103e-07,1.958104e-07,1.958106e-07,1.958108e-07,1.958109e-07,1.958111e-07,1.958113e-07,1.958114e-07,1.958116e-07,1.958118e-07,1.958119e-07,1.958121e-07,1.958123e-07,1.958124e-07,1.958126e-07,1.958128e-07,1.958129e-07,1.958131e-07,1.958133e-07,1.958134e-07,1.958136e-07,1.958138e-07,1.958139e-07,1.958141e-07,1.958143e-07,1.958144e-07,1.958146e-07,1.958148e-07,1.958149e-07,1.958151e-07,1.958153e-07,1.958154e-07,1.958156e-07,1.958158e-07,1.958159e-07,1.958161e-07,1.958163e-07,1.958164e-07,1.958166e-07,1.958168e-07,1.958169e-07,1.958171e-07,1.958173e-07,1.958174e-07,1.958176e-07,1.958178e-07,1.958179e-07,1.958181e-07,1.958183e-07,1.958184e-07,1.958186e-07,1.958188e-07,1.958189e-07,1.958191e-07,1.958193e-07,1.958194e-07,1.958196e-07,1.958198e-07,1.958199e-07,1.958201e-07,1.958203e-07,1.958204e-07,1.958206e-07,1.958208e-07,1.958209e-07,1.958211e-07,1.958213e-07,1.958214e-07,1.958216e-07,1.958218e-07,1.958219e-07,1.958221e-07,1.958223e-07,1.958224e-07,1.958226e-07,1.958228e-07,1.958229e-07,1.958231e-07,1.958233e-07,1.958234e-07,1.958236e-07,1.958238e-07,1.958240e-07,1.958241e-07,1.958243e-07,1.958245e-07,1.958246e-07,1.958248e-07,1.958250e-07,1.958251e-07,1.958253e-07,1.958255e-07,1.958256e-07,1.958258e-07,1.958260e-07,1.958261e-07,1.958263e-07,1.958265e-07,1.958266e-07,1.958268e-07,1.958270e-07,1.958271e-07,1.958273e-07,1.958275e-07,1.958276e-07,1.958278e-07,1.958280e-07,1.958281e-07,1.958283e-07,1.958285e-07,1.958286e-07,1.958288e-07,1.958290e-07,1.958291e-07,1.958293e-07,1.958295e-07,1.958296e-07,1.958298e-07,1.958300e-07,1.958301e-07,1.958303e-07,1.958305e-07,1.958306e-07,1.958308e-07,1.958310e-07,1.958311e-07,1.958313e-07,1.958315e-07,1.958316e-07,1.958318e-07,1.958320e-07,1.958321e-07,1.958323e-07,1.958325e-07,1.958326e-07,1.958328e-07,1.958330e-07,1.958331e-07,1.958333e-07,1.958335e-07,1.958336e-07,1.958338e-07,1.958340e-07,1.958341e-07,1.958343e-07,1.958345e-07,1.958346e-07,1.958348e-07,1.958350e-07,1.958351e-07,1.958353e-07,1.958355e-07,1.958356e-07,1.958358e-07,1.958360e-07,1.958361e-07,1.958363e-07,1.958365e-07,1.958366e-07,1.958368e-07,1.958370e-07,1.958371e-07,1.958373e-07,1.958375e-07,1.958376e-07,1.958378e-07,1.958380e-07,1.958381e-07,1.958383e-07,1.958385e-07,1.958386e-07,1.958388e-07,1.958390e-07,1.958391e-07,1.958393e-07,1.958395e-07,1.958396e-07,1.958398e-07,1.958400e-07,1.958401e-07,1.958403e-07,1.958405e-07,1.958406e-07,1.958408e-07,1.958410e-07,1.958411e-07,1.958413e-07,1.958415e-07,1.958416e-07,1.958418e-07,1.958420e-07,1.958421e-07,1.958423e-07,1.958425e-07,1.958426e-07,1.958428e-07,1.958430e-07,1.958431e-07,1.958433e-07,1.958435e-07,1.958436e-07,1.958438e-07,1.958440e-07,1.958441e-07,1.958443e-07,1.958445e-07,1.958446e-07,1.958448e-07,1.958450e-07,1.958451e-07,1.958453e-07,1.958455e-07,1.958456e-07,1.958458e-07,1.958460e-07,1.958461e-07,1.958463e-07,1.958465e-07,1.958466e-07,1.958468e-07,1.958470e-07,1.958471e-07,1.958473e-07,1.958475e-07,1.958476e-07,1.958478e-07,1.958480e-07,1.958481e-07,1.958483e-07,1.958485e-07,1.958486e-07,1.958488e-07,1.958490e-07,1.958491e-07,1.958493e-07,1.958495e-07,1.958496e-07,1.958498e-07,1.958500e-07,1.958501e-07,1.958503e-07,1.958505e-07,1.958506e-07,1.958508e-07,1.958510e-07,1.958511e-07,1.958513e-07,1.958515e-07,1.958516e-07,1.958518e-07,1.958520e-07,1.958521e-07,1.958523e-07,1.958524e-07,1.958526e-07,1.958528e-07,1.958529e-07,1.958531e-07,1.958533e-07,1.958534e-07,1.958536e-07,1.958538e-07,1.958539e-07,1.958541e-07,1.958543e-07,1.958544e-07,1.958546e-07,1.958548e-07,1.958549e-07,1.958551e-07,1.958553e-07,1.958554e-07,1.958556e-07,1.958558e-07,1.958559e-07,1.958561e-07,1.958563e-07,1.958564e-07,1.958566e-07,1.958568e-07,1.958569e-07,1.958571e-07,1.958573e-07,1.958574e-07,1.958576e-07,1.958578e-07,1.958579e-07,1.958581e-07,1.958583e-07,1.958584e-07,1.958586e-07,1.958588e-07,1.958589e-07,1.958591e-07,1.958593e-07,1.958594e-07,1.958596e-07,1.958598e-07,1.958599e-07,1.958601e-07,1.958603e-07,1.958604e-07,1.958606e-07,1.958608e-07,1.958609e-07,1.958611e-07,1.958613e-07,1.958614e-07,1.958616e-07,1.958618e-07,1.958619e-07,1.958621e-07,1.958623e-07,1.958624e-07,1.958626e-07,1.958628e-07,1.958629e-07,1.958631e-07,1.958633e-07,1.958634e-07,1.958636e-07,1.958638e-07,1.958639e-07,1.958641e-07,1.958643e-07,1.958644e-07,1.958646e-07,1.958648e-07,1.958649e-07,1.958651e-07,1.958653e-07,1.958654e-07,1.958656e-07,1.958658e-07,1.958659e-07,1.958661e-07,1.958663e-07,1.958664e-07,1.958666e-07,1.958668e-07,1.958669e-07,1.958671e-07,1.958673e-07,1.958674e-07,1.958676e-07,1.958678e-07,1.958679e-07,1.958681e-07,1.958683e-07,1.958684e-07,1.958686e-07,1.958688e-07,1.958689e-07,1.958691e-07,1.958692e-07,1.958694e-07,1.958696e-07,1.958697e-07,1.958699e-07,1.958701e-07,1.958702e-07,1.958704e-07,1.958706e-07,1.958707e-07,1.958709e-07,1.958711e-07,1.958712e-07,1.958714e-07,1.958716e-07,1.958717e-07,1.958719e-07,1.958721e-07,1.958722e-07,1.958724e-07,1.958726e-07,1.958727e-07,1.958729e-07,1.958731e-07,1.958732e-07,1.958734e-07,1.958736e-07,1.958737e-07,1.958739e-07,1.958741e-07,1.958742e-07,1.958744e-07,1.958746e-07,1.958747e-07,1.958749e-07,1.958751e-07,1.958752e-07,1.958754e-07,1.958756e-07,1.958757e-07,1.958759e-07,1.958761e-07,1.958762e-07,1.958764e-07,1.958766e-07,1.958767e-07,1.958769e-07,1.958771e-07,1.958772e-07,1.958774e-07,1.958776e-07,1.958777e-07,1.958779e-07,1.958781e-07,1.958782e-07,1.958784e-07,1.958786e-07,1.958787e-07,1.958789e-07,1.958791e-07,1.958792e-07,1.958794e-07,1.958796e-07,1.958797e-07,1.958799e-07,1.958800e-07,1.958802e-07,1.958804e-07,1.958805e-07,1.958807e-07,1.958809e-07,1.958810e-07,1.958812e-07,1.958814e-07,1.958815e-07,1.958817e-07,1.958819e-07,1.958820e-07,1.958822e-07,1.958824e-07,1.958825e-07,1.958827e-07,1.958829e-07,1.958830e-07,1.958832e-07,1.958834e-07,1.958835e-07,1.958837e-07,1.958839e-07,1.958840e-07,1.958842e-07,1.958844e-07,1.958845e-07,1.958847e-07,1.958849e-07,1.958850e-07,1.958852e-07,1.958854e-07,1.958855e-07,1.958857e-07,1.958859e-07,1.958860e-07,1.958862e-07,1.958864e-07,1.958865e-07,1.958867e-07,1.958869e-07,1.958870e-07,1.958872e-07,1.958874e-07,1.958875e-07,1.958877e-07,1.958879e-07,1.958880e-07,1.958882e-07,1.958883e-07,1.958885e-07,1.958887e-07,1.958888e-07,1.958890e-07,1.958892e-07,1.958893e-07,1.958895e-07,1.958897e-07,1.958898e-07,1.958900e-07,1.958902e-07,1.958903e-07,1.958905e-07,1.958907e-07,1.958908e-07,1.958910e-07,1.958912e-07,1.958913e-07,1.958915e-07,1.958917e-07,1.958918e-07,1.958920e-07,1.958922e-07,1.958923e-07,1.958925e-07,1.958927e-07,1.958928e-07,1.958930e-07,1.958932e-07,1.958933e-07,1.958935e-07,1.958937e-07,1.958938e-07,1.958940e-07,1.958942e-07,1.958943e-07,1.958945e-07,1.958947e-07,1.958948e-07,1.958950e-07,1.958952e-07,1.958953e-07,1.958955e-07,1.958956e-07,1.958958e-07,1.958960e-07,1.958961e-07,1.958963e-07,1.958965e-07,1.958966e-07,1.958968e-07,1.958970e-07,1.958971e-07,1.958973e-07,1.958975e-07,1.958976e-07,1.958978e-07,1.958980e-07,1.958981e-07,1.958983e-07,1.958985e-07,1.958986e-07,1.958988e-07,1.958990e-07,1.958991e-07,1.958993e-07,1.958995e-07,1.958996e-07,1.958998e-07,1.959000e-07,1.959001e-07,1.959003e-07,1.959005e-07,1.959006e-07,1.959008e-07,1.959010e-07,1.959011e-07,1.959013e-07,1.959015e-07,1.959016e-07,1.959018e-07,1.959019e-07,1.959021e-07,1.959023e-07,1.959024e-07,1.959026e-07,1.959028e-07,1.959029e-07,1.959031e-07,1.959033e-07,1.959034e-07,1.959036e-07,1.959038e-07,1.959039e-07,1.959041e-07,1.959043e-07,1.959044e-07,1.959046e-07,1.959048e-07,1.959049e-07,1.959051e-07,1.959053e-07,1.959054e-07,1.959056e-07,1.959058e-07,1.959059e-07,1.959061e-07,1.959063e-07,1.959064e-07,1.959066e-07,1.959068e-07,1.959069e-07,1.959071e-07,1.959073e-07,1.959074e-07,1.959076e-07,1.959077e-07,1.959079e-07,1.959081e-07,1.959082e-07,1.959084e-07,1.959086e-07,1.959087e-07,1.959089e-07,1.959091e-07,1.959092e-07,1.959094e-07,1.959096e-07,1.959097e-07,1.959099e-07,1.959101e-07,1.959102e-07,1.959104e-07,1.959106e-07,1.959107e-07,1.959109e-07,1.959111e-07,1.959112e-07,1.959114e-07,1.959116e-07,1.959117e-07,1.959119e-07,1.959121e-07,1.959122e-07,1.959124e-07,1.959126e-07,1.959127e-07,1.959129e-07,1.959131e-07,1.959132e-07,1.959134e-07,1.959135e-07,1.959137e-07,1.959139e-07,1.959140e-07,1.959142e-07,1.959144e-07,1.959145e-07,1.959147e-07,1.959149e-07,1.959150e-07,1.959152e-07,1.959154e-07,1.959155e-07,1.959157e-07,1.959159e-07,1.959160e-07,1.959162e-07,1.959164e-07,1.959165e-07,1.959167e-07,1.959169e-07,1.959170e-07,1.959172e-07,1.959174e-07,1.959175e-07,1.959177e-07,1.959179e-07,1.959180e-07,1.959182e-07,1.959183e-07,1.959185e-07,1.959187e-07,1.959188e-07,1.959190e-07,1.959192e-07,1.959193e-07,1.959195e-07,1.959197e-07,1.959198e-07,1.959200e-07,1.959202e-07,1.959203e-07,1.959205e-07,1.959207e-07,1.959208e-07,1.959210e-07,1.959212e-07,1.959213e-07,1.959215e-07,1.959217e-07,1.959218e-07,1.959220e-07,1.959222e-07,1.959223e-07,1.959225e-07,1.959227e-07,1.959228e-07,1.959230e-07,1.959231e-07,1.959233e-07,1.959235e-07,1.959236e-07,1.959238e-07,1.959240e-07,1.959241e-07,1.959243e-07,1.959245e-07,1.959246e-07,1.959248e-07,1.959250e-07,1.959251e-07,1.959253e-07,1.959255e-07,1.959256e-07,1.959258e-07,1.959260e-07,1.959261e-07,1.959263e-07,1.959265e-07,1.959266e-07,1.959268e-07,1.959270e-07,1.959271e-07,1.959273e-07,1.959274e-07,1.959276e-07,1.959278e-07,1.959279e-07,1.959281e-07,1.959283e-07,1.959284e-07,1.959286e-07,1.959288e-07,1.959289e-07,1.959291e-07,1.959293e-07,1.959294e-07,1.959296e-07,1.959298e-07,1.959299e-07,1.959301e-07,1.959303e-07,1.959304e-07,1.959306e-07,1.959308e-07,1.959309e-07,1.959311e-07,1.959313e-07,1.959314e-07,1.959316e-07,1.959317e-07,1.959319e-07,1.959321e-07,1.959322e-07,1.959324e-07,1.959326e-07,1.959327e-07,1.959329e-07,1.959331e-07,1.959332e-07,1.959334e-07,1.959336e-07,1.959337e-07,1.959339e-07,1.959341e-07,1.959342e-07,1.959344e-07,1.959346e-07,1.959347e-07,1.959349e-07,1.959351e-07,1.959352e-07,1.959354e-07,1.959356e-07,1.959357e-07,1.959359e-07,1.959360e-07,1.959362e-07,1.959364e-07,1.959365e-07,1.959367e-07,1.959369e-07,1.959370e-07,1.959372e-07,1.959374e-07,1.959375e-07,1.959377e-07,1.959379e-07,1.959380e-07,1.959382e-07,1.959384e-07,1.959385e-07,1.959387e-07,1.959389e-07,1.959390e-07,1.959392e-07,1.959394e-07,1.959395e-07,1.959397e-07,1.959398e-07,1.959400e-07,1.959402e-07,1.959403e-07,1.959405e-07,1.959407e-07,1.959408e-07,1.959410e-07,1.959412e-07,1.959413e-07,1.959415e-07,1.959417e-07,1.959418e-07,1.959420e-07,1.959422e-07,1.959423e-07,1.959425e-07,1.959427e-07,1.959428e-07,1.959430e-07,1.959432e-07,1.959433e-07,1.959435e-07,1.959436e-07,1.959438e-07,1.959440e-07,1.959441e-07,1.959443e-07,1.959445e-07,1.959446e-07,1.959448e-07,1.959450e-07,1.959451e-07,1.959453e-07,1.959455e-07,1.959456e-07,1.959458e-07,1.959460e-07,1.959461e-07,1.959463e-07,1.959465e-07,1.959466e-07,1.959468e-07,1.959469e-07,1.959471e-07,1.959473e-07,1.959474e-07,1.959476e-07,1.959478e-07,1.959479e-07,1.959481e-07,1.959483e-07,1.959484e-07,1.959486e-07,1.959488e-07,1.959489e-07,1.959491e-07,1.959493e-07,1.959494e-07,1.959496e-07,1.959498e-07,1.959499e-07,1.959501e-07,1.959503e-07,1.959504e-07,1.959506e-07,1.959507e-07,1.959509e-07,1.959511e-07,1.959512e-07,1.959514e-07,1.959516e-07,1.959517e-07,1.959519e-07,1.959521e-07,1.959522e-07,1.959524e-07,1.959526e-07,1.959527e-07,1.959529e-07,1.959531e-07,1.959532e-07,1.959534e-07,1.959536e-07,1.959537e-07,1.959539e-07,1.959540e-07,1.959542e-07,1.959544e-07,1.959545e-07,1.959547e-07,1.959549e-07,1.959550e-07,1.959552e-07,1.959554e-07,1.959555e-07,1.959557e-07,1.959559e-07,1.959560e-07,1.959562e-07,1.959564e-07,1.959565e-07,1.959567e-07,1.959569e-07,1.959570e-07,1.959572e-07,1.959573e-07,1.959575e-07,1.959577e-07,1.959578e-07,1.959580e-07,1.959582e-07,1.959583e-07,1.959585e-07,1.959587e-07,1.959588e-07,1.959590e-07,1.959592e-07,1.959593e-07,1.959595e-07,1.959597e-07,1.959598e-07,1.959600e-07,1.959602e-07,1.959603e-07,1.959605e-07,1.959606e-07,1.959608e-07,1.959610e-07,1.959611e-07,1.959613e-07,1.959615e-07,1.959616e-07,1.959618e-07,1.959620e-07,1.959621e-07,1.959623e-07,1.959625e-07,1.959626e-07,1.959628e-07,1.959630e-07,1.959631e-07,1.959633e-07,1.959634e-07,1.959636e-07,1.959638e-07,1.959639e-07,1.959641e-07,1.959643e-07,1.959644e-07,1.959646e-07,1.959648e-07,1.959649e-07,1.959651e-07,1.959653e-07,1.959654e-07,1.959656e-07,1.959658e-07,1.959659e-07,1.959661e-07,1.959663e-07,1.959664e-07,1.959666e-07,1.959667e-07,1.959669e-07,1.959671e-07,1.959672e-07,1.959674e-07,1.959676e-07,1.959677e-07,1.959679e-07,1.959681e-07,1.959682e-07,1.959684e-07,1.959686e-07,1.959687e-07,1.959689e-07,1.959691e-07,1.959692e-07,1.959694e-07,1.959695e-07,1.959697e-07,1.959699e-07,1.959700e-07,1.959702e-07,1.959704e-07,1.959705e-07,1.959707e-07,1.959709e-07,1.959710e-07,1.959712e-07,1.959714e-07,1.959715e-07,1.959717e-07,1.959719e-07,1.959720e-07,1.959722e-07,1.959724e-07,1.959725e-07,1.959727e-07,1.959728e-07,1.959730e-07,1.959732e-07,1.959733e-07,1.959735e-07,1.959737e-07,1.959738e-07,1.959740e-07,1.959742e-07,1.959743e-07,1.959745e-07,1.959747e-07,1.959748e-07,1.959750e-07,1.959752e-07,1.959753e-07,1.959755e-07,1.959756e-07,1.959758e-07,1.959760e-07,1.959761e-07,1.959763e-07,1.959765e-07,1.959766e-07,1.959768e-07,1.959770e-07,1.959771e-07,1.959773e-07,1.959775e-07,1.959776e-07,1.959778e-07,1.959780e-07,1.959781e-07,1.959783e-07,1.959784e-07,1.959786e-07,1.959788e-07,1.959789e-07,1.959791e-07,1.959793e-07,1.959794e-07,1.959796e-07,1.959798e-07,1.959799e-07,1.959801e-07,1.959803e-07,1.959804e-07,1.959806e-07,1.959808e-07,1.959809e-07,1.959811e-07,1.959812e-07,1.959814e-07,1.959816e-07,1.959817e-07,1.959819e-07,1.959821e-07,1.959822e-07,1.959824e-07,1.959826e-07,1.959827e-07,1.959829e-07,1.959831e-07,1.959832e-07,1.959834e-07,1.959835e-07,1.959837e-07,1.959839e-07,1.959840e-07,1.959842e-07,1.959844e-07,1.959845e-07,1.959847e-07,1.959849e-07,1.959850e-07,1.959852e-07,1.959854e-07,1.959855e-07,1.959857e-07,1.959859e-07,1.959860e-07,1.959862e-07,1.959863e-07,1.959865e-07,1.959867e-07,1.959868e-07,1.959870e-07,1.959872e-07,1.959873e-07,1.959875e-07,1.959877e-07,1.959878e-07,1.959880e-07,1.959882e-07,1.959883e-07,1.959885e-07,1.959887e-07,1.959888e-07,1.959890e-07,1.959891e-07,1.959893e-07,1.959895e-07,1.959896e-07,1.959898e-07,1.959900e-07,1.959901e-07,1.959903e-07,1.959905e-07,1.959906e-07,1.959908e-07,1.959910e-07,1.959911e-07,1.959913e-07,1.959914e-07,1.959916e-07,1.959918e-07,1.959919e-07,1.959921e-07,1.959923e-07,1.959924e-07,1.959926e-07,1.959928e-07,1.959929e-07,1.959931e-07,1.959933e-07,1.959934e-07,1.959936e-07,1.959937e-07,1.959939e-07,1.959941e-07,1.959942e-07,1.959944e-07,1.959946e-07,1.959947e-07,1.959949e-07,1.959951e-07,1.959952e-07,1.959954e-07,1.959956e-07,1.959957e-07,1.959959e-07,1.959961e-07,1.959962e-07,1.959964e-07,1.959965e-07,1.959967e-07,1.959969e-07,1.959970e-07,1.959972e-07,1.959974e-07,1.959975e-07,1.959977e-07,1.959979e-07,1.959980e-07,1.959982e-07,1.959984e-07,1.959985e-07,1.959987e-07,1.959988e-07,1.959990e-07,1.959992e-07,1.959993e-07,1.959995e-07,1.959997e-07,1.959998e-07,1.960000e-07,1.960002e-07,1.960003e-07,1.960005e-07,1.960007e-07,1.960008e-07,1.960010e-07,1.960011e-07,1.960013e-07,1.960015e-07,1.960016e-07,1.960018e-07,1.960020e-07,1.960021e-07,1.960023e-07,1.960025e-07,1.960026e-07,1.960028e-07,1.960030e-07,1.960031e-07,1.960033e-07,1.960034e-07,1.960036e-07,1.960038e-07,1.960039e-07,1.960041e-07,1.960043e-07,1.960044e-07,1.960046e-07,1.960048e-07,1.960049e-07,1.960051e-07,1.960053e-07,1.960054e-07,1.960056e-07,1.960057e-07,1.960059e-07,1.960061e-07,1.960062e-07,1.960064e-07,1.960066e-07,1.960067e-07,1.960069e-07,1.960071e-07,1.960072e-07,1.960074e-07,1.960076e-07,1.960077e-07,1.960079e-07,1.960080e-07,1.960082e-07,1.960084e-07,1.960085e-07,1.960087e-07,1.960089e-07,1.960090e-07,1.960092e-07,1.960094e-07,1.960095e-07,1.960097e-07,1.960099e-07,1.960100e-07,1.960102e-07,1.960103e-07,1.960105e-07,1.960107e-07,1.960108e-07,1.960110e-07,1.960112e-07,1.960113e-07,1.960115e-07,1.960117e-07,1.960118e-07,1.960120e-07,1.960122e-07,1.960123e-07,1.960125e-07,1.960126e-07,1.960128e-07,1.960130e-07,1.960131e-07,1.960133e-07,1.960135e-07,1.960136e-07,1.960138e-07,1.960140e-07,1.960141e-07,1.960143e-07,1.960145e-07,1.960146e-07,1.960148e-07,1.960149e-07,1.960151e-07,1.960153e-07,1.960154e-07,1.960156e-07,1.960158e-07,1.960159e-07,1.960161e-07,1.960163e-07,1.960164e-07,1.960166e-07,1.960168e-07,1.960169e-07,1.960171e-07,1.960172e-07,1.960174e-07,1.960176e-07,1.960177e-07,1.960179e-07,1.960181e-07,1.960182e-07,1.960184e-07,1.960186e-07,1.960187e-07,1.960189e-07,1.960190e-07,1.960192e-07,1.960194e-07,1.960195e-07,1.960197e-07,1.960199e-07,1.960200e-07,1.960202e-07,1.960204e-07,1.960205e-07,1.960207e-07,1.960209e-07,1.960210e-07,1.960212e-07,1.960213e-07,1.960215e-07,1.960217e-07,1.960218e-07,1.960220e-07,1.960222e-07,1.960223e-07,1.960225e-07,1.960227e-07,1.960228e-07,1.960230e-07,1.960232e-07,1.960233e-07,1.960235e-07,1.960236e-07,1.960238e-07,1.960240e-07,1.960241e-07,1.960243e-07,1.960245e-07,1.960246e-07,1.960248e-07,1.960250e-07,1.960251e-07,1.960253e-07,1.960254e-07,1.960256e-07,1.960258e-07,1.960259e-07,1.960261e-07,1.960263e-07,1.960264e-07,1.960266e-07,1.960268e-07,1.960269e-07,1.960271e-07,1.960273e-07,1.960274e-07,1.960276e-07,1.960277e-07,1.960279e-07,1.960281e-07,1.960282e-07,1.960284e-07,1.960286e-07,1.960287e-07,1.960289e-07,1.960291e-07,1.960292e-07,1.960294e-07,1.960295e-07,1.960297e-07,1.960299e-07,1.960300e-07,1.960302e-07,1.960304e-07,1.960305e-07,1.960307e-07,1.960309e-07,1.960310e-07,1.960312e-07,1.960314e-07,1.960315e-07,1.960317e-07,1.960318e-07,1.960320e-07,1.960322e-07,1.960323e-07,1.960325e-07,1.960327e-07,1.960328e-07,1.960330e-07,1.960332e-07,1.960333e-07,1.960335e-07,1.960336e-07,1.960338e-07,1.960340e-07,1.960341e-07,1.960343e-07,1.960345e-07,1.960346e-07,1.960348e-07,1.960350e-07,1.960351e-07,1.960353e-07,1.960354e-07,1.960356e-07,1.960358e-07,1.960359e-07,1.960361e-07,1.960363e-07,1.960364e-07,1.960366e-07,1.960368e-07,1.960369e-07,1.960371e-07,1.960373e-07,1.960374e-07,1.960376e-07,1.960377e-07,1.960379e-07,1.960381e-07,1.960382e-07,1.960384e-07,1.960386e-07,1.960387e-07,1.960389e-07,1.960391e-07,1.960392e-07,1.960394e-07,1.960395e-07,1.960397e-07,1.960399e-07,1.960400e-07,1.960402e-07,1.960404e-07,1.960405e-07,1.960407e-07,1.960409e-07,1.960410e-07,1.960412e-07,1.960413e-07,1.960415e-07,1.960417e-07,1.960418e-07,1.960420e-07,1.960422e-07,1.960423e-07,1.960425e-07,1.960427e-07,1.960428e-07,1.960430e-07,1.960431e-07,1.960433e-07,1.960435e-07,1.960436e-07,1.960438e-07,1.960440e-07,1.960441e-07,1.960443e-07,1.960445e-07,1.960446e-07,1.960448e-07,1.960450e-07,1.960451e-07,1.960453e-07,1.960454e-07,1.960456e-07,1.960458e-07,1.960459e-07,1.960461e-07,1.960463e-07,1.960464e-07,1.960466e-07,1.960468e-07,1.960469e-07,1.960471e-07,1.960472e-07,1.960474e-07,1.960476e-07,1.960477e-07,1.960479e-07,1.960481e-07,1.960482e-07,1.960484e-07,1.960486e-07,1.960487e-07,1.960489e-07,1.960490e-07,1.960492e-07,1.960494e-07,1.960495e-07,1.960497e-07,1.960499e-07,1.960500e-07,1.960502e-07,1.960504e-07,1.960505e-07,1.960507e-07,1.960508e-07,1.960510e-07,1.960512e-07,1.960513e-07,1.960515e-07,1.960517e-07,1.960518e-07,1.960520e-07,1.960522e-07,1.960523e-07,1.960525e-07,1.960526e-07,1.960528e-07,1.960530e-07,1.960531e-07,1.960533e-07,1.960535e-07,1.960536e-07,1.960538e-07,1.960540e-07,1.960541e-07,1.960543e-07,1.960544e-07,1.960546e-07,1.960548e-07,1.960549e-07,1.960551e-07,1.960553e-07,1.960554e-07,1.960556e-07,1.960558e-07,1.960559e-07,1.960561e-07,1.960562e-07,1.960564e-07,1.960566e-07,1.960567e-07,1.960569e-07,1.960571e-07,1.960572e-07,1.960574e-07,1.960576e-07,1.960577e-07,1.960579e-07,1.960580e-07,1.960582e-07,1.960584e-07,1.960585e-07,1.960587e-07,1.960589e-07,1.960590e-07,1.960592e-07,1.960594e-07,1.960595e-07,1.960597e-07,1.960598e-07,1.960600e-07,1.960602e-07,1.960603e-07,1.960605e-07,1.960607e-07,1.960608e-07,1.960610e-07,1.960611e-07,1.960613e-07,1.960615e-07,1.960616e-07,1.960618e-07,1.960620e-07,1.960621e-07,1.960623e-07,1.960625e-07,1.960626e-07,1.960628e-07,1.960629e-07,1.960631e-07,1.960633e-07,1.960634e-07,1.960636e-07,1.960638e-07,1.960639e-07,1.960641e-07,1.960643e-07,1.960644e-07,1.960646e-07,1.960647e-07,1.960649e-07,1.960651e-07,1.960652e-07,1.960654e-07,1.960656e-07,1.960657e-07,1.960659e-07,1.960661e-07,1.960662e-07,1.960664e-07,1.960665e-07,1.960667e-07,1.960669e-07,1.960670e-07,1.960672e-07,1.960674e-07,1.960675e-07,1.960677e-07,1.960679e-07,1.960680e-07,1.960682e-07,1.960683e-07,1.960685e-07,1.960687e-07,1.960688e-07,1.960690e-07,1.960692e-07,1.960693e-07,1.960695e-07,1.960696e-07,1.960698e-07,1.960700e-07,1.960701e-07,1.960703e-07,1.960705e-07,1.960706e-07,1.960708e-07,1.960710e-07,1.960711e-07,1.960713e-07,1.960714e-07,1.960716e-07,1.960718e-07,1.960719e-07,1.960721e-07,1.960723e-07,1.960724e-07,1.960726e-07,1.960728e-07,1.960729e-07,1.960731e-07,1.960732e-07,1.960734e-07,1.960736e-07,1.960737e-07,1.960739e-07,1.960741e-07,1.960742e-07,1.960744e-07,1.960746e-07,1.960747e-07,1.960749e-07,1.960750e-07,1.960752e-07,1.960754e-07,1.960755e-07,1.960757e-07,1.960759e-07,1.960760e-07,1.960762e-07,1.960763e-07,1.960765e-07,1.960767e-07,1.960768e-07,1.960770e-07,1.960772e-07,1.960773e-07,1.960775e-07,1.960777e-07,1.960778e-07,1.960780e-07,1.960781e-07,1.960783e-07,1.960785e-07,1.960786e-07,1.960788e-07,1.960790e-07,1.960791e-07,1.960793e-07,1.960794e-07,1.960796e-07,1.960798e-07,1.960799e-07,1.960801e-07,1.960803e-07,1.960804e-07,1.960806e-07,1.960808e-07,1.960809e-07,1.960811e-07,1.960812e-07,1.960814e-07,1.960816e-07,1.960817e-07,1.960819e-07,1.960821e-07,1.960822e-07,1.960824e-07,1.960826e-07,1.960827e-07,1.960829e-07,1.960830e-07,1.960832e-07,1.960834e-07,1.960835e-07,1.960837e-07,1.960839e-07,1.960840e-07,1.960842e-07,1.960843e-07,1.960845e-07,1.960847e-07,1.960848e-07,1.960850e-07,1.960852e-07,1.960853e-07,1.960855e-07,1.960857e-07,1.960858e-07,1.960860e-07,1.960861e-07,1.960863e-07,1.960865e-07,1.960866e-07,1.960868e-07,1.960870e-07,1.960871e-07,1.960873e-07,1.960874e-07,1.960876e-07,1.960878e-07,1.960879e-07,1.960881e-07,1.960883e-07,1.960884e-07,1.960886e-07,1.960888e-07,1.960889e-07,1.960891e-07,1.960892e-07,1.960894e-07,1.960896e-07,1.960897e-07,1.960899e-07,1.960901e-07,1.960902e-07,1.960904e-07,1.960905e-07,1.960907e-07,1.960909e-07,1.960910e-07,1.960912e-07,1.960914e-07,1.960915e-07,1.960917e-07,1.960919e-07,1.960920e-07,1.960922e-07,1.960923e-07,1.960925e-07,1.960927e-07,1.960928e-07,1.960930e-07,1.960932e-07,1.960933e-07,1.960935e-07,1.960936e-07,1.960938e-07,1.960940e-07,1.960941e-07,1.960943e-07,1.960945e-07,1.960946e-07,1.960948e-07,1.960949e-07,1.960951e-07,1.960953e-07,1.960954e-07,1.960956e-07,1.960958e-07,1.960959e-07,1.960961e-07,1.960963e-07,1.960964e-07,1.960966e-07,1.960967e-07,1.960969e-07,1.960971e-07,1.960972e-07,1.960974e-07,1.960976e-07,1.960977e-07,1.960979e-07,1.960980e-07,1.960982e-07,1.960984e-07,1.960985e-07,1.960987e-07,1.960989e-07,1.960990e-07,1.960992e-07,1.960994e-07,1.960995e-07,1.960997e-07,1.960998e-07,1.961000e-07,1.961002e-07,1.961003e-07,1.961005e-07,1.961007e-07,1.961008e-07,1.961010e-07,1.961011e-07,1.961013e-07,1.961015e-07,1.961016e-07,1.961018e-07,1.961020e-07,1.961021e-07,1.961023e-07,1.961024e-07,1.961026e-07,1.961028e-07,1.961029e-07,1.961031e-07,1.961033e-07,1.961034e-07,1.961036e-07,1.961038e-07,1.961039e-07,1.961041e-07,1.961042e-07,1.961044e-07,1.961046e-07,1.961047e-07,1.961049e-07,1.961051e-07,1.961052e-07,1.961054e-07,1.961055e-07,1.961057e-07,1.961059e-07,1.961060e-07,1.961062e-07,1.961064e-07,1.961065e-07,1.961067e-07,1.961068e-07,1.961070e-07,1.961072e-07,1.961073e-07,1.961075e-07,1.961077e-07,1.961078e-07,1.961080e-07,1.961081e-07,1.961083e-07,1.961085e-07,1.961086e-07,1.961088e-07,1.961090e-07,1.961091e-07,1.961093e-07,1.961095e-07,1.961096e-07,1.961098e-07,1.961099e-07,1.961101e-07,1.961103e-07,1.961104e-07,1.961106e-07,1.961108e-07,1.961109e-07,1.961111e-07,1.961112e-07,1.961114e-07,1.961116e-07,1.961117e-07,1.961119e-07,1.961121e-07,1.961122e-07,1.961124e-07,1.961125e-07,1.961127e-07,1.961129e-07,1.961130e-07,1.961132e-07,1.961134e-07,1.961135e-07,1.961137e-07,1.961138e-07,1.961140e-07,1.961142e-07,1.961143e-07,1.961145e-07,1.961147e-07,1.961148e-07,1.961150e-07,1.961151e-07,1.961153e-07,1.961155e-07,1.961156e-07,1.961158e-07,1.961160e-07,1.961161e-07,1.961163e-07,1.961165e-07,1.961166e-07,1.961168e-07,1.961169e-07,1.961171e-07,1.961173e-07,1.961174e-07,1.961176e-07,1.961178e-07,1.961179e-07,1.961181e-07,1.961182e-07,1.961184e-07,1.961186e-07,1.961187e-07,1.961189e-07,1.961191e-07,1.961192e-07,1.961194e-07,1.961195e-07,1.961197e-07,1.961199e-07,1.961200e-07,1.961202e-07,1.961204e-07,1.961205e-07,1.961207e-07,1.961208e-07,1.961210e-07,1.961212e-07,1.961213e-07,1.961215e-07,1.961217e-07,1.961218e-07,1.961220e-07,1.961221e-07,1.961223e-07,1.961225e-07,1.961226e-07,1.961228e-07,1.961230e-07,1.961231e-07,1.961233e-07,1.961234e-07,1.961236e-07,1.961238e-07,1.961239e-07,1.961241e-07,1.961243e-07,1.961244e-07,1.961246e-07,1.961247e-07,1.961249e-07,1.961251e-07,1.961252e-07,1.961254e-07,1.961256e-07,1.961257e-07,1.961259e-07,1.961260e-07,1.961262e-07,1.961264e-07,1.961265e-07,1.961267e-07,1.961269e-07,1.961270e-07,1.961272e-07,1.961274e-07,1.961275e-07,1.961277e-07,1.961278e-07,1.961280e-07,1.961282e-07,1.961283e-07,1.961285e-07,1.961287e-07,1.961288e-07,1.961290e-07,1.961291e-07,1.961293e-07,1.961295e-07,1.961296e-07,1.961298e-07,1.961300e-07,1.961301e-07,1.961303e-07,1.961304e-07,1.961306e-07,1.961308e-07,1.961309e-07,1.961311e-07,1.961313e-07,1.961314e-07,1.961316e-07,1.961317e-07,1.961319e-07,1.961321e-07,1.961322e-07,1.961324e-07,1.961326e-07,1.961327e-07,1.961329e-07,1.961330e-07,1.961332e-07,1.961334e-07,1.961335e-07,1.961337e-07,1.961339e-07,1.961340e-07,1.961342e-07,1.961343e-07,1.961345e-07,1.961347e-07,1.961348e-07,1.961350e-07,1.961352e-07,1.961353e-07,1.961355e-07,1.961356e-07,1.961358e-07,1.961360e-07,1.961361e-07,1.961363e-07,1.961365e-07,1.961366e-07,1.961368e-07,1.961369e-07,1.961371e-07,1.961373e-07,1.961374e-07,1.961376e-07,1.961378e-07,1.961379e-07,1.961381e-07,1.961382e-07,1.961384e-07,1.961386e-07,1.961387e-07,1.961389e-07,1.961391e-07,1.961392e-07,1.961394e-07,1.961395e-07,1.961397e-07,1.961399e-07,1.961400e-07,1.961402e-07,1.961404e-07,1.961405e-07,1.961407e-07,1.961408e-07,1.961410e-07,1.961412e-07,1.961413e-07,1.961415e-07,1.961417e-07,1.961418e-07,1.961420e-07,1.961421e-07,1.961423e-07,1.961425e-07,1.961426e-07,1.961428e-07,1.961429e-07,1.961431e-07,1.961433e-07,1.961434e-07,1.961436e-07,1.961438e-07,1.961439e-07,1.961441e-07,1.961442e-07,1.961444e-07,1.961446e-07,1.961447e-07,1.961449e-07,1.961451e-07,1.961452e-07,1.961454e-07,1.961455e-07,1.961457e-07,1.961459e-07,1.961460e-07,1.961462e-07,1.961464e-07,1.961465e-07,1.961467e-07,1.961468e-07,1.961470e-07,1.961472e-07,1.961473e-07,1.961475e-07,1.961477e-07,1.961478e-07,1.961480e-07,1.961481e-07,1.961483e-07,1.961485e-07,1.961486e-07,1.961488e-07,1.961490e-07,1.961491e-07,1.961493e-07,1.961494e-07,1.961496e-07,1.961498e-07,1.961499e-07,1.961501e-07,1.961503e-07,1.961504e-07,1.961506e-07,1.961507e-07,1.961509e-07,1.961511e-07,1.961512e-07,1.961514e-07,1.961516e-07,1.961517e-07,1.961519e-07,1.961520e-07,1.961522e-07,1.961524e-07,1.961525e-07,1.961527e-07,1.961529e-07,1.961530e-07,1.961532e-07,1.961533e-07,1.961535e-07,1.961537e-07,1.961538e-07,1.961540e-07,1.961541e-07,1.961543e-07,1.961545e-07,1.961546e-07,1.961548e-07,1.961550e-07,1.961551e-07,1.961553e-07,1.961554e-07,1.961556e-07,1.961558e-07,1.961559e-07,1.961561e-07,1.961563e-07,1.961564e-07,1.961566e-07,1.961567e-07,1.961569e-07,1.961571e-07,1.961572e-07,1.961574e-07,1.961576e-07,1.961577e-07,1.961579e-07,1.961580e-07,1.961582e-07,1.961584e-07,1.961585e-07,1.961587e-07,1.961589e-07,1.961590e-07,1.961592e-07,1.961593e-07,1.961595e-07,1.961597e-07,1.961598e-07,1.961600e-07,1.961601e-07,1.961603e-07,1.961605e-07,1.961606e-07,1.961608e-07,1.961610e-07,1.961611e-07,1.961613e-07,1.961614e-07,1.961616e-07,1.961618e-07,1.961619e-07,1.961621e-07,1.961623e-07,1.961624e-07,1.961626e-07,1.961627e-07,1.961629e-07,1.961631e-07,1.961632e-07,1.961634e-07,1.961636e-07,1.961637e-07,1.961639e-07,1.961640e-07,1.961642e-07,1.961644e-07,1.961645e-07,1.961647e-07,1.961649e-07,1.961650e-07,1.961652e-07,1.961653e-07,1.961655e-07,1.961657e-07,1.961658e-07,1.961660e-07,1.961661e-07,1.961663e-07,1.961665e-07,1.961666e-07,1.961668e-07,1.961670e-07,1.961671e-07,1.961673e-07,1.961674e-07,1.961676e-07,1.961678e-07,1.961679e-07,1.961681e-07,1.961683e-07,1.961684e-07,1.961686e-07,1.961687e-07,1.961689e-07,1.961691e-07,1.961692e-07,1.961694e-07,1.961695e-07,1.961697e-07,1.961699e-07,1.961700e-07,1.961702e-07,1.961704e-07,1.961705e-07,1.961707e-07,1.961708e-07,1.961710e-07,1.961712e-07,1.961713e-07,1.961715e-07,1.961717e-07,1.961718e-07,1.961720e-07,1.961721e-07,1.961723e-07,1.961725e-07,1.961726e-07,1.961728e-07,1.961730e-07,1.961731e-07,1.961733e-07,1.961734e-07,1.961736e-07,1.961738e-07,1.961739e-07,1.961741e-07,1.961742e-07,1.961744e-07,1.961746e-07,1.961747e-07,1.961749e-07,1.961751e-07,1.961752e-07,1.961754e-07,1.961755e-07,1.961757e-07,1.961759e-07,1.961760e-07,1.961762e-07,1.961764e-07,1.961765e-07,1.961767e-07,1.961768e-07,1.961770e-07,1.961772e-07,1.961773e-07,1.961775e-07,1.961776e-07,1.961778e-07,1.961780e-07,1.961781e-07,1.961783e-07,1.961785e-07,1.961786e-07,1.961788e-07,1.961789e-07,1.961791e-07,1.961793e-07,1.961794e-07,1.961796e-07,1.961798e-07,1.961799e-07,1.961801e-07,1.961802e-07,1.961804e-07,1.961806e-07,1.961807e-07,1.961809e-07,1.961810e-07,1.961812e-07,1.961814e-07,1.961815e-07,1.961817e-07,1.961819e-07,1.961820e-07,1.961822e-07,1.961823e-07,1.961825e-07,1.961827e-07,1.961828e-07,1.961830e-07,1.961832e-07,1.961833e-07,1.961835e-07,1.961836e-07,1.961838e-07,1.961840e-07,1.961841e-07,1.961843e-07,1.961844e-07,1.961846e-07,1.961848e-07,1.961849e-07,1.961851e-07,1.961853e-07,1.961854e-07,1.961856e-07,1.961857e-07,1.961859e-07,1.961861e-07,1.961862e-07,1.961864e-07,1.961865e-07,1.961867e-07,1.961869e-07,1.961870e-07,1.961872e-07,1.961874e-07,1.961875e-07,1.961877e-07,1.961878e-07,1.961880e-07,1.961882e-07,1.961883e-07,1.961885e-07,1.961887e-07,1.961888e-07,1.961890e-07,1.961891e-07,1.961893e-07,1.961895e-07,1.961896e-07,1.961898e-07,1.961899e-07,1.961901e-07,1.961903e-07,1.961904e-07,1.961906e-07,1.961908e-07,1.961909e-07,1.961911e-07,1.961912e-07,1.961914e-07,1.961916e-07,1.961917e-07,1.961919e-07,1.961920e-07,1.961922e-07,1.961924e-07,1.961925e-07,1.961927e-07,1.961929e-07,1.961930e-07,1.961932e-07,1.961933e-07,1.961935e-07,1.961937e-07,1.961938e-07,1.961940e-07,1.961941e-07,1.961943e-07,1.961945e-07,1.961946e-07,1.961948e-07,1.961950e-07,1.961951e-07,1.961953e-07,1.961954e-07,1.961956e-07,1.961958e-07,1.961959e-07,1.961961e-07,1.961963e-07,1.961964e-07,1.961966e-07,1.961967e-07,1.961969e-07,1.961971e-07,1.961972e-07,1.961974e-07,1.961975e-07,1.961977e-07,1.961979e-07,1.961980e-07,1.961982e-07,1.961984e-07,1.961985e-07,1.961987e-07,1.961988e-07,1.961990e-07,1.961992e-07,1.961993e-07,1.961995e-07,1.961996e-07,1.961998e-07,1.962000e-07,1.962001e-07,1.962003e-07,1.962005e-07,1.962006e-07,1.962008e-07,1.962009e-07,1.962011e-07,1.962013e-07,1.962014e-07,1.962016e-07,1.962017e-07,1.962019e-07,1.962021e-07,1.962022e-07,1.962024e-07,1.962026e-07,1.962027e-07,1.962029e-07,1.962030e-07,1.962032e-07,1.962034e-07,1.962035e-07,1.962037e-07,1.962038e-07,1.962040e-07,1.962042e-07,1.962043e-07,1.962045e-07,1.962047e-07,1.962048e-07,1.962050e-07,1.962051e-07,1.962053e-07,1.962055e-07,1.962056e-07,1.962058e-07,1.962059e-07,1.962061e-07,1.962063e-07,1.962064e-07,1.962066e-07,1.962068e-07,1.962069e-07,1.962071e-07,1.962072e-07,1.962074e-07,1.962076e-07,1.962077e-07,1.962079e-07,1.962080e-07,1.962082e-07,1.962084e-07,1.962085e-07,1.962087e-07,1.962089e-07,1.962090e-07,1.962092e-07,1.962093e-07,1.962095e-07,1.962097e-07,1.962098e-07,1.962100e-07,1.962101e-07,1.962103e-07,1.962105e-07,1.962106e-07,1.962108e-07,1.962110e-07,1.962111e-07,1.962113e-07,1.962114e-07,1.962116e-07,1.962118e-07,1.962119e-07,1.962121e-07,1.962122e-07,1.962124e-07,1.962126e-07,1.962127e-07,1.962129e-07,1.962131e-07,1.962132e-07,1.962134e-07,1.962135e-07,1.962137e-07,1.962139e-07,1.962140e-07,1.962142e-07,1.962143e-07,1.962145e-07,1.962147e-07,1.962148e-07,1.962150e-07,1.962151e-07,1.962153e-07,1.962155e-07,1.962156e-07,1.962158e-07,1.962160e-07,1.962161e-07,1.962163e-07,1.962164e-07,1.962166e-07,1.962168e-07,1.962169e-07,1.962171e-07,1.962172e-07,1.962174e-07,1.962176e-07,1.962177e-07,1.962179e-07,1.962181e-07,1.962182e-07,1.962184e-07,1.962185e-07,1.962187e-07,1.962189e-07,1.962190e-07,1.962192e-07,1.962193e-07,1.962195e-07,1.962197e-07,1.962198e-07,1.962200e-07,1.962202e-07,1.962203e-07,1.962205e-07,1.962206e-07,1.962208e-07,1.962210e-07,1.962211e-07,1.962213e-07,1.962214e-07,1.962216e-07,1.962218e-07,1.962219e-07,1.962221e-07,1.962222e-07,1.962224e-07,1.962226e-07,1.962227e-07,1.962229e-07,1.962231e-07,1.962232e-07,1.962234e-07,1.962235e-07,1.962237e-07,1.962239e-07,1.962240e-07,1.962242e-07,1.962243e-07,1.962245e-07,1.962247e-07,1.962248e-07,1.962250e-07,1.962251e-07,1.962253e-07,1.962255e-07,1.962256e-07,1.962258e-07,1.962260e-07,1.962261e-07,1.962263e-07,1.962264e-07,1.962266e-07,1.962268e-07,1.962269e-07,1.962271e-07,1.962272e-07,1.962274e-07,1.962276e-07,1.962277e-07,1.962279e-07,1.962281e-07,1.962282e-07,1.962284e-07,1.962285e-07,1.962287e-07,1.962289e-07,1.962290e-07,1.962292e-07,1.962293e-07,1.962295e-07,1.962297e-07,1.962298e-07,1.962300e-07,1.962301e-07,1.962303e-07,1.962305e-07,1.962306e-07,1.962308e-07,1.962310e-07,1.962311e-07,1.962313e-07,1.962314e-07,1.962316e-07,1.962318e-07,1.962319e-07,1.962321e-07,1.962322e-07,1.962324e-07,1.962326e-07,1.962327e-07,1.962329e-07,1.962330e-07,1.962332e-07,1.962334e-07,1.962335e-07,1.962337e-07,1.962339e-07,1.962340e-07,1.962342e-07,1.962343e-07,1.962345e-07,1.962347e-07,1.962348e-07,1.962350e-07,1.962351e-07,1.962353e-07,1.962355e-07,1.962356e-07,1.962358e-07,1.962359e-07,1.962361e-07,1.962363e-07,1.962364e-07,1.962366e-07,1.962368e-07,1.962369e-07,1.962371e-07,1.962372e-07,1.962374e-07,1.962376e-07,1.962377e-07,1.962379e-07,1.962380e-07,1.962382e-07,1.962384e-07,1.962385e-07,1.962387e-07,1.962388e-07,1.962390e-07,1.962392e-07,1.962393e-07,1.962395e-07,1.962397e-07,1.962398e-07,1.962400e-07,1.962401e-07,1.962403e-07,1.962405e-07,1.962406e-07,1.962408e-07,1.962409e-07,1.962411e-07,1.962413e-07,1.962414e-07,1.962416e-07,1.962417e-07,1.962419e-07,1.962421e-07,1.962422e-07,1.962424e-07,1.962426e-07,1.962427e-07,1.962429e-07,1.962430e-07,1.962432e-07,1.962434e-07,1.962435e-07,1.962437e-07,1.962438e-07,1.962440e-07,1.962442e-07,1.962443e-07,1.962445e-07,1.962446e-07,1.962448e-07,1.962450e-07,1.962451e-07,1.962453e-07,1.962454e-07,1.962456e-07,1.962458e-07,1.962459e-07,1.962461e-07,1.962463e-07,1.962464e-07,1.962466e-07,1.962467e-07,1.962469e-07,1.962471e-07,1.962472e-07,1.962474e-07,1.962475e-07,1.962477e-07,1.962479e-07,1.962480e-07,1.962482e-07,1.962483e-07,1.962485e-07,1.962487e-07,1.962488e-07,1.962490e-07,1.962492e-07,1.962493e-07,1.962495e-07,1.962496e-07,1.962498e-07,1.962500e-07,1.962501e-07,1.962503e-07,1.962504e-07,1.962506e-07,1.962508e-07,1.962509e-07,1.962511e-07,1.962512e-07,1.962514e-07,1.962516e-07,1.962517e-07,1.962519e-07,1.962520e-07,1.962522e-07,1.962524e-07,1.962525e-07,1.962527e-07,1.962529e-07,1.962530e-07,1.962532e-07,1.962533e-07,1.962535e-07,1.962537e-07,1.962538e-07,1.962540e-07,1.962541e-07,1.962543e-07,1.962545e-07,1.962546e-07,1.962548e-07,1.962549e-07,1.962551e-07,1.962553e-07,1.962554e-07,1.962556e-07,1.962557e-07,1.962559e-07,1.962561e-07,1.962562e-07,1.962564e-07,1.962566e-07,1.962567e-07,1.962569e-07,1.962570e-07,1.962572e-07,1.962574e-07,1.962575e-07,1.962577e-07,1.962578e-07,1.962580e-07,1.962582e-07,1.962583e-07,1.962585e-07,1.962586e-07,1.962588e-07,1.962590e-07,1.962591e-07,1.962593e-07,1.962594e-07,1.962596e-07,1.962598e-07,1.962599e-07,1.962601e-07,1.962602e-07,1.962604e-07,1.962606e-07,1.962607e-07,1.962609e-07,1.962611e-07,1.962612e-07,1.962614e-07,1.962615e-07,1.962617e-07,1.962619e-07,1.962620e-07,1.962622e-07,1.962623e-07,1.962625e-07,1.962627e-07,1.962628e-07,1.962630e-07,1.962631e-07,1.962633e-07,1.962635e-07,1.962636e-07,1.962638e-07,1.962639e-07,1.962641e-07,1.962643e-07,1.962644e-07,1.962646e-07,1.962647e-07,1.962649e-07,1.962651e-07,1.962652e-07,1.962654e-07,1.962656e-07,1.962657e-07,1.962659e-07,1.962660e-07,1.962662e-07,1.962664e-07,1.962665e-07,1.962667e-07,1.962668e-07,1.962670e-07,1.962672e-07,1.962673e-07,1.962675e-07,1.962676e-07,1.962678e-07,1.962680e-07,1.962681e-07,1.962683e-07,1.962684e-07,1.962686e-07,1.962688e-07,1.962689e-07,1.962691e-07,1.962692e-07,1.962694e-07,1.962696e-07,1.962697e-07,1.962699e-07,1.962701e-07,1.962702e-07,1.962704e-07,1.962705e-07,1.962707e-07,1.962709e-07,1.962710e-07,1.962712e-07,1.962713e-07,1.962715e-07,1.962717e-07,1.962718e-07,1.962720e-07,1.962721e-07,1.962723e-07,1.962725e-07,1.962726e-07,1.962728e-07,1.962729e-07,1.962731e-07,1.962733e-07,1.962734e-07,1.962736e-07,1.962737e-07,1.962739e-07,1.962741e-07,1.962742e-07,1.962744e-07,1.962745e-07,1.962747e-07,1.962749e-07,1.962750e-07,1.962752e-07,1.962754e-07,1.962755e-07,1.962757e-07,1.962758e-07,1.962760e-07,1.962762e-07,1.962763e-07,1.962765e-07,1.962766e-07,1.962768e-07,1.962770e-07,1.962771e-07,1.962773e-07,1.962774e-07,1.962776e-07,1.962778e-07,1.962779e-07,1.962781e-07,1.962782e-07,1.962784e-07,1.962786e-07,1.962787e-07,1.962789e-07,1.962790e-07,1.962792e-07,1.962794e-07,1.962795e-07,1.962797e-07,1.962798e-07,1.962800e-07,1.962802e-07,1.962803e-07,1.962805e-07,1.962806e-07,1.962808e-07,1.962810e-07,1.962811e-07,1.962813e-07,1.962815e-07,1.962816e-07,1.962818e-07,1.962819e-07,1.962821e-07,1.962823e-07,1.962824e-07,1.962826e-07,1.962827e-07,1.962829e-07,1.962831e-07,1.962832e-07,1.962834e-07,1.962835e-07,1.962837e-07,1.962839e-07,1.962840e-07,1.962842e-07,1.962843e-07,1.962845e-07,1.962847e-07,1.962848e-07,1.962850e-07,1.962851e-07,1.962853e-07,1.962855e-07,1.962856e-07,1.962858e-07,1.962859e-07,1.962861e-07,1.962863e-07,1.962864e-07,1.962866e-07,1.962867e-07,1.962869e-07,1.962871e-07,1.962872e-07,1.962874e-07,1.962875e-07,1.962877e-07,1.962879e-07,1.962880e-07,1.962882e-07,1.962883e-07,1.962885e-07,1.962887e-07,1.962888e-07,1.962890e-07,1.962892e-07,1.962893e-07,1.962895e-07,1.962896e-07,1.962898e-07,1.962900e-07,1.962901e-07,1.962903e-07,1.962904e-07,1.962906e-07,1.962908e-07,1.962909e-07,1.962911e-07,1.962912e-07,1.962914e-07,1.962916e-07,1.962917e-07,1.962919e-07,1.962920e-07,1.962922e-07,1.962924e-07,1.962925e-07,1.962927e-07,1.962928e-07,1.962930e-07,1.962932e-07,1.962933e-07,1.962935e-07,1.962936e-07,1.962938e-07,1.962940e-07,1.962941e-07,1.962943e-07,1.962944e-07,1.962946e-07,1.962948e-07,1.962949e-07,1.962951e-07,1.962952e-07,1.962954e-07,1.962956e-07,1.962957e-07,1.962959e-07,1.962960e-07,1.962962e-07,1.962964e-07,1.962965e-07,1.962967e-07,1.962968e-07,1.962970e-07,1.962972e-07,1.962973e-07,1.962975e-07,1.962976e-07,1.962978e-07,1.962980e-07,1.962981e-07,1.962983e-07,1.962984e-07,1.962986e-07,1.962988e-07,1.962989e-07,1.962991e-07,1.962992e-07,1.962994e-07,1.962996e-07,1.962997e-07,1.962999e-07,1.963001e-07,1.963002e-07,1.963004e-07,1.963005e-07,1.963007e-07,1.963009e-07,1.963010e-07,1.963012e-07,1.963013e-07,1.963015e-07,1.963017e-07,1.963018e-07,1.963020e-07,1.963021e-07,1.963023e-07,1.963025e-07,1.963026e-07,1.963028e-07,1.963029e-07,1.963031e-07,1.963033e-07,1.963034e-07,1.963036e-07,1.963037e-07,1.963039e-07,1.963041e-07,1.963042e-07,1.963044e-07,1.963045e-07,1.963047e-07,1.963049e-07,1.963050e-07,1.963052e-07,1.963053e-07,1.963055e-07,1.963057e-07,1.963058e-07,1.963060e-07,1.963061e-07,1.963063e-07,1.963065e-07,1.963066e-07,1.963068e-07,1.963069e-07,1.963071e-07,1.963073e-07,1.963074e-07,1.963076e-07,1.963077e-07,1.963079e-07,1.963081e-07,1.963082e-07,1.963084e-07,1.963085e-07,1.963087e-07,1.963089e-07,1.963090e-07,1.963092e-07,1.963093e-07,1.963095e-07,1.963097e-07,1.963098e-07,1.963100e-07,1.963101e-07,1.963103e-07,1.963105e-07,1.963106e-07,1.963108e-07,1.963109e-07,1.963111e-07,1.963113e-07,1.963114e-07,1.963116e-07,1.963117e-07,1.963119e-07,1.963121e-07,1.963122e-07,1.963124e-07,1.963125e-07,1.963127e-07,1.963129e-07,1.963130e-07,1.963132e-07,1.963133e-07,1.963135e-07,1.963137e-07,1.963138e-07,1.963140e-07,1.963141e-07,1.963143e-07,1.963145e-07,1.963146e-07,1.963148e-07,1.963149e-07,1.963151e-07,1.963153e-07,1.963154e-07,1.963156e-07,1.963157e-07,1.963159e-07,1.963161e-07,1.963162e-07,1.963164e-07,1.963165e-07,1.963167e-07,1.963169e-07,1.963170e-07,1.963172e-07,1.963173e-07,1.963175e-07,1.963177e-07,1.963178e-07,1.963180e-07,1.963181e-07,1.963183e-07,1.963185e-07,1.963186e-07,1.963188e-07,1.963189e-07,1.963191e-07,1.963193e-07,1.963194e-07,1.963196e-07,1.963197e-07,1.963199e-07,1.963201e-07,1.963202e-07,1.963204e-07,1.963205e-07,1.963207e-07,1.963209e-07,1.963210e-07,1.963212e-07,1.963213e-07,1.963215e-07,1.963217e-07,1.963218e-07,1.963220e-07,1.963221e-07,1.963223e-07,1.963225e-07,1.963226e-07,1.963228e-07,1.963229e-07,1.963231e-07,1.963233e-07,1.963234e-07,1.963236e-07,1.963237e-07,1.963239e-07,1.963241e-07,1.963242e-07,1.963244e-07,1.963245e-07,1.963247e-07,1.963249e-07,1.963250e-07,1.963252e-07,1.963253e-07,1.963255e-07,1.963257e-07,1.963258e-07,1.963260e-07,1.963261e-07,1.963263e-07,1.963265e-07,1.963266e-07,1.963268e-07,1.963269e-07,1.963271e-07,1.963273e-07,1.963274e-07,1.963276e-07,1.963277e-07,1.963279e-07,1.963281e-07,1.963282e-07,1.963284e-07,1.963285e-07,1.963287e-07,1.963289e-07,1.963290e-07,1.963292e-07,1.963293e-07,1.963295e-07,1.963297e-07,1.963298e-07,1.963300e-07,1.963301e-07,1.963303e-07,1.963305e-07,1.963306e-07,1.963308e-07,1.963309e-07,1.963311e-07,1.963313e-07,1.963314e-07,1.963316e-07,1.963317e-07,1.963319e-07,1.963320e-07,1.963322e-07,1.963324e-07,1.963325e-07,1.963327e-07,1.963328e-07,1.963330e-07,1.963332e-07,1.963333e-07,1.963335e-07,1.963336e-07,1.963338e-07,1.963340e-07,1.963341e-07,1.963343e-07,1.963344e-07,1.963346e-07,1.963348e-07,1.963349e-07,1.963351e-07,1.963352e-07,1.963354e-07,1.963356e-07,1.963357e-07,1.963359e-07,1.963360e-07,1.963362e-07,1.963364e-07,1.963365e-07,1.963367e-07,1.963368e-07,1.963370e-07,1.963372e-07,1.963373e-07,1.963375e-07,1.963376e-07,1.963378e-07,1.963380e-07,1.963381e-07,1.963383e-07,1.963384e-07,1.963386e-07,1.963388e-07,1.963389e-07,1.963391e-07,1.963392e-07,1.963394e-07,1.963396e-07,1.963397e-07,1.963399e-07,1.963400e-07,1.963402e-07,1.963404e-07,1.963405e-07,1.963407e-07,1.963408e-07,1.963410e-07,1.963412e-07,1.963413e-07,1.963415e-07,1.963416e-07,1.963418e-07,1.963420e-07,1.963421e-07,1.963423e-07,1.963424e-07,1.963426e-07,1.963428e-07,1.963429e-07,1.963431e-07,1.963432e-07,1.963434e-07,1.963435e-07,1.963437e-07,1.963439e-07,1.963440e-07,1.963442e-07,1.963443e-07,1.963445e-07,1.963447e-07,1.963448e-07,1.963450e-07,1.963451e-07,1.963453e-07,1.963455e-07,1.963456e-07,1.963458e-07,1.963459e-07,1.963461e-07,1.963463e-07,1.963464e-07,1.963466e-07,1.963467e-07,1.963469e-07,1.963471e-07,1.963472e-07,1.963474e-07,1.963475e-07,1.963477e-07,1.963479e-07,1.963480e-07,1.963482e-07,1.963483e-07,1.963485e-07,1.963487e-07,1.963488e-07,1.963490e-07,1.963491e-07,1.963493e-07,1.963495e-07,1.963496e-07,1.963498e-07,1.963499e-07,1.963501e-07,1.963503e-07,1.963504e-07,1.963506e-07,1.963507e-07,1.963509e-07,1.963510e-07,1.963512e-07,1.963514e-07,1.963515e-07,1.963517e-07,1.963518e-07,1.963520e-07,1.963522e-07,1.963523e-07,1.963525e-07,1.963526e-07,1.963528e-07,1.963530e-07,1.963531e-07,1.963533e-07,1.963534e-07,1.963536e-07,1.963538e-07,1.963539e-07,1.963541e-07,1.963542e-07,1.963544e-07,1.963546e-07,1.963547e-07,1.963549e-07,1.963550e-07,1.963552e-07,1.963554e-07,1.963555e-07,1.963557e-07,1.963558e-07,1.963560e-07,1.963562e-07,1.963563e-07,1.963565e-07,1.963566e-07,1.963568e-07,1.963569e-07,1.963571e-07,1.963573e-07,1.963574e-07,1.963576e-07,1.963577e-07,1.963579e-07,1.963581e-07,1.963582e-07,1.963584e-07,1.963585e-07,1.963587e-07,1.963589e-07,1.963590e-07,1.963592e-07,1.963593e-07,1.963595e-07,1.963597e-07,1.963598e-07,1.963600e-07,1.963601e-07,1.963603e-07,1.963605e-07,1.963606e-07,1.963608e-07,1.963609e-07,1.963611e-07,1.963613e-07,1.963614e-07,1.963616e-07,1.963617e-07,1.963619e-07,1.963620e-07,1.963622e-07,1.963624e-07,1.963625e-07,1.963627e-07,1.963628e-07,1.963630e-07,1.963632e-07,1.963633e-07,1.963635e-07,1.963636e-07,1.963638e-07,1.963640e-07,1.963641e-07,1.963643e-07,1.963644e-07,1.963646e-07,1.963648e-07,1.963649e-07,1.963651e-07,1.963652e-07,1.963654e-07,1.963656e-07,1.963657e-07,1.963659e-07,1.963660e-07,1.963662e-07,1.963664e-07,1.963665e-07,1.963667e-07,1.963668e-07,1.963670e-07,1.963671e-07,1.963673e-07,1.963675e-07,1.963676e-07,1.963678e-07,1.963679e-07,1.963681e-07,1.963683e-07,1.963684e-07,1.963686e-07,1.963687e-07,1.963689e-07,1.963691e-07,1.963692e-07,1.963694e-07,1.963695e-07,1.963697e-07,1.963699e-07,1.963700e-07,1.963702e-07,1.963703e-07,1.963705e-07,1.963707e-07,1.963708e-07,1.963710e-07,1.963711e-07,1.963713e-07,1.963714e-07,1.963716e-07,1.963718e-07,1.963719e-07,1.963721e-07,1.963722e-07,1.963724e-07,1.963726e-07,1.963727e-07,1.963729e-07,1.963730e-07,1.963732e-07,1.963734e-07,1.963735e-07,1.963737e-07,1.963738e-07,1.963740e-07,1.963742e-07,1.963743e-07,1.963745e-07,1.963746e-07,1.963748e-07,1.963750e-07,1.963751e-07,1.963753e-07,1.963754e-07,1.963756e-07,1.963757e-07,1.963759e-07,1.963761e-07,1.963762e-07,1.963764e-07,1.963765e-07,1.963767e-07,1.963769e-07,1.963770e-07,1.963772e-07,1.963773e-07,1.963775e-07,1.963777e-07,1.963778e-07,1.963780e-07,1.963781e-07,1.963783e-07,1.963785e-07,1.963786e-07,1.963788e-07,1.963789e-07,1.963791e-07,1.963792e-07,1.963794e-07,1.963796e-07,1.963797e-07,1.963799e-07,1.963800e-07,1.963802e-07,1.963804e-07,1.963805e-07,1.963807e-07,1.963808e-07,1.963810e-07,1.963812e-07,1.963813e-07,1.963815e-07,1.963816e-07,1.963818e-07,1.963820e-07,1.963821e-07,1.963823e-07,1.963824e-07,1.963826e-07,1.963827e-07,1.963829e-07,1.963831e-07,1.963832e-07,1.963834e-07,1.963835e-07,1.963837e-07,1.963839e-07,1.963840e-07,1.963842e-07,1.963843e-07,1.963845e-07,1.963847e-07,1.963848e-07,1.963850e-07,1.963851e-07,1.963853e-07,1.963855e-07,1.963856e-07,1.963858e-07,1.963859e-07,1.963861e-07,1.963862e-07,1.963864e-07,1.963866e-07,1.963867e-07,1.963869e-07,1.963870e-07,1.963872e-07,1.963874e-07,1.963875e-07,1.963877e-07,1.963878e-07,1.963880e-07,1.963882e-07,1.963883e-07,1.963885e-07,1.963886e-07,1.963888e-07,1.963890e-07,1.963891e-07,1.963893e-07,1.963894e-07,1.963896e-07,1.963897e-07,1.963899e-07,1.963901e-07,1.963902e-07,1.963904e-07,1.963905e-07,1.963907e-07,1.963909e-07,1.963910e-07,1.963912e-07,1.963913e-07,1.963915e-07,1.963917e-07,1.963918e-07,1.963920e-07,1.963921e-07,1.963923e-07,1.963925e-07,1.963926e-07,1.963928e-07,1.963929e-07,1.963931e-07,1.963932e-07,1.963934e-07,1.963936e-07,1.963937e-07,1.963939e-07,1.963940e-07,1.963942e-07,1.963944e-07,1.963945e-07,1.963947e-07,1.963948e-07,1.963950e-07,1.963952e-07,1.963953e-07,1.963955e-07,1.963956e-07,1.963958e-07,1.963959e-07,1.963961e-07,1.963963e-07,1.963964e-07,1.963966e-07,1.963967e-07,1.963969e-07,1.963971e-07,1.963972e-07,1.963974e-07,1.963975e-07,1.963977e-07,1.963979e-07,1.963980e-07,1.963982e-07,1.963983e-07,1.963985e-07,1.963986e-07,1.963988e-07,1.963990e-07,1.963991e-07,1.963993e-07,1.963994e-07,1.963996e-07,1.963998e-07,1.963999e-07,1.964001e-07,1.964002e-07,1.964004e-07,1.964006e-07,1.964007e-07,1.964009e-07,1.964010e-07,1.964012e-07,1.964013e-07,1.964015e-07,1.964017e-07,1.964018e-07,1.964020e-07,1.964021e-07,1.964023e-07,1.964025e-07,1.964026e-07,1.964028e-07,1.964029e-07,1.964031e-07,1.964033e-07,1.964034e-07,1.964036e-07,1.964037e-07,1.964039e-07,1.964040e-07,1.964042e-07,1.964044e-07,1.964045e-07,1.964047e-07,1.964048e-07,1.964050e-07,1.964052e-07,1.964053e-07,1.964055e-07,1.964056e-07,1.964058e-07,1.964060e-07,1.964061e-07,1.964063e-07,1.964064e-07,1.964066e-07,1.964067e-07,1.964069e-07,1.964071e-07,1.964072e-07,1.964074e-07,1.964075e-07,1.964077e-07,1.964079e-07,1.964080e-07,1.964082e-07,1.964083e-07,1.964085e-07,1.964087e-07,1.964088e-07,1.964090e-07,1.964091e-07,1.964093e-07,1.964094e-07,1.964096e-07,1.964098e-07,1.964099e-07,1.964101e-07,1.964102e-07,1.964104e-07,1.964106e-07,1.964107e-07,1.964109e-07,1.964110e-07,1.964112e-07,1.964114e-07,1.964115e-07,1.964117e-07,1.964118e-07,1.964120e-07,1.964121e-07,1.964123e-07,1.964125e-07,1.964126e-07,1.964128e-07,1.964129e-07,1.964131e-07,1.964133e-07,1.964134e-07,1.964136e-07,1.964137e-07,1.964139e-07,1.964140e-07,1.964142e-07,1.964144e-07,1.964145e-07,1.964147e-07,1.964148e-07,1.964150e-07,1.964152e-07,1.964153e-07,1.964155e-07,1.964156e-07,1.964158e-07,1.964160e-07,1.964161e-07,1.964163e-07,1.964164e-07,1.964166e-07,1.964167e-07,1.964169e-07,1.964171e-07,1.964172e-07,1.964174e-07,1.964175e-07,1.964177e-07,1.964179e-07,1.964180e-07,1.964182e-07,1.964183e-07,1.964185e-07,1.964186e-07,1.964188e-07,1.964190e-07,1.964191e-07,1.964193e-07,1.964194e-07,1.964196e-07,1.964198e-07,1.964199e-07,1.964201e-07,1.964202e-07,1.964204e-07,1.964206e-07,1.964207e-07,1.964209e-07,1.964210e-07,1.964212e-07,1.964213e-07,1.964215e-07,1.964217e-07,1.964218e-07,1.964220e-07,1.964221e-07,1.964223e-07,1.964225e-07,1.964226e-07,1.964228e-07,1.964229e-07,1.964231e-07,1.964232e-07,1.964234e-07,1.964236e-07,1.964237e-07,1.964239e-07,1.964240e-07,1.964242e-07,1.964244e-07,1.964245e-07,1.964247e-07,1.964248e-07,1.964250e-07,1.964251e-07,1.964253e-07,1.964255e-07,1.964256e-07,1.964258e-07,1.964259e-07,1.964261e-07,1.964263e-07,1.964264e-07,1.964266e-07,1.964267e-07,1.964269e-07,1.964271e-07,1.964272e-07,1.964274e-07,1.964275e-07,1.964277e-07,1.964278e-07,1.964280e-07,1.964282e-07,1.964283e-07,1.964285e-07,1.964286e-07,1.964288e-07,1.964290e-07,1.964291e-07,1.964293e-07,1.964294e-07,1.964296e-07,1.964297e-07,1.964299e-07,1.964301e-07,1.964302e-07,1.964304e-07,1.964305e-07,1.964307e-07,1.964309e-07,1.964310e-07,1.964312e-07,1.964313e-07,1.964315e-07,1.964316e-07,1.964318e-07,1.964320e-07,1.964321e-07,1.964323e-07,1.964324e-07,1.964326e-07,1.964328e-07,1.964329e-07,1.964331e-07,1.964332e-07,1.964334e-07,1.964335e-07,1.964337e-07,1.964339e-07,1.964340e-07,1.964342e-07,1.964343e-07,1.964345e-07,1.964347e-07,1.964348e-07,1.964350e-07,1.964351e-07,1.964353e-07,1.964354e-07,1.964356e-07,1.964358e-07,1.964359e-07,1.964361e-07,1.964362e-07,1.964364e-07,1.964366e-07,1.964367e-07,1.964369e-07,1.964370e-07,1.964372e-07,1.964373e-07,1.964375e-07,1.964377e-07,1.964378e-07,1.964380e-07,1.964381e-07,1.964383e-07,1.964385e-07,1.964386e-07,1.964388e-07,1.964389e-07,1.964391e-07,1.964392e-07,1.964394e-07,1.964396e-07,1.964397e-07,1.964399e-07,1.964400e-07,1.964402e-07,1.964404e-07,1.964405e-07,1.964407e-07,1.964408e-07,1.964410e-07,1.964411e-07,1.964413e-07,1.964415e-07,1.964416e-07,1.964418e-07,1.964419e-07,1.964421e-07,1.964423e-07,1.964424e-07,1.964426e-07,1.964427e-07,1.964429e-07,1.964430e-07,1.964432e-07,1.964434e-07,1.964435e-07,1.964437e-07,1.964438e-07,1.964440e-07,1.964442e-07,1.964443e-07,1.964445e-07,1.964446e-07,1.964448e-07,1.964449e-07,1.964451e-07,1.964453e-07,1.964454e-07,1.964456e-07,1.964457e-07,1.964459e-07,1.964461e-07,1.964462e-07,1.964464e-07,1.964465e-07,1.964467e-07,1.964468e-07,1.964470e-07,1.964472e-07,1.964473e-07,1.964475e-07,1.964476e-07,1.964478e-07,1.964480e-07,1.964481e-07,1.964483e-07,1.964484e-07,1.964486e-07,1.964487e-07,1.964489e-07,1.964491e-07,1.964492e-07,1.964494e-07,1.964495e-07,1.964497e-07,1.964499e-07,1.964500e-07,1.964502e-07,1.964503e-07,1.964505e-07,1.964506e-07,1.964508e-07,1.964510e-07,1.964511e-07,1.964513e-07,1.964514e-07,1.964516e-07,1.964518e-07,1.964519e-07,1.964521e-07,1.964522e-07,1.964524e-07,1.964525e-07,1.964527e-07,1.964529e-07,1.964530e-07,1.964532e-07,1.964533e-07,1.964535e-07,1.964536e-07,1.964538e-07,1.964540e-07,1.964541e-07,1.964543e-07,1.964544e-07,1.964546e-07,1.964548e-07,1.964549e-07,1.964551e-07,1.964552e-07,1.964554e-07,1.964555e-07,1.964557e-07,1.964559e-07,1.964560e-07,1.964562e-07,1.964563e-07,1.964565e-07,1.964567e-07,1.964568e-07,1.964570e-07,1.964571e-07,1.964573e-07,1.964574e-07,1.964576e-07,1.964578e-07,1.964579e-07,1.964581e-07,1.964582e-07,1.964584e-07,1.964585e-07,1.964587e-07,1.964589e-07,1.964590e-07,1.964592e-07,1.964593e-07,1.964595e-07,1.964597e-07,1.964598e-07,1.964600e-07,1.964601e-07,1.964603e-07,1.964604e-07,1.964606e-07,1.964608e-07,1.964609e-07,1.964611e-07,1.964612e-07,1.964614e-07,1.964616e-07,1.964617e-07,1.964619e-07,1.964620e-07,1.964622e-07,1.964623e-07,1.964625e-07,1.964627e-07,1.964628e-07,1.964630e-07,1.964631e-07,1.964633e-07,1.964634e-07,1.964636e-07,1.964638e-07,1.964639e-07,1.964641e-07,1.964642e-07,1.964644e-07,1.964646e-07,1.964647e-07,1.964649e-07,1.964650e-07,1.964652e-07,1.964653e-07,1.964655e-07,1.964657e-07,1.964658e-07,1.964660e-07,1.964661e-07,1.964663e-07,1.964664e-07,1.964666e-07,1.964668e-07,1.964669e-07,1.964671e-07,1.964672e-07,1.964674e-07,1.964676e-07,1.964677e-07,1.964679e-07,1.964680e-07,1.964682e-07,1.964683e-07,1.964685e-07,1.964687e-07,1.964688e-07,1.964690e-07,1.964691e-07,1.964693e-07,1.964695e-07,1.964696e-07,1.964698e-07,1.964699e-07,1.964701e-07,1.964702e-07,1.964704e-07,1.964706e-07,1.964707e-07,1.964709e-07,1.964710e-07,1.964712e-07,1.964713e-07,1.964715e-07,1.964717e-07,1.964718e-07,1.964720e-07,1.964721e-07,1.964723e-07,1.964725e-07,1.964726e-07,1.964728e-07,1.964729e-07,1.964731e-07,1.964732e-07,1.964734e-07,1.964736e-07,1.964737e-07,1.964739e-07,1.964740e-07,1.964742e-07,1.964743e-07,1.964745e-07,1.964747e-07,1.964748e-07,1.964750e-07,1.964751e-07,1.964753e-07,1.964754e-07,1.964756e-07,1.964758e-07,1.964759e-07,1.964761e-07,1.964762e-07,1.964764e-07,1.964766e-07,1.964767e-07,1.964769e-07,1.964770e-07,1.964772e-07,1.964773e-07,1.964775e-07,1.964777e-07,1.964778e-07,1.964780e-07,1.964781e-07,1.964783e-07,1.964784e-07,1.964786e-07,1.964788e-07,1.964789e-07,1.964791e-07,1.964792e-07,1.964794e-07,1.964796e-07,1.964797e-07,1.964799e-07,1.964800e-07,1.964802e-07,1.964803e-07,1.964805e-07,1.964807e-07,1.964808e-07,1.964810e-07,1.964811e-07,1.964813e-07,1.964814e-07,1.964816e-07,1.964818e-07,1.964819e-07,1.964821e-07,1.964822e-07,1.964824e-07,1.964825e-07,1.964827e-07,1.964829e-07,1.964830e-07,1.964832e-07,1.964833e-07,1.964835e-07,1.964837e-07,1.964838e-07,1.964840e-07,1.964841e-07,1.964843e-07,1.964844e-07,1.964846e-07,1.964848e-07,1.964849e-07,1.964851e-07,1.964852e-07,1.964854e-07,1.964855e-07,1.964857e-07,1.964859e-07,1.964860e-07,1.964862e-07,1.964863e-07,1.964865e-07,1.964867e-07,1.964868e-07,1.964870e-07,1.964871e-07,1.964873e-07,1.964874e-07,1.964876e-07,1.964878e-07,1.964879e-07,1.964881e-07,1.964882e-07,1.964884e-07,1.964885e-07,1.964887e-07,1.964889e-07,1.964890e-07,1.964892e-07,1.964893e-07,1.964895e-07,1.964896e-07,1.964898e-07,1.964900e-07,1.964901e-07,1.964903e-07,1.964904e-07,1.964906e-07,1.964907e-07,1.964909e-07,1.964911e-07,1.964912e-07,1.964914e-07,1.964915e-07,1.964917e-07,1.964919e-07,1.964920e-07,1.964922e-07,1.964923e-07,1.964925e-07,1.964926e-07,1.964928e-07,1.964930e-07,1.964931e-07,1.964933e-07,1.964934e-07,1.964936e-07,1.964937e-07,1.964939e-07,1.964941e-07,1.964942e-07,1.964944e-07,1.964945e-07,1.964947e-07,1.964948e-07,1.964950e-07,1.964952e-07,1.964953e-07,1.964955e-07,1.964956e-07,1.964958e-07,1.964960e-07,1.964961e-07,1.964963e-07,1.964964e-07,1.964966e-07,1.964967e-07,1.964969e-07,1.964971e-07,1.964972e-07,1.964974e-07,1.964975e-07,1.964977e-07,1.964978e-07,1.964980e-07,1.964982e-07,1.964983e-07,1.964985e-07,1.964986e-07,1.964988e-07,1.964989e-07,1.964991e-07,1.964993e-07,1.964994e-07,1.964996e-07,1.964997e-07,1.964999e-07,1.965000e-07,1.965002e-07,1.965004e-07,1.965005e-07,1.965007e-07,1.965008e-07,1.965010e-07,1.965011e-07,1.965013e-07,1.965015e-07,1.965016e-07,1.965018e-07,1.965019e-07,1.965021e-07,1.965023e-07,1.965024e-07,1.965026e-07,1.965027e-07,1.965029e-07,1.965030e-07,1.965032e-07,1.965034e-07,1.965035e-07,1.965037e-07,1.965038e-07,1.965040e-07,1.965041e-07,1.965043e-07,1.965045e-07,1.965046e-07,1.965048e-07,1.965049e-07,1.965051e-07,1.965052e-07,1.965054e-07,1.965056e-07,1.965057e-07,1.965059e-07,1.965060e-07,1.965062e-07,1.965063e-07,1.965065e-07,1.965067e-07,1.965068e-07,1.965070e-07,1.965071e-07,1.965073e-07,1.965074e-07,1.965076e-07,1.965078e-07,1.965079e-07,1.965081e-07,1.965082e-07,1.965084e-07,1.965085e-07,1.965087e-07,1.965089e-07,1.965090e-07,1.965092e-07,1.965093e-07,1.965095e-07,1.965096e-07,1.965098e-07,1.965100e-07,1.965101e-07,1.965103e-07,1.965104e-07,1.965106e-07,1.965108e-07,1.965109e-07,1.965111e-07,1.965112e-07,1.965114e-07,1.965115e-07,1.965117e-07,1.965119e-07,1.965120e-07,1.965122e-07,1.965123e-07,1.965125e-07,1.965126e-07,1.965128e-07,1.965130e-07,1.965131e-07,1.965133e-07,1.965134e-07,1.965136e-07,1.965137e-07,1.965139e-07,1.965141e-07,1.965142e-07,1.965144e-07,1.965145e-07,1.965147e-07,1.965148e-07,1.965150e-07,1.965152e-07,1.965153e-07,1.965155e-07,1.965156e-07,1.965158e-07,1.965159e-07,1.965161e-07,1.965163e-07,1.965164e-07,1.965166e-07,1.965167e-07,1.965169e-07,1.965170e-07,1.965172e-07,1.965174e-07,1.965175e-07,1.965177e-07,1.965178e-07,1.965180e-07,1.965181e-07,1.965183e-07,1.965185e-07,1.965186e-07,1.965188e-07,1.965189e-07,1.965191e-07,1.965192e-07,1.965194e-07,1.965196e-07,1.965197e-07,1.965199e-07,1.965200e-07,1.965202e-07,1.965203e-07,1.965205e-07,1.965207e-07,1.965208e-07,1.965210e-07,1.965211e-07,1.965213e-07,1.965214e-07,1.965216e-07,1.965218e-07,1.965219e-07,1.965221e-07,1.965222e-07,1.965224e-07,1.965225e-07,1.965227e-07,1.965229e-07,1.965230e-07,1.965232e-07,1.965233e-07,1.965235e-07,1.965236e-07,1.965238e-07,1.965240e-07,1.965241e-07,1.965243e-07,1.965244e-07,1.965246e-07,1.965247e-07,1.965249e-07,1.965251e-07,1.965252e-07,1.965254e-07,1.965255e-07,1.965257e-07,1.965258e-07,1.965260e-07,1.965262e-07,1.965263e-07,1.965265e-07,1.965266e-07,1.965268e-07,1.965269e-07,1.965271e-07,1.965273e-07,1.965274e-07,1.965276e-07,1.965277e-07,1.965279e-07,1.965280e-07,1.965282e-07,1.965284e-07,1.965285e-07,1.965287e-07,1.965288e-07,1.965290e-07,1.965291e-07,1.965293e-07,1.965295e-07,1.965296e-07,1.965298e-07,1.965299e-07,1.965301e-07,1.965302e-07,1.965304e-07,1.965306e-07,1.965307e-07,1.965309e-07,1.965310e-07,1.965312e-07,1.965313e-07,1.965315e-07,1.965317e-07,1.965318e-07,1.965320e-07,1.965321e-07,1.965323e-07,1.965324e-07,1.965326e-07,1.965328e-07,1.965329e-07,1.965331e-07,1.965332e-07,1.965334e-07,1.965335e-07,1.965337e-07,1.965339e-07,1.965340e-07,1.965342e-07,1.965343e-07,1.965345e-07,1.965346e-07,1.965348e-07,1.965350e-07,1.965351e-07,1.965353e-07,1.965354e-07,1.965356e-07,1.965357e-07,1.965359e-07,1.965361e-07,1.965362e-07,1.965364e-07,1.965365e-07,1.965367e-07,1.965368e-07,1.965370e-07,1.965372e-07,1.965373e-07,1.965375e-07,1.965376e-07,1.965378e-07,1.965379e-07,1.965381e-07,1.965383e-07,1.965384e-07,1.965386e-07,1.965387e-07,1.965389e-07,1.965390e-07,1.965392e-07,1.965394e-07,1.965395e-07,1.965397e-07,1.965398e-07,1.965400e-07,1.965401e-07,1.965403e-07,1.965405e-07,1.965406e-07,1.965408e-07,1.965409e-07,1.965411e-07,1.965412e-07,1.965414e-07,1.965416e-07,1.965417e-07,1.965419e-07,1.965420e-07,1.965422e-07,1.965423e-07,1.965425e-07,1.965427e-07,1.965428e-07,1.965430e-07,1.965431e-07,1.965433e-07,1.965434e-07,1.965436e-07,1.965438e-07,1.965439e-07,1.965441e-07,1.965442e-07,1.965444e-07,1.965445e-07,1.965447e-07,1.965448e-07,1.965450e-07,1.965452e-07,1.965453e-07,1.965455e-07,1.965456e-07,1.965458e-07,1.965459e-07,1.965461e-07,1.965463e-07,1.965464e-07,1.965466e-07,1.965467e-07,1.965469e-07,1.965470e-07,1.965472e-07,1.965474e-07,1.965475e-07,1.965477e-07,1.965478e-07,1.965480e-07,1.965481e-07,1.965483e-07,1.965485e-07,1.965486e-07,1.965488e-07,1.965489e-07,1.965491e-07,1.965492e-07,1.965494e-07,1.965496e-07,1.965497e-07,1.965499e-07,1.965500e-07,1.965502e-07,1.965503e-07,1.965505e-07,1.965507e-07,1.965508e-07,1.965510e-07,1.965511e-07,1.965513e-07,1.965514e-07,1.965516e-07,1.965518e-07,1.965519e-07,1.965521e-07,1.965522e-07,1.965524e-07,1.965525e-07,1.965527e-07,1.965528e-07,1.965530e-07,1.965532e-07,1.965533e-07,1.965535e-07,1.965536e-07,1.965538e-07,1.965539e-07,1.965541e-07,1.965543e-07,1.965544e-07,1.965546e-07,1.965547e-07,1.965549e-07,1.965550e-07,1.965552e-07,1.965554e-07,1.965555e-07,1.965557e-07,1.965558e-07,1.965560e-07,1.965561e-07,1.965563e-07,1.965565e-07,1.965566e-07,1.965568e-07,1.965569e-07,1.965571e-07,1.965572e-07,1.965574e-07,1.965576e-07,1.965577e-07,1.965579e-07,1.965580e-07,1.965582e-07,1.965583e-07,1.965585e-07,1.965586e-07,1.965588e-07,1.965590e-07,1.965591e-07,1.965593e-07,1.965594e-07,1.965596e-07,1.965597e-07,1.965599e-07,1.965601e-07,1.965602e-07,1.965604e-07,1.965605e-07,1.965607e-07,1.965608e-07,1.965610e-07,1.965612e-07,1.965613e-07,1.965615e-07,1.965616e-07,1.965618e-07,1.965619e-07,1.965621e-07,1.965623e-07,1.965624e-07,1.965626e-07,1.965627e-07,1.965629e-07,1.965630e-07,1.965632e-07,1.965633e-07,1.965635e-07,1.965637e-07,1.965638e-07,1.965640e-07,1.965641e-07,1.965643e-07,1.965644e-07,1.965646e-07,1.965648e-07,1.965649e-07,1.965651e-07,1.965652e-07,1.965654e-07,1.965655e-07,1.965657e-07,1.965659e-07,1.965660e-07,1.965662e-07,1.965663e-07,1.965665e-07,1.965666e-07,1.965668e-07,1.965670e-07,1.965671e-07,1.965673e-07,1.965674e-07,1.965676e-07,1.965677e-07,1.965679e-07,1.965680e-07,1.965682e-07,1.965684e-07,1.965685e-07,1.965687e-07,1.965688e-07,1.965690e-07,1.965691e-07,1.965693e-07,1.965695e-07,1.965696e-07,1.965698e-07,1.965699e-07,1.965701e-07,1.965702e-07,1.965704e-07,1.965706e-07,1.965707e-07,1.965709e-07,1.965710e-07,1.965712e-07,1.965713e-07,1.965715e-07,1.965716e-07,1.965718e-07,1.965720e-07,1.965721e-07,1.965723e-07,1.965724e-07,1.965726e-07,1.965727e-07,1.965729e-07,1.965731e-07,1.965732e-07,1.965734e-07,1.965735e-07,1.965737e-07,1.965738e-07,1.965740e-07,1.965742e-07,1.965743e-07,1.965745e-07,1.965746e-07,1.965748e-07,1.965749e-07,1.965751e-07,1.965752e-07,1.965754e-07,1.965756e-07,1.965757e-07,1.965759e-07,1.965760e-07,1.965762e-07,1.965763e-07,1.965765e-07,1.965767e-07,1.965768e-07,1.965770e-07,1.965771e-07,1.965773e-07,1.965774e-07,1.965776e-07,1.965778e-07,1.965779e-07,1.965781e-07,1.965782e-07,1.965784e-07,1.965785e-07,1.965787e-07,1.965788e-07,1.965790e-07,1.965792e-07,1.965793e-07,1.965795e-07,1.965796e-07,1.965798e-07,1.965799e-07,1.965801e-07,1.965803e-07,1.965804e-07,1.965806e-07,1.965807e-07,1.965809e-07,1.965810e-07,1.965812e-07,1.965814e-07,1.965815e-07,1.965817e-07,1.965818e-07,1.965820e-07,1.965821e-07,1.965823e-07,1.965824e-07,1.965826e-07,1.965828e-07,1.965829e-07,1.965831e-07,1.965832e-07,1.965834e-07,1.965835e-07,1.965837e-07,1.965839e-07,1.965840e-07,1.965842e-07,1.965843e-07,1.965845e-07,1.965846e-07,1.965848e-07,1.965849e-07,1.965851e-07,1.965853e-07,1.965854e-07,1.965856e-07,1.965857e-07,1.965859e-07,1.965860e-07,1.965862e-07,1.965864e-07,1.965865e-07,1.965867e-07,1.965868e-07,1.965870e-07,1.965871e-07,1.965873e-07,1.965874e-07,1.965876e-07,1.965878e-07,1.965879e-07,1.965881e-07,1.965882e-07,1.965884e-07,1.965885e-07,1.965887e-07,1.965889e-07,1.965890e-07,1.965892e-07,1.965893e-07,1.965895e-07,1.965896e-07,1.965898e-07,1.965900e-07,1.965901e-07,1.965903e-07,1.965904e-07,1.965906e-07,1.965907e-07,1.965909e-07,1.965910e-07,1.965912e-07,1.965914e-07,1.965915e-07,1.965917e-07,1.965918e-07,1.965920e-07,1.965921e-07,1.965923e-07,1.965925e-07,1.965926e-07,1.965928e-07,1.965929e-07,1.965931e-07,1.965932e-07,1.965934e-07,1.965935e-07,1.965937e-07,1.965939e-07,1.965940e-07,1.965942e-07,1.965943e-07,1.965945e-07,1.965946e-07,1.965948e-07,1.965950e-07,1.965951e-07,1.965953e-07,1.965954e-07,1.965956e-07,1.965957e-07,1.965959e-07,1.965960e-07,1.965962e-07,1.965964e-07,1.965965e-07,1.965967e-07,1.965968e-07,1.965970e-07,1.965971e-07,1.965973e-07,1.965975e-07,1.965976e-07,1.965978e-07,1.965979e-07,1.965981e-07,1.965982e-07,1.965984e-07,1.965985e-07,1.965987e-07,1.965989e-07,1.965990e-07,1.965992e-07,1.965993e-07,1.965995e-07,1.965996e-07,1.965998e-07,1.965999e-07,1.966001e-07,1.966003e-07,1.966004e-07,1.966006e-07,1.966007e-07,1.966009e-07,1.966010e-07,1.966012e-07,1.966014e-07,1.966015e-07,1.966017e-07,1.966018e-07,1.966020e-07,1.966021e-07,1.966023e-07,1.966024e-07,1.966026e-07,1.966028e-07,1.966029e-07,1.966031e-07,1.966032e-07,1.966034e-07,1.966035e-07,1.966037e-07,1.966039e-07,1.966040e-07,1.966042e-07,1.966043e-07,1.966045e-07,1.966046e-07,1.966048e-07,1.966049e-07,1.966051e-07,1.966053e-07,1.966054e-07,1.966056e-07,1.966057e-07,1.966059e-07,1.966060e-07,1.966062e-07,1.966064e-07,1.966065e-07,1.966067e-07,1.966068e-07,1.966070e-07,1.966071e-07,1.966073e-07,1.966074e-07,1.966076e-07,1.966078e-07,1.966079e-07,1.966081e-07,1.966082e-07,1.966084e-07,1.966085e-07,1.966087e-07,1.966088e-07,1.966090e-07,1.966092e-07,1.966093e-07,1.966095e-07,1.966096e-07,1.966098e-07,1.966099e-07,1.966101e-07,1.966103e-07,1.966104e-07,1.966106e-07,1.966107e-07,1.966109e-07,1.966110e-07,1.966112e-07,1.966113e-07,1.966115e-07,1.966117e-07,1.966118e-07,1.966120e-07,1.966121e-07,1.966123e-07,1.966124e-07,1.966126e-07,1.966127e-07,1.966129e-07,1.966131e-07,1.966132e-07,1.966134e-07,1.966135e-07,1.966137e-07,1.966138e-07,1.966140e-07,1.966142e-07,1.966143e-07,1.966145e-07,1.966146e-07,1.966148e-07,1.966149e-07,1.966151e-07,1.966152e-07,1.966154e-07,1.966156e-07,1.966157e-07,1.966159e-07,1.966160e-07,1.966162e-07,1.966163e-07,1.966165e-07,1.966166e-07,1.966168e-07,1.966170e-07,1.966171e-07,1.966173e-07,1.966174e-07,1.966176e-07,1.966177e-07,1.966179e-07,1.966181e-07,1.966182e-07,1.966184e-07,1.966185e-07,1.966187e-07,1.966188e-07,1.966190e-07,1.966191e-07,1.966193e-07,1.966195e-07,1.966196e-07,1.966198e-07,1.966199e-07,1.966201e-07,1.966202e-07,1.966204e-07,1.966205e-07,1.966207e-07,1.966209e-07,1.966210e-07,1.966212e-07,1.966213e-07,1.966215e-07,1.966216e-07,1.966218e-07,1.966219e-07,1.966221e-07,1.966223e-07,1.966224e-07,1.966226e-07,1.966227e-07,1.966229e-07,1.966230e-07,1.966232e-07,1.966234e-07,1.966235e-07,1.966237e-07,1.966238e-07,1.966240e-07,1.966241e-07,1.966243e-07,1.966244e-07,1.966246e-07,1.966248e-07,1.966249e-07,1.966251e-07,1.966252e-07,1.966254e-07,1.966255e-07,1.966257e-07,1.966258e-07,1.966260e-07,1.966262e-07,1.966263e-07,1.966265e-07,1.966266e-07,1.966268e-07,1.966269e-07,1.966271e-07,1.966272e-07,1.966274e-07,1.966276e-07,1.966277e-07,1.966279e-07,1.966280e-07,1.966282e-07,1.966283e-07,1.966285e-07,1.966286e-07,1.966288e-07,1.966290e-07,1.966291e-07,1.966293e-07,1.966294e-07,1.966296e-07,1.966297e-07,1.966299e-07,1.966301e-07,1.966302e-07,1.966304e-07,1.966305e-07,1.966307e-07,1.966308e-07,1.966310e-07,1.966311e-07,1.966313e-07,1.966315e-07,1.966316e-07,1.966318e-07,1.966319e-07,1.966321e-07,1.966322e-07,1.966324e-07,1.966325e-07,1.966327e-07,1.966329e-07,1.966330e-07,1.966332e-07,1.966333e-07,1.966335e-07,1.966336e-07,1.966338e-07,1.966339e-07,1.966341e-07,1.966343e-07,1.966344e-07,1.966346e-07,1.966347e-07,1.966349e-07,1.966350e-07,1.966352e-07,1.966353e-07,1.966355e-07,1.966357e-07,1.966358e-07,1.966360e-07,1.966361e-07,1.966363e-07,1.966364e-07,1.966366e-07,1.966367e-07,1.966369e-07,1.966371e-07,1.966372e-07,1.966374e-07,1.966375e-07,1.966377e-07,1.966378e-07,1.966380e-07,1.966381e-07,1.966383e-07,1.966385e-07,1.966386e-07,1.966388e-07,1.966389e-07,1.966391e-07,1.966392e-07,1.966394e-07,1.966395e-07,1.966397e-07,1.966399e-07,1.966400e-07,1.966402e-07,1.966403e-07,1.966405e-07,1.966406e-07,1.966408e-07,1.966409e-07,1.966411e-07,1.966413e-07,1.966414e-07,1.966416e-07,1.966417e-07,1.966419e-07,1.966420e-07,1.966422e-07,1.966423e-07,1.966425e-07,1.966427e-07,1.966428e-07,1.966430e-07,1.966431e-07,1.966433e-07,1.966434e-07,1.966436e-07,1.966438e-07,1.966439e-07,1.966441e-07,1.966442e-07,1.966444e-07,1.966445e-07,1.966447e-07,1.966448e-07,1.966450e-07,1.966452e-07,1.966453e-07,1.966455e-07,1.966456e-07,1.966458e-07,1.966459e-07,1.966461e-07,1.966462e-07,1.966464e-07,1.966466e-07,1.966467e-07,1.966469e-07,1.966470e-07,1.966472e-07,1.966473e-07,1.966475e-07,1.966476e-07,1.966478e-07,1.966480e-07,1.966481e-07,1.966483e-07,1.966484e-07,1.966486e-07,1.966487e-07,1.966489e-07,1.966490e-07,1.966492e-07,1.966493e-07,1.966495e-07,1.966497e-07,1.966498e-07,1.966500e-07,1.966501e-07,1.966503e-07,1.966504e-07,1.966506e-07,1.966507e-07,1.966509e-07,1.966511e-07,1.966512e-07,1.966514e-07,1.966515e-07,1.966517e-07,1.966518e-07,1.966520e-07,1.966521e-07,1.966523e-07,1.966525e-07,1.966526e-07,1.966528e-07,1.966529e-07,1.966531e-07,1.966532e-07,1.966534e-07,1.966535e-07,1.966537e-07,1.966539e-07,1.966540e-07,1.966542e-07,1.966543e-07,1.966545e-07,1.966546e-07,1.966548e-07,1.966549e-07,1.966551e-07,1.966553e-07,1.966554e-07,1.966556e-07,1.966557e-07,1.966559e-07,1.966560e-07,1.966562e-07,1.966563e-07,1.966565e-07,1.966567e-07,1.966568e-07,1.966570e-07,1.966571e-07,1.966573e-07,1.966574e-07,1.966576e-07,1.966577e-07,1.966579e-07,1.966581e-07,1.966582e-07,1.966584e-07,1.966585e-07,1.966587e-07,1.966588e-07,1.966590e-07,1.966591e-07,1.966593e-07,1.966595e-07,1.966596e-07,1.966598e-07,1.966599e-07,1.966601e-07,1.966602e-07,1.966604e-07,1.966605e-07,1.966607e-07,1.966609e-07,1.966610e-07,1.966612e-07,1.966613e-07,1.966615e-07,1.966616e-07,1.966618e-07,1.966619e-07,1.966621e-07,1.966622e-07,1.966624e-07,1.966626e-07,1.966627e-07,1.966629e-07,1.966630e-07,1.966632e-07,1.966633e-07,1.966635e-07,1.966636e-07,1.966638e-07,1.966640e-07,1.966641e-07,1.966643e-07,1.966644e-07,1.966646e-07,1.966647e-07,1.966649e-07,1.966650e-07,1.966652e-07,1.966654e-07,1.966655e-07,1.966657e-07,1.966658e-07,1.966660e-07,1.966661e-07,1.966663e-07,1.966664e-07,1.966666e-07,1.966668e-07,1.966669e-07,1.966671e-07,1.966672e-07,1.966674e-07,1.966675e-07,1.966677e-07,1.966678e-07,1.966680e-07,1.966682e-07,1.966683e-07,1.966685e-07,1.966686e-07,1.966688e-07,1.966689e-07,1.966691e-07,1.966692e-07,1.966694e-07,1.966695e-07,1.966697e-07,1.966699e-07,1.966700e-07,1.966702e-07,1.966703e-07,1.966705e-07,1.966706e-07,1.966708e-07,1.966709e-07,1.966711e-07,1.966713e-07,1.966714e-07,1.966716e-07,1.966717e-07,1.966719e-07,1.966720e-07,1.966722e-07,1.966723e-07,1.966725e-07,1.966727e-07,1.966728e-07,1.966730e-07,1.966731e-07,1.966733e-07,1.966734e-07,1.966736e-07,1.966737e-07,1.966739e-07,1.966740e-07,1.966742e-07,1.966744e-07,1.966745e-07,1.966747e-07,1.966748e-07,1.966750e-07,1.966751e-07,1.966753e-07,1.966754e-07,1.966756e-07,1.966758e-07,1.966759e-07,1.966761e-07,1.966762e-07,1.966764e-07,1.966765e-07,1.966767e-07,1.966768e-07,1.966770e-07,1.966772e-07,1.966773e-07,1.966775e-07,1.966776e-07,1.966778e-07,1.966779e-07,1.966781e-07,1.966782e-07,1.966784e-07,1.966785e-07,1.966787e-07,1.966789e-07,1.966790e-07,1.966792e-07,1.966793e-07,1.966795e-07,1.966796e-07,1.966798e-07,1.966799e-07,1.966801e-07,1.966803e-07,1.966804e-07,1.966806e-07,1.966807e-07,1.966809e-07,1.966810e-07,1.966812e-07,1.966813e-07,1.966815e-07,1.966817e-07,1.966818e-07,1.966820e-07,1.966821e-07,1.966823e-07,1.966824e-07,1.966826e-07,1.966827e-07,1.966829e-07,1.966830e-07,1.966832e-07,1.966834e-07,1.966835e-07,1.966837e-07,1.966838e-07,1.966840e-07,1.966841e-07,1.966843e-07,1.966844e-07,1.966846e-07,1.966848e-07,1.966849e-07,1.966851e-07,1.966852e-07,1.966854e-07,1.966855e-07,1.966857e-07,1.966858e-07,1.966860e-07,1.966861e-07,1.966863e-07,1.966865e-07,1.966866e-07,1.966868e-07,1.966869e-07,1.966871e-07,1.966872e-07,1.966874e-07,1.966875e-07,1.966877e-07,1.966879e-07,1.966880e-07,1.966882e-07,1.966883e-07,1.966885e-07,1.966886e-07,1.966888e-07,1.966889e-07,1.966891e-07,1.966892e-07,1.966894e-07,1.966896e-07,1.966897e-07,1.966899e-07,1.966900e-07,1.966902e-07,1.966903e-07,1.966905e-07,1.966906e-07,1.966908e-07,1.966910e-07,1.966911e-07,1.966913e-07,1.966914e-07,1.966916e-07,1.966917e-07,1.966919e-07,1.966920e-07,1.966922e-07,1.966923e-07,1.966925e-07,1.966927e-07,1.966928e-07,1.966930e-07,1.966931e-07,1.966933e-07,1.966934e-07,1.966936e-07,1.966937e-07,1.966939e-07,1.966941e-07,1.966942e-07,1.966944e-07,1.966945e-07,1.966947e-07,1.966948e-07,1.966950e-07,1.966951e-07,1.966953e-07,1.966954e-07,1.966956e-07,1.966958e-07,1.966959e-07,1.966961e-07,1.966962e-07,1.966964e-07,1.966965e-07,1.966967e-07,1.966968e-07,1.966970e-07,1.966971e-07,1.966973e-07,1.966975e-07,1.966976e-07,1.966978e-07,1.966979e-07,1.966981e-07,1.966982e-07,1.966984e-07,1.966985e-07,1.966987e-07,1.966989e-07,1.966990e-07,1.966992e-07,1.966993e-07,1.966995e-07,1.966996e-07,1.966998e-07,1.966999e-07,1.967001e-07,1.967002e-07,1.967004e-07,1.967006e-07,1.967007e-07,1.967009e-07,1.967010e-07,1.967012e-07,1.967013e-07,1.967015e-07,1.967016e-07,1.967018e-07,1.967019e-07,1.967021e-07,1.967023e-07,1.967024e-07,1.967026e-07,1.967027e-07,1.967029e-07,1.967030e-07,1.967032e-07,1.967033e-07,1.967035e-07,1.967037e-07,1.967038e-07,1.967040e-07,1.967041e-07,1.967043e-07,1.967044e-07,1.967046e-07,1.967047e-07,1.967049e-07,1.967050e-07,1.967052e-07,1.967054e-07,1.967055e-07,1.967057e-07,1.967058e-07,1.967060e-07,1.967061e-07,1.967063e-07,1.967064e-07,1.967066e-07,1.967067e-07,1.967069e-07,1.967071e-07,1.967072e-07,1.967074e-07,1.967075e-07,1.967077e-07,1.967078e-07,1.967080e-07,1.967081e-07,1.967083e-07,1.967084e-07,1.967086e-07,1.967088e-07,1.967089e-07,1.967091e-07,1.967092e-07,1.967094e-07,1.967095e-07,1.967097e-07,1.967098e-07,1.967100e-07,1.967102e-07,1.967103e-07,1.967105e-07,1.967106e-07,1.967108e-07,1.967109e-07,1.967111e-07,1.967112e-07,1.967114e-07,1.967115e-07,1.967117e-07,1.967119e-07,1.967120e-07,1.967122e-07,1.967123e-07,1.967125e-07,1.967126e-07,1.967128e-07,1.967129e-07,1.967131e-07,1.967132e-07,1.967134e-07,1.967136e-07,1.967137e-07,1.967139e-07,1.967140e-07,1.967142e-07,1.967143e-07,1.967145e-07,1.967146e-07,1.967148e-07,1.967149e-07,1.967151e-07,1.967153e-07,1.967154e-07,1.967156e-07,1.967157e-07,1.967159e-07,1.967160e-07,1.967162e-07,1.967163e-07,1.967165e-07,1.967166e-07,1.967168e-07,1.967170e-07,1.967171e-07,1.967173e-07,1.967174e-07,1.967176e-07,1.967177e-07,1.967179e-07,1.967180e-07,1.967182e-07,1.967183e-07,1.967185e-07,1.967187e-07,1.967188e-07,1.967190e-07,1.967191e-07,1.967193e-07,1.967194e-07,1.967196e-07,1.967197e-07,1.967199e-07,1.967200e-07,1.967202e-07,1.967204e-07,1.967205e-07,1.967207e-07,1.967208e-07,1.967210e-07,1.967211e-07,1.967213e-07,1.967214e-07,1.967216e-07,1.967217e-07,1.967219e-07,1.967221e-07,1.967222e-07,1.967224e-07,1.967225e-07,1.967227e-07,1.967228e-07,1.967230e-07,1.967231e-07,1.967233e-07,1.967234e-07,1.967236e-07,1.967238e-07,1.967239e-07,1.967241e-07,1.967242e-07,1.967244e-07,1.967245e-07,1.967247e-07,1.967248e-07,1.967250e-07,1.967251e-07,1.967253e-07,1.967255e-07,1.967256e-07,1.967258e-07,1.967259e-07,1.967261e-07,1.967262e-07,1.967264e-07,1.967265e-07,1.967267e-07,1.967268e-07,1.967270e-07,1.967272e-07,1.967273e-07,1.967275e-07,1.967276e-07,1.967278e-07,1.967279e-07,1.967281e-07,1.967282e-07,1.967284e-07,1.967285e-07,1.967287e-07,1.967289e-07,1.967290e-07,1.967292e-07,1.967293e-07,1.967295e-07,1.967296e-07,1.967298e-07,1.967299e-07,1.967301e-07,1.967302e-07,1.967304e-07,1.967306e-07,1.967307e-07,1.967309e-07,1.967310e-07,1.967312e-07,1.967313e-07,1.967315e-07,1.967316e-07,1.967318e-07,1.967319e-07,1.967321e-07,1.967323e-07,1.967324e-07,1.967326e-07,1.967327e-07,1.967329e-07,1.967330e-07,1.967332e-07,1.967333e-07,1.967335e-07,1.967336e-07,1.967338e-07,1.967340e-07,1.967341e-07,1.967343e-07,1.967344e-07,1.967346e-07,1.967347e-07,1.967349e-07,1.967350e-07,1.967352e-07,1.967353e-07,1.967355e-07,1.967356e-07,1.967358e-07,1.967360e-07,1.967361e-07,1.967363e-07,1.967364e-07,1.967366e-07,1.967367e-07,1.967369e-07,1.967370e-07,1.967372e-07,1.967373e-07,1.967375e-07,1.967377e-07,1.967378e-07,1.967380e-07,1.967381e-07,1.967383e-07,1.967384e-07,1.967386e-07,1.967387e-07,1.967389e-07,1.967390e-07,1.967392e-07,1.967394e-07,1.967395e-07,1.967397e-07,1.967398e-07,1.967400e-07,1.967401e-07,1.967403e-07,1.967404e-07,1.967406e-07,1.967407e-07,1.967409e-07,1.967411e-07,1.967412e-07,1.967414e-07,1.967415e-07,1.967417e-07,1.967418e-07,1.967420e-07,1.967421e-07,1.967423e-07,1.967424e-07,1.967426e-07,1.967427e-07,1.967429e-07,1.967431e-07,1.967432e-07,1.967434e-07,1.967435e-07,1.967437e-07,1.967438e-07,1.967440e-07,1.967441e-07,1.967443e-07,1.967444e-07,1.967446e-07,1.967448e-07,1.967449e-07,1.967451e-07,1.967452e-07,1.967454e-07,1.967455e-07,1.967457e-07,1.967458e-07,1.967460e-07,1.967461e-07,1.967463e-07,1.967465e-07,1.967466e-07,1.967468e-07,1.967469e-07,1.967471e-07,1.967472e-07,1.967474e-07,1.967475e-07,1.967477e-07,1.967478e-07,1.967480e-07,1.967481e-07,1.967483e-07,1.967485e-07,1.967486e-07,1.967488e-07,1.967489e-07,1.967491e-07,1.967492e-07,1.967494e-07,1.967495e-07,1.967497e-07,1.967498e-07,1.967500e-07,1.967502e-07,1.967503e-07,1.967505e-07,1.967506e-07,1.967508e-07,1.967509e-07,1.967511e-07,1.967512e-07,1.967514e-07,1.967515e-07,1.967517e-07,1.967518e-07,1.967520e-07,1.967522e-07,1.967523e-07,1.967525e-07,1.967526e-07,1.967528e-07,1.967529e-07,1.967531e-07,1.967532e-07,1.967534e-07,1.967535e-07,1.967537e-07,1.967539e-07,1.967540e-07,1.967542e-07,1.967543e-07,1.967545e-07,1.967546e-07,1.967548e-07,1.967549e-07,1.967551e-07,1.967552e-07,1.967554e-07,1.967555e-07,1.967557e-07,1.967559e-07,1.967560e-07,1.967562e-07,1.967563e-07,1.967565e-07,1.967566e-07,1.967568e-07,1.967569e-07,1.967571e-07,1.967572e-07,1.967574e-07,1.967575e-07,1.967577e-07,1.967579e-07,1.967580e-07,1.967582e-07,1.967583e-07,1.967585e-07,1.967586e-07,1.967588e-07,1.967589e-07,1.967591e-07,1.967592e-07,1.967594e-07,1.967596e-07,1.967597e-07,1.967599e-07,1.967600e-07,1.967602e-07,1.967603e-07,1.967605e-07,1.967606e-07,1.967608e-07,1.967609e-07,1.967611e-07,1.967612e-07,1.967614e-07,1.967616e-07,1.967617e-07,1.967619e-07,1.967620e-07,1.967622e-07,1.967623e-07,1.967625e-07,1.967626e-07,1.967628e-07,1.967629e-07,1.967631e-07,1.967632e-07,1.967634e-07,1.967636e-07,1.967637e-07,1.967639e-07,1.967640e-07,1.967642e-07,1.967643e-07,1.967645e-07,1.967646e-07,1.967648e-07,1.967649e-07,1.967651e-07,1.967653e-07,1.967654e-07,1.967656e-07,1.967657e-07,1.967659e-07,1.967660e-07,1.967662e-07,1.967663e-07,1.967665e-07,1.967666e-07,1.967668e-07,1.967669e-07,1.967671e-07,1.967673e-07,1.967674e-07,1.967676e-07,1.967677e-07,1.967679e-07,1.967680e-07,1.967682e-07,1.967683e-07,1.967685e-07,1.967686e-07,1.967688e-07,1.967689e-07,1.967691e-07,1.967693e-07,1.967694e-07,1.967696e-07,1.967697e-07,1.967699e-07,1.967700e-07,1.967702e-07,1.967703e-07,1.967705e-07,1.967706e-07,1.967708e-07,1.967709e-07,1.967711e-07,1.967713e-07,1.967714e-07,1.967716e-07,1.967717e-07,1.967719e-07,1.967720e-07,1.967722e-07,1.967723e-07,1.967725e-07,1.967726e-07,1.967728e-07,1.967729e-07,1.967731e-07,1.967733e-07,1.967734e-07,1.967736e-07,1.967737e-07,1.967739e-07,1.967740e-07,1.967742e-07,1.967743e-07,1.967745e-07,1.967746e-07,1.967748e-07,1.967749e-07,1.967751e-07,1.967753e-07,1.967754e-07,1.967756e-07,1.967757e-07,1.967759e-07,1.967760e-07,1.967762e-07,1.967763e-07,1.967765e-07,1.967766e-07,1.967768e-07,1.967769e-07,1.967771e-07,1.967773e-07,1.967774e-07,1.967776e-07,1.967777e-07,1.967779e-07,1.967780e-07,1.967782e-07,1.967783e-07,1.967785e-07,1.967786e-07,1.967788e-07,1.967789e-07,1.967791e-07,1.967793e-07,1.967794e-07,1.967796e-07,1.967797e-07,1.967799e-07,1.967800e-07,1.967802e-07,1.967803e-07,1.967805e-07,1.967806e-07,1.967808e-07,1.967809e-07,1.967811e-07,1.967813e-07,1.967814e-07,1.967816e-07,1.967817e-07,1.967819e-07,1.967820e-07,1.967822e-07,1.967823e-07,1.967825e-07,1.967826e-07,1.967828e-07,1.967829e-07,1.967831e-07,1.967833e-07,1.967834e-07,1.967836e-07,1.967837e-07,1.967839e-07,1.967840e-07,1.967842e-07,1.967843e-07,1.967845e-07,1.967846e-07,1.967848e-07,1.967849e-07,1.967851e-07,1.967853e-07,1.967854e-07,1.967856e-07,1.967857e-07,1.967859e-07,1.967860e-07,1.967862e-07,1.967863e-07,1.967865e-07,1.967866e-07,1.967868e-07,1.967869e-07,1.967871e-07,1.967872e-07,1.967874e-07,1.967876e-07,1.967877e-07,1.967879e-07,1.967880e-07,1.967882e-07,1.967883e-07,1.967885e-07,1.967886e-07,1.967888e-07,1.967889e-07,1.967891e-07,1.967892e-07,1.967894e-07,1.967896e-07,1.967897e-07,1.967899e-07,1.967900e-07,1.967902e-07,1.967903e-07,1.967905e-07,1.967906e-07,1.967908e-07,1.967909e-07,1.967911e-07,1.967912e-07,1.967914e-07,1.967916e-07,1.967917e-07,1.967919e-07,1.967920e-07,1.967922e-07,1.967923e-07,1.967925e-07,1.967926e-07,1.967928e-07,1.967929e-07,1.967931e-07,1.967932e-07,1.967934e-07,1.967935e-07,1.967937e-07,1.967939e-07,1.967940e-07,1.967942e-07,1.967943e-07,1.967945e-07,1.967946e-07,1.967948e-07,1.967949e-07,1.967951e-07,1.967952e-07,1.967954e-07,1.967955e-07,1.967957e-07,1.967959e-07,1.967960e-07,1.967962e-07,1.967963e-07,1.967965e-07,1.967966e-07,1.967968e-07,1.967969e-07,1.967971e-07,1.967972e-07,1.967974e-07,1.967975e-07,1.967977e-07,1.967978e-07,1.967980e-07,1.967982e-07,1.967983e-07,1.967985e-07,1.967986e-07,1.967988e-07,1.967989e-07,1.967991e-07,1.967992e-07,1.967994e-07,1.967995e-07,1.967997e-07,1.967998e-07,1.968000e-07,1.968002e-07,1.968003e-07,1.968005e-07,1.968006e-07,1.968008e-07,1.968009e-07,1.968011e-07,1.968012e-07,1.968014e-07,1.968015e-07,1.968017e-07,1.968018e-07,1.968020e-07,1.968021e-07,1.968023e-07,1.968025e-07,1.968026e-07,1.968028e-07,1.968029e-07,1.968031e-07,1.968032e-07,1.968034e-07,1.968035e-07,1.968037e-07,1.968038e-07,1.968040e-07,1.968041e-07,1.968043e-07,1.968044e-07,1.968046e-07,1.968048e-07,1.968049e-07,1.968051e-07,1.968052e-07,1.968054e-07,1.968055e-07,1.968057e-07,1.968058e-07,1.968060e-07,1.968061e-07,1.968063e-07,1.968064e-07,1.968066e-07,1.968068e-07,1.968069e-07,1.968071e-07,1.968072e-07,1.968074e-07,1.968075e-07,1.968077e-07,1.968078e-07,1.968080e-07,1.968081e-07,1.968083e-07,1.968084e-07,1.968086e-07,1.968087e-07,1.968089e-07,1.968091e-07,1.968092e-07,1.968094e-07,1.968095e-07,1.968097e-07,1.968098e-07,1.968100e-07,1.968101e-07,1.968103e-07,1.968104e-07,1.968106e-07,1.968107e-07,1.968109e-07,1.968110e-07,1.968112e-07,1.968114e-07,1.968115e-07,1.968117e-07,1.968118e-07,1.968120e-07,1.968121e-07,1.968123e-07,1.968124e-07,1.968126e-07,1.968127e-07,1.968129e-07,1.968130e-07,1.968132e-07,1.968133e-07,1.968135e-07,1.968137e-07,1.968138e-07,1.968140e-07,1.968141e-07,1.968143e-07,1.968144e-07,1.968146e-07,1.968147e-07,1.968149e-07,1.968150e-07,1.968152e-07,1.968153e-07,1.968155e-07,1.968156e-07,1.968158e-07,1.968160e-07,1.968161e-07,1.968163e-07,1.968164e-07,1.968166e-07,1.968167e-07,1.968169e-07,1.968170e-07,1.968172e-07,1.968173e-07,1.968175e-07,1.968176e-07,1.968178e-07,1.968179e-07,1.968181e-07,1.968183e-07,1.968184e-07,1.968186e-07,1.968187e-07,1.968189e-07,1.968190e-07,1.968192e-07,1.968193e-07,1.968195e-07,1.968196e-07,1.968198e-07,1.968199e-07,1.968201e-07,1.968202e-07,1.968204e-07,1.968206e-07,1.968207e-07,1.968209e-07,1.968210e-07,1.968212e-07,1.968213e-07,1.968215e-07,1.968216e-07,1.968218e-07,1.968219e-07,1.968221e-07,1.968222e-07,1.968224e-07,1.968225e-07,1.968227e-07,1.968229e-07,1.968230e-07,1.968232e-07,1.968233e-07,1.968235e-07,1.968236e-07,1.968238e-07,1.968239e-07,1.968241e-07,1.968242e-07,1.968244e-07,1.968245e-07,1.968247e-07,1.968248e-07,1.968250e-07,1.968251e-07,1.968253e-07,1.968255e-07,1.968256e-07,1.968258e-07,1.968259e-07,1.968261e-07,1.968262e-07,1.968264e-07,1.968265e-07,1.968267e-07,1.968268e-07,1.968270e-07,1.968271e-07,1.968273e-07,1.968274e-07,1.968276e-07,1.968278e-07,1.968279e-07,1.968281e-07,1.968282e-07,1.968284e-07,1.968285e-07,1.968287e-07,1.968288e-07,1.968290e-07,1.968291e-07,1.968293e-07,1.968294e-07,1.968296e-07,1.968297e-07,1.968299e-07,1.968301e-07,1.968302e-07,1.968304e-07,1.968305e-07,1.968307e-07,1.968308e-07,1.968310e-07,1.968311e-07,1.968313e-07,1.968314e-07,1.968316e-07,1.968317e-07,1.968319e-07,1.968320e-07,1.968322e-07,1.968323e-07,1.968325e-07,1.968327e-07,1.968328e-07,1.968330e-07,1.968331e-07,1.968333e-07,1.968334e-07,1.968336e-07,1.968337e-07,1.968339e-07,1.968340e-07,1.968342e-07,1.968343e-07,1.968345e-07,1.968346e-07,1.968348e-07,1.968349e-07,1.968351e-07,1.968353e-07,1.968354e-07,1.968356e-07,1.968357e-07,1.968359e-07,1.968360e-07,1.968362e-07,1.968363e-07,1.968365e-07,1.968366e-07,1.968368e-07,1.968369e-07,1.968371e-07,1.968372e-07,1.968374e-07,1.968376e-07,1.968377e-07,1.968379e-07,1.968380e-07,1.968382e-07,1.968383e-07,1.968385e-07,1.968386e-07,1.968388e-07,1.968389e-07,1.968391e-07,1.968392e-07,1.968394e-07,1.968395e-07,1.968397e-07,1.968398e-07,1.968400e-07,1.968402e-07,1.968403e-07,1.968405e-07,1.968406e-07,1.968408e-07,1.968409e-07,1.968411e-07,1.968412e-07,1.968414e-07,1.968415e-07,1.968417e-07,1.968418e-07,1.968420e-07,1.968421e-07,1.968423e-07,1.968424e-07,1.968426e-07,1.968428e-07,1.968429e-07,1.968431e-07,1.968432e-07,1.968434e-07,1.968435e-07,1.968437e-07,1.968438e-07,1.968440e-07,1.968441e-07,1.968443e-07,1.968444e-07,1.968446e-07,1.968447e-07,1.968449e-07,1.968450e-07,1.968452e-07,1.968454e-07,1.968455e-07,1.968457e-07,1.968458e-07,1.968460e-07,1.968461e-07,1.968463e-07,1.968464e-07,1.968466e-07,1.968467e-07,1.968469e-07,1.968470e-07,1.968472e-07,1.968473e-07,1.968475e-07,1.968476e-07,1.968478e-07,1.968480e-07,1.968481e-07,1.968483e-07,1.968484e-07,1.968486e-07,1.968487e-07,1.968489e-07,1.968490e-07,1.968492e-07,1.968493e-07,1.968495e-07,1.968496e-07,1.968498e-07,1.968499e-07,1.968501e-07,1.968502e-07,1.968504e-07,1.968506e-07,1.968507e-07,1.968509e-07,1.968510e-07,1.968512e-07,1.968513e-07,1.968515e-07,1.968516e-07,1.968518e-07,1.968519e-07,1.968521e-07,1.968522e-07,1.968524e-07,1.968525e-07,1.968527e-07,1.968528e-07,1.968530e-07,1.968532e-07,1.968533e-07,1.968535e-07,1.968536e-07,1.968538e-07,1.968539e-07,1.968541e-07,1.968542e-07,1.968544e-07,1.968545e-07,1.968547e-07,1.968548e-07,1.968550e-07,1.968551e-07,1.968553e-07,1.968554e-07,1.968556e-07,1.968557e-07,1.968559e-07,1.968561e-07,1.968562e-07,1.968564e-07,1.968565e-07,1.968567e-07,1.968568e-07,1.968570e-07,1.968571e-07,1.968573e-07,1.968574e-07,1.968576e-07,1.968577e-07,1.968579e-07,1.968580e-07,1.968582e-07,1.968583e-07,1.968585e-07,1.968587e-07,1.968588e-07,1.968590e-07,1.968591e-07,1.968593e-07,1.968594e-07,1.968596e-07,1.968597e-07,1.968599e-07,1.968600e-07,1.968602e-07,1.968603e-07,1.968605e-07,1.968606e-07,1.968608e-07,1.968609e-07,1.968611e-07,1.968612e-07,1.968614e-07,1.968616e-07,1.968617e-07,1.968619e-07,1.968620e-07,1.968622e-07,1.968623e-07,1.968625e-07,1.968626e-07,1.968628e-07,1.968629e-07,1.968631e-07,1.968632e-07,1.968634e-07,1.968635e-07,1.968637e-07,1.968638e-07,1.968640e-07,1.968641e-07,1.968643e-07,1.968645e-07,1.968646e-07,1.968648e-07,1.968649e-07,1.968651e-07,1.968652e-07,1.968654e-07,1.968655e-07,1.968657e-07,1.968658e-07,1.968660e-07,1.968661e-07,1.968663e-07,1.968664e-07,1.968666e-07,1.968667e-07,1.968669e-07,1.968670e-07,1.968672e-07,1.968674e-07,1.968675e-07,1.968677e-07,1.968678e-07,1.968680e-07,1.968681e-07,1.968683e-07,1.968684e-07,1.968686e-07,1.968687e-07,1.968689e-07,1.968690e-07,1.968692e-07,1.968693e-07,1.968695e-07,1.968696e-07,1.968698e-07,1.968699e-07,1.968701e-07,1.968703e-07,1.968704e-07,1.968706e-07,1.968707e-07,1.968709e-07,1.968710e-07,1.968712e-07,1.968713e-07,1.968715e-07,1.968716e-07,1.968718e-07,1.968719e-07,1.968721e-07,1.968722e-07,1.968724e-07,1.968725e-07,1.968727e-07,1.968728e-07,1.968730e-07,1.968732e-07,1.968733e-07,1.968735e-07,1.968736e-07,1.968738e-07,1.968739e-07,1.968741e-07,1.968742e-07,1.968744e-07,1.968745e-07,1.968747e-07,1.968748e-07,1.968750e-07,1.968751e-07,1.968753e-07,1.968754e-07,1.968756e-07,1.968757e-07,1.968759e-07,1.968761e-07,1.968762e-07,1.968764e-07,1.968765e-07,1.968767e-07,1.968768e-07,1.968770e-07,1.968771e-07,1.968773e-07,1.968774e-07,1.968776e-07,1.968777e-07,1.968779e-07,1.968780e-07,1.968782e-07,1.968783e-07,1.968785e-07,1.968786e-07,1.968788e-07,1.968789e-07,1.968791e-07,1.968793e-07,1.968794e-07,1.968796e-07,1.968797e-07,1.968799e-07,1.968800e-07,1.968802e-07,1.968803e-07,1.968805e-07,1.968806e-07,1.968808e-07,1.968809e-07,1.968811e-07,1.968812e-07,1.968814e-07,1.968815e-07,1.968817e-07,1.968818e-07,1.968820e-07,1.968822e-07,1.968823e-07,1.968825e-07,1.968826e-07,1.968828e-07,1.968829e-07,1.968831e-07,1.968832e-07,1.968834e-07,1.968835e-07,1.968837e-07,1.968838e-07,1.968840e-07,1.968841e-07,1.968843e-07,1.968844e-07,1.968846e-07,1.968847e-07,1.968849e-07,1.968850e-07,1.968852e-07,1.968854e-07,1.968855e-07,1.968857e-07,1.968858e-07,1.968860e-07,1.968861e-07,1.968863e-07,1.968864e-07,1.968866e-07,1.968867e-07,1.968869e-07,1.968870e-07,1.968872e-07,1.968873e-07,1.968875e-07,1.968876e-07,1.968878e-07,1.968879e-07,1.968881e-07,1.968882e-07,1.968884e-07,1.968886e-07,1.968887e-07,1.968889e-07,1.968890e-07,1.968892e-07,1.968893e-07,1.968895e-07,1.968896e-07,1.968898e-07,1.968899e-07,1.968901e-07,1.968902e-07,1.968904e-07,1.968905e-07,1.968907e-07,1.968908e-07,1.968910e-07,1.968911e-07,1.968913e-07,1.968914e-07,1.968916e-07,1.968918e-07,1.968919e-07,1.968921e-07,1.968922e-07,1.968924e-07,1.968925e-07,1.968927e-07,1.968928e-07,1.968930e-07,1.968931e-07,1.968933e-07,1.968934e-07,1.968936e-07,1.968937e-07,1.968939e-07,1.968940e-07,1.968942e-07,1.968943e-07,1.968945e-07,1.968946e-07,1.968948e-07,1.968950e-07,1.968951e-07,1.968953e-07,1.968954e-07,1.968956e-07,1.968957e-07,1.968959e-07,1.968960e-07,1.968962e-07,1.968963e-07,1.968965e-07,1.968966e-07,1.968968e-07,1.968969e-07,1.968971e-07,1.968972e-07,1.968974e-07,1.968975e-07,1.968977e-07,1.968978e-07,1.968980e-07,1.968981e-07,1.968983e-07,1.968985e-07,1.968986e-07,1.968988e-07,1.968989e-07,1.968991e-07,1.968992e-07,1.968994e-07,1.968995e-07,1.968997e-07,1.968998e-07,1.969000e-07,1.969001e-07,1.969003e-07,1.969004e-07,1.969006e-07,1.969007e-07,1.969009e-07,1.969010e-07,1.969012e-07,1.969013e-07,1.969015e-07,1.969016e-07,1.969018e-07,1.969020e-07,1.969021e-07,1.969023e-07,1.969024e-07,1.969026e-07,1.969027e-07,1.969029e-07,1.969030e-07,1.969032e-07,1.969033e-07,1.969035e-07,1.969036e-07,1.969038e-07,1.969039e-07,1.969041e-07,1.969042e-07,1.969044e-07,1.969045e-07,1.969047e-07,1.969048e-07,1.969050e-07,1.969051e-07,1.969053e-07,1.969055e-07,1.969056e-07,1.969058e-07,1.969059e-07,1.969061e-07,1.969062e-07,1.969064e-07,1.969065e-07,1.969067e-07,1.969068e-07,1.969070e-07,1.969071e-07,1.969073e-07,1.969074e-07,1.969076e-07,1.969077e-07,1.969079e-07,1.969080e-07,1.969082e-07,1.969083e-07,1.969085e-07,1.969086e-07,1.969088e-07,1.969090e-07,1.969091e-07,1.969093e-07,1.969094e-07,1.969096e-07,1.969097e-07,1.969099e-07,1.969100e-07,1.969102e-07,1.969103e-07,1.969105e-07,1.969106e-07,1.969108e-07,1.969109e-07,1.969111e-07,1.969112e-07,1.969114e-07,1.969115e-07,1.969117e-07,1.969118e-07,1.969120e-07,1.969121e-07,1.969123e-07,1.969124e-07,1.969126e-07,1.969128e-07,1.969129e-07,1.969131e-07,1.969132e-07,1.969134e-07,1.969135e-07,1.969137e-07,1.969138e-07,1.969140e-07,1.969141e-07,1.969143e-07,1.969144e-07,1.969146e-07,1.969147e-07,1.969149e-07,1.969150e-07,1.969152e-07,1.969153e-07,1.969155e-07,1.969156e-07,1.969158e-07,1.969159e-07,1.969161e-07,1.969163e-07,1.969164e-07,1.969166e-07,1.969167e-07,1.969169e-07,1.969170e-07,1.969172e-07,1.969173e-07,1.969175e-07,1.969176e-07,1.969178e-07,1.969179e-07,1.969181e-07,1.969182e-07,1.969184e-07,1.969185e-07,1.969187e-07,1.969188e-07,1.969190e-07,1.969191e-07,1.969193e-07,1.969194e-07,1.969196e-07,1.969197e-07,1.969199e-07,1.969200e-07,1.969202e-07,1.969204e-07,1.969205e-07,1.969207e-07,1.969208e-07,1.969210e-07,1.969211e-07,1.969213e-07,1.969214e-07,1.969216e-07,1.969217e-07,1.969219e-07,1.969220e-07,1.969222e-07,1.969223e-07,1.969225e-07,1.969226e-07,1.969228e-07,1.969229e-07,1.969231e-07,1.969232e-07,1.969234e-07,1.969235e-07,1.969237e-07,1.969238e-07,1.969240e-07,1.969242e-07,1.969243e-07,1.969245e-07,1.969246e-07,1.969248e-07,1.969249e-07,1.969251e-07,1.969252e-07,1.969254e-07,1.969255e-07,1.969257e-07,1.969258e-07,1.969260e-07,1.969261e-07,1.969263e-07,1.969264e-07,1.969266e-07,1.969267e-07,1.969269e-07,1.969270e-07,1.969272e-07,1.969273e-07,1.969275e-07,1.969276e-07,1.969278e-07,1.969279e-07,1.969281e-07,1.969283e-07,1.969284e-07,1.969286e-07,1.969287e-07,1.969289e-07,1.969290e-07,1.969292e-07,1.969293e-07,1.969295e-07,1.969296e-07,1.969298e-07,1.969299e-07,1.969301e-07,1.969302e-07,1.969304e-07,1.969305e-07,1.969307e-07,1.969308e-07,1.969310e-07,1.969311e-07,1.969313e-07,1.969314e-07,1.969316e-07,1.969317e-07,1.969319e-07,1.969320e-07,1.969322e-07,1.969324e-07,1.969325e-07,1.969327e-07,1.969328e-07,1.969330e-07,1.969331e-07,1.969333e-07,1.969334e-07,1.969336e-07,1.969337e-07,1.969339e-07,1.969340e-07,1.969342e-07,1.969343e-07,1.969345e-07,1.969346e-07,1.969348e-07,1.969349e-07,1.969351e-07,1.969352e-07,1.969354e-07,1.969355e-07,1.969357e-07,1.969358e-07,1.969360e-07,1.969361e-07,1.969363e-07,1.969364e-07,1.969366e-07,1.969368e-07,1.969369e-07,1.969371e-07,1.969372e-07,1.969374e-07,1.969375e-07,1.969377e-07,1.969378e-07,1.969380e-07,1.969381e-07,1.969383e-07,1.969384e-07,1.969386e-07,1.969387e-07,1.969389e-07,1.969390e-07,1.969392e-07,1.969393e-07,1.969395e-07,1.969396e-07,1.969398e-07,1.969399e-07,1.969401e-07,1.969402e-07,1.969404e-07,1.969405e-07,1.969407e-07,1.969408e-07,1.969410e-07,1.969412e-07,1.969413e-07,1.969415e-07,1.969416e-07,1.969418e-07,1.969419e-07,1.969421e-07,1.969422e-07,1.969424e-07,1.969425e-07,1.969427e-07,1.969428e-07,1.969430e-07,1.969431e-07,1.969433e-07,1.969434e-07,1.969436e-07,1.969437e-07,1.969439e-07,1.969440e-07,1.969442e-07,1.969443e-07,1.969445e-07,1.969446e-07,1.969448e-07,1.969449e-07,1.969451e-07,1.969452e-07,1.969454e-07,1.969456e-07,1.969457e-07,1.969459e-07,1.969460e-07,1.969462e-07,1.969463e-07,1.969465e-07,1.969466e-07,1.969468e-07,1.969469e-07,1.969471e-07,1.969472e-07,1.969474e-07,1.969475e-07,1.969477e-07,1.969478e-07,1.969480e-07,1.969481e-07,1.969483e-07,1.969484e-07,1.969486e-07,1.969487e-07,1.969489e-07,1.969490e-07,1.969492e-07,1.969493e-07,1.969495e-07,1.969496e-07,1.969498e-07,1.969499e-07,1.969501e-07,1.969503e-07,1.969504e-07,1.969506e-07,1.969507e-07,1.969509e-07,1.969510e-07,1.969512e-07,1.969513e-07,1.969515e-07,1.969516e-07,1.969518e-07,1.969519e-07,1.969521e-07,1.969522e-07,1.969524e-07,1.969525e-07,1.969527e-07,1.969528e-07,1.969530e-07,1.969531e-07,1.969533e-07,1.969534e-07,1.969536e-07,1.969537e-07,1.969539e-07,1.969540e-07,1.969542e-07,1.969543e-07,1.969545e-07,1.969546e-07,1.969548e-07,1.969549e-07,1.969551e-07,1.969553e-07,1.969554e-07,1.969556e-07,1.969557e-07,1.969559e-07,1.969560e-07,1.969562e-07,1.969563e-07,1.969565e-07,1.969566e-07,1.969568e-07,1.969569e-07,1.969571e-07,1.969572e-07,1.969574e-07,1.969575e-07,1.969577e-07,1.969578e-07,1.969580e-07,1.969581e-07,1.969583e-07,1.969584e-07,1.969586e-07,1.969587e-07,1.969589e-07,1.969590e-07,1.969592e-07,1.969593e-07,1.969595e-07,1.969596e-07,1.969598e-07,1.969599e-07,1.969601e-07,1.969602e-07,1.969604e-07,1.969606e-07,1.969607e-07,1.969609e-07,1.969610e-07,1.969612e-07,1.969613e-07,1.969615e-07,1.969616e-07,1.969618e-07,1.969619e-07,1.969621e-07,1.969622e-07,1.969624e-07,1.969625e-07,1.969627e-07,1.969628e-07,1.969630e-07,1.969631e-07,1.969633e-07,1.969634e-07,1.969636e-07,1.969637e-07,1.969639e-07,1.969640e-07,1.969642e-07,1.969643e-07,1.969645e-07,1.969646e-07,1.969648e-07,1.969649e-07,1.969651e-07,1.969652e-07,1.969654e-07,1.969655e-07,1.969657e-07,1.969659e-07,1.969660e-07,1.969662e-07,1.969663e-07,1.969665e-07,1.969666e-07,1.969668e-07,1.969669e-07,1.969671e-07,1.969672e-07,1.969674e-07,1.969675e-07,1.969677e-07,1.969678e-07,1.969680e-07,1.969681e-07,1.969683e-07,1.969684e-07,1.969686e-07,1.969687e-07,1.969689e-07,1.969690e-07,1.969692e-07,1.969693e-07,1.969695e-07,1.969696e-07,1.969698e-07,1.969699e-07,1.969701e-07,1.969702e-07,1.969704e-07,1.969705e-07,1.969707e-07,1.969708e-07,1.969710e-07,1.969711e-07,1.969713e-07,1.969715e-07,1.969716e-07,1.969718e-07,1.969719e-07,1.969721e-07,1.969722e-07,1.969724e-07,1.969725e-07,1.969727e-07,1.969728e-07,1.969730e-07,1.969731e-07,1.969733e-07,1.969734e-07,1.969736e-07,1.969737e-07,1.969739e-07,1.969740e-07,1.969742e-07,1.969743e-07,1.969745e-07,1.969746e-07,1.969748e-07,1.969749e-07,1.969751e-07,1.969752e-07,1.969754e-07,1.969755e-07,1.969757e-07,1.969758e-07,1.969760e-07,1.969761e-07,1.969763e-07,1.969764e-07,1.969766e-07,1.969767e-07,1.969769e-07,1.969770e-07,1.969772e-07,1.969773e-07,1.969775e-07,1.969777e-07,1.969778e-07,1.969780e-07,1.969781e-07,1.969783e-07,1.969784e-07,1.969786e-07,1.969787e-07,1.969789e-07,1.969790e-07,1.969792e-07,1.969793e-07,1.969795e-07,1.969796e-07,1.969798e-07,1.969799e-07,1.969801e-07,1.969802e-07,1.969804e-07,1.969805e-07,1.969807e-07,1.969808e-07,1.969810e-07,1.969811e-07,1.969813e-07,1.969814e-07,1.969816e-07,1.969817e-07,1.969819e-07,1.969820e-07,1.969822e-07,1.969823e-07,1.969825e-07,1.969826e-07,1.969828e-07,1.969829e-07,1.969831e-07,1.969832e-07,1.969834e-07,1.969835e-07,1.969837e-07,1.969838e-07,1.969840e-07,1.969842e-07,1.969843e-07,1.969845e-07,1.969846e-07,1.969848e-07,1.969849e-07,1.969851e-07,1.969852e-07,1.969854e-07,1.969855e-07,1.969857e-07,1.969858e-07,1.969860e-07,1.969861e-07,1.969863e-07,1.969864e-07,1.969866e-07,1.969867e-07,1.969869e-07,1.969870e-07,1.969872e-07,1.969873e-07,1.969875e-07,1.969876e-07,1.969878e-07,1.969879e-07,1.969881e-07,1.969882e-07,1.969884e-07,1.969885e-07,1.969887e-07,1.969888e-07,1.969890e-07,1.969891e-07,1.969893e-07,1.969894e-07,1.969896e-07,1.969897e-07,1.969899e-07,1.969900e-07,1.969902e-07,1.969903e-07,1.969905e-07,1.969906e-07,1.969908e-07,1.969910e-07,1.969911e-07,1.969913e-07,1.969914e-07,1.969916e-07,1.969917e-07,1.969919e-07,1.969920e-07,1.969922e-07,1.969923e-07,1.969925e-07,1.969926e-07,1.969928e-07,1.969929e-07,1.969931e-07,1.969932e-07,1.969934e-07,1.969935e-07,1.969937e-07,1.969938e-07,1.969940e-07,1.969941e-07,1.969943e-07,1.969944e-07,1.969946e-07,1.969947e-07,1.969949e-07,1.969950e-07,1.969952e-07,1.969953e-07,1.969955e-07,1.969956e-07,1.969958e-07,1.969959e-07,1.969961e-07,1.969962e-07,1.969964e-07,1.969965e-07,1.969967e-07,1.969968e-07,1.969970e-07,1.969971e-07,1.969973e-07,1.969974e-07,1.969976e-07,1.969977e-07,1.969979e-07,1.969980e-07,1.969982e-07,1.969983e-07,1.969985e-07,1.969987e-07,1.969988e-07,1.969990e-07,1.969991e-07,1.969993e-07,1.969994e-07,1.969996e-07,1.969997e-07,1.969999e-07,1.970000e-07,1.970002e-07,1.970003e-07,1.970005e-07,1.970006e-07,1.970008e-07,1.970009e-07,1.970011e-07,1.970012e-07,1.970014e-07,1.970015e-07,1.970017e-07,1.970018e-07,1.970020e-07,1.970021e-07,1.970023e-07,1.970024e-07,1.970026e-07,1.970027e-07,1.970029e-07,1.970030e-07,1.970032e-07,1.970033e-07,1.970035e-07,1.970036e-07,1.970038e-07,1.970039e-07,1.970041e-07,1.970042e-07,1.970044e-07,1.970045e-07,1.970047e-07,1.970048e-07,1.970050e-07,1.970051e-07,1.970053e-07,1.970054e-07,1.970056e-07,1.970057e-07,1.970059e-07,1.970060e-07,1.970062e-07,1.970063e-07,1.970065e-07,1.970066e-07,1.970068e-07,1.970069e-07,1.970071e-07,1.970073e-07,1.970074e-07,1.970076e-07,1.970077e-07,1.970079e-07,1.970080e-07,1.970082e-07,1.970083e-07,1.970085e-07,1.970086e-07,1.970088e-07,1.970089e-07,1.970091e-07,1.970092e-07,1.970094e-07,1.970095e-07,1.970097e-07,1.970098e-07,1.970100e-07,1.970101e-07,1.970103e-07,1.970104e-07,1.970106e-07,1.970107e-07,1.970109e-07,1.970110e-07,1.970112e-07,1.970113e-07,1.970115e-07,1.970116e-07,1.970118e-07,1.970119e-07,1.970121e-07,1.970122e-07,1.970124e-07,1.970125e-07,1.970127e-07,1.970128e-07,1.970130e-07,1.970131e-07,1.970133e-07,1.970134e-07,1.970136e-07,1.970137e-07,1.970139e-07,1.970140e-07,1.970142e-07,1.970143e-07,1.970145e-07,1.970146e-07,1.970148e-07,1.970149e-07,1.970151e-07,1.970152e-07,1.970154e-07,1.970155e-07,1.970157e-07,1.970158e-07,1.970160e-07,1.970161e-07,1.970163e-07,1.970164e-07,1.970166e-07,1.970168e-07,1.970169e-07,1.970171e-07,1.970172e-07,1.970174e-07,1.970175e-07,1.970177e-07,1.970178e-07,1.970180e-07,1.970181e-07,1.970183e-07,1.970184e-07,1.970186e-07,1.970187e-07,1.970189e-07,1.970190e-07,1.970192e-07,1.970193e-07,1.970195e-07,1.970196e-07,1.970198e-07,1.970199e-07,1.970201e-07,1.970202e-07,1.970204e-07,1.970205e-07,1.970207e-07,1.970208e-07,1.970210e-07,1.970211e-07,1.970213e-07,1.970214e-07,1.970216e-07,1.970217e-07,1.970219e-07,1.970220e-07,1.970222e-07,1.970223e-07,1.970225e-07,1.970226e-07,1.970228e-07,1.970229e-07,1.970231e-07,1.970232e-07,1.970234e-07,1.970235e-07,1.970237e-07,1.970238e-07,1.970240e-07,1.970241e-07,1.970243e-07,1.970244e-07,1.970246e-07,1.970247e-07,1.970249e-07,1.970250e-07,1.970252e-07,1.970253e-07,1.970255e-07,1.970256e-07,1.970258e-07,1.970259e-07,1.970261e-07,1.970262e-07,1.970264e-07,1.970265e-07,1.970267e-07,1.970268e-07,1.970270e-07,1.970271e-07,1.970273e-07,1.970274e-07,1.970276e-07,1.970277e-07,1.970279e-07,1.970280e-07,1.970282e-07,1.970283e-07,1.970285e-07,1.970286e-07,1.970288e-07,1.970290e-07,1.970291e-07,1.970293e-07,1.970294e-07,1.970296e-07,1.970297e-07,1.970299e-07,1.970300e-07,1.970302e-07,1.970303e-07,1.970305e-07,1.970306e-07,1.970308e-07,1.970309e-07,1.970311e-07,1.970312e-07,1.970314e-07,1.970315e-07,1.970317e-07,1.970318e-07,1.970320e-07,1.970321e-07,1.970323e-07,1.970324e-07,1.970326e-07,1.970327e-07,1.970329e-07,1.970330e-07,1.970332e-07,1.970333e-07,1.970335e-07,1.970336e-07,1.970338e-07,1.970339e-07,1.970341e-07,1.970342e-07,1.970344e-07,1.970345e-07,1.970347e-07,1.970348e-07,1.970350e-07,1.970351e-07,1.970353e-07,1.970354e-07,1.970356e-07,1.970357e-07,1.970359e-07,1.970360e-07,1.970362e-07,1.970363e-07,1.970365e-07,1.970366e-07,1.970368e-07,1.970369e-07,1.970371e-07,1.970372e-07,1.970374e-07,1.970375e-07,1.970377e-07,1.970378e-07,1.970380e-07,1.970381e-07,1.970383e-07,1.970384e-07,1.970386e-07,1.970387e-07,1.970389e-07,1.970390e-07,1.970392e-07,1.970393e-07,1.970395e-07,1.970396e-07,1.970398e-07,1.970399e-07,1.970401e-07,1.970402e-07,1.970404e-07,1.970405e-07,1.970407e-07,1.970408e-07,1.970410e-07,1.970411e-07,1.970413e-07,1.970414e-07,1.970416e-07,1.970417e-07,1.970419e-07,1.970420e-07,1.970422e-07,1.970423e-07,1.970425e-07,1.970426e-07,1.970428e-07,1.970429e-07,1.970431e-07,1.970432e-07,1.970434e-07,1.970435e-07,1.970437e-07,1.970438e-07,1.970440e-07,1.970441e-07,1.970443e-07,1.970444e-07,1.970446e-07,1.970447e-07,1.970449e-07,1.970450e-07,1.970452e-07,1.970453e-07,1.970455e-07,1.970457e-07,1.970458e-07,1.970460e-07,1.970461e-07,1.970463e-07,1.970464e-07,1.970466e-07,1.970467e-07,1.970469e-07,1.970470e-07,1.970472e-07,1.970473e-07,1.970475e-07,1.970476e-07,1.970478e-07,1.970479e-07,1.970481e-07,1.970482e-07,1.970484e-07,1.970485e-07,1.970487e-07,1.970488e-07,1.970490e-07,1.970491e-07,1.970493e-07,1.970494e-07,1.970496e-07,1.970497e-07,1.970499e-07,1.970500e-07,1.970502e-07,1.970503e-07,1.970505e-07,1.970506e-07,1.970508e-07,1.970509e-07,1.970511e-07,1.970512e-07,1.970514e-07,1.970515e-07,1.970517e-07,1.970518e-07,1.970520e-07,1.970521e-07,1.970523e-07,1.970524e-07,1.970526e-07,1.970527e-07,1.970529e-07,1.970530e-07,1.970532e-07,1.970533e-07,1.970535e-07,1.970536e-07,1.970538e-07,1.970539e-07,1.970541e-07,1.970542e-07,1.970544e-07,1.970545e-07,1.970547e-07,1.970548e-07,1.970550e-07,1.970551e-07,1.970553e-07,1.970554e-07,1.970556e-07,1.970557e-07,1.970559e-07,1.970560e-07,1.970562e-07,1.970563e-07,1.970565e-07,1.970566e-07,1.970568e-07,1.970569e-07,1.970571e-07,1.970572e-07,1.970574e-07,1.970575e-07,1.970577e-07,1.970578e-07,1.970580e-07,1.970581e-07,1.970583e-07,1.970584e-07,1.970586e-07,1.970587e-07,1.970589e-07,1.970590e-07,1.970592e-07,1.970593e-07,1.970595e-07,1.970596e-07,1.970598e-07,1.970599e-07,1.970601e-07,1.970602e-07,1.970604e-07,1.970605e-07,1.970607e-07,1.970608e-07,1.970610e-07,1.970611e-07,1.970613e-07,1.970614e-07,1.970616e-07,1.970617e-07,1.970619e-07,1.970620e-07,1.970622e-07,1.970623e-07,1.970625e-07,1.970626e-07,1.970628e-07,1.970629e-07,1.970631e-07,1.970632e-07,1.970634e-07,1.970635e-07,1.970637e-07,1.970638e-07,1.970640e-07,1.970641e-07,1.970643e-07,1.970644e-07,1.970646e-07,1.970647e-07,1.970649e-07,1.970650e-07,1.970652e-07,1.970653e-07,1.970655e-07,1.970656e-07,1.970658e-07,1.970659e-07,1.970661e-07,1.970662e-07,1.970664e-07,1.970665e-07,1.970667e-07,1.970668e-07,1.970670e-07,1.970671e-07,1.970673e-07,1.970674e-07,1.970676e-07,1.970677e-07,1.970679e-07,1.970680e-07,1.970682e-07,1.970683e-07,1.970685e-07,1.970686e-07,1.970688e-07,1.970689e-07,1.970691e-07,1.970692e-07,1.970694e-07,1.970695e-07,1.970697e-07,1.970698e-07,1.970700e-07,1.970701e-07,1.970703e-07,1.970704e-07,1.970706e-07,1.970707e-07,1.970709e-07,1.970710e-07,1.970712e-07,1.970713e-07,1.970715e-07,1.970716e-07,1.970718e-07,1.970719e-07,1.970721e-07,1.970722e-07,1.970724e-07,1.970725e-07,1.970727e-07,1.970728e-07,1.970730e-07,1.970731e-07,1.970733e-07,1.970734e-07,1.970736e-07,1.970737e-07,1.970739e-07,1.970740e-07,1.970742e-07,1.970743e-07,1.970745e-07,1.970746e-07,1.970748e-07,1.970749e-07,1.970751e-07,1.970752e-07,1.970754e-07,1.970755e-07,1.970757e-07,1.970758e-07,1.970760e-07,1.970761e-07,1.970763e-07,1.970764e-07,1.970766e-07,1.970767e-07,1.970769e-07,1.970770e-07,1.970772e-07,1.970773e-07,1.970775e-07,1.970776e-07,1.970778e-07,1.970779e-07,1.970781e-07,1.970782e-07,1.970784e-07,1.970785e-07,1.970787e-07,1.970788e-07,1.970790e-07,1.970791e-07,1.970793e-07,1.970794e-07,1.970796e-07,1.970797e-07,1.970799e-07,1.970800e-07,1.970802e-07,1.970803e-07,1.970805e-07,1.970806e-07,1.970808e-07,1.970809e-07,1.970811e-07,1.970812e-07,1.970814e-07,1.970815e-07,1.970817e-07,1.970818e-07,1.970820e-07,1.970821e-07,1.970823e-07,1.970824e-07,1.970826e-07,1.970827e-07,1.970829e-07,1.970830e-07,1.970832e-07,1.970833e-07,1.970835e-07,1.970836e-07,1.970838e-07,1.970839e-07,1.970841e-07,1.970842e-07,1.970844e-07,1.970845e-07,1.970847e-07,1.970848e-07,1.970850e-07,1.970851e-07,1.970853e-07,1.970854e-07,1.970856e-07,1.970857e-07,1.970859e-07,1.970860e-07,1.970862e-07,1.970863e-07,1.970865e-07,1.970866e-07,1.970868e-07,1.970869e-07,1.970871e-07,1.970872e-07,1.970874e-07,1.970875e-07,1.970877e-07,1.970878e-07,1.970880e-07,1.970881e-07,1.970883e-07,1.970884e-07,1.970886e-07,1.970887e-07,1.970889e-07,1.970890e-07,1.970892e-07,1.970893e-07,1.970895e-07,1.970896e-07,1.970898e-07,1.970899e-07,1.970901e-07,1.970902e-07,1.970904e-07,1.970905e-07,1.970907e-07,1.970908e-07,1.970910e-07,1.970911e-07,1.970913e-07,1.970914e-07,1.970916e-07,1.970917e-07,1.970919e-07,1.970920e-07,1.970922e-07,1.970923e-07,1.970925e-07,1.970926e-07,1.970928e-07,1.970929e-07,1.970931e-07,1.970932e-07,1.970934e-07,1.970935e-07,1.970937e-07,1.970938e-07,1.970940e-07,1.970941e-07,1.970943e-07,1.970944e-07,1.970946e-07,1.970947e-07,1.970949e-07,1.970950e-07,1.970952e-07,1.970953e-07,1.970955e-07,1.970956e-07,1.970958e-07,1.970959e-07,1.970961e-07,1.970962e-07,1.970964e-07,1.970965e-07,1.970967e-07,1.970968e-07,1.970970e-07,1.970971e-07,1.970973e-07,1.970974e-07,1.970976e-07,1.970977e-07,1.970979e-07,1.970980e-07,1.970982e-07,1.970983e-07,1.970984e-07,1.970986e-07,1.970987e-07,1.970989e-07,1.970990e-07,1.970992e-07,1.970993e-07,1.970995e-07,1.970996e-07,1.970998e-07,1.970999e-07,1.971001e-07,1.971002e-07,1.971004e-07,1.971005e-07,1.971007e-07,1.971008e-07,1.971010e-07,1.971011e-07,1.971013e-07,1.971014e-07,1.971016e-07,1.971017e-07,1.971019e-07,1.971020e-07,1.971022e-07,1.971023e-07,1.971025e-07,1.971026e-07,1.971028e-07,1.971029e-07,1.971031e-07,1.971032e-07,1.971034e-07,1.971035e-07,1.971037e-07,1.971038e-07,1.971040e-07,1.971041e-07,1.971043e-07,1.971044e-07,1.971046e-07,1.971047e-07,1.971049e-07,1.971050e-07,1.971052e-07,1.971053e-07,1.971055e-07,1.971056e-07,1.971058e-07,1.971059e-07,1.971061e-07,1.971062e-07,1.971064e-07,1.971065e-07,1.971067e-07,1.971068e-07,1.971070e-07,1.971071e-07,1.971073e-07,1.971074e-07,1.971076e-07,1.971077e-07,1.971079e-07,1.971080e-07,1.971082e-07,1.971083e-07,1.971085e-07,1.971086e-07,1.971088e-07,1.971089e-07,1.971091e-07,1.971092e-07,1.971094e-07,1.971095e-07,1.971097e-07,1.971098e-07,1.971100e-07,1.971101e-07,1.971103e-07,1.971104e-07,1.971106e-07,1.971107e-07,1.971109e-07,1.971110e-07,1.971112e-07,1.971113e-07,1.971115e-07,1.971116e-07,1.971118e-07,1.971119e-07,1.971121e-07,1.971122e-07,1.971124e-07,1.971125e-07,1.971127e-07,1.971128e-07,1.971130e-07,1.971131e-07,1.971133e-07,1.971134e-07,1.971136e-07,1.971137e-07,1.971139e-07,1.971140e-07,1.971142e-07,1.971143e-07,1.971145e-07,1.971146e-07,1.971148e-07,1.971149e-07,1.971151e-07,1.971152e-07,1.971153e-07,1.971155e-07,1.971156e-07,1.971158e-07,1.971159e-07,1.971161e-07,1.971162e-07,1.971164e-07,1.971165e-07,1.971167e-07,1.971168e-07,1.971170e-07,1.971171e-07,1.971173e-07,1.971174e-07,1.971176e-07,1.971177e-07,1.971179e-07,1.971180e-07,1.971182e-07,1.971183e-07,1.971185e-07,1.971186e-07,1.971188e-07,1.971189e-07,1.971191e-07,1.971192e-07,1.971194e-07,1.971195e-07,1.971197e-07,1.971198e-07,1.971200e-07,1.971201e-07,1.971203e-07,1.971204e-07,1.971206e-07,1.971207e-07,1.971209e-07,1.971210e-07,1.971212e-07,1.971213e-07,1.971215e-07,1.971216e-07,1.971218e-07,1.971219e-07,1.971221e-07,1.971222e-07,1.971224e-07,1.971225e-07,1.971227e-07,1.971228e-07,1.971230e-07,1.971231e-07,1.971233e-07,1.971234e-07,1.971236e-07,1.971237e-07,1.971239e-07,1.971240e-07,1.971242e-07,1.971243e-07,1.971245e-07,1.971246e-07,1.971248e-07,1.971249e-07,1.971251e-07,1.971252e-07,1.971254e-07,1.971255e-07,1.971257e-07,1.971258e-07,1.971260e-07,1.971261e-07,1.971263e-07,1.971264e-07,1.971266e-07,1.971267e-07,1.971269e-07,1.971270e-07,1.971271e-07,1.971273e-07,1.971274e-07,1.971276e-07,1.971277e-07,1.971279e-07,1.971280e-07,1.971282e-07,1.971283e-07,1.971285e-07,1.971286e-07,1.971288e-07,1.971289e-07,1.971291e-07,1.971292e-07,1.971294e-07,1.971295e-07,1.971297e-07,1.971298e-07,1.971300e-07,1.971301e-07,1.971303e-07,1.971304e-07,1.971306e-07,1.971307e-07,1.971309e-07,1.971310e-07,1.971312e-07,1.971313e-07,1.971315e-07,1.971316e-07,1.971318e-07,1.971319e-07,1.971321e-07,1.971322e-07,1.971324e-07,1.971325e-07,1.971327e-07,1.971328e-07,1.971330e-07,1.971331e-07,1.971333e-07,1.971334e-07,1.971336e-07,1.971337e-07,1.971339e-07,1.971340e-07,1.971342e-07,1.971343e-07,1.971345e-07,1.971346e-07,1.971348e-07,1.971349e-07,1.971351e-07,1.971352e-07,1.971354e-07,1.971355e-07,1.971357e-07,1.971358e-07,1.971360e-07,1.971361e-07,1.971363e-07,1.971364e-07,1.971366e-07,1.971367e-07,1.971368e-07,1.971370e-07,1.971371e-07,1.971373e-07,1.971374e-07,1.971376e-07,1.971377e-07,1.971379e-07,1.971380e-07,1.971382e-07,1.971383e-07,1.971385e-07,1.971386e-07,1.971388e-07,1.971389e-07,1.971391e-07,1.971392e-07,1.971394e-07,1.971395e-07,1.971397e-07,1.971398e-07,1.971400e-07,1.971401e-07,1.971403e-07,1.971404e-07,1.971406e-07,1.971407e-07,1.971409e-07,1.971410e-07,1.971412e-07,1.971413e-07,1.971415e-07,1.971416e-07,1.971418e-07,1.971419e-07,1.971421e-07,1.971422e-07,1.971424e-07,1.971425e-07,1.971427e-07,1.971428e-07,1.971430e-07,1.971431e-07,1.971433e-07,1.971434e-07,1.971436e-07,1.971437e-07,1.971439e-07,1.971440e-07,1.971442e-07,1.971443e-07,1.971445e-07,1.971446e-07,1.971448e-07,1.971449e-07,1.971451e-07,1.971452e-07,1.971453e-07,1.971455e-07,1.971456e-07,1.971458e-07,1.971459e-07,1.971461e-07,1.971462e-07,1.971464e-07,1.971465e-07,1.971467e-07,1.971468e-07,1.971470e-07,1.971471e-07,1.971473e-07,1.971474e-07,1.971476e-07,1.971477e-07,1.971479e-07,1.971480e-07,1.971482e-07,1.971483e-07,1.971485e-07,1.971486e-07,1.971488e-07,1.971489e-07,1.971491e-07,1.971492e-07,1.971494e-07,1.971495e-07,1.971497e-07,1.971498e-07,1.971500e-07,1.971501e-07,1.971503e-07,1.971504e-07,1.971506e-07,1.971507e-07,1.971509e-07,1.971510e-07,1.971512e-07,1.971513e-07,1.971515e-07,1.971516e-07,1.971518e-07,1.971519e-07,1.971521e-07,1.971522e-07,1.971524e-07,1.971525e-07,1.971527e-07,1.971528e-07,1.971529e-07,1.971531e-07,1.971532e-07,1.971534e-07,1.971535e-07,1.971537e-07,1.971538e-07,1.971540e-07,1.971541e-07,1.971543e-07,1.971544e-07,1.971546e-07,1.971547e-07,1.971549e-07,1.971550e-07,1.971552e-07,1.971553e-07,1.971555e-07,1.971556e-07,1.971558e-07,1.971559e-07,1.971561e-07,1.971562e-07,1.971564e-07,1.971565e-07,1.971567e-07,1.971568e-07,1.971570e-07,1.971571e-07,1.971573e-07,1.971574e-07,1.971576e-07,1.971577e-07,1.971579e-07,1.971580e-07,1.971582e-07,1.971583e-07,1.971585e-07,1.971586e-07,1.971588e-07,1.971589e-07,1.971591e-07,1.971592e-07,1.971594e-07,1.971595e-07,1.971597e-07,1.971598e-07,1.971599e-07,1.971601e-07,1.971602e-07,1.971604e-07,1.971605e-07,1.971607e-07,1.971608e-07,1.971610e-07,1.971611e-07,1.971613e-07,1.971614e-07,1.971616e-07,1.971617e-07,1.971619e-07,1.971620e-07,1.971622e-07,1.971623e-07,1.971625e-07,1.971626e-07,1.971628e-07,1.971629e-07,1.971631e-07,1.971632e-07,1.971634e-07,1.971635e-07,1.971637e-07,1.971638e-07,1.971640e-07,1.971641e-07,1.971643e-07,1.971644e-07,1.971646e-07,1.971647e-07,1.971649e-07,1.971650e-07,1.971652e-07,1.971653e-07,1.971655e-07,1.971656e-07,1.971658e-07,1.971659e-07,1.971661e-07,1.971662e-07,1.971663e-07,1.971665e-07,1.971666e-07,1.971668e-07,1.971669e-07,1.971671e-07,1.971672e-07,1.971674e-07,1.971675e-07,1.971677e-07,1.971678e-07,1.971680e-07,1.971681e-07,1.971683e-07,1.971684e-07,1.971686e-07,1.971687e-07,1.971689e-07,1.971690e-07,1.971692e-07,1.971693e-07,1.971695e-07,1.971696e-07,1.971698e-07,1.971699e-07,1.971701e-07,1.971702e-07,1.971704e-07,1.971705e-07,1.971707e-07,1.971708e-07,1.971710e-07,1.971711e-07,1.971713e-07,1.971714e-07,1.971716e-07,1.971717e-07,1.971719e-07,1.971720e-07,1.971721e-07,1.971723e-07,1.971724e-07,1.971726e-07,1.971727e-07,1.971729e-07,1.971730e-07,1.971732e-07,1.971733e-07,1.971735e-07,1.971736e-07,1.971738e-07,1.971739e-07,1.971741e-07,1.971742e-07,1.971744e-07,1.971745e-07,1.971747e-07,1.971748e-07,1.971750e-07,1.971751e-07,1.971753e-07,1.971754e-07,1.971756e-07,1.971757e-07,1.971759e-07,1.971760e-07,1.971762e-07,1.971763e-07,1.971765e-07,1.971766e-07,1.971768e-07,1.971769e-07,1.971771e-07,1.971772e-07,1.971774e-07,1.971775e-07,1.971777e-07,1.971778e-07,1.971779e-07,1.971781e-07,1.971782e-07,1.971784e-07,1.971785e-07,1.971787e-07,1.971788e-07,1.971790e-07,1.971791e-07,1.971793e-07,1.971794e-07,1.971796e-07,1.971797e-07,1.971799e-07,1.971800e-07,1.971802e-07,1.971803e-07,1.971805e-07,1.971806e-07,1.971808e-07,1.971809e-07,1.971811e-07,1.971812e-07,1.971814e-07,1.971815e-07,1.971817e-07,1.971818e-07,1.971820e-07,1.971821e-07,1.971823e-07,1.971824e-07,1.971826e-07,1.971827e-07,1.971829e-07,1.971830e-07,1.971831e-07,1.971833e-07,1.971834e-07,1.971836e-07,1.971837e-07,1.971839e-07,1.971840e-07,1.971842e-07,1.971843e-07,1.971845e-07,1.971846e-07,1.971848e-07,1.971849e-07,1.971851e-07,1.971852e-07,1.971854e-07,1.971855e-07,1.971857e-07,1.971858e-07,1.971860e-07,1.971861e-07,1.971863e-07,1.971864e-07,1.971866e-07,1.971867e-07,1.971869e-07,1.971870e-07,1.971872e-07,1.971873e-07,1.971875e-07,1.971876e-07,1.971878e-07,1.971879e-07,1.971881e-07,1.971882e-07,1.971883e-07,1.971885e-07,1.971886e-07,1.971888e-07,1.971889e-07,1.971891e-07,1.971892e-07,1.971894e-07,1.971895e-07,1.971897e-07,1.971898e-07,1.971900e-07,1.971901e-07,1.971903e-07,1.971904e-07,1.971906e-07,1.971907e-07,1.971909e-07,1.971910e-07,1.971912e-07,1.971913e-07,1.971915e-07,1.971916e-07,1.971918e-07,1.971919e-07,1.971921e-07,1.971922e-07,1.971924e-07,1.971925e-07,1.971927e-07,1.971928e-07,1.971930e-07,1.971931e-07,1.971932e-07,1.971934e-07,1.971935e-07,1.971937e-07,1.971938e-07,1.971940e-07,1.971941e-07,1.971943e-07,1.971944e-07,1.971946e-07,1.971947e-07,1.971949e-07,1.971950e-07,1.971952e-07,1.971953e-07,1.971955e-07,1.971956e-07,1.971958e-07,1.971959e-07,1.971961e-07,1.971962e-07,1.971964e-07,1.971965e-07,1.971967e-07,1.971968e-07,1.971970e-07,1.971971e-07,1.971973e-07,1.971974e-07,1.971976e-07,1.971977e-07,1.971979e-07,1.971980e-07,1.971981e-07,1.971983e-07,1.971984e-07,1.971986e-07,1.971987e-07,1.971989e-07,1.971990e-07,1.971992e-07,1.971993e-07,1.971995e-07,1.971996e-07,1.971998e-07,1.971999e-07,1.972001e-07,1.972002e-07,1.972004e-07,1.972005e-07,1.972007e-07,1.972008e-07,1.972010e-07,1.972011e-07,1.972013e-07,1.972014e-07,1.972016e-07,1.972017e-07,1.972019e-07,1.972020e-07,1.972022e-07,1.972023e-07,1.972024e-07,1.972026e-07,1.972027e-07,1.972029e-07,1.972030e-07,1.972032e-07,1.972033e-07,1.972035e-07,1.972036e-07,1.972038e-07,1.972039e-07,1.972041e-07,1.972042e-07,1.972044e-07,1.972045e-07,1.972047e-07,1.972048e-07,1.972050e-07,1.972051e-07,1.972053e-07,1.972054e-07,1.972056e-07,1.972057e-07,1.972059e-07,1.972060e-07,1.972062e-07,1.972063e-07,1.972065e-07,1.972066e-07,1.972068e-07,1.972069e-07,1.972070e-07,1.972072e-07,1.972073e-07,1.972075e-07,1.972076e-07,1.972078e-07,1.972079e-07,1.972081e-07,1.972082e-07,1.972084e-07,1.972085e-07,1.972087e-07,1.972088e-07,1.972090e-07,1.972091e-07,1.972093e-07,1.972094e-07,1.972096e-07,1.972097e-07,1.972099e-07,1.972100e-07,1.972102e-07,1.972103e-07,1.972105e-07,1.972106e-07,1.972108e-07,1.972109e-07,1.972110e-07,1.972112e-07,1.972113e-07,1.972115e-07,1.972116e-07,1.972118e-07,1.972119e-07,1.972121e-07,1.972122e-07,1.972124e-07,1.972125e-07,1.972127e-07,1.972128e-07,1.972130e-07,1.972131e-07,1.972133e-07,1.972134e-07,1.972136e-07,1.972137e-07,1.972139e-07,1.972140e-07,1.972142e-07,1.972143e-07,1.972145e-07,1.972146e-07,1.972148e-07,1.972149e-07,1.972151e-07,1.972152e-07,1.972153e-07,1.972155e-07,1.972156e-07,1.972158e-07,1.972159e-07,1.972161e-07,1.972162e-07,1.972164e-07,1.972165e-07,1.972167e-07,1.972168e-07,1.972170e-07,1.972171e-07,1.972173e-07,1.972174e-07,1.972176e-07,1.972177e-07,1.972179e-07,1.972180e-07,1.972182e-07,1.972183e-07,1.972185e-07,1.972186e-07,1.972188e-07,1.972189e-07,1.972191e-07,1.972192e-07,1.972193e-07,1.972195e-07,1.972196e-07,1.972198e-07,1.972199e-07,1.972201e-07,1.972202e-07,1.972204e-07,1.972205e-07,1.972207e-07,1.972208e-07,1.972210e-07,1.972211e-07,1.972213e-07,1.972214e-07,1.972216e-07,1.972217e-07,1.972219e-07,1.972220e-07,1.972222e-07,1.972223e-07,1.972225e-07,1.972226e-07,1.972228e-07,1.972229e-07,1.972231e-07,1.972232e-07,1.972233e-07,1.972235e-07,1.972236e-07,1.972238e-07,1.972239e-07,1.972241e-07,1.972242e-07,1.972244e-07,1.972245e-07,1.972247e-07,1.972248e-07,1.972250e-07,1.972251e-07,1.972253e-07,1.972254e-07,1.972256e-07,1.972257e-07,1.972259e-07,1.972260e-07,1.972262e-07,1.972263e-07,1.972265e-07,1.972266e-07,1.972268e-07,1.972269e-07,1.972270e-07,1.972272e-07,1.972273e-07,1.972275e-07,1.972276e-07,1.972278e-07,1.972279e-07,1.972281e-07,1.972282e-07,1.972284e-07,1.972285e-07,1.972287e-07,1.972288e-07,1.972290e-07,1.972291e-07,1.972293e-07,1.972294e-07,1.972296e-07,1.972297e-07,1.972299e-07,1.972300e-07,1.972302e-07,1.972303e-07,1.972305e-07,1.972306e-07,1.972307e-07,1.972309e-07,1.972310e-07,1.972312e-07,1.972313e-07,1.972315e-07,1.972316e-07,1.972318e-07,1.972319e-07,1.972321e-07,1.972322e-07,1.972324e-07,1.972325e-07,1.972327e-07,1.972328e-07,1.972330e-07,1.972331e-07,1.972333e-07,1.972334e-07,1.972336e-07,1.972337e-07,1.972339e-07,1.972340e-07,1.972342e-07,1.972343e-07,1.972344e-07,1.972346e-07,1.972347e-07,1.972349e-07,1.972350e-07,1.972352e-07,1.972353e-07,1.972355e-07,1.972356e-07,1.972358e-07,1.972359e-07,1.972361e-07,1.972362e-07,1.972364e-07,1.972365e-07,1.972367e-07,1.972368e-07,1.972370e-07,1.972371e-07,1.972373e-07,1.972374e-07,1.972376e-07,1.972377e-07,1.972378e-07,1.972380e-07,1.972381e-07,1.972383e-07,1.972384e-07,1.972386e-07,1.972387e-07,1.972389e-07,1.972390e-07,1.972392e-07,1.972393e-07,1.972395e-07,1.972396e-07,1.972398e-07,1.972399e-07,1.972401e-07,1.972402e-07,1.972404e-07,1.972405e-07,1.972407e-07,1.972408e-07,1.972410e-07,1.972411e-07,1.972412e-07,1.972414e-07,1.972415e-07,1.972417e-07,1.972418e-07,1.972420e-07,1.972421e-07,1.972423e-07,1.972424e-07,1.972426e-07,1.972427e-07,1.972429e-07,1.972430e-07,1.972432e-07,1.972433e-07,1.972435e-07,1.972436e-07,1.972438e-07,1.972439e-07,1.972441e-07,1.972442e-07,1.972444e-07,1.972445e-07,1.972446e-07,1.972448e-07,1.972449e-07,1.972451e-07,1.972452e-07,1.972454e-07,1.972455e-07,1.972457e-07,1.972458e-07,1.972460e-07,1.972461e-07,1.972463e-07,1.972464e-07,1.972466e-07,1.972467e-07,1.972469e-07,1.972470e-07,1.972472e-07,1.972473e-07,1.972475e-07,1.972476e-07,1.972478e-07,1.972479e-07,1.972480e-07,1.972482e-07,1.972483e-07,1.972485e-07,1.972486e-07,1.972488e-07,1.972489e-07,1.972491e-07,1.972492e-07,1.972494e-07,1.972495e-07,1.972497e-07,1.972498e-07,1.972500e-07,1.972501e-07,1.972503e-07,1.972504e-07,1.972506e-07,1.972507e-07,1.972509e-07,1.972510e-07,1.972512e-07,1.972513e-07,1.972514e-07,1.972516e-07,1.972517e-07,1.972519e-07,1.972520e-07,1.972522e-07,1.972523e-07,1.972525e-07,1.972526e-07,1.972528e-07,1.972529e-07,1.972531e-07,1.972532e-07,1.972534e-07,1.972535e-07,1.972537e-07,1.972538e-07,1.972540e-07,1.972541e-07,1.972543e-07,1.972544e-07,1.972545e-07,1.972547e-07,1.972548e-07,1.972550e-07,1.972551e-07,1.972553e-07,1.972554e-07,1.972556e-07,1.972557e-07,1.972559e-07,1.972560e-07,1.972562e-07,1.972563e-07,1.972565e-07,1.972566e-07,1.972568e-07,1.972569e-07,1.972571e-07,1.972572e-07,1.972574e-07,1.972575e-07,1.972576e-07,1.972578e-07,1.972579e-07,1.972581e-07,1.972582e-07,1.972584e-07,1.972585e-07,1.972587e-07,1.972588e-07,1.972590e-07,1.972591e-07,1.972593e-07,1.972594e-07,1.972596e-07,1.972597e-07,1.972599e-07,1.972600e-07,1.972602e-07,1.972603e-07,1.972605e-07,1.972606e-07,1.972607e-07,1.972609e-07,1.972610e-07,1.972612e-07,1.972613e-07,1.972615e-07,1.972616e-07,1.972618e-07,1.972619e-07,1.972621e-07,1.972622e-07,1.972624e-07,1.972625e-07,1.972627e-07,1.972628e-07,1.972630e-07,1.972631e-07,1.972633e-07,1.972634e-07,1.972636e-07,1.972637e-07,1.972638e-07,1.972640e-07,1.972641e-07,1.972643e-07,1.972644e-07,1.972646e-07,1.972647e-07,1.972649e-07,1.972650e-07,1.972652e-07,1.972653e-07,1.972655e-07,1.972656e-07,1.972658e-07,1.972659e-07,1.972661e-07,1.972662e-07,1.972664e-07,1.972665e-07,1.972667e-07,1.972668e-07,1.972669e-07,1.972671e-07,1.972672e-07,1.972674e-07,1.972675e-07,1.972677e-07,1.972678e-07,1.972680e-07,1.972681e-07,1.972683e-07,1.972684e-07,1.972686e-07,1.972687e-07,1.972689e-07,1.972690e-07,1.972692e-07,1.972693e-07,1.972695e-07,1.972696e-07,1.972697e-07,1.972699e-07,1.972700e-07,1.972702e-07,1.972703e-07,1.972705e-07,1.972706e-07,1.972708e-07,1.972709e-07,1.972711e-07,1.972712e-07,1.972714e-07,1.972715e-07,1.972717e-07,1.972718e-07,1.972720e-07,1.972721e-07,1.972723e-07,1.972724e-07,1.972726e-07,1.972727e-07,1.972728e-07,1.972730e-07,1.972731e-07,1.972733e-07,1.972734e-07,1.972736e-07,1.972737e-07,1.972739e-07,1.972740e-07,1.972742e-07,1.972743e-07,1.972745e-07,1.972746e-07,1.972748e-07,1.972749e-07,1.972751e-07,1.972752e-07,1.972754e-07,1.972755e-07,1.972756e-07,1.972758e-07,1.972759e-07,1.972761e-07,1.972762e-07,1.972764e-07,1.972765e-07,1.972767e-07,1.972768e-07,1.972770e-07,1.972771e-07,1.972773e-07,1.972774e-07,1.972776e-07,1.972777e-07,1.972779e-07,1.972780e-07,1.972782e-07,1.972783e-07,1.972784e-07,1.972786e-07,1.972787e-07,1.972789e-07,1.972790e-07,1.972792e-07,1.972793e-07,1.972795e-07,1.972796e-07,1.972798e-07,1.972799e-07,1.972801e-07,1.972802e-07,1.972804e-07,1.972805e-07,1.972807e-07,1.972808e-07,1.972810e-07,1.972811e-07,1.972812e-07,1.972814e-07,1.972815e-07,1.972817e-07,1.972818e-07,1.972820e-07,1.972821e-07,1.972823e-07,1.972824e-07,1.972826e-07,1.972827e-07,1.972829e-07,1.972830e-07,1.972832e-07,1.972833e-07,1.972835e-07,1.972836e-07,1.972838e-07,1.972839e-07,1.972840e-07,1.972842e-07,1.972843e-07,1.972845e-07,1.972846e-07,1.972848e-07,1.972849e-07,1.972851e-07,1.972852e-07,1.972854e-07,1.972855e-07,1.972857e-07,1.972858e-07,1.972860e-07,1.972861e-07,1.972863e-07,1.972864e-07,1.972866e-07,1.972867e-07,1.972868e-07,1.972870e-07,1.972871e-07,1.972873e-07,1.972874e-07,1.972876e-07,1.972877e-07,1.972879e-07,1.972880e-07,1.972882e-07,1.972883e-07,1.972885e-07,1.972886e-07,1.972888e-07,1.972889e-07,1.972891e-07,1.972892e-07,1.972893e-07,1.972895e-07,1.972896e-07,1.972898e-07,1.972899e-07,1.972901e-07,1.972902e-07,1.972904e-07,1.972905e-07,1.972907e-07,1.972908e-07,1.972910e-07,1.972911e-07,1.972913e-07,1.972914e-07,1.972916e-07,1.972917e-07,1.972919e-07,1.972920e-07,1.972921e-07,1.972923e-07,1.972924e-07,1.972926e-07,1.972927e-07,1.972929e-07,1.972930e-07,1.972932e-07,1.972933e-07,1.972935e-07,1.972936e-07,1.972938e-07,1.972939e-07,1.972941e-07,1.972942e-07,1.972944e-07,1.972945e-07,1.972946e-07,1.972948e-07,1.972949e-07,1.972951e-07,1.972952e-07,1.972954e-07,1.972955e-07,1.972957e-07,1.972958e-07,1.972960e-07,1.972961e-07,1.972963e-07,1.972964e-07,1.972966e-07,1.972967e-07,1.972969e-07,1.972970e-07,1.972971e-07,1.972973e-07,1.972974e-07,1.972976e-07,1.972977e-07,1.972979e-07,1.972980e-07,1.972982e-07,1.972983e-07,1.972985e-07,1.972986e-07,1.972988e-07,1.972989e-07,1.972991e-07,1.972992e-07,1.972994e-07,1.972995e-07,1.972997e-07,1.972998e-07,1.972999e-07,1.973001e-07,1.973002e-07,1.973004e-07,1.973005e-07,1.973007e-07,1.973008e-07,1.973010e-07,1.973011e-07,1.973013e-07,1.973014e-07,1.973016e-07,1.973017e-07,1.973019e-07,1.973020e-07,1.973022e-07,1.973023e-07,1.973024e-07,1.973026e-07,1.973027e-07,1.973029e-07,1.973030e-07,1.973032e-07,1.973033e-07,1.973035e-07,1.973036e-07,1.973038e-07,1.973039e-07,1.973041e-07,1.973042e-07,1.973044e-07,1.973045e-07,1.973047e-07,1.973048e-07,1.973049e-07,1.973051e-07,1.973052e-07,1.973054e-07,1.973055e-07,1.973057e-07,1.973058e-07,1.973060e-07,1.973061e-07,1.973063e-07,1.973064e-07,1.973066e-07,1.973067e-07,1.973069e-07,1.973070e-07,1.973072e-07,1.973073e-07,1.973074e-07,1.973076e-07,1.973077e-07,1.973079e-07,1.973080e-07,1.973082e-07,1.973083e-07,1.973085e-07,1.973086e-07,1.973088e-07,1.973089e-07,1.973091e-07,1.973092e-07,1.973094e-07,1.973095e-07,1.973097e-07,1.973098e-07,1.973099e-07,1.973101e-07,1.973102e-07,1.973104e-07,1.973105e-07,1.973107e-07,1.973108e-07,1.973110e-07,1.973111e-07,1.973113e-07,1.973114e-07,1.973116e-07,1.973117e-07,1.973119e-07,1.973120e-07,1.973121e-07,1.973123e-07,1.973124e-07,1.973126e-07,1.973127e-07,1.973129e-07,1.973130e-07,1.973132e-07,1.973133e-07,1.973135e-07,1.973136e-07,1.973138e-07,1.973139e-07,1.973141e-07,1.973142e-07,1.973144e-07,1.973145e-07,1.973146e-07,1.973148e-07,1.973149e-07,1.973151e-07,1.973152e-07,1.973154e-07,1.973155e-07,1.973157e-07,1.973158e-07,1.973160e-07,1.973161e-07,1.973163e-07,1.973164e-07,1.973166e-07,1.973167e-07,1.973169e-07,1.973170e-07,1.973171e-07,1.973173e-07,1.973174e-07,1.973176e-07,1.973177e-07,1.973179e-07,1.973180e-07,1.973182e-07,1.973183e-07,1.973185e-07,1.973186e-07,1.973188e-07,1.973189e-07,1.973191e-07,1.973192e-07,1.973193e-07,1.973195e-07,1.973196e-07,1.973198e-07,1.973199e-07,1.973201e-07,1.973202e-07,1.973204e-07,1.973205e-07,1.973207e-07,1.973208e-07,1.973210e-07,1.973211e-07,1.973213e-07,1.973214e-07,1.973216e-07,1.973217e-07,1.973218e-07,1.973220e-07,1.973221e-07,1.973223e-07,1.973224e-07,1.973226e-07,1.973227e-07,1.973229e-07,1.973230e-07,1.973232e-07,1.973233e-07,1.973235e-07,1.973236e-07,1.973238e-07,1.973239e-07,1.973240e-07,1.973242e-07,1.973243e-07,1.973245e-07,1.973246e-07,1.973248e-07,1.973249e-07,1.973251e-07,1.973252e-07,1.973254e-07,1.973255e-07,1.973257e-07,1.973258e-07,1.973260e-07,1.973261e-07,1.973262e-07,1.973264e-07,1.973265e-07,1.973267e-07,1.973268e-07,1.973270e-07,1.973271e-07,1.973273e-07,1.973274e-07,1.973276e-07,1.973277e-07,1.973279e-07,1.973280e-07,1.973282e-07,1.973283e-07,1.973284e-07,1.973286e-07,1.973287e-07,1.973289e-07,1.973290e-07,1.973292e-07,1.973293e-07,1.973295e-07,1.973296e-07,1.973298e-07,1.973299e-07,1.973301e-07,1.973302e-07,1.973304e-07,1.973305e-07,1.973307e-07,1.973308e-07,1.973309e-07,1.973311e-07,1.973312e-07,1.973314e-07,1.973315e-07,1.973317e-07,1.973318e-07,1.973320e-07,1.973321e-07,1.973323e-07,1.973324e-07,1.973326e-07,1.973327e-07,1.973329e-07,1.973330e-07,1.973331e-07,1.973333e-07,1.973334e-07,1.973336e-07,1.973337e-07,1.973339e-07,1.973340e-07,1.973342e-07,1.973343e-07,1.973345e-07,1.973346e-07,1.973348e-07,1.973349e-07,1.973351e-07,1.973352e-07,1.973353e-07,1.973355e-07,1.973356e-07,1.973358e-07,1.973359e-07,1.973361e-07,1.973362e-07,1.973364e-07,1.973365e-07,1.973367e-07,1.973368e-07,1.973370e-07,1.973371e-07,1.973373e-07,1.973374e-07,1.973375e-07,1.973377e-07,1.973378e-07,1.973380e-07,1.973381e-07,1.973383e-07,1.973384e-07,1.973386e-07,1.973387e-07,1.973389e-07,1.973390e-07,1.973392e-07,1.973393e-07,1.973395e-07,1.973396e-07,1.973397e-07,1.973399e-07,1.973400e-07,1.973402e-07,1.973403e-07,1.973405e-07,1.973406e-07,1.973408e-07,1.973409e-07,1.973411e-07,1.973412e-07,1.973414e-07,1.973415e-07,1.973416e-07,1.973418e-07,1.973419e-07,1.973421e-07,1.973422e-07,1.973424e-07,1.973425e-07,1.973427e-07,1.973428e-07,1.973430e-07,1.973431e-07,1.973433e-07,1.973434e-07,1.973436e-07,1.973437e-07,1.973438e-07,1.973440e-07,1.973441e-07,1.973443e-07,1.973444e-07,1.973446e-07,1.973447e-07,1.973449e-07,1.973450e-07,1.973452e-07,1.973453e-07,1.973455e-07,1.973456e-07,1.973458e-07,1.973459e-07,1.973460e-07,1.973462e-07,1.973463e-07,1.973465e-07,1.973466e-07,1.973468e-07,1.973469e-07,1.973471e-07,1.973472e-07,1.973474e-07,1.973475e-07,1.973477e-07,1.973478e-07,1.973480e-07,1.973481e-07,1.973482e-07,1.973484e-07,1.973485e-07,1.973487e-07,1.973488e-07,1.973490e-07,1.973491e-07,1.973493e-07,1.973494e-07,1.973496e-07,1.973497e-07,1.973499e-07,1.973500e-07,1.973501e-07,1.973503e-07,1.973504e-07,1.973506e-07,1.973507e-07,1.973509e-07,1.973510e-07,1.973512e-07,1.973513e-07,1.973515e-07,1.973516e-07,1.973518e-07,1.973519e-07,1.973521e-07,1.973522e-07,1.973523e-07,1.973525e-07,1.973526e-07,1.973528e-07,1.973529e-07,1.973531e-07,1.973532e-07,1.973534e-07,1.973535e-07,1.973537e-07,1.973538e-07,1.973540e-07,1.973541e-07,1.973542e-07,1.973544e-07,1.973545e-07,1.973547e-07,1.973548e-07,1.973550e-07,1.973551e-07,1.973553e-07,1.973554e-07,1.973556e-07,1.973557e-07,1.973559e-07,1.973560e-07,1.973562e-07,1.973563e-07,1.973564e-07,1.973566e-07,1.973567e-07,1.973569e-07,1.973570e-07,1.973572e-07,1.973573e-07,1.973575e-07,1.973576e-07,1.973578e-07,1.973579e-07,1.973581e-07,1.973582e-07,1.973583e-07,1.973585e-07,1.973586e-07,1.973588e-07,1.973589e-07,1.973591e-07,1.973592e-07,1.973594e-07,1.973595e-07,1.973597e-07,1.973598e-07,1.973600e-07,1.973601e-07,1.973603e-07,1.973604e-07,1.973605e-07,1.973607e-07,1.973608e-07,1.973610e-07,1.973611e-07,1.973613e-07,1.973614e-07,1.973616e-07,1.973617e-07,1.973619e-07,1.973620e-07,1.973622e-07,1.973623e-07,1.973624e-07,1.973626e-07,1.973627e-07,1.973629e-07,1.973630e-07,1.973632e-07,1.973633e-07,1.973635e-07,1.973636e-07,1.973638e-07,1.973639e-07,1.973641e-07,1.973642e-07,1.973643e-07,1.973645e-07,1.973646e-07,1.973648e-07,1.973649e-07,1.973651e-07,1.973652e-07,1.973654e-07,1.973655e-07,1.973657e-07,1.973658e-07,1.973660e-07,1.973661e-07,1.973663e-07,1.973664e-07,1.973665e-07,1.973667e-07,1.973668e-07,1.973670e-07,1.973671e-07,1.973673e-07,1.973674e-07,1.973676e-07,1.973677e-07,1.973679e-07,1.973680e-07,1.973682e-07,1.973683e-07,1.973684e-07,1.973686e-07,1.973687e-07,1.973689e-07,1.973690e-07,1.973692e-07,1.973693e-07,1.973695e-07,1.973696e-07,1.973698e-07,1.973699e-07,1.973701e-07,1.973702e-07,1.973703e-07,1.973705e-07,1.973706e-07,1.973708e-07,1.973709e-07,1.973711e-07,1.973712e-07,1.973714e-07,1.973715e-07,1.973717e-07,1.973718e-07,1.973720e-07,1.973721e-07,1.973722e-07,1.973724e-07,1.973725e-07,1.973727e-07,1.973728e-07,1.973730e-07,1.973731e-07,1.973733e-07,1.973734e-07,1.973736e-07,1.973737e-07,1.973739e-07,1.973740e-07,1.973741e-07,1.973743e-07,1.973744e-07,1.973746e-07,1.973747e-07,1.973749e-07,1.973750e-07,1.973752e-07,1.973753e-07,1.973755e-07,1.973756e-07,1.973758e-07,1.973759e-07,1.973760e-07,1.973762e-07,1.973763e-07,1.973765e-07,1.973766e-07,1.973768e-07,1.973769e-07,1.973771e-07,1.973772e-07,1.973774e-07,1.973775e-07,1.973777e-07,1.973778e-07,1.973779e-07,1.973781e-07,1.973782e-07,1.973784e-07,1.973785e-07,1.973787e-07,1.973788e-07,1.973790e-07,1.973791e-07,1.973793e-07,1.973794e-07,1.973796e-07,1.973797e-07,1.973798e-07,1.973800e-07,1.973801e-07,1.973803e-07,1.973804e-07,1.973806e-07,1.973807e-07,1.973809e-07,1.973810e-07,1.973812e-07,1.973813e-07,1.973815e-07,1.973816e-07,1.973817e-07,1.973819e-07,1.973820e-07,1.973822e-07,1.973823e-07,1.973825e-07,1.973826e-07,1.973828e-07,1.973829e-07,1.973831e-07,1.973832e-07,1.973834e-07,1.973835e-07,1.973836e-07,1.973838e-07,1.973839e-07,1.973841e-07,1.973842e-07,1.973844e-07,1.973845e-07,1.973847e-07,1.973848e-07,1.973850e-07,1.973851e-07,1.973853e-07,1.973854e-07,1.973855e-07,1.973857e-07,1.973858e-07,1.973860e-07,1.973861e-07,1.973863e-07,1.973864e-07,1.973866e-07,1.973867e-07,1.973869e-07,1.973870e-07,1.973871e-07,1.973873e-07,1.973874e-07,1.973876e-07,1.973877e-07,1.973879e-07,1.973880e-07,1.973882e-07,1.973883e-07,1.973885e-07,1.973886e-07,1.973888e-07,1.973889e-07,1.973890e-07,1.973892e-07,1.973893e-07,1.973895e-07,1.973896e-07,1.973898e-07,1.973899e-07,1.973901e-07,1.973902e-07,1.973904e-07,1.973905e-07,1.973907e-07,1.973908e-07,1.973909e-07,1.973911e-07,1.973912e-07,1.973914e-07,1.973915e-07,1.973917e-07,1.973918e-07,1.973920e-07,1.973921e-07,1.973923e-07,1.973924e-07,1.973926e-07,1.973927e-07,1.973928e-07,1.973930e-07,1.973931e-07,1.973933e-07,1.973934e-07,1.973936e-07,1.973937e-07,1.973939e-07,1.973940e-07,1.973942e-07,1.973943e-07,1.973944e-07,1.973946e-07,1.973947e-07,1.973949e-07,1.973950e-07,1.973952e-07,1.973953e-07,1.973955e-07,1.973956e-07,1.973958e-07,1.973959e-07,1.973961e-07,1.973962e-07,1.973963e-07,1.973965e-07,1.973966e-07,1.973968e-07,1.973969e-07,1.973971e-07,1.973972e-07,1.973974e-07,1.973975e-07,1.973977e-07,1.973978e-07,1.973979e-07,1.973981e-07,1.973982e-07,1.973984e-07,1.973985e-07,1.973987e-07,1.973988e-07,1.973990e-07,1.973991e-07,1.973993e-07,1.973994e-07,1.973996e-07,1.973997e-07,1.973998e-07,1.974000e-07,1.974001e-07,1.974003e-07,1.974004e-07,1.974006e-07,1.974007e-07,1.974009e-07,1.974010e-07,1.974012e-07,1.974013e-07,1.974015e-07,1.974016e-07,1.974017e-07,1.974019e-07,1.974020e-07,1.974022e-07,1.974023e-07,1.974025e-07,1.974026e-07,1.974028e-07,1.974029e-07,1.974031e-07,1.974032e-07,1.974033e-07,1.974035e-07,1.974036e-07,1.974038e-07,1.974039e-07,1.974041e-07,1.974042e-07,1.974044e-07,1.974045e-07,1.974047e-07,1.974048e-07,1.974049e-07,1.974051e-07,1.974052e-07,1.974054e-07,1.974055e-07,1.974057e-07,1.974058e-07,1.974060e-07,1.974061e-07,1.974063e-07,1.974064e-07,1.974066e-07,1.974067e-07,1.974068e-07,1.974070e-07,1.974071e-07,1.974073e-07,1.974074e-07,1.974076e-07,1.974077e-07,1.974079e-07,1.974080e-07,1.974082e-07,1.974083e-07,1.974084e-07,1.974086e-07,1.974087e-07,1.974089e-07,1.974090e-07,1.974092e-07,1.974093e-07,1.974095e-07,1.974096e-07,1.974098e-07,1.974099e-07,1.974101e-07,1.974102e-07,1.974103e-07,1.974105e-07,1.974106e-07,1.974108e-07,1.974109e-07,1.974111e-07,1.974112e-07,1.974114e-07,1.974115e-07,1.974117e-07,1.974118e-07,1.974119e-07,1.974121e-07,1.974122e-07,1.974124e-07,1.974125e-07,1.974127e-07,1.974128e-07,1.974130e-07,1.974131e-07,1.974133e-07,1.974134e-07,1.974135e-07,1.974137e-07,1.974138e-07,1.974140e-07,1.974141e-07,1.974143e-07,1.974144e-07,1.974146e-07,1.974147e-07,1.974149e-07,1.974150e-07,1.974152e-07,1.974153e-07,1.974154e-07,1.974156e-07,1.974157e-07,1.974159e-07,1.974160e-07,1.974162e-07,1.974163e-07,1.974165e-07,1.974166e-07,1.974168e-07,1.974169e-07,1.974170e-07,1.974172e-07,1.974173e-07,1.974175e-07,1.974176e-07,1.974178e-07,1.974179e-07,1.974181e-07,1.974182e-07,1.974184e-07,1.974185e-07,1.974186e-07,1.974188e-07,1.974189e-07,1.974191e-07,1.974192e-07,1.974194e-07,1.974195e-07,1.974197e-07,1.974198e-07,1.974200e-07,1.974201e-07,1.974202e-07,1.974204e-07,1.974205e-07,1.974207e-07,1.974208e-07,1.974210e-07,1.974211e-07,1.974213e-07,1.974214e-07,1.974216e-07,1.974217e-07,1.974219e-07,1.974220e-07,1.974221e-07,1.974223e-07,1.974224e-07,1.974226e-07,1.974227e-07,1.974229e-07,1.974230e-07,1.974232e-07,1.974233e-07,1.974235e-07,1.974236e-07,1.974237e-07,1.974239e-07,1.974240e-07,1.974242e-07,1.974243e-07,1.974245e-07,1.974246e-07,1.974248e-07,1.974249e-07,1.974251e-07,1.974252e-07,1.974253e-07,1.974255e-07,1.974256e-07,1.974258e-07,1.974259e-07,1.974261e-07,1.974262e-07,1.974264e-07,1.974265e-07,1.974267e-07,1.974268e-07,1.974269e-07,1.974271e-07,1.974272e-07,1.974274e-07,1.974275e-07,1.974277e-07,1.974278e-07,1.974280e-07,1.974281e-07,1.974283e-07,1.974284e-07,1.974285e-07,1.974287e-07,1.974288e-07,1.974290e-07,1.974291e-07,1.974293e-07,1.974294e-07,1.974296e-07,1.974297e-07,1.974299e-07,1.974300e-07,1.974301e-07,1.974303e-07,1.974304e-07,1.974306e-07,1.974307e-07,1.974309e-07,1.974310e-07,1.974312e-07,1.974313e-07,1.974315e-07,1.974316e-07,1.974317e-07,1.974319e-07,1.974320e-07,1.974322e-07,1.974323e-07,1.974325e-07,1.974326e-07,1.974328e-07,1.974329e-07,1.974331e-07,1.974332e-07,1.974333e-07,1.974335e-07,1.974336e-07,1.974338e-07,1.974339e-07,1.974341e-07,1.974342e-07,1.974344e-07,1.974345e-07,1.974347e-07,1.974348e-07,1.974349e-07,1.974351e-07,1.974352e-07,1.974354e-07,1.974355e-07,1.974357e-07,1.974358e-07,1.974360e-07,1.974361e-07,1.974363e-07,1.974364e-07,1.974365e-07,1.974367e-07,1.974368e-07,1.974370e-07,1.974371e-07,1.974373e-07,1.974374e-07,1.974376e-07,1.974377e-07,1.974379e-07,1.974380e-07,1.974381e-07,1.974383e-07,1.974384e-07,1.974386e-07,1.974387e-07,1.974389e-07,1.974390e-07,1.974392e-07,1.974393e-07,1.974395e-07,1.974396e-07,1.974397e-07,1.974399e-07,1.974400e-07,1.974402e-07,1.974403e-07,1.974405e-07,1.974406e-07,1.974408e-07,1.974409e-07,1.974411e-07,1.974412e-07,1.974413e-07,1.974415e-07,1.974416e-07,1.974418e-07,1.974419e-07,1.974421e-07,1.974422e-07,1.974424e-07,1.974425e-07,1.974427e-07,1.974428e-07,1.974429e-07,1.974431e-07,1.974432e-07,1.974434e-07,1.974435e-07,1.974437e-07,1.974438e-07,1.974440e-07,1.974441e-07,1.974442e-07,1.974444e-07,1.974445e-07,1.974447e-07,1.974448e-07,1.974450e-07,1.974451e-07,1.974453e-07,1.974454e-07,1.974456e-07,1.974457e-07,1.974458e-07,1.974460e-07,1.974461e-07,1.974463e-07,1.974464e-07,1.974466e-07,1.974467e-07,1.974469e-07,1.974470e-07,1.974472e-07,1.974473e-07,1.974474e-07,1.974476e-07,1.974477e-07,1.974479e-07,1.974480e-07,1.974482e-07,1.974483e-07,1.974485e-07,1.974486e-07,1.974488e-07,1.974489e-07,1.974490e-07,1.974492e-07,1.974493e-07,1.974495e-07,1.974496e-07,1.974498e-07,1.974499e-07,1.974501e-07,1.974502e-07,1.974504e-07,1.974505e-07,1.974506e-07,1.974508e-07,1.974509e-07,1.974511e-07,1.974512e-07,1.974514e-07,1.974515e-07,1.974517e-07,1.974518e-07,1.974519e-07,1.974521e-07,1.974522e-07,1.974524e-07,1.974525e-07,1.974527e-07,1.974528e-07,1.974530e-07,1.974531e-07,1.974533e-07,1.974534e-07,1.974535e-07,1.974537e-07,1.974538e-07,1.974540e-07,1.974541e-07,1.974543e-07,1.974544e-07,1.974546e-07,1.974547e-07,1.974549e-07,1.974550e-07,1.974551e-07,1.974553e-07,1.974554e-07,1.974556e-07,1.974557e-07,1.974559e-07,1.974560e-07,1.974562e-07,1.974563e-07,1.974564e-07,1.974566e-07,1.974567e-07,1.974569e-07,1.974570e-07,1.974572e-07,1.974573e-07,1.974575e-07,1.974576e-07,1.974578e-07,1.974579e-07,1.974580e-07,1.974582e-07,1.974583e-07,1.974585e-07,1.974586e-07,1.974588e-07,1.974589e-07,1.974591e-07,1.974592e-07,1.974594e-07,1.974595e-07,1.974596e-07,1.974598e-07,1.974599e-07,1.974601e-07,1.974602e-07,1.974604e-07,1.974605e-07,1.974607e-07,1.974608e-07,1.974609e-07,1.974611e-07,1.974612e-07,1.974614e-07,1.974615e-07,1.974617e-07,1.974618e-07,1.974620e-07,1.974621e-07,1.974623e-07,1.974624e-07,1.974625e-07,1.974627e-07,1.974628e-07,1.974630e-07,1.974631e-07,1.974633e-07,1.974634e-07,1.974636e-07,1.974637e-07,1.974638e-07,1.974640e-07,1.974641e-07,1.974643e-07,1.974644e-07,1.974646e-07,1.974647e-07,1.974649e-07,1.974650e-07,1.974652e-07,1.974653e-07,1.974654e-07,1.974656e-07,1.974657e-07,1.974659e-07,1.974660e-07,1.974662e-07,1.974663e-07,1.974665e-07,1.974666e-07,1.974667e-07,1.974669e-07,1.974670e-07,1.974672e-07,1.974673e-07,1.974675e-07,1.974676e-07,1.974678e-07,1.974679e-07,1.974681e-07,1.974682e-07,1.974683e-07,1.974685e-07,1.974686e-07,1.974688e-07,1.974689e-07,1.974691e-07,1.974692e-07,1.974694e-07,1.974695e-07,1.974696e-07,1.974698e-07,1.974699e-07,1.974701e-07,1.974702e-07,1.974704e-07,1.974705e-07,1.974707e-07,1.974708e-07,1.974710e-07,1.974711e-07,1.974712e-07,1.974714e-07,1.974715e-07,1.974717e-07,1.974718e-07,1.974720e-07,1.974721e-07,1.974723e-07,1.974724e-07,1.974725e-07,1.974727e-07,1.974728e-07,1.974730e-07,1.974731e-07,1.974733e-07,1.974734e-07,1.974736e-07,1.974737e-07,1.974739e-07,1.974740e-07,1.974741e-07,1.974743e-07,1.974744e-07,1.974746e-07,1.974747e-07,1.974749e-07,1.974750e-07,1.974752e-07,1.974753e-07,1.974754e-07,1.974756e-07,1.974757e-07,1.974759e-07,1.974760e-07,1.974762e-07,1.974763e-07,1.974765e-07,1.974766e-07,1.974768e-07,1.974769e-07,1.974770e-07,1.974772e-07,1.974773e-07,1.974775e-07,1.974776e-07,1.974778e-07,1.974779e-07,1.974781e-07,1.974782e-07,1.974783e-07,1.974785e-07,1.974786e-07,1.974788e-07,1.974789e-07,1.974791e-07,1.974792e-07,1.974794e-07,1.974795e-07,1.974797e-07,1.974798e-07,1.974799e-07,1.974801e-07,1.974802e-07,1.974804e-07,1.974805e-07,1.974807e-07,1.974808e-07,1.974810e-07,1.974811e-07,1.974812e-07,1.974814e-07,1.974815e-07,1.974817e-07,1.974818e-07,1.974820e-07,1.974821e-07,1.974823e-07,1.974824e-07,1.974825e-07,1.974827e-07,1.974828e-07,1.974830e-07,1.974831e-07,1.974833e-07,1.974834e-07,1.974836e-07,1.974837e-07,1.974839e-07,1.974840e-07,1.974841e-07,1.974843e-07,1.974844e-07,1.974846e-07,1.974847e-07,1.974849e-07,1.974850e-07,1.974852e-07,1.974853e-07,1.974854e-07,1.974856e-07,1.974857e-07,1.974859e-07,1.974860e-07,1.974862e-07,1.974863e-07,1.974865e-07,1.974866e-07,1.974867e-07,1.974869e-07,1.974870e-07,1.974872e-07,1.974873e-07,1.974875e-07,1.974876e-07,1.974878e-07,1.974879e-07,1.974880e-07,1.974882e-07,1.974883e-07,1.974885e-07,1.974886e-07,1.974888e-07,1.974889e-07,1.974891e-07,1.974892e-07,1.974894e-07,1.974895e-07,1.974896e-07,1.974898e-07,1.974899e-07,1.974901e-07,1.974902e-07,1.974904e-07,1.974905e-07,1.974907e-07,1.974908e-07,1.974909e-07,1.974911e-07,1.974912e-07,1.974914e-07,1.974915e-07,1.974917e-07,1.974918e-07,1.974920e-07,1.974921e-07,1.974922e-07,1.974924e-07,1.974925e-07,1.974927e-07,1.974928e-07,1.974930e-07,1.974931e-07,1.974933e-07,1.974934e-07,1.974935e-07,1.974937e-07,1.974938e-07,1.974940e-07,1.974941e-07,1.974943e-07,1.974944e-07,1.974946e-07,1.974947e-07,1.974949e-07,1.974950e-07,1.974951e-07,1.974953e-07,1.974954e-07,1.974956e-07,1.974957e-07,1.974959e-07,1.974960e-07,1.974962e-07,1.974963e-07,1.974964e-07,1.974966e-07,1.974967e-07,1.974969e-07,1.974970e-07,1.974972e-07,1.974973e-07,1.974975e-07,1.974976e-07,1.974977e-07,1.974979e-07,1.974980e-07,1.974982e-07,1.974983e-07,1.974985e-07,1.974986e-07,1.974988e-07,1.974989e-07,1.974990e-07,1.974992e-07,1.974993e-07,1.974995e-07,1.974996e-07,1.974998e-07,1.974999e-07,1.975001e-07,1.975002e-07,1.975003e-07,1.975005e-07,1.975006e-07,1.975008e-07,1.975009e-07,1.975011e-07,1.975012e-07,1.975014e-07,1.975015e-07,1.975016e-07,1.975018e-07,1.975019e-07,1.975021e-07,1.975022e-07,1.975024e-07,1.975025e-07,1.975027e-07,1.975028e-07,1.975030e-07,1.975031e-07,1.975032e-07,1.975034e-07,1.975035e-07,1.975037e-07,1.975038e-07,1.975040e-07,1.975041e-07,1.975043e-07,1.975044e-07,1.975045e-07,1.975047e-07,1.975048e-07,1.975050e-07,1.975051e-07,1.975053e-07,1.975054e-07,1.975056e-07,1.975057e-07,1.975058e-07,1.975060e-07,1.975061e-07,1.975063e-07,1.975064e-07,1.975066e-07,1.975067e-07,1.975069e-07,1.975070e-07,1.975071e-07,1.975073e-07,1.975074e-07,1.975076e-07,1.975077e-07,1.975079e-07,1.975080e-07,1.975082e-07,1.975083e-07,1.975084e-07,1.975086e-07,1.975087e-07,1.975089e-07,1.975090e-07,1.975092e-07,1.975093e-07,1.975095e-07,1.975096e-07,1.975097e-07,1.975099e-07,1.975100e-07,1.975102e-07,1.975103e-07,1.975105e-07,1.975106e-07,1.975108e-07,1.975109e-07,1.975110e-07,1.975112e-07,1.975113e-07,1.975115e-07,1.975116e-07,1.975118e-07,1.975119e-07,1.975121e-07,1.975122e-07,1.975123e-07,1.975125e-07,1.975126e-07,1.975128e-07,1.975129e-07,1.975131e-07,1.975132e-07,1.975134e-07,1.975135e-07,1.975136e-07,1.975138e-07,1.975139e-07,1.975141e-07,1.975142e-07,1.975144e-07,1.975145e-07,1.975147e-07,1.975148e-07,1.975149e-07,1.975151e-07,1.975152e-07,1.975154e-07,1.975155e-07,1.975157e-07,1.975158e-07,1.975160e-07,1.975161e-07,1.975162e-07,1.975164e-07,1.975165e-07,1.975167e-07,1.975168e-07,1.975170e-07,1.975171e-07,1.975173e-07,1.975174e-07,1.975175e-07,1.975177e-07,1.975178e-07,1.975180e-07,1.975181e-07,1.975183e-07,1.975184e-07,1.975186e-07,1.975187e-07,1.975188e-07,1.975190e-07,1.975191e-07,1.975193e-07,1.975194e-07,1.975196e-07,1.975197e-07,1.975199e-07,1.975200e-07,1.975201e-07,1.975203e-07,1.975204e-07,1.975206e-07,1.975207e-07,1.975209e-07,1.975210e-07,1.975212e-07,1.975213e-07,1.975214e-07,1.975216e-07,1.975217e-07,1.975219e-07,1.975220e-07,1.975222e-07,1.975223e-07,1.975225e-07,1.975226e-07,1.975227e-07,1.975229e-07,1.975230e-07,1.975232e-07,1.975233e-07,1.975235e-07,1.975236e-07,1.975238e-07,1.975239e-07,1.975240e-07,1.975242e-07,1.975243e-07,1.975245e-07,1.975246e-07,1.975248e-07,1.975249e-07,1.975251e-07,1.975252e-07,1.975253e-07,1.975255e-07,1.975256e-07,1.975258e-07,1.975259e-07,1.975261e-07,1.975262e-07,1.975263e-07,1.975265e-07,1.975266e-07,1.975268e-07,1.975269e-07,1.975271e-07,1.975272e-07,1.975274e-07,1.975275e-07,1.975276e-07,1.975278e-07,1.975279e-07,1.975281e-07,1.975282e-07,1.975284e-07,1.975285e-07,1.975287e-07,1.975288e-07,1.975289e-07,1.975291e-07,1.975292e-07,1.975294e-07,1.975295e-07,1.975297e-07,1.975298e-07,1.975300e-07,1.975301e-07,1.975302e-07,1.975304e-07,1.975305e-07,1.975307e-07,1.975308e-07,1.975310e-07,1.975311e-07,1.975313e-07,1.975314e-07,1.975315e-07,1.975317e-07,1.975318e-07,1.975320e-07,1.975321e-07,1.975323e-07,1.975324e-07,1.975326e-07,1.975327e-07,1.975328e-07,1.975330e-07,1.975331e-07,1.975333e-07,1.975334e-07,1.975336e-07,1.975337e-07,1.975339e-07,1.975340e-07,1.975341e-07,1.975343e-07,1.975344e-07,1.975346e-07,1.975347e-07,1.975349e-07,1.975350e-07,1.975351e-07,1.975353e-07,1.975354e-07,1.975356e-07,1.975357e-07,1.975359e-07,1.975360e-07,1.975362e-07,1.975363e-07,1.975364e-07,1.975366e-07,1.975367e-07,1.975369e-07,1.975370e-07,1.975372e-07,1.975373e-07,1.975375e-07,1.975376e-07,1.975377e-07,1.975379e-07,1.975380e-07,1.975382e-07,1.975383e-07,1.975385e-07,1.975386e-07,1.975388e-07,1.975389e-07,1.975390e-07,1.975392e-07,1.975393e-07,1.975395e-07,1.975396e-07,1.975398e-07,1.975399e-07,1.975400e-07,1.975402e-07,1.975403e-07,1.975405e-07,1.975406e-07,1.975408e-07,1.975409e-07,1.975411e-07,1.975412e-07,1.975413e-07,1.975415e-07,1.975416e-07,1.975418e-07,1.975419e-07,1.975421e-07,1.975422e-07,1.975424e-07,1.975425e-07,1.975426e-07,1.975428e-07,1.975429e-07,1.975431e-07,1.975432e-07,1.975434e-07,1.975435e-07,1.975437e-07,1.975438e-07,1.975439e-07,1.975441e-07,1.975442e-07,1.975444e-07,1.975445e-07,1.975447e-07,1.975448e-07,1.975449e-07,1.975451e-07,1.975452e-07,1.975454e-07,1.975455e-07,1.975457e-07,1.975458e-07,1.975460e-07,1.975461e-07,1.975462e-07,1.975464e-07,1.975465e-07,1.975467e-07,1.975468e-07,1.975470e-07,1.975471e-07,1.975473e-07,1.975474e-07,1.975475e-07,1.975477e-07,1.975478e-07,1.975480e-07,1.975481e-07,1.975483e-07,1.975484e-07,1.975485e-07,1.975487e-07,1.975488e-07,1.975490e-07,1.975491e-07,1.975493e-07,1.975494e-07,1.975496e-07,1.975497e-07,1.975498e-07,1.975500e-07,1.975501e-07,1.975503e-07,1.975504e-07,1.975506e-07,1.975507e-07,1.975509e-07,1.975510e-07,1.975511e-07,1.975513e-07,1.975514e-07,1.975516e-07,1.975517e-07,1.975519e-07,1.975520e-07,1.975521e-07,1.975523e-07,1.975524e-07,1.975526e-07,1.975527e-07,1.975529e-07,1.975530e-07,1.975532e-07,1.975533e-07,1.975534e-07,1.975536e-07,1.975537e-07,1.975539e-07,1.975540e-07,1.975542e-07,1.975543e-07,1.975545e-07,1.975546e-07,1.975547e-07,1.975549e-07,1.975550e-07,1.975552e-07,1.975553e-07,1.975555e-07,1.975556e-07,1.975557e-07,1.975559e-07,1.975560e-07,1.975562e-07,1.975563e-07,1.975565e-07,1.975566e-07,1.975568e-07,1.975569e-07,1.975570e-07,1.975572e-07,1.975573e-07,1.975575e-07,1.975576e-07,1.975578e-07,1.975579e-07,1.975581e-07,1.975582e-07,1.975583e-07,1.975585e-07,1.975586e-07,1.975588e-07,1.975589e-07,1.975591e-07,1.975592e-07,1.975593e-07,1.975595e-07,1.975596e-07,1.975598e-07,1.975599e-07,1.975601e-07,1.975602e-07,1.975604e-07,1.975605e-07,1.975606e-07,1.975608e-07,1.975609e-07,1.975611e-07,1.975612e-07,1.975614e-07,1.975615e-07,1.975616e-07,1.975618e-07,1.975619e-07,1.975621e-07,1.975622e-07,1.975624e-07,1.975625e-07,1.975627e-07,1.975628e-07,1.975629e-07,1.975631e-07,1.975632e-07,1.975634e-07,1.975635e-07,1.975637e-07,1.975638e-07,1.975639e-07,1.975641e-07,1.975642e-07,1.975644e-07,1.975645e-07,1.975647e-07,1.975648e-07,1.975650e-07,1.975651e-07,1.975652e-07,1.975654e-07,1.975655e-07,1.975657e-07,1.975658e-07,1.975660e-07,1.975661e-07,1.975663e-07,1.975664e-07,1.975665e-07,1.975667e-07,1.975668e-07,1.975670e-07,1.975671e-07,1.975673e-07,1.975674e-07,1.975675e-07,1.975677e-07,1.975678e-07,1.975680e-07,1.975681e-07,1.975683e-07,1.975684e-07,1.975686e-07,1.975687e-07,1.975688e-07,1.975690e-07,1.975691e-07,1.975693e-07,1.975694e-07,1.975696e-07,1.975697e-07,1.975698e-07,1.975700e-07,1.975701e-07,1.975703e-07,1.975704e-07,1.975706e-07,1.975707e-07,1.975709e-07,1.975710e-07,1.975711e-07,1.975713e-07,1.975714e-07,1.975716e-07,1.975717e-07,1.975719e-07,1.975720e-07,1.975721e-07,1.975723e-07,1.975724e-07,1.975726e-07,1.975727e-07,1.975729e-07,1.975730e-07,1.975732e-07,1.975733e-07,1.975734e-07,1.975736e-07,1.975737e-07,1.975739e-07,1.975740e-07,1.975742e-07,1.975743e-07,1.975744e-07,1.975746e-07,1.975747e-07,1.975749e-07,1.975750e-07,1.975752e-07,1.975753e-07,1.975755e-07,1.975756e-07,1.975757e-07,1.975759e-07,1.975760e-07,1.975762e-07,1.975763e-07,1.975765e-07,1.975766e-07,1.975767e-07,1.975769e-07,1.975770e-07,1.975772e-07,1.975773e-07,1.975775e-07,1.975776e-07,1.975777e-07,1.975779e-07,1.975780e-07,1.975782e-07,1.975783e-07,1.975785e-07,1.975786e-07,1.975788e-07,1.975789e-07,1.975790e-07,1.975792e-07,1.975793e-07,1.975795e-07,1.975796e-07,1.975798e-07,1.975799e-07,1.975800e-07,1.975802e-07,1.975803e-07,1.975805e-07,1.975806e-07,1.975808e-07,1.975809e-07,1.975811e-07,1.975812e-07,1.975813e-07,1.975815e-07,1.975816e-07,1.975818e-07,1.975819e-07,1.975821e-07,1.975822e-07,1.975823e-07,1.975825e-07,1.975826e-07,1.975828e-07,1.975829e-07,1.975831e-07,1.975832e-07,1.975834e-07,1.975835e-07,1.975836e-07,1.975838e-07,1.975839e-07,1.975841e-07,1.975842e-07,1.975844e-07,1.975845e-07,1.975846e-07,1.975848e-07,1.975849e-07,1.975851e-07,1.975852e-07,1.975854e-07,1.975855e-07,1.975856e-07,1.975858e-07,1.975859e-07,1.975861e-07,1.975862e-07,1.975864e-07,1.975865e-07,1.975867e-07,1.975868e-07,1.975869e-07,1.975871e-07,1.975872e-07,1.975874e-07,1.975875e-07,1.975877e-07,1.975878e-07,1.975879e-07,1.975881e-07,1.975882e-07,1.975884e-07,1.975885e-07,1.975887e-07,1.975888e-07,1.975889e-07,1.975891e-07,1.975892e-07,1.975894e-07,1.975895e-07,1.975897e-07,1.975898e-07,1.975900e-07,1.975901e-07,1.975902e-07,1.975904e-07,1.975905e-07,1.975907e-07,1.975908e-07,1.975910e-07,1.975911e-07,1.975912e-07,1.975914e-07,1.975915e-07,1.975917e-07,1.975918e-07,1.975920e-07,1.975921e-07,1.975922e-07,1.975924e-07,1.975925e-07,1.975927e-07,1.975928e-07,1.975930e-07,1.975931e-07,1.975933e-07,1.975934e-07,1.975935e-07,1.975937e-07,1.975938e-07,1.975940e-07,1.975941e-07,1.975943e-07,1.975944e-07,1.975945e-07,1.975947e-07,1.975948e-07,1.975950e-07,1.975951e-07,1.975953e-07,1.975954e-07,1.975955e-07,1.975957e-07,1.975958e-07,1.975960e-07,1.975961e-07,1.975963e-07,1.975964e-07,1.975966e-07,1.975967e-07,1.975968e-07,1.975970e-07,1.975971e-07,1.975973e-07,1.975974e-07,1.975976e-07,1.975977e-07,1.975978e-07,1.975980e-07,1.975981e-07,1.975983e-07,1.975984e-07,1.975986e-07,1.975987e-07,1.975988e-07,1.975990e-07,1.975991e-07,1.975993e-07,1.975994e-07,1.975996e-07,1.975997e-07,1.975999e-07,1.976000e-07,1.976001e-07,1.976003e-07,1.976004e-07,1.976006e-07,1.976007e-07,1.976009e-07,1.976010e-07,1.976011e-07,1.976013e-07,1.976014e-07,1.976016e-07,1.976017e-07,1.976019e-07,1.976020e-07,1.976021e-07,1.976023e-07,1.976024e-07,1.976026e-07,1.976027e-07,1.976029e-07,1.976030e-07,1.976031e-07,1.976033e-07,1.976034e-07,1.976036e-07,1.976037e-07,1.976039e-07,1.976040e-07,1.976042e-07,1.976043e-07,1.976044e-07,1.976046e-07,1.976047e-07,1.976049e-07,1.976050e-07,1.976052e-07,1.976053e-07,1.976054e-07,1.976056e-07,1.976057e-07,1.976059e-07,1.976060e-07,1.976062e-07,1.976063e-07,1.976064e-07,1.976066e-07,1.976067e-07,1.976069e-07,1.976070e-07,1.976072e-07,1.976073e-07,1.976074e-07,1.976076e-07,1.976077e-07,1.976079e-07,1.976080e-07,1.976082e-07,1.976083e-07,1.976085e-07,1.976086e-07,1.976087e-07,1.976089e-07,1.976090e-07,1.976092e-07,1.976093e-07,1.976095e-07,1.976096e-07,1.976097e-07,1.976099e-07,1.976100e-07,1.976102e-07,1.976103e-07,1.976105e-07,1.976106e-07,1.976107e-07,1.976109e-07,1.976110e-07,1.976112e-07,1.976113e-07,1.976115e-07,1.976116e-07,1.976117e-07,1.976119e-07,1.976120e-07,1.976122e-07,1.976123e-07,1.976125e-07,1.976126e-07,1.976128e-07,1.976129e-07,1.976130e-07,1.976132e-07,1.976133e-07,1.976135e-07,1.976136e-07,1.976138e-07,1.976139e-07,1.976140e-07,1.976142e-07,1.976143e-07,1.976145e-07,1.976146e-07,1.976148e-07,1.976149e-07,1.976150e-07,1.976152e-07,1.976153e-07,1.976155e-07,1.976156e-07,1.976158e-07,1.976159e-07,1.976160e-07,1.976162e-07,1.976163e-07,1.976165e-07,1.976166e-07,1.976168e-07,1.976169e-07,1.976170e-07,1.976172e-07,1.976173e-07,1.976175e-07,1.976176e-07,1.976178e-07,1.976179e-07,1.976180e-07,1.976182e-07,1.976183e-07,1.976185e-07,1.976186e-07,1.976188e-07,1.976189e-07,1.976191e-07,1.976192e-07,1.976193e-07,1.976195e-07,1.976196e-07,1.976198e-07,1.976199e-07,1.976201e-07,1.976202e-07,1.976203e-07,1.976205e-07,1.976206e-07,1.976208e-07,1.976209e-07,1.976211e-07,1.976212e-07,1.976213e-07,1.976215e-07,1.976216e-07,1.976218e-07,1.976219e-07,1.976221e-07,1.976222e-07,1.976223e-07,1.976225e-07,1.976226e-07,1.976228e-07,1.976229e-07,1.976231e-07,1.976232e-07,1.976233e-07,1.976235e-07,1.976236e-07,1.976238e-07,1.976239e-07,1.976241e-07,1.976242e-07,1.976243e-07,1.976245e-07,1.976246e-07,1.976248e-07,1.976249e-07,1.976251e-07,1.976252e-07,1.976253e-07,1.976255e-07,1.976256e-07,1.976258e-07,1.976259e-07,1.976261e-07,1.976262e-07,1.976263e-07,1.976265e-07,1.976266e-07,1.976268e-07,1.976269e-07,1.976271e-07,1.976272e-07,1.976274e-07,1.976275e-07,1.976276e-07,1.976278e-07,1.976279e-07,1.976281e-07,1.976282e-07,1.976284e-07,1.976285e-07,1.976286e-07,1.976288e-07,1.976289e-07,1.976291e-07,1.976292e-07,1.976294e-07,1.976295e-07,1.976296e-07,1.976298e-07,1.976299e-07,1.976301e-07,1.976302e-07,1.976304e-07,1.976305e-07,1.976306e-07,1.976308e-07,1.976309e-07,1.976311e-07,1.976312e-07,1.976314e-07,1.976315e-07,1.976316e-07,1.976318e-07,1.976319e-07,1.976321e-07,1.976322e-07,1.976324e-07,1.976325e-07,1.976326e-07,1.976328e-07,1.976329e-07,1.976331e-07,1.976332e-07,1.976334e-07,1.976335e-07,1.976336e-07,1.976338e-07,1.976339e-07,1.976341e-07,1.976342e-07,1.976344e-07,1.976345e-07,1.976346e-07,1.976348e-07,1.976349e-07,1.976351e-07,1.976352e-07,1.976354e-07,1.976355e-07,1.976356e-07,1.976358e-07,1.976359e-07,1.976361e-07,1.976362e-07,1.976364e-07,1.976365e-07,1.976366e-07,1.976368e-07,1.976369e-07,1.976371e-07,1.976372e-07,1.976374e-07,1.976375e-07,1.976376e-07,1.976378e-07,1.976379e-07,1.976381e-07,1.976382e-07,1.976384e-07,1.976385e-07,1.976386e-07,1.976388e-07,1.976389e-07,1.976391e-07,1.976392e-07,1.976394e-07,1.976395e-07,1.976396e-07,1.976398e-07,1.976399e-07,1.976401e-07,1.976402e-07,1.976404e-07,1.976405e-07,1.976406e-07,1.976408e-07,1.976409e-07,1.976411e-07,1.976412e-07,1.976414e-07,1.976415e-07,1.976416e-07,1.976418e-07,1.976419e-07,1.976421e-07,1.976422e-07,1.976424e-07,1.976425e-07,1.976426e-07,1.976428e-07,1.976429e-07,1.976431e-07,1.976432e-07,1.976434e-07,1.976435e-07,1.976436e-07,1.976438e-07,1.976439e-07,1.976441e-07,1.976442e-07,1.976444e-07,1.976445e-07,1.976446e-07,1.976448e-07,1.976449e-07,1.976451e-07,1.976452e-07,1.976454e-07,1.976455e-07,1.976456e-07,1.976458e-07,1.976459e-07,1.976461e-07,1.976462e-07,1.976464e-07,1.976465e-07,1.976466e-07,1.976468e-07,1.976469e-07,1.976471e-07,1.976472e-07,1.976474e-07,1.976475e-07,1.976476e-07,1.976478e-07,1.976479e-07,1.976481e-07,1.976482e-07,1.976484e-07,1.976485e-07,1.976486e-07,1.976488e-07,1.976489e-07,1.976491e-07,1.976492e-07,1.976494e-07,1.976495e-07,1.976496e-07,1.976498e-07,1.976499e-07,1.976501e-07,1.976502e-07,1.976504e-07,1.976505e-07,1.976506e-07,1.976508e-07,1.976509e-07,1.976511e-07,1.976512e-07,1.976514e-07,1.976515e-07,1.976516e-07,1.976518e-07,1.976519e-07,1.976521e-07,1.976522e-07,1.976524e-07,1.976525e-07,1.976526e-07,1.976528e-07,1.976529e-07,1.976531e-07,1.976532e-07,1.976534e-07,1.976535e-07,1.976536e-07,1.976538e-07,1.976539e-07,1.976541e-07,1.976542e-07,1.976544e-07,1.976545e-07,1.976546e-07,1.976548e-07,1.976549e-07,1.976551e-07,1.976552e-07,1.976554e-07,1.976555e-07,1.976556e-07,1.976558e-07,1.976559e-07,1.976561e-07,1.976562e-07,1.976564e-07,1.976565e-07,1.976566e-07,1.976568e-07,1.976569e-07,1.976571e-07,1.976572e-07,1.976574e-07,1.976575e-07,1.976576e-07,1.976578e-07,1.976579e-07,1.976581e-07,1.976582e-07,1.976584e-07,1.976585e-07,1.976586e-07,1.976588e-07,1.976589e-07,1.976591e-07,1.976592e-07,1.976594e-07,1.976595e-07,1.976596e-07,1.976598e-07,1.976599e-07,1.976601e-07,1.976602e-07,1.976603e-07,1.976605e-07,1.976606e-07,1.976608e-07,1.976609e-07,1.976611e-07,1.976612e-07,1.976613e-07,1.976615e-07,1.976616e-07,1.976618e-07,1.976619e-07,1.976621e-07,1.976622e-07,1.976623e-07,1.976625e-07,1.976626e-07,1.976628e-07,1.976629e-07,1.976631e-07,1.976632e-07,1.976633e-07,1.976635e-07,1.976636e-07,1.976638e-07,1.976639e-07,1.976641e-07,1.976642e-07,1.976643e-07,1.976645e-07,1.976646e-07,1.976648e-07,1.976649e-07,1.976651e-07,1.976652e-07,1.976653e-07,1.976655e-07,1.976656e-07,1.976658e-07,1.976659e-07,1.976661e-07,1.976662e-07,1.976663e-07,1.976665e-07,1.976666e-07,1.976668e-07,1.976669e-07,1.976671e-07,1.976672e-07,1.976673e-07,1.976675e-07,1.976676e-07,1.976678e-07,1.976679e-07,1.976681e-07,1.976682e-07,1.976683e-07,1.976685e-07,1.976686e-07,1.976688e-07,1.976689e-07,1.976690e-07,1.976692e-07,1.976693e-07,1.976695e-07,1.976696e-07,1.976698e-07,1.976699e-07,1.976700e-07,1.976702e-07,1.976703e-07,1.976705e-07,1.976706e-07,1.976708e-07,1.976709e-07,1.976710e-07,1.976712e-07,1.976713e-07,1.976715e-07,1.976716e-07,1.976718e-07,1.976719e-07,1.976720e-07,1.976722e-07,1.976723e-07,1.976725e-07,1.976726e-07,1.976728e-07,1.976729e-07,1.976730e-07,1.976732e-07,1.976733e-07,1.976735e-07,1.976736e-07,1.976738e-07,1.976739e-07,1.976740e-07,1.976742e-07,1.976743e-07,1.976745e-07,1.976746e-07,1.976747e-07,1.976749e-07,1.976750e-07,1.976752e-07,1.976753e-07,1.976755e-07,1.976756e-07,1.976757e-07,1.976759e-07,1.976760e-07,1.976762e-07,1.976763e-07,1.976765e-07,1.976766e-07,1.976767e-07,1.976769e-07,1.976770e-07,1.976772e-07,1.976773e-07,1.976775e-07,1.976776e-07,1.976777e-07,1.976779e-07,1.976780e-07,1.976782e-07,1.976783e-07,1.976785e-07,1.976786e-07,1.976787e-07,1.976789e-07,1.976790e-07,1.976792e-07,1.976793e-07,1.976794e-07,1.976796e-07,1.976797e-07,1.976799e-07,1.976800e-07,1.976802e-07,1.976803e-07,1.976804e-07,1.976806e-07,1.976807e-07,1.976809e-07,1.976810e-07,1.976812e-07,1.976813e-07,1.976814e-07,1.976816e-07,1.976817e-07,1.976819e-07,1.976820e-07,1.976822e-07,1.976823e-07,1.976824e-07,1.976826e-07,1.976827e-07,1.976829e-07,1.976830e-07,1.976832e-07,1.976833e-07,1.976834e-07,1.976836e-07,1.976837e-07,1.976839e-07,1.976840e-07,1.976841e-07,1.976843e-07,1.976844e-07,1.976846e-07,1.976847e-07,1.976849e-07,1.976850e-07,1.976851e-07,1.976853e-07,1.976854e-07,1.976856e-07,1.976857e-07,1.976859e-07,1.976860e-07,1.976861e-07,1.976863e-07,1.976864e-07,1.976866e-07,1.976867e-07,1.976869e-07,1.976870e-07,1.976871e-07,1.976873e-07,1.976874e-07,1.976876e-07,1.976877e-07,1.976878e-07,1.976880e-07,1.976881e-07,1.976883e-07,1.976884e-07,1.976886e-07,1.976887e-07,1.976888e-07,1.976890e-07,1.976891e-07,1.976893e-07,1.976894e-07,1.976896e-07,1.976897e-07,1.976898e-07,1.976900e-07,1.976901e-07,1.976903e-07,1.976904e-07,1.976906e-07,1.976907e-07,1.976908e-07,1.976910e-07,1.976911e-07,1.976913e-07,1.976914e-07,1.976915e-07,1.976917e-07,1.976918e-07,1.976920e-07,1.976921e-07,1.976923e-07,1.976924e-07,1.976925e-07,1.976927e-07,1.976928e-07,1.976930e-07,1.976931e-07,1.976933e-07,1.976934e-07,1.976935e-07,1.976937e-07,1.976938e-07,1.976940e-07,1.976941e-07,1.976943e-07,1.976944e-07,1.976945e-07,1.976947e-07,1.976948e-07,1.976950e-07,1.976951e-07,1.976952e-07,1.976954e-07,1.976955e-07,1.976957e-07,1.976958e-07,1.976960e-07,1.976961e-07,1.976962e-07,1.976964e-07,1.976965e-07,1.976967e-07,1.976968e-07,1.976970e-07,1.976971e-07,1.976972e-07,1.976974e-07,1.976975e-07,1.976977e-07,1.976978e-07,1.976979e-07,1.976981e-07,1.976982e-07,1.976984e-07,1.976985e-07,1.976987e-07,1.976988e-07,1.976989e-07,1.976991e-07,1.976992e-07,1.976994e-07,1.976995e-07,1.976997e-07,1.976998e-07,1.976999e-07,1.977001e-07,1.977002e-07,1.977004e-07,1.977005e-07,1.977007e-07,1.977008e-07,1.977009e-07,1.977011e-07,1.977012e-07,1.977014e-07,1.977015e-07,1.977016e-07,1.977018e-07,1.977019e-07,1.977021e-07,1.977022e-07,1.977024e-07,1.977025e-07,1.977026e-07,1.977028e-07,1.977029e-07,1.977031e-07,1.977032e-07,1.977034e-07,1.977035e-07,1.977036e-07,1.977038e-07,1.977039e-07,1.977041e-07,1.977042e-07,1.977043e-07,1.977045e-07,1.977046e-07,1.977048e-07,1.977049e-07,1.977051e-07,1.977052e-07,1.977053e-07,1.977055e-07,1.977056e-07,1.977058e-07,1.977059e-07,1.977061e-07,1.977062e-07,1.977063e-07,1.977065e-07,1.977066e-07,1.977068e-07,1.977069e-07,1.977070e-07,1.977072e-07,1.977073e-07,1.977075e-07,1.977076e-07,1.977078e-07,1.977079e-07,1.977080e-07,1.977082e-07,1.977083e-07,1.977085e-07,1.977086e-07,1.977088e-07,1.977089e-07,1.977090e-07,1.977092e-07,1.977093e-07,1.977095e-07,1.977096e-07,1.977097e-07,1.977099e-07,1.977100e-07,1.977102e-07,1.977103e-07,1.977105e-07,1.977106e-07,1.977107e-07,1.977109e-07,1.977110e-07,1.977112e-07,1.977113e-07,1.977115e-07,1.977116e-07,1.977117e-07,1.977119e-07,1.977120e-07,1.977122e-07,1.977123e-07,1.977124e-07,1.977126e-07,1.977127e-07,1.977129e-07,1.977130e-07,1.977132e-07,1.977133e-07,1.977134e-07,1.977136e-07,1.977137e-07,1.977139e-07,1.977140e-07,1.977141e-07,1.977143e-07,1.977144e-07,1.977146e-07,1.977147e-07,1.977149e-07,1.977150e-07,1.977151e-07,1.977153e-07,1.977154e-07,1.977156e-07,1.977157e-07,1.977159e-07,1.977160e-07,1.977161e-07,1.977163e-07,1.977164e-07,1.977166e-07,1.977167e-07,1.977168e-07,1.977170e-07,1.977171e-07,1.977173e-07,1.977174e-07,1.977176e-07,1.977177e-07,1.977178e-07,1.977180e-07,1.977181e-07,1.977183e-07,1.977184e-07,1.977185e-07,1.977187e-07,1.977188e-07,1.977190e-07,1.977191e-07,1.977193e-07,1.977194e-07,1.977195e-07,1.977197e-07,1.977198e-07,1.977200e-07,1.977201e-07,1.977203e-07,1.977204e-07,1.977205e-07,1.977207e-07,1.977208e-07,1.977210e-07,1.977211e-07,1.977212e-07,1.977214e-07,1.977215e-07,1.977217e-07,1.977218e-07,1.977220e-07,1.977221e-07,1.977222e-07,1.977224e-07,1.977225e-07,1.977227e-07,1.977228e-07,1.977229e-07,1.977231e-07,1.977232e-07,1.977234e-07,1.977235e-07,1.977237e-07,1.977238e-07,1.977239e-07,1.977241e-07,1.977242e-07,1.977244e-07,1.977245e-07,1.977247e-07,1.977248e-07,1.977249e-07,1.977251e-07,1.977252e-07,1.977254e-07,1.977255e-07,1.977256e-07,1.977258e-07,1.977259e-07,1.977261e-07,1.977262e-07,1.977264e-07,1.977265e-07,1.977266e-07,1.977268e-07,1.977269e-07,1.977271e-07,1.977272e-07,1.977273e-07,1.977275e-07,1.977276e-07,1.977278e-07,1.977279e-07,1.977281e-07,1.977282e-07,1.977283e-07,1.977285e-07,1.977286e-07,1.977288e-07,1.977289e-07,1.977290e-07,1.977292e-07,1.977293e-07,1.977295e-07,1.977296e-07,1.977298e-07,1.977299e-07,1.977300e-07,1.977302e-07,1.977303e-07,1.977305e-07,1.977306e-07,1.977308e-07,1.977309e-07,1.977310e-07,1.977312e-07,1.977313e-07,1.977315e-07,1.977316e-07,1.977317e-07,1.977319e-07,1.977320e-07,1.977322e-07,1.977323e-07,1.977325e-07,1.977326e-07,1.977327e-07,1.977329e-07,1.977330e-07,1.977332e-07,1.977333e-07,1.977334e-07,1.977336e-07,1.977337e-07,1.977339e-07,1.977340e-07,1.977342e-07,1.977343e-07,1.977344e-07,1.977346e-07,1.977347e-07,1.977349e-07,1.977350e-07,1.977351e-07,1.977353e-07,1.977354e-07,1.977356e-07,1.977357e-07,1.977359e-07,1.977360e-07,1.977361e-07,1.977363e-07,1.977364e-07,1.977366e-07,1.977367e-07,1.977368e-07,1.977370e-07,1.977371e-07,1.977373e-07,1.977374e-07,1.977376e-07,1.977377e-07,1.977378e-07,1.977380e-07,1.977381e-07,1.977383e-07,1.977384e-07,1.977385e-07,1.977387e-07,1.977388e-07,1.977390e-07,1.977391e-07,1.977393e-07,1.977394e-07,1.977395e-07,1.977397e-07,1.977398e-07,1.977400e-07,1.977401e-07,1.977402e-07,1.977404e-07,1.977405e-07,1.977407e-07,1.977408e-07,1.977410e-07,1.977411e-07,1.977412e-07,1.977414e-07,1.977415e-07,1.977417e-07,1.977418e-07,1.977419e-07,1.977421e-07,1.977422e-07,1.977424e-07,1.977425e-07,1.977427e-07,1.977428e-07,1.977429e-07,1.977431e-07,1.977432e-07,1.977434e-07,1.977435e-07,1.977436e-07,1.977438e-07,1.977439e-07,1.977441e-07,1.977442e-07,1.977444e-07,1.977445e-07,1.977446e-07,1.977448e-07,1.977449e-07,1.977451e-07,1.977452e-07,1.977453e-07,1.977455e-07,1.977456e-07,1.977458e-07,1.977459e-07,1.977461e-07,1.977462e-07,1.977463e-07,1.977465e-07,1.977466e-07,1.977468e-07,1.977469e-07,1.977470e-07,1.977472e-07,1.977473e-07,1.977475e-07,1.977476e-07,1.977478e-07,1.977479e-07,1.977480e-07,1.977482e-07,1.977483e-07,1.977485e-07,1.977486e-07,1.977487e-07,1.977489e-07,1.977490e-07,1.977492e-07,1.977493e-07,1.977495e-07,1.977496e-07,1.977497e-07,1.977499e-07,1.977500e-07,1.977502e-07,1.977503e-07,1.977504e-07,1.977506e-07,1.977507e-07,1.977509e-07,1.977510e-07,1.977512e-07,1.977513e-07,1.977514e-07,1.977516e-07,1.977517e-07,1.977519e-07,1.977520e-07,1.977521e-07,1.977523e-07,1.977524e-07,1.977526e-07,1.977527e-07,1.977528e-07,1.977530e-07,1.977531e-07,1.977533e-07,1.977534e-07,1.977536e-07,1.977537e-07,1.977538e-07,1.977540e-07,1.977541e-07,1.977543e-07,1.977544e-07,1.977545e-07,1.977547e-07,1.977548e-07,1.977550e-07,1.977551e-07,1.977553e-07,1.977554e-07,1.977555e-07,1.977557e-07,1.977558e-07,1.977560e-07,1.977561e-07,1.977562e-07,1.977564e-07,1.977565e-07,1.977567e-07,1.977568e-07,1.977570e-07,1.977571e-07,1.977572e-07,1.977574e-07,1.977575e-07,1.977577e-07,1.977578e-07,1.977579e-07,1.977581e-07,1.977582e-07,1.977584e-07,1.977585e-07,1.977587e-07,1.977588e-07,1.977589e-07,1.977591e-07,1.977592e-07,1.977594e-07,1.977595e-07,1.977596e-07,1.977598e-07,1.977599e-07,1.977601e-07,1.977602e-07,1.977603e-07,1.977605e-07,1.977606e-07,1.977608e-07,1.977609e-07,1.977611e-07,1.977612e-07,1.977613e-07,1.977615e-07,1.977616e-07,1.977618e-07,1.977619e-07,1.977620e-07,1.977622e-07,1.977623e-07,1.977625e-07,1.977626e-07,1.977628e-07,1.977629e-07,1.977630e-07,1.977632e-07,1.977633e-07,1.977635e-07,1.977636e-07,1.977637e-07,1.977639e-07,1.977640e-07,1.977642e-07,1.977643e-07,1.977644e-07,1.977646e-07,1.977647e-07,1.977649e-07,1.977650e-07,1.977652e-07,1.977653e-07,1.977654e-07,1.977656e-07,1.977657e-07,1.977659e-07,1.977660e-07,1.977661e-07,1.977663e-07,1.977664e-07,1.977666e-07,1.977667e-07,1.977669e-07,1.977670e-07,1.977671e-07,1.977673e-07,1.977674e-07,1.977676e-07,1.977677e-07,1.977678e-07,1.977680e-07,1.977681e-07,1.977683e-07,1.977684e-07,1.977685e-07,1.977687e-07,1.977688e-07,1.977690e-07,1.977691e-07,1.977693e-07,1.977694e-07,1.977695e-07,1.977697e-07,1.977698e-07,1.977700e-07,1.977701e-07,1.977702e-07,1.977704e-07,1.977705e-07,1.977707e-07,1.977708e-07,1.977710e-07,1.977711e-07,1.977712e-07,1.977714e-07,1.977715e-07,1.977717e-07,1.977718e-07,1.977719e-07,1.977721e-07,1.977722e-07,1.977724e-07,1.977725e-07,1.977726e-07,1.977728e-07,1.977729e-07,1.977731e-07,1.977732e-07,1.977734e-07,1.977735e-07,1.977736e-07,1.977738e-07,1.977739e-07,1.977741e-07,1.977742e-07,1.977743e-07,1.977745e-07,1.977746e-07,1.977748e-07,1.977749e-07,1.977750e-07,1.977752e-07,1.977753e-07,1.977755e-07,1.977756e-07,1.977758e-07,1.977759e-07,1.977760e-07,1.977762e-07,1.977763e-07,1.977765e-07,1.977766e-07,1.977767e-07,1.977769e-07,1.977770e-07,1.977772e-07,1.977773e-07,1.977775e-07,1.977776e-07,1.977777e-07,1.977779e-07,1.977780e-07,1.977782e-07,1.977783e-07,1.977784e-07,1.977786e-07,1.977787e-07,1.977789e-07,1.977790e-07,1.977791e-07,1.977793e-07,1.977794e-07,1.977796e-07,1.977797e-07,1.977799e-07,1.977800e-07,1.977801e-07,1.977803e-07,1.977804e-07,1.977806e-07,1.977807e-07,1.977808e-07,1.977810e-07,1.977811e-07,1.977813e-07,1.977814e-07,1.977815e-07,1.977817e-07,1.977818e-07,1.977820e-07,1.977821e-07,1.977823e-07,1.977824e-07,1.977825e-07,1.977827e-07,1.977828e-07,1.977830e-07,1.977831e-07,1.977832e-07,1.977834e-07,1.977835e-07,1.977837e-07,1.977838e-07,1.977839e-07,1.977841e-07,1.977842e-07,1.977844e-07,1.977845e-07,1.977847e-07,1.977848e-07,1.977849e-07,1.977851e-07,1.977852e-07,1.977854e-07,1.977855e-07,1.977856e-07,1.977858e-07,1.977859e-07,1.977861e-07,1.977862e-07,1.977863e-07,1.977865e-07,1.977866e-07,1.977868e-07,1.977869e-07,1.977871e-07,1.977872e-07,1.977873e-07,1.977875e-07,1.977876e-07,1.977878e-07,1.977879e-07,1.977880e-07,1.977882e-07,1.977883e-07,1.977885e-07,1.977886e-07,1.977887e-07,1.977889e-07,1.977890e-07,1.977892e-07,1.977893e-07,1.977894e-07,1.977896e-07,1.977897e-07,1.977899e-07,1.977900e-07,1.977902e-07,1.977903e-07,1.977904e-07,1.977906e-07,1.977907e-07,1.977909e-07,1.977910e-07,1.977911e-07,1.977913e-07,1.977914e-07,1.977916e-07,1.977917e-07,1.977918e-07,1.977920e-07,1.977921e-07,1.977923e-07,1.977924e-07,1.977926e-07,1.977927e-07,1.977928e-07,1.977930e-07,1.977931e-07,1.977933e-07,1.977934e-07,1.977935e-07,1.977937e-07,1.977938e-07,1.977940e-07,1.977941e-07,1.977942e-07,1.977944e-07,1.977945e-07,1.977947e-07,1.977948e-07,1.977949e-07,1.977951e-07,1.977952e-07,1.977954e-07,1.977955e-07,1.977957e-07,1.977958e-07,1.977959e-07,1.977961e-07,1.977962e-07,1.977964e-07,1.977965e-07,1.977966e-07,1.977968e-07,1.977969e-07,1.977971e-07,1.977972e-07,1.977973e-07,1.977975e-07,1.977976e-07,1.977978e-07,1.977979e-07,1.977981e-07,1.977982e-07,1.977983e-07,1.977985e-07,1.977986e-07,1.977988e-07,1.977989e-07,1.977990e-07,1.977992e-07,1.977993e-07,1.977995e-07,1.977996e-07,1.977997e-07,1.977999e-07,1.978000e-07,1.978002e-07,1.978003e-07,1.978004e-07,1.978006e-07,1.978007e-07,1.978009e-07,1.978010e-07,1.978012e-07,1.978013e-07,1.978014e-07,1.978016e-07,1.978017e-07,1.978019e-07,1.978020e-07,1.978021e-07,1.978023e-07,1.978024e-07,1.978026e-07,1.978027e-07,1.978028e-07,1.978030e-07,1.978031e-07,1.978033e-07,1.978034e-07,1.978035e-07,1.978037e-07,1.978038e-07,1.978040e-07,1.978041e-07,1.978043e-07,1.978044e-07,1.978045e-07,1.978047e-07,1.978048e-07,1.978050e-07,1.978051e-07,1.978052e-07,1.978054e-07,1.978055e-07,1.978057e-07,1.978058e-07,1.978059e-07,1.978061e-07,1.978062e-07,1.978064e-07,1.978065e-07,1.978066e-07,1.978068e-07,1.978069e-07,1.978071e-07,1.978072e-07,1.978074e-07,1.978075e-07,1.978076e-07,1.978078e-07,1.978079e-07,1.978081e-07,1.978082e-07,1.978083e-07,1.978085e-07,1.978086e-07,1.978088e-07,1.978089e-07,1.978090e-07,1.978092e-07,1.978093e-07,1.978095e-07,1.978096e-07,1.978097e-07,1.978099e-07,1.978100e-07,1.978102e-07,1.978103e-07,1.978105e-07,1.978106e-07,1.978107e-07,1.978109e-07,1.978110e-07,1.978112e-07,1.978113e-07,1.978114e-07,1.978116e-07,1.978117e-07,1.978119e-07,1.978120e-07,1.978121e-07,1.978123e-07,1.978124e-07,1.978126e-07,1.978127e-07,1.978128e-07,1.978130e-07,1.978131e-07,1.978133e-07,1.978134e-07,1.978136e-07,1.978137e-07,1.978138e-07,1.978140e-07,1.978141e-07,1.978143e-07,1.978144e-07,1.978145e-07,1.978147e-07,1.978148e-07,1.978150e-07,1.978151e-07,1.978152e-07,1.978154e-07,1.978155e-07,1.978157e-07,1.978158e-07,1.978159e-07,1.978161e-07,1.978162e-07,1.978164e-07,1.978165e-07,1.978166e-07,1.978168e-07,1.978169e-07,1.978171e-07,1.978172e-07,1.978174e-07,1.978175e-07,1.978176e-07,1.978178e-07,1.978179e-07,1.978181e-07,1.978182e-07,1.978183e-07,1.978185e-07,1.978186e-07,1.978188e-07,1.978189e-07,1.978190e-07,1.978192e-07,1.978193e-07,1.978195e-07,1.978196e-07,1.978197e-07,1.978199e-07,1.978200e-07,1.978202e-07,1.978203e-07,1.978204e-07,1.978206e-07,1.978207e-07,1.978209e-07,1.978210e-07,1.978212e-07,1.978213e-07,1.978214e-07,1.978216e-07,1.978217e-07,1.978219e-07,1.978220e-07,1.978221e-07,1.978223e-07,1.978224e-07,1.978226e-07,1.978227e-07,1.978228e-07,1.978230e-07,1.978231e-07,1.978233e-07,1.978234e-07,1.978235e-07,1.978237e-07,1.978238e-07,1.978240e-07,1.978241e-07,1.978242e-07,1.978244e-07,1.978245e-07,1.978247e-07,1.978248e-07,1.978249e-07,1.978251e-07,1.978252e-07,1.978254e-07,1.978255e-07,1.978257e-07,1.978258e-07,1.978259e-07,1.978261e-07,1.978262e-07,1.978264e-07,1.978265e-07,1.978266e-07,1.978268e-07,1.978269e-07,1.978271e-07,1.978272e-07,1.978273e-07,1.978275e-07,1.978276e-07,1.978278e-07,1.978279e-07,1.978280e-07,1.978282e-07,1.978283e-07,1.978285e-07,1.978286e-07,1.978287e-07,1.978289e-07,1.978290e-07,1.978292e-07,1.978293e-07,1.978294e-07,1.978296e-07,1.978297e-07,1.978299e-07,1.978300e-07,1.978302e-07,1.978303e-07,1.978304e-07,1.978306e-07,1.978307e-07,1.978309e-07,1.978310e-07,1.978311e-07,1.978313e-07,1.978314e-07,1.978316e-07,1.978317e-07,1.978318e-07,1.978320e-07,1.978321e-07,1.978323e-07,1.978324e-07,1.978325e-07,1.978327e-07,1.978328e-07,1.978330e-07,1.978331e-07,1.978332e-07,1.978334e-07,1.978335e-07,1.978337e-07,1.978338e-07,1.978339e-07,1.978341e-07,1.978342e-07,1.978344e-07,1.978345e-07,1.978347e-07,1.978348e-07,1.978349e-07,1.978351e-07,1.978352e-07,1.978354e-07,1.978355e-07,1.978356e-07,1.978358e-07,1.978359e-07,1.978361e-07,1.978362e-07,1.978363e-07,1.978365e-07,1.978366e-07,1.978368e-07,1.978369e-07,1.978370e-07,1.978372e-07,1.978373e-07,1.978375e-07,1.978376e-07,1.978377e-07,1.978379e-07,1.978380e-07,1.978382e-07,1.978383e-07,1.978384e-07,1.978386e-07,1.978387e-07,1.978389e-07,1.978390e-07,1.978391e-07,1.978393e-07,1.978394e-07,1.978396e-07,1.978397e-07,1.978398e-07,1.978400e-07,1.978401e-07,1.978403e-07,1.978404e-07,1.978406e-07,1.978407e-07,1.978408e-07,1.978410e-07,1.978411e-07,1.978413e-07,1.978414e-07,1.978415e-07,1.978417e-07,1.978418e-07,1.978420e-07,1.978421e-07,1.978422e-07,1.978424e-07,1.978425e-07,1.978427e-07,1.978428e-07,1.978429e-07,1.978431e-07,1.978432e-07,1.978434e-07,1.978435e-07,1.978436e-07,1.978438e-07,1.978439e-07,1.978441e-07,1.978442e-07,1.978443e-07,1.978445e-07,1.978446e-07,1.978448e-07,1.978449e-07,1.978450e-07,1.978452e-07,1.978453e-07,1.978455e-07,1.978456e-07,1.978457e-07,1.978459e-07,1.978460e-07,1.978462e-07,1.978463e-07,1.978465e-07,1.978466e-07,1.978467e-07,1.978469e-07,1.978470e-07,1.978472e-07,1.978473e-07,1.978474e-07,1.978476e-07,1.978477e-07,1.978479e-07,1.978480e-07,1.978481e-07,1.978483e-07,1.978484e-07,1.978486e-07,1.978487e-07,1.978488e-07,1.978490e-07,1.978491e-07,1.978493e-07,1.978494e-07,1.978495e-07,1.978497e-07,1.978498e-07,1.978500e-07,1.978501e-07,1.978502e-07,1.978504e-07,1.978505e-07,1.978507e-07,1.978508e-07,1.978509e-07,1.978511e-07,1.978512e-07,1.978514e-07,1.978515e-07,1.978516e-07,1.978518e-07,1.978519e-07,1.978521e-07,1.978522e-07,1.978523e-07,1.978525e-07,1.978526e-07,1.978528e-07,1.978529e-07,1.978530e-07,1.978532e-07,1.978533e-07,1.978535e-07,1.978536e-07,1.978537e-07,1.978539e-07,1.978540e-07,1.978542e-07,1.978543e-07,1.978545e-07,1.978546e-07,1.978547e-07,1.978549e-07,1.978550e-07,1.978552e-07,1.978553e-07,1.978554e-07,1.978556e-07,1.978557e-07,1.978559e-07,1.978560e-07,1.978561e-07,1.978563e-07,1.978564e-07,1.978566e-07,1.978567e-07,1.978568e-07,1.978570e-07,1.978571e-07,1.978573e-07,1.978574e-07,1.978575e-07,1.978577e-07,1.978578e-07,1.978580e-07,1.978581e-07,1.978582e-07,1.978584e-07,1.978585e-07,1.978587e-07,1.978588e-07,1.978589e-07,1.978591e-07,1.978592e-07,1.978594e-07,1.978595e-07,1.978596e-07,1.978598e-07,1.978599e-07,1.978601e-07,1.978602e-07,1.978603e-07,1.978605e-07,1.978606e-07,1.978608e-07,1.978609e-07,1.978610e-07,1.978612e-07,1.978613e-07,1.978615e-07,1.978616e-07,1.978617e-07,1.978619e-07,1.978620e-07,1.978622e-07,1.978623e-07,1.978624e-07,1.978626e-07,1.978627e-07,1.978629e-07,1.978630e-07,1.978631e-07,1.978633e-07,1.978634e-07,1.978636e-07,1.978637e-07,1.978638e-07,1.978640e-07,1.978641e-07,1.978643e-07,1.978644e-07,1.978645e-07,1.978647e-07,1.978648e-07,1.978650e-07,1.978651e-07,1.978652e-07,1.978654e-07,1.978655e-07,1.978657e-07,1.978658e-07,1.978660e-07,1.978661e-07,1.978662e-07,1.978664e-07,1.978665e-07,1.978667e-07,1.978668e-07,1.978669e-07,1.978671e-07,1.978672e-07,1.978674e-07,1.978675e-07,1.978676e-07,1.978678e-07,1.978679e-07,1.978681e-07,1.978682e-07,1.978683e-07,1.978685e-07,1.978686e-07,1.978688e-07,1.978689e-07,1.978690e-07,1.978692e-07,1.978693e-07,1.978695e-07,1.978696e-07,1.978697e-07,1.978699e-07,1.978700e-07,1.978702e-07,1.978703e-07,1.978704e-07,1.978706e-07,1.978707e-07,1.978709e-07,1.978710e-07,1.978711e-07,1.978713e-07,1.978714e-07,1.978716e-07,1.978717e-07,1.978718e-07,1.978720e-07,1.978721e-07,1.978723e-07,1.978724e-07,1.978725e-07,1.978727e-07,1.978728e-07,1.978730e-07,1.978731e-07,1.978732e-07,1.978734e-07,1.978735e-07,1.978737e-07,1.978738e-07,1.978739e-07,1.978741e-07,1.978742e-07,1.978744e-07,1.978745e-07,1.978746e-07,1.978748e-07,1.978749e-07,1.978751e-07,1.978752e-07,1.978753e-07,1.978755e-07,1.978756e-07,1.978758e-07,1.978759e-07,1.978760e-07,1.978762e-07,1.978763e-07,1.978765e-07,1.978766e-07,1.978767e-07,1.978769e-07,1.978770e-07,1.978772e-07,1.978773e-07,1.978774e-07,1.978776e-07,1.978777e-07,1.978779e-07,1.978780e-07,1.978781e-07,1.978783e-07,1.978784e-07,1.978786e-07,1.978787e-07,1.978788e-07,1.978790e-07,1.978791e-07,1.978793e-07,1.978794e-07,1.978795e-07,1.978797e-07,1.978798e-07,1.978800e-07,1.978801e-07,1.978802e-07,1.978804e-07,1.978805e-07,1.978807e-07,1.978808e-07,1.978809e-07,1.978811e-07,1.978812e-07,1.978814e-07,1.978815e-07,1.978816e-07,1.978818e-07,1.978819e-07,1.978821e-07,1.978822e-07,1.978823e-07,1.978825e-07,1.978826e-07,1.978828e-07,1.978829e-07,1.978830e-07,1.978832e-07,1.978833e-07,1.978835e-07,1.978836e-07,1.978837e-07,1.978839e-07,1.978840e-07,1.978842e-07,1.978843e-07,1.978844e-07,1.978846e-07,1.978847e-07,1.978849e-07,1.978850e-07,1.978851e-07,1.978853e-07,1.978854e-07,1.978856e-07,1.978857e-07,1.978858e-07,1.978860e-07,1.978861e-07,1.978863e-07,1.978864e-07,1.978865e-07,1.978867e-07,1.978868e-07,1.978870e-07,1.978871e-07,1.978872e-07,1.978874e-07,1.978875e-07,1.978877e-07,1.978878e-07,1.978879e-07,1.978881e-07,1.978882e-07,1.978884e-07,1.978885e-07,1.978886e-07,1.978888e-07,1.978889e-07,1.978891e-07,1.978892e-07,1.978893e-07,1.978895e-07,1.978896e-07,1.978898e-07,1.978899e-07,1.978900e-07,1.978902e-07,1.978903e-07,1.978905e-07,1.978906e-07,1.978907e-07,1.978909e-07,1.978910e-07,1.978912e-07,1.978913e-07,1.978914e-07,1.978916e-07,1.978917e-07,1.978919e-07,1.978920e-07,1.978921e-07,1.978923e-07,1.978924e-07,1.978926e-07,1.978927e-07,1.978928e-07,1.978930e-07,1.978931e-07,1.978933e-07,1.978934e-07,1.978935e-07,1.978937e-07,1.978938e-07,1.978940e-07,1.978941e-07,1.978942e-07,1.978944e-07,1.978945e-07,1.978947e-07,1.978948e-07,1.978949e-07,1.978951e-07,1.978952e-07,1.978953e-07,1.978955e-07,1.978956e-07,1.978958e-07,1.978959e-07,1.978960e-07,1.978962e-07,1.978963e-07,1.978965e-07,1.978966e-07,1.978967e-07,1.978969e-07,1.978970e-07,1.978972e-07,1.978973e-07,1.978974e-07,1.978976e-07,1.978977e-07,1.978979e-07,1.978980e-07,1.978981e-07,1.978983e-07,1.978984e-07,1.978986e-07,1.978987e-07,1.978988e-07,1.978990e-07,1.978991e-07,1.978993e-07,1.978994e-07,1.978995e-07,1.978997e-07,1.978998e-07,1.979000e-07,1.979001e-07,1.979002e-07,1.979004e-07,1.979005e-07,1.979007e-07,1.979008e-07,1.979009e-07,1.979011e-07,1.979012e-07,1.979014e-07,1.979015e-07,1.979016e-07,1.979018e-07,1.979019e-07,1.979021e-07,1.979022e-07,1.979023e-07,1.979025e-07,1.979026e-07,1.979028e-07,1.979029e-07,1.979030e-07,1.979032e-07,1.979033e-07,1.979035e-07,1.979036e-07,1.979037e-07,1.979039e-07,1.979040e-07,1.979042e-07,1.979043e-07,1.979044e-07,1.979046e-07,1.979047e-07,1.979049e-07,1.979050e-07,1.979051e-07,1.979053e-07,1.979054e-07,1.979056e-07,1.979057e-07,1.979058e-07,1.979060e-07,1.979061e-07,1.979063e-07,1.979064e-07,1.979065e-07,1.979067e-07,1.979068e-07,1.979069e-07,1.979071e-07,1.979072e-07,1.979074e-07,1.979075e-07,1.979076e-07,1.979078e-07,1.979079e-07,1.979081e-07,1.979082e-07,1.979083e-07,1.979085e-07,1.979086e-07,1.979088e-07,1.979089e-07,1.979090e-07,1.979092e-07,1.979093e-07,1.979095e-07,1.979096e-07,1.979097e-07,1.979099e-07,1.979100e-07,1.979102e-07,1.979103e-07,1.979104e-07,1.979106e-07,1.979107e-07,1.979109e-07,1.979110e-07,1.979111e-07,1.979113e-07,1.979114e-07,1.979116e-07,1.979117e-07,1.979118e-07,1.979120e-07,1.979121e-07,1.979123e-07,1.979124e-07,1.979125e-07,1.979127e-07,1.979128e-07,1.979130e-07,1.979131e-07,1.979132e-07,1.979134e-07,1.979135e-07,1.979137e-07,1.979138e-07,1.979139e-07,1.979141e-07,1.979142e-07,1.979143e-07,1.979145e-07,1.979146e-07,1.979148e-07,1.979149e-07,1.979150e-07,1.979152e-07,1.979153e-07,1.979155e-07,1.979156e-07,1.979157e-07,1.979159e-07,1.979160e-07,1.979162e-07,1.979163e-07,1.979164e-07,1.979166e-07,1.979167e-07,1.979169e-07,1.979170e-07,1.979171e-07,1.979173e-07,1.979174e-07,1.979176e-07,1.979177e-07,1.979178e-07,1.979180e-07,1.979181e-07,1.979183e-07,1.979184e-07,1.979185e-07,1.979187e-07,1.979188e-07,1.979190e-07,1.979191e-07,1.979192e-07,1.979194e-07,1.979195e-07,1.979197e-07,1.979198e-07,1.979199e-07,1.979201e-07,1.979202e-07,1.979204e-07,1.979205e-07,1.979206e-07,1.979208e-07,1.979209e-07,1.979210e-07,1.979212e-07,1.979213e-07,1.979215e-07,1.979216e-07,1.979217e-07,1.979219e-07,1.979220e-07,1.979222e-07,1.979223e-07,1.979224e-07,1.979226e-07,1.979227e-07,1.979229e-07,1.979230e-07,1.979231e-07,1.979233e-07,1.979234e-07,1.979236e-07,1.979237e-07,1.979238e-07,1.979240e-07,1.979241e-07,1.979243e-07,1.979244e-07,1.979245e-07,1.979247e-07,1.979248e-07,1.979250e-07,1.979251e-07,1.979252e-07,1.979254e-07,1.979255e-07,1.979257e-07,1.979258e-07,1.979259e-07,1.979261e-07,1.979262e-07,1.979263e-07,1.979265e-07,1.979266e-07,1.979268e-07,1.979269e-07,1.979270e-07,1.979272e-07,1.979273e-07,1.979275e-07,1.979276e-07,1.979277e-07,1.979279e-07,1.979280e-07,1.979282e-07,1.979283e-07,1.979284e-07,1.979286e-07,1.979287e-07,1.979289e-07,1.979290e-07,1.979291e-07,1.979293e-07,1.979294e-07,1.979296e-07,1.979297e-07,1.979298e-07,1.979300e-07,1.979301e-07,1.979303e-07,1.979304e-07,1.979305e-07,1.979307e-07,1.979308e-07,1.979309e-07,1.979311e-07,1.979312e-07,1.979314e-07,1.979315e-07,1.979316e-07,1.979318e-07,1.979319e-07,1.979321e-07,1.979322e-07,1.979323e-07,1.979325e-07,1.979326e-07,1.979328e-07,1.979329e-07,1.979330e-07,1.979332e-07,1.979333e-07,1.979335e-07,1.979336e-07,1.979337e-07,1.979339e-07,1.979340e-07,1.979342e-07,1.979343e-07,1.979344e-07,1.979346e-07,1.979347e-07,1.979349e-07,1.979350e-07,1.979351e-07,1.979353e-07,1.979354e-07,1.979355e-07,1.979357e-07,1.979358e-07,1.979360e-07,1.979361e-07,1.979362e-07,1.979364e-07,1.979365e-07,1.979367e-07,1.979368e-07,1.979369e-07,1.979371e-07,1.979372e-07,1.979374e-07,1.979375e-07,1.979376e-07,1.979378e-07,1.979379e-07,1.979381e-07,1.979382e-07,1.979383e-07,1.979385e-07,1.979386e-07,1.979388e-07,1.979389e-07,1.979390e-07,1.979392e-07,1.979393e-07,1.979394e-07,1.979396e-07,1.979397e-07,1.979399e-07,1.979400e-07,1.979401e-07,1.979403e-07,1.979404e-07,1.979406e-07,1.979407e-07,1.979408e-07,1.979410e-07,1.979411e-07,1.979413e-07,1.979414e-07,1.979415e-07,1.979417e-07,1.979418e-07,1.979420e-07,1.979421e-07,1.979422e-07,1.979424e-07,1.979425e-07,1.979427e-07,1.979428e-07,1.979429e-07,1.979431e-07,1.979432e-07,1.979433e-07,1.979435e-07,1.979436e-07,1.979438e-07,1.979439e-07,1.979440e-07,1.979442e-07,1.979443e-07,1.979445e-07,1.979446e-07,1.979447e-07,1.979449e-07,1.979450e-07,1.979452e-07,1.979453e-07,1.979454e-07,1.979456e-07,1.979457e-07,1.979459e-07,1.979460e-07,1.979461e-07,1.979463e-07,1.979464e-07,1.979466e-07,1.979467e-07,1.979468e-07,1.979470e-07,1.979471e-07,1.979472e-07,1.979474e-07,1.979475e-07,1.979477e-07,1.979478e-07,1.979479e-07,1.979481e-07,1.979482e-07,1.979484e-07,1.979485e-07,1.979486e-07,1.979488e-07,1.979489e-07,1.979491e-07,1.979492e-07,1.979493e-07,1.979495e-07,1.979496e-07,1.979498e-07,1.979499e-07,1.979500e-07,1.979502e-07,1.979503e-07,1.979504e-07,1.979506e-07,1.979507e-07,1.979509e-07,1.979510e-07,1.979511e-07,1.979513e-07,1.979514e-07,1.979516e-07,1.979517e-07,1.979518e-07,1.979520e-07,1.979521e-07,1.979523e-07,1.979524e-07,1.979525e-07,1.979527e-07,1.979528e-07,1.979530e-07,1.979531e-07,1.979532e-07,1.979534e-07,1.979535e-07,1.979536e-07,1.979538e-07,1.979539e-07,1.979541e-07,1.979542e-07,1.979543e-07,1.979545e-07,1.979546e-07,1.979548e-07,1.979549e-07,1.979550e-07,1.979552e-07,1.979553e-07,1.979555e-07,1.979556e-07,1.979557e-07,1.979559e-07,1.979560e-07,1.979562e-07,1.979563e-07,1.979564e-07,1.979566e-07,1.979567e-07,1.979568e-07,1.979570e-07,1.979571e-07,1.979573e-07,1.979574e-07,1.979575e-07,1.979577e-07,1.979578e-07,1.979580e-07,1.979581e-07,1.979582e-07,1.979584e-07,1.979585e-07,1.979587e-07,1.979588e-07,1.979589e-07,1.979591e-07,1.979592e-07,1.979594e-07,1.979595e-07,1.979596e-07,1.979598e-07,1.979599e-07,1.979600e-07,1.979602e-07,1.979603e-07,1.979605e-07,1.979606e-07,1.979607e-07,1.979609e-07,1.979610e-07,1.979612e-07,1.979613e-07,1.979614e-07,1.979616e-07,1.979617e-07,1.979619e-07,1.979620e-07,1.979621e-07,1.979623e-07,1.979624e-07,1.979625e-07,1.979627e-07,1.979628e-07,1.979630e-07,1.979631e-07,1.979632e-07,1.979634e-07,1.979635e-07,1.979637e-07,1.979638e-07,1.979639e-07,1.979641e-07,1.979642e-07,1.979644e-07,1.979645e-07,1.979646e-07,1.979648e-07,1.979649e-07,1.979651e-07,1.979652e-07,1.979653e-07,1.979655e-07,1.979656e-07,1.979657e-07,1.979659e-07,1.979660e-07,1.979662e-07,1.979663e-07,1.979664e-07,1.979666e-07,1.979667e-07,1.979669e-07,1.979670e-07,1.979671e-07,1.979673e-07,1.979674e-07,1.979676e-07,1.979677e-07,1.979678e-07,1.979680e-07,1.979681e-07,1.979682e-07,1.979684e-07,1.979685e-07,1.979687e-07,1.979688e-07,1.979689e-07,1.979691e-07,1.979692e-07,1.979694e-07,1.979695e-07,1.979696e-07,1.979698e-07,1.979699e-07,1.979701e-07,1.979702e-07,1.979703e-07,1.979705e-07,1.979706e-07,1.979707e-07,1.979709e-07,1.979710e-07,1.979712e-07,1.979713e-07,1.979714e-07,1.979716e-07,1.979717e-07,1.979719e-07,1.979720e-07,1.979721e-07,1.979723e-07,1.979724e-07,1.979726e-07,1.979727e-07,1.979728e-07,1.979730e-07,1.979731e-07,1.979732e-07,1.979734e-07,1.979735e-07,1.979737e-07,1.979738e-07,1.979739e-07,1.979741e-07,1.979742e-07,1.979744e-07,1.979745e-07,1.979746e-07,1.979748e-07,1.979749e-07,1.979751e-07,1.979752e-07,1.979753e-07,1.979755e-07,1.979756e-07,1.979757e-07,1.979759e-07,1.979760e-07,1.979762e-07,1.979763e-07,1.979764e-07,1.979766e-07,1.979767e-07,1.979769e-07,1.979770e-07,1.979771e-07,1.979773e-07,1.979774e-07,1.979776e-07,1.979777e-07,1.979778e-07,1.979780e-07,1.979781e-07,1.979782e-07,1.979784e-07,1.979785e-07,1.979787e-07,1.979788e-07,1.979789e-07,1.979791e-07,1.979792e-07,1.979794e-07,1.979795e-07,1.979796e-07,1.979798e-07,1.979799e-07,1.979801e-07,1.979802e-07,1.979803e-07,1.979805e-07,1.979806e-07,1.979807e-07,1.979809e-07,1.979810e-07,1.979812e-07,1.979813e-07,1.979814e-07,1.979816e-07,1.979817e-07,1.979819e-07,1.979820e-07,1.979821e-07,1.979823e-07,1.979824e-07,1.979826e-07,1.979827e-07,1.979828e-07,1.979830e-07,1.979831e-07,1.979832e-07,1.979834e-07,1.979835e-07,1.979837e-07,1.979838e-07,1.979839e-07,1.979841e-07,1.979842e-07,1.979844e-07,1.979845e-07,1.979846e-07,1.979848e-07,1.979849e-07,1.979850e-07,1.979852e-07,1.979853e-07,1.979855e-07,1.979856e-07,1.979857e-07,1.979859e-07,1.979860e-07,1.979862e-07,1.979863e-07,1.979864e-07,1.979866e-07,1.979867e-07,1.979869e-07,1.979870e-07,1.979871e-07,1.979873e-07,1.979874e-07,1.979875e-07,1.979877e-07,1.979878e-07,1.979880e-07,1.979881e-07,1.979882e-07,1.979884e-07,1.979885e-07,1.979887e-07,1.979888e-07,1.979889e-07,1.979891e-07,1.979892e-07,1.979893e-07,1.979895e-07,1.979896e-07,1.979898e-07,1.979899e-07,1.979900e-07,1.979902e-07,1.979903e-07,1.979905e-07,1.979906e-07,1.979907e-07,1.979909e-07,1.979910e-07,1.979912e-07,1.979913e-07,1.979914e-07,1.979916e-07,1.979917e-07,1.979918e-07,1.979920e-07,1.979921e-07,1.979923e-07,1.979924e-07,1.979925e-07,1.979927e-07,1.979928e-07,1.979930e-07,1.979931e-07,1.979932e-07,1.979934e-07,1.979935e-07,1.979936e-07,1.979938e-07,1.979939e-07,1.979941e-07,1.979942e-07,1.979943e-07,1.979945e-07,1.979946e-07,1.979948e-07,1.979949e-07,1.979950e-07,1.979952e-07,1.979953e-07,1.979955e-07,1.979956e-07,1.979957e-07,1.979959e-07,1.979960e-07,1.979961e-07,1.979963e-07,1.979964e-07,1.979966e-07,1.979967e-07,1.979968e-07,1.979970e-07,1.979971e-07,1.979973e-07,1.979974e-07,1.979975e-07,1.979977e-07,1.979978e-07,1.979979e-07,1.979981e-07,1.979982e-07,1.979984e-07,1.979985e-07,1.979986e-07,1.979988e-07,1.979989e-07,1.979991e-07,1.979992e-07,1.979993e-07,1.979995e-07,1.979996e-07,1.979997e-07,1.979999e-07,1.980000e-07,1.980002e-07,1.980003e-07,1.980004e-07,1.980006e-07,1.980007e-07,1.980009e-07,1.980010e-07,1.980011e-07,1.980013e-07,1.980014e-07,1.980015e-07,1.980017e-07,1.980018e-07,1.980020e-07,1.980021e-07,1.980022e-07,1.980024e-07,1.980025e-07,1.980027e-07,1.980028e-07,1.980029e-07,1.980031e-07,1.980032e-07,1.980033e-07,1.980035e-07,1.980036e-07,1.980038e-07,1.980039e-07,1.980040e-07,1.980042e-07,1.980043e-07,1.980045e-07,1.980046e-07,1.980047e-07,1.980049e-07,1.980050e-07,1.980052e-07,1.980053e-07,1.980054e-07,1.980056e-07,1.980057e-07,1.980058e-07,1.980060e-07,1.980061e-07,1.980063e-07,1.980064e-07,1.980065e-07,1.980067e-07,1.980068e-07,1.980070e-07,1.980071e-07,1.980072e-07,1.980074e-07,1.980075e-07,1.980076e-07,1.980078e-07,1.980079e-07,1.980081e-07,1.980082e-07,1.980083e-07,1.980085e-07,1.980086e-07,1.980088e-07,1.980089e-07,1.980090e-07,1.980092e-07,1.980093e-07,1.980094e-07,1.980096e-07,1.980097e-07,1.980099e-07,1.980100e-07,1.980101e-07,1.980103e-07,1.980104e-07,1.980106e-07,1.980107e-07,1.980108e-07,1.980110e-07,1.980111e-07,1.980112e-07,1.980114e-07,1.980115e-07,1.980117e-07,1.980118e-07,1.980119e-07,1.980121e-07,1.980122e-07,1.980124e-07,1.980125e-07,1.980126e-07,1.980128e-07,1.980129e-07,1.980130e-07,1.980132e-07,1.980133e-07,1.980135e-07,1.980136e-07,1.980137e-07,1.980139e-07,1.980140e-07,1.980142e-07,1.980143e-07,1.980144e-07,1.980146e-07,1.980147e-07,1.980148e-07,1.980150e-07,1.980151e-07,1.980153e-07,1.980154e-07,1.980155e-07,1.980157e-07,1.980158e-07,1.980159e-07,1.980161e-07,1.980162e-07,1.980164e-07,1.980165e-07,1.980166e-07,1.980168e-07,1.980169e-07,1.980171e-07,1.980172e-07,1.980173e-07,1.980175e-07,1.980176e-07,1.980177e-07,1.980179e-07,1.980180e-07,1.980182e-07,1.980183e-07,1.980184e-07,1.980186e-07,1.980187e-07,1.980189e-07,1.980190e-07,1.980191e-07,1.980193e-07,1.980194e-07,1.980195e-07,1.980197e-07,1.980198e-07,1.980200e-07,1.980201e-07,1.980202e-07,1.980204e-07,1.980205e-07,1.980207e-07,1.980208e-07,1.980209e-07,1.980211e-07,1.980212e-07,1.980213e-07,1.980215e-07,1.980216e-07,1.980218e-07,1.980219e-07,1.980220e-07,1.980222e-07,1.980223e-07,1.980225e-07,1.980226e-07,1.980227e-07,1.980229e-07,1.980230e-07,1.980231e-07,1.980233e-07,1.980234e-07,1.980236e-07,1.980237e-07,1.980238e-07,1.980240e-07,1.980241e-07,1.980243e-07,1.980244e-07,1.980245e-07,1.980247e-07,1.980248e-07,1.980249e-07,1.980251e-07,1.980252e-07,1.980254e-07,1.980255e-07,1.980256e-07,1.980258e-07,1.980259e-07,1.980260e-07,1.980262e-07,1.980263e-07,1.980265e-07,1.980266e-07,1.980267e-07,1.980269e-07,1.980270e-07,1.980272e-07,1.980273e-07,1.980274e-07,1.980276e-07,1.980277e-07,1.980278e-07,1.980280e-07,1.980281e-07,1.980283e-07,1.980284e-07,1.980285e-07,1.980287e-07,1.980288e-07,1.980290e-07,1.980291e-07,1.980292e-07,1.980294e-07,1.980295e-07,1.980296e-07,1.980298e-07,1.980299e-07,1.980301e-07,1.980302e-07,1.980303e-07,1.980305e-07,1.980306e-07,1.980307e-07,1.980309e-07,1.980310e-07,1.980312e-07,1.980313e-07,1.980314e-07,1.980316e-07,1.980317e-07,1.980319e-07,1.980320e-07,1.980321e-07,1.980323e-07,1.980324e-07,1.980325e-07,1.980327e-07,1.980328e-07,1.980330e-07,1.980331e-07,1.980332e-07,1.980334e-07,1.980335e-07,1.980337e-07,1.980338e-07,1.980339e-07,1.980341e-07,1.980342e-07,1.980343e-07,1.980345e-07,1.980346e-07,1.980348e-07,1.980349e-07,1.980350e-07,1.980352e-07,1.980353e-07,1.980354e-07,1.980356e-07,1.980357e-07,1.980359e-07,1.980360e-07,1.980361e-07,1.980363e-07,1.980364e-07,1.980366e-07,1.980367e-07,1.980368e-07,1.980370e-07,1.980371e-07,1.980372e-07,1.980374e-07,1.980375e-07,1.980377e-07,1.980378e-07,1.980379e-07,1.980381e-07,1.980382e-07,1.980383e-07,1.980385e-07,1.980386e-07,1.980388e-07,1.980389e-07,1.980390e-07,1.980392e-07,1.980393e-07,1.980395e-07,1.980396e-07,1.980397e-07,1.980399e-07,1.980400e-07,1.980401e-07,1.980403e-07,1.980404e-07,1.980406e-07,1.980407e-07,1.980408e-07,1.980410e-07,1.980411e-07,1.980412e-07,1.980414e-07,1.980415e-07,1.980417e-07,1.980418e-07,1.980419e-07,1.980421e-07,1.980422e-07,1.980424e-07,1.980425e-07,1.980426e-07,1.980428e-07,1.980429e-07,1.980430e-07,1.980432e-07,1.980433e-07,1.980435e-07,1.980436e-07,1.980437e-07,1.980439e-07,1.980440e-07,1.980441e-07,1.980443e-07,1.980444e-07,1.980446e-07,1.980447e-07,1.980448e-07,1.980450e-07,1.980451e-07,1.980453e-07,1.980454e-07,1.980455e-07,1.980457e-07,1.980458e-07,1.980459e-07,1.980461e-07,1.980462e-07,1.980464e-07,1.980465e-07,1.980466e-07,1.980468e-07,1.980469e-07,1.980470e-07,1.980472e-07,1.980473e-07,1.980475e-07,1.980476e-07,1.980477e-07,1.980479e-07,1.980480e-07,1.980481e-07,1.980483e-07,1.980484e-07,1.980486e-07,1.980487e-07,1.980488e-07,1.980490e-07,1.980491e-07,1.980493e-07,1.980494e-07,1.980495e-07,1.980497e-07,1.980498e-07,1.980499e-07,1.980501e-07,1.980502e-07,1.980504e-07,1.980505e-07,1.980506e-07,1.980508e-07,1.980509e-07,1.980510e-07,1.980512e-07,1.980513e-07,1.980515e-07,1.980516e-07,1.980517e-07,1.980519e-07,1.980520e-07,1.980522e-07,1.980523e-07,1.980524e-07,1.980526e-07,1.980527e-07,1.980528e-07,1.980530e-07,1.980531e-07,1.980533e-07,1.980534e-07,1.980535e-07,1.980537e-07,1.980538e-07,1.980539e-07,1.980541e-07,1.980542e-07,1.980544e-07,1.980545e-07,1.980546e-07,1.980548e-07,1.980549e-07,1.980550e-07,1.980552e-07,1.980553e-07,1.980555e-07,1.980556e-07,1.980557e-07,1.980559e-07,1.980560e-07,1.980562e-07,1.980563e-07,1.980564e-07,1.980566e-07,1.980567e-07,1.980568e-07,1.980570e-07,1.980571e-07,1.980573e-07,1.980574e-07,1.980575e-07,1.980577e-07,1.980578e-07,1.980579e-07,1.980581e-07,1.980582e-07,1.980584e-07,1.980585e-07,1.980586e-07,1.980588e-07,1.980589e-07,1.980590e-07,1.980592e-07,1.980593e-07,1.980595e-07,1.980596e-07,1.980597e-07,1.980599e-07,1.980600e-07,1.980602e-07,1.980603e-07,1.980604e-07,1.980606e-07,1.980607e-07,1.980608e-07,1.980610e-07,1.980611e-07,1.980613e-07,1.980614e-07,1.980615e-07,1.980617e-07,1.980618e-07,1.980619e-07,1.980621e-07,1.980622e-07,1.980624e-07,1.980625e-07,1.980626e-07,1.980628e-07,1.980629e-07,1.980630e-07,1.980632e-07,1.980633e-07,1.980635e-07,1.980636e-07,1.980637e-07,1.980639e-07,1.980640e-07,1.980641e-07,1.980643e-07,1.980644e-07,1.980646e-07,1.980647e-07,1.980648e-07,1.980650e-07,1.980651e-07,1.980653e-07,1.980654e-07,1.980655e-07,1.980657e-07,1.980658e-07,1.980659e-07,1.980661e-07,1.980662e-07,1.980664e-07,1.980665e-07,1.980666e-07,1.980668e-07,1.980669e-07,1.980670e-07,1.980672e-07,1.980673e-07,1.980675e-07,1.980676e-07,1.980677e-07,1.980679e-07,1.980680e-07,1.980681e-07,1.980683e-07,1.980684e-07,1.980686e-07,1.980687e-07,1.980688e-07,1.980690e-07,1.980691e-07,1.980692e-07,1.980694e-07,1.980695e-07,1.980697e-07,1.980698e-07,1.980699e-07,1.980701e-07,1.980702e-07,1.980703e-07,1.980705e-07,1.980706e-07,1.980708e-07,1.980709e-07,1.980710e-07,1.980712e-07,1.980713e-07,1.980714e-07,1.980716e-07,1.980717e-07,1.980719e-07,1.980720e-07,1.980721e-07,1.980723e-07,1.980724e-07,1.980726e-07,1.980727e-07,1.980728e-07,1.980730e-07,1.980731e-07,1.980732e-07,1.980734e-07,1.980735e-07,1.980737e-07,1.980738e-07,1.980739e-07,1.980741e-07,1.980742e-07,1.980743e-07,1.980745e-07,1.980746e-07,1.980748e-07,1.980749e-07,1.980750e-07,1.980752e-07,1.980753e-07,1.980754e-07,1.980756e-07,1.980757e-07,1.980759e-07,1.980760e-07,1.980761e-07,1.980763e-07,1.980764e-07,1.980765e-07,1.980767e-07,1.980768e-07,1.980770e-07,1.980771e-07,1.980772e-07,1.980774e-07,1.980775e-07,1.980776e-07,1.980778e-07,1.980779e-07,1.980781e-07,1.980782e-07,1.980783e-07,1.980785e-07,1.980786e-07,1.980787e-07,1.980789e-07,1.980790e-07,1.980792e-07,1.980793e-07,1.980794e-07,1.980796e-07,1.980797e-07,1.980798e-07,1.980800e-07,1.980801e-07,1.980803e-07,1.980804e-07,1.980805e-07,1.980807e-07,1.980808e-07,1.980809e-07,1.980811e-07,1.980812e-07,1.980814e-07,1.980815e-07,1.980816e-07,1.980818e-07,1.980819e-07,1.980821e-07,1.980822e-07,1.980823e-07,1.980825e-07,1.980826e-07,1.980827e-07,1.980829e-07,1.980830e-07,1.980832e-07,1.980833e-07,1.980834e-07,1.980836e-07,1.980837e-07,1.980838e-07,1.980840e-07,1.980841e-07,1.980843e-07,1.980844e-07,1.980845e-07,1.980847e-07,1.980848e-07,1.980849e-07,1.980851e-07,1.980852e-07,1.980854e-07,1.980855e-07,1.980856e-07,1.980858e-07,1.980859e-07,1.980860e-07,1.980862e-07,1.980863e-07,1.980865e-07,1.980866e-07,1.980867e-07,1.980869e-07,1.980870e-07,1.980871e-07,1.980873e-07,1.980874e-07,1.980876e-07,1.980877e-07,1.980878e-07,1.980880e-07,1.980881e-07,1.980882e-07,1.980884e-07,1.980885e-07,1.980887e-07,1.980888e-07,1.980889e-07,1.980891e-07,1.980892e-07,1.980893e-07,1.980895e-07,1.980896e-07,1.980898e-07,1.980899e-07,1.980900e-07,1.980902e-07,1.980903e-07,1.980904e-07,1.980906e-07,1.980907e-07,1.980909e-07,1.980910e-07,1.980911e-07,1.980913e-07,1.980914e-07,1.980915e-07,1.980917e-07,1.980918e-07,1.980920e-07,1.980921e-07,1.980922e-07,1.980924e-07,1.980925e-07,1.980926e-07,1.980928e-07,1.980929e-07,1.980931e-07,1.980932e-07,1.980933e-07,1.980935e-07,1.980936e-07,1.980937e-07,1.980939e-07,1.980940e-07,1.980942e-07,1.980943e-07,1.980944e-07,1.980946e-07,1.980947e-07,1.980948e-07,1.980950e-07,1.980951e-07,1.980953e-07,1.980954e-07,1.980955e-07,1.980957e-07,1.980958e-07,1.980959e-07,1.980961e-07,1.980962e-07,1.980964e-07,1.980965e-07,1.980966e-07,1.980968e-07,1.980969e-07,1.980970e-07,1.980972e-07,1.980973e-07,1.980975e-07,1.980976e-07,1.980977e-07,1.980979e-07,1.980980e-07,1.980981e-07,1.980983e-07,1.980984e-07,1.980986e-07,1.980987e-07,1.980988e-07,1.980990e-07,1.980991e-07,1.980992e-07,1.980994e-07,1.980995e-07,1.980997e-07,1.980998e-07,1.980999e-07,1.981001e-07,1.981002e-07,1.981003e-07,1.981005e-07,1.981006e-07,1.981008e-07,1.981009e-07,1.981010e-07,1.981012e-07,1.981013e-07,1.981014e-07,1.981016e-07,1.981017e-07,1.981018e-07,1.981020e-07,1.981021e-07,1.981023e-07,1.981024e-07,1.981025e-07,1.981027e-07,1.981028e-07,1.981029e-07,1.981031e-07,1.981032e-07,1.981034e-07,1.981035e-07,1.981036e-07,1.981038e-07,1.981039e-07,1.981040e-07,1.981042e-07,1.981043e-07,1.981045e-07,1.981046e-07,1.981047e-07,1.981049e-07,1.981050e-07,1.981051e-07,1.981053e-07,1.981054e-07,1.981056e-07,1.981057e-07,1.981058e-07,1.981060e-07,1.981061e-07,1.981062e-07,1.981064e-07,1.981065e-07,1.981067e-07,1.981068e-07,1.981069e-07,1.981071e-07,1.981072e-07,1.981073e-07,1.981075e-07,1.981076e-07,1.981078e-07,1.981079e-07,1.981080e-07,1.981082e-07,1.981083e-07,1.981084e-07,1.981086e-07,1.981087e-07,1.981089e-07,1.981090e-07,1.981091e-07,1.981093e-07,1.981094e-07,1.981095e-07,1.981097e-07,1.981098e-07,1.981100e-07,1.981101e-07,1.981102e-07,1.981104e-07,1.981105e-07,1.981106e-07,1.981108e-07,1.981109e-07,1.981111e-07,1.981112e-07,1.981113e-07,1.981115e-07,1.981116e-07,1.981117e-07,1.981119e-07,1.981120e-07,1.981121e-07,1.981123e-07,1.981124e-07,1.981126e-07,1.981127e-07,1.981128e-07,1.981130e-07,1.981131e-07,1.981132e-07,1.981134e-07,1.981135e-07,1.981137e-07,1.981138e-07,1.981139e-07,1.981141e-07,1.981142e-07,1.981143e-07,1.981145e-07,1.981146e-07,1.981148e-07,1.981149e-07,1.981150e-07,1.981152e-07,1.981153e-07,1.981154e-07,1.981156e-07,1.981157e-07,1.981159e-07,1.981160e-07,1.981161e-07,1.981163e-07,1.981164e-07,1.981165e-07,1.981167e-07,1.981168e-07,1.981170e-07,1.981171e-07,1.981172e-07,1.981174e-07,1.981175e-07,1.981176e-07,1.981178e-07,1.981179e-07,1.981180e-07,1.981182e-07,1.981183e-07,1.981185e-07,1.981186e-07,1.981187e-07,1.981189e-07,1.981190e-07,1.981191e-07,1.981193e-07,1.981194e-07,1.981196e-07,1.981197e-07,1.981198e-07,1.981200e-07,1.981201e-07,1.981202e-07,1.981204e-07,1.981205e-07,1.981207e-07,1.981208e-07,1.981209e-07,1.981211e-07,1.981212e-07,1.981213e-07,1.981215e-07,1.981216e-07,1.981218e-07,1.981219e-07,1.981220e-07,1.981222e-07,1.981223e-07,1.981224e-07,1.981226e-07,1.981227e-07,1.981228e-07,1.981230e-07,1.981231e-07,1.981233e-07,1.981234e-07,1.981235e-07,1.981237e-07,1.981238e-07,1.981239e-07,1.981241e-07,1.981242e-07,1.981244e-07,1.981245e-07,1.981246e-07,1.981248e-07,1.981249e-07,1.981250e-07,1.981252e-07,1.981253e-07,1.981255e-07,1.981256e-07,1.981257e-07,1.981259e-07,1.981260e-07,1.981261e-07,1.981263e-07,1.981264e-07,1.981266e-07,1.981267e-07,1.981268e-07,1.981270e-07,1.981271e-07,1.981272e-07,1.981274e-07,1.981275e-07,1.981276e-07,1.981278e-07,1.981279e-07,1.981281e-07,1.981282e-07,1.981283e-07,1.981285e-07,1.981286e-07,1.981287e-07,1.981289e-07,1.981290e-07,1.981292e-07,1.981293e-07,1.981294e-07,1.981296e-07,1.981297e-07,1.981298e-07,1.981300e-07,1.981301e-07,1.981303e-07,1.981304e-07,1.981305e-07,1.981307e-07,1.981308e-07,1.981309e-07,1.981311e-07,1.981312e-07,1.981313e-07,1.981315e-07,1.981316e-07,1.981318e-07,1.981319e-07,1.981320e-07,1.981322e-07,1.981323e-07,1.981324e-07,1.981326e-07,1.981327e-07,1.981329e-07,1.981330e-07,1.981331e-07,1.981333e-07,1.981334e-07,1.981335e-07,1.981337e-07,1.981338e-07,1.981340e-07,1.981341e-07,1.981342e-07,1.981344e-07,1.981345e-07,1.981346e-07,1.981348e-07,1.981349e-07,1.981350e-07,1.981352e-07,1.981353e-07,1.981355e-07,1.981356e-07,1.981357e-07,1.981359e-07,1.981360e-07,1.981361e-07,1.981363e-07,1.981364e-07,1.981366e-07,1.981367e-07,1.981368e-07,1.981370e-07,1.981371e-07,1.981372e-07,1.981374e-07,1.981375e-07,1.981377e-07,1.981378e-07,1.981379e-07,1.981381e-07,1.981382e-07,1.981383e-07,1.981385e-07,1.981386e-07,1.981387e-07,1.981389e-07,1.981390e-07,1.981392e-07,1.981393e-07,1.981394e-07,1.981396e-07,1.981397e-07,1.981398e-07,1.981400e-07,1.981401e-07,1.981403e-07,1.981404e-07,1.981405e-07,1.981407e-07,1.981408e-07,1.981409e-07,1.981411e-07,1.981412e-07,1.981413e-07,1.981415e-07,1.981416e-07,1.981418e-07,1.981419e-07,1.981420e-07,1.981422e-07,1.981423e-07,1.981424e-07,1.981426e-07,1.981427e-07,1.981429e-07,1.981430e-07,1.981431e-07,1.981433e-07,1.981434e-07,1.981435e-07,1.981437e-07,1.981438e-07,1.981439e-07,1.981441e-07,1.981442e-07,1.981444e-07,1.981445e-07,1.981446e-07,1.981448e-07,1.981449e-07,1.981450e-07,1.981452e-07,1.981453e-07,1.981455e-07,1.981456e-07,1.981457e-07,1.981459e-07,1.981460e-07,1.981461e-07,1.981463e-07,1.981464e-07,1.981465e-07,1.981467e-07,1.981468e-07,1.981470e-07,1.981471e-07,1.981472e-07,1.981474e-07,1.981475e-07,1.981476e-07,1.981478e-07,1.981479e-07,1.981481e-07,1.981482e-07,1.981483e-07,1.981485e-07,1.981486e-07,1.981487e-07,1.981489e-07,1.981490e-07,1.981491e-07,1.981493e-07,1.981494e-07,1.981496e-07,1.981497e-07,1.981498e-07,1.981500e-07,1.981501e-07,1.981502e-07,1.981504e-07,1.981505e-07,1.981507e-07,1.981508e-07,1.981509e-07,1.981511e-07,1.981512e-07,1.981513e-07,1.981515e-07,1.981516e-07,1.981517e-07,1.981519e-07,1.981520e-07,1.981522e-07,1.981523e-07,1.981524e-07,1.981526e-07,1.981527e-07,1.981528e-07,1.981530e-07,1.981531e-07,1.981533e-07,1.981534e-07,1.981535e-07,1.981537e-07,1.981538e-07,1.981539e-07,1.981541e-07,1.981542e-07,1.981543e-07,1.981545e-07,1.981546e-07,1.981548e-07,1.981549e-07,1.981550e-07,1.981552e-07,1.981553e-07,1.981554e-07,1.981556e-07,1.981557e-07,1.981559e-07,1.981560e-07,1.981561e-07,1.981563e-07,1.981564e-07,1.981565e-07,1.981567e-07,1.981568e-07,1.981569e-07,1.981571e-07,1.981572e-07,1.981574e-07,1.981575e-07,1.981576e-07,1.981578e-07,1.981579e-07,1.981580e-07,1.981582e-07,1.981583e-07,1.981584e-07,1.981586e-07,1.981587e-07,1.981589e-07,1.981590e-07,1.981591e-07,1.981593e-07,1.981594e-07,1.981595e-07,1.981597e-07,1.981598e-07,1.981600e-07,1.981601e-07,1.981602e-07,1.981604e-07,1.981605e-07,1.981606e-07,1.981608e-07,1.981609e-07,1.981610e-07,1.981612e-07,1.981613e-07,1.981615e-07,1.981616e-07,1.981617e-07,1.981619e-07,1.981620e-07,1.981621e-07,1.981623e-07,1.981624e-07,1.981625e-07,1.981627e-07,1.981628e-07,1.981630e-07,1.981631e-07,1.981632e-07,1.981634e-07,1.981635e-07,1.981636e-07,1.981638e-07,1.981639e-07,1.981641e-07,1.981642e-07,1.981643e-07,1.981645e-07,1.981646e-07,1.981647e-07,1.981649e-07,1.981650e-07,1.981651e-07,1.981653e-07,1.981654e-07,1.981656e-07,1.981657e-07,1.981658e-07,1.981660e-07,1.981661e-07,1.981662e-07,1.981664e-07,1.981665e-07,1.981666e-07,1.981668e-07,1.981669e-07,1.981671e-07,1.981672e-07,1.981673e-07,1.981675e-07,1.981676e-07,1.981677e-07,1.981679e-07,1.981680e-07,1.981682e-07,1.981683e-07,1.981684e-07,1.981686e-07,1.981687e-07,1.981688e-07,1.981690e-07,1.981691e-07,1.981692e-07,1.981694e-07,1.981695e-07,1.981697e-07,1.981698e-07,1.981699e-07,1.981701e-07,1.981702e-07,1.981703e-07,1.981705e-07,1.981706e-07,1.981707e-07,1.981709e-07,1.981710e-07,1.981712e-07,1.981713e-07,1.981714e-07,1.981716e-07,1.981717e-07,1.981718e-07,1.981720e-07,1.981721e-07,1.981722e-07,1.981724e-07,1.981725e-07,1.981727e-07,1.981728e-07,1.981729e-07,1.981731e-07,1.981732e-07,1.981733e-07,1.981735e-07,1.981736e-07,1.981738e-07,1.981739e-07,1.981740e-07,1.981742e-07,1.981743e-07,1.981744e-07,1.981746e-07,1.981747e-07,1.981748e-07,1.981750e-07,1.981751e-07,1.981753e-07,1.981754e-07,1.981755e-07,1.981757e-07,1.981758e-07,1.981759e-07,1.981761e-07,1.981762e-07,1.981763e-07,1.981765e-07,1.981766e-07,1.981768e-07,1.981769e-07,1.981770e-07,1.981772e-07,1.981773e-07,1.981774e-07,1.981776e-07,1.981777e-07,1.981778e-07,1.981780e-07,1.981781e-07,1.981783e-07,1.981784e-07,1.981785e-07,1.981787e-07,1.981788e-07,1.981789e-07,1.981791e-07,1.981792e-07,1.981793e-07,1.981795e-07,1.981796e-07,1.981798e-07,1.981799e-07,1.981800e-07,1.981802e-07,1.981803e-07,1.981804e-07,1.981806e-07,1.981807e-07,1.981808e-07,1.981810e-07,1.981811e-07,1.981813e-07,1.981814e-07,1.981815e-07,1.981817e-07,1.981818e-07,1.981819e-07,1.981821e-07,1.981822e-07,1.981823e-07,1.981825e-07,1.981826e-07,1.981828e-07,1.981829e-07,1.981830e-07,1.981832e-07,1.981833e-07,1.981834e-07,1.981836e-07,1.981837e-07,1.981839e-07,1.981840e-07,1.981841e-07,1.981843e-07,1.981844e-07,1.981845e-07,1.981847e-07,1.981848e-07,1.981849e-07,1.981851e-07,1.981852e-07,1.981854e-07,1.981855e-07,1.981856e-07,1.981858e-07,1.981859e-07,1.981860e-07,1.981862e-07,1.981863e-07,1.981864e-07,1.981866e-07,1.981867e-07,1.981869e-07,1.981870e-07,1.981871e-07,1.981873e-07,1.981874e-07,1.981875e-07,1.981877e-07,1.981878e-07,1.981879e-07,1.981881e-07,1.981882e-07,1.981884e-07,1.981885e-07,1.981886e-07,1.981888e-07,1.981889e-07,1.981890e-07,1.981892e-07,1.981893e-07,1.981894e-07,1.981896e-07,1.981897e-07,1.981899e-07,1.981900e-07,1.981901e-07,1.981903e-07,1.981904e-07,1.981905e-07,1.981907e-07,1.981908e-07,1.981909e-07,1.981911e-07,1.981912e-07,1.981914e-07,1.981915e-07,1.981916e-07,1.981918e-07,1.981919e-07,1.981920e-07,1.981922e-07,1.981923e-07,1.981924e-07,1.981926e-07,1.981927e-07,1.981929e-07,1.981930e-07,1.981931e-07,1.981933e-07,1.981934e-07,1.981935e-07,1.981937e-07,1.981938e-07,1.981939e-07,1.981941e-07,1.981942e-07,1.981944e-07,1.981945e-07,1.981946e-07,1.981948e-07,1.981949e-07,1.981950e-07,1.981952e-07,1.981953e-07,1.981954e-07,1.981956e-07,1.981957e-07,1.981958e-07,1.981960e-07,1.981961e-07,1.981963e-07,1.981964e-07,1.981965e-07,1.981967e-07,1.981968e-07,1.981969e-07,1.981971e-07,1.981972e-07,1.981973e-07,1.981975e-07,1.981976e-07,1.981978e-07,1.981979e-07,1.981980e-07,1.981982e-07,1.981983e-07,1.981984e-07,1.981986e-07,1.981987e-07,1.981988e-07,1.981990e-07,1.981991e-07,1.981993e-07,1.981994e-07,1.981995e-07,1.981997e-07,1.981998e-07,1.981999e-07,1.982001e-07,1.982002e-07,1.982003e-07,1.982005e-07,1.982006e-07,1.982008e-07,1.982009e-07,1.982010e-07,1.982012e-07,1.982013e-07,1.982014e-07,1.982016e-07,1.982017e-07,1.982018e-07,1.982020e-07,1.982021e-07,1.982023e-07,1.982024e-07,1.982025e-07,1.982027e-07,1.982028e-07,1.982029e-07,1.982031e-07,1.982032e-07,1.982033e-07,1.982035e-07,1.982036e-07,1.982038e-07,1.982039e-07,1.982040e-07,1.982042e-07,1.982043e-07,1.982044e-07,1.982046e-07,1.982047e-07,1.982048e-07,1.982050e-07,1.982051e-07,1.982052e-07,1.982054e-07,1.982055e-07,1.982057e-07,1.982058e-07,1.982059e-07,1.982061e-07,1.982062e-07,1.982063e-07,1.982065e-07,1.982066e-07,1.982067e-07,1.982069e-07,1.982070e-07,1.982072e-07,1.982073e-07,1.982074e-07,1.982076e-07,1.982077e-07,1.982078e-07,1.982080e-07,1.982081e-07,1.982082e-07,1.982084e-07,1.982085e-07,1.982087e-07,1.982088e-07,1.982089e-07,1.982091e-07,1.982092e-07,1.982093e-07,1.982095e-07,1.982096e-07,1.982097e-07,1.982099e-07,1.982100e-07,1.982101e-07,1.982103e-07,1.982104e-07,1.982106e-07,1.982107e-07,1.982108e-07,1.982110e-07,1.982111e-07,1.982112e-07,1.982114e-07,1.982115e-07,1.982116e-07,1.982118e-07,1.982119e-07,1.982121e-07,1.982122e-07,1.982123e-07,1.982125e-07,1.982126e-07,1.982127e-07,1.982129e-07,1.982130e-07,1.982131e-07,1.982133e-07,1.982134e-07,1.982136e-07,1.982137e-07,1.982138e-07,1.982140e-07,1.982141e-07,1.982142e-07,1.982144e-07,1.982145e-07,1.982146e-07,1.982148e-07,1.982149e-07,1.982150e-07,1.982152e-07,1.982153e-07,1.982155e-07,1.982156e-07,1.982157e-07,1.982159e-07,1.982160e-07,1.982161e-07,1.982163e-07,1.982164e-07,1.982165e-07,1.982167e-07,1.982168e-07,1.982170e-07,1.982171e-07,1.982172e-07,1.982174e-07,1.982175e-07,1.982176e-07,1.982178e-07,1.982179e-07,1.982180e-07,1.982182e-07,1.982183e-07,1.982184e-07,1.982186e-07,1.982187e-07,1.982189e-07,1.982190e-07,1.982191e-07,1.982193e-07,1.982194e-07,1.982195e-07,1.982197e-07,1.982198e-07,1.982199e-07,1.982201e-07,1.982202e-07,1.982204e-07,1.982205e-07,1.982206e-07,1.982208e-07,1.982209e-07,1.982210e-07,1.982212e-07,1.982213e-07,1.982214e-07,1.982216e-07,1.982217e-07,1.982218e-07,1.982220e-07,1.982221e-07,1.982223e-07,1.982224e-07,1.982225e-07,1.982227e-07,1.982228e-07,1.982229e-07,1.982231e-07,1.982232e-07,1.982233e-07,1.982235e-07,1.982236e-07,1.982238e-07,1.982239e-07,1.982240e-07,1.982242e-07,1.982243e-07,1.982244e-07,1.982246e-07,1.982247e-07,1.982248e-07,1.982250e-07,1.982251e-07,1.982252e-07,1.982254e-07,1.982255e-07,1.982257e-07,1.982258e-07,1.982259e-07,1.982261e-07,1.982262e-07,1.982263e-07,1.982265e-07,1.982266e-07,1.982267e-07,1.982269e-07,1.982270e-07,1.982272e-07,1.982273e-07,1.982274e-07,1.982276e-07,1.982277e-07,1.982278e-07,1.982280e-07,1.982281e-07,1.982282e-07,1.982284e-07,1.982285e-07,1.982286e-07,1.982288e-07,1.982289e-07,1.982291e-07,1.982292e-07,1.982293e-07,1.982295e-07,1.982296e-07,1.982297e-07,1.982299e-07,1.982300e-07,1.982301e-07,1.982303e-07,1.982304e-07,1.982305e-07,1.982307e-07,1.982308e-07,1.982310e-07,1.982311e-07,1.982312e-07,1.982314e-07,1.982315e-07,1.982316e-07,1.982318e-07,1.982319e-07,1.982320e-07,1.982322e-07,1.982323e-07,1.982325e-07,1.982326e-07,1.982327e-07,1.982329e-07,1.982330e-07,1.982331e-07,1.982333e-07,1.982334e-07,1.982335e-07,1.982337e-07,1.982338e-07,1.982339e-07,1.982341e-07,1.982342e-07,1.982344e-07,1.982345e-07,1.982346e-07,1.982348e-07,1.982349e-07,1.982350e-07,1.982352e-07,1.982353e-07,1.982354e-07,1.982356e-07,1.982357e-07,1.982358e-07,1.982360e-07,1.982361e-07,1.982363e-07,1.982364e-07,1.982365e-07,1.982367e-07,1.982368e-07,1.982369e-07,1.982371e-07,1.982372e-07,1.982373e-07,1.982375e-07,1.982376e-07,1.982377e-07,1.982379e-07,1.982380e-07,1.982382e-07,1.982383e-07,1.982384e-07,1.982386e-07,1.982387e-07,1.982388e-07,1.982390e-07,1.982391e-07,1.982392e-07,1.982394e-07,1.982395e-07,1.982396e-07,1.982398e-07,1.982399e-07,1.982401e-07,1.982402e-07,1.982403e-07,1.982405e-07,1.982406e-07,1.982407e-07,1.982409e-07,1.982410e-07,1.982411e-07,1.982413e-07,1.982414e-07,1.982415e-07,1.982417e-07,1.982418e-07,1.982420e-07,1.982421e-07,1.982422e-07,1.982424e-07,1.982425e-07,1.982426e-07,1.982428e-07,1.982429e-07,1.982430e-07,1.982432e-07,1.982433e-07,1.982435e-07,1.982436e-07,1.982437e-07,1.982439e-07,1.982440e-07,1.982441e-07,1.982443e-07,1.982444e-07,1.982445e-07,1.982447e-07,1.982448e-07,1.982449e-07,1.982451e-07,1.982452e-07,1.982454e-07,1.982455e-07,1.982456e-07,1.982458e-07,1.982459e-07,1.982460e-07,1.982462e-07,1.982463e-07,1.982464e-07,1.982466e-07,1.982467e-07,1.982468e-07,1.982470e-07,1.982471e-07,1.982472e-07,1.982474e-07,1.982475e-07,1.982477e-07,1.982478e-07,1.982479e-07,1.982481e-07,1.982482e-07,1.982483e-07,1.982485e-07,1.982486e-07,1.982487e-07,1.982489e-07,1.982490e-07,1.982491e-07,1.982493e-07,1.982494e-07,1.982496e-07,1.982497e-07,1.982498e-07,1.982500e-07,1.982501e-07,1.982502e-07,1.982504e-07,1.982505e-07,1.982506e-07,1.982508e-07,1.982509e-07,1.982510e-07,1.982512e-07,1.982513e-07,1.982515e-07,1.982516e-07,1.982517e-07,1.982519e-07,1.982520e-07,1.982521e-07,1.982523e-07,1.982524e-07,1.982525e-07,1.982527e-07,1.982528e-07,1.982529e-07,1.982531e-07,1.982532e-07,1.982534e-07,1.982535e-07,1.982536e-07,1.982538e-07,1.982539e-07,1.982540e-07,1.982542e-07,1.982543e-07,1.982544e-07,1.982546e-07,1.982547e-07,1.982548e-07,1.982550e-07,1.982551e-07,1.982553e-07,1.982554e-07,1.982555e-07,1.982557e-07,1.982558e-07,1.982559e-07,1.982561e-07,1.982562e-07,1.982563e-07,1.982565e-07,1.982566e-07,1.982567e-07,1.982569e-07,1.982570e-07,1.982572e-07,1.982573e-07,1.982574e-07,1.982576e-07,1.982577e-07,1.982578e-07,1.982580e-07,1.982581e-07,1.982582e-07,1.982584e-07,1.982585e-07,1.982586e-07,1.982588e-07,1.982589e-07,1.982590e-07,1.982592e-07,1.982593e-07,1.982595e-07,1.982596e-07,1.982597e-07,1.982599e-07,1.982600e-07,1.982601e-07,1.982603e-07,1.982604e-07,1.982605e-07,1.982607e-07,1.982608e-07,1.982609e-07,1.982611e-07,1.982612e-07,1.982614e-07,1.982615e-07,1.982616e-07,1.982618e-07,1.982619e-07,1.982620e-07,1.982622e-07,1.982623e-07,1.982624e-07,1.982626e-07,1.982627e-07,1.982628e-07,1.982630e-07,1.982631e-07,1.982632e-07,1.982634e-07,1.982635e-07,1.982637e-07,1.982638e-07,1.982639e-07,1.982641e-07,1.982642e-07,1.982643e-07,1.982645e-07,1.982646e-07,1.982647e-07,1.982649e-07,1.982650e-07,1.982651e-07,1.982653e-07,1.982654e-07,1.982656e-07,1.982657e-07,1.982658e-07,1.982660e-07,1.982661e-07,1.982662e-07,1.982664e-07,1.982665e-07,1.982666e-07,1.982668e-07,1.982669e-07,1.982670e-07,1.982672e-07,1.982673e-07,1.982674e-07,1.982676e-07,1.982677e-07,1.982679e-07,1.982680e-07,1.982681e-07,1.982683e-07,1.982684e-07,1.982685e-07,1.982687e-07,1.982688e-07,1.982689e-07,1.982691e-07,1.982692e-07,1.982693e-07,1.982695e-07,1.982696e-07,1.982698e-07,1.982699e-07,1.982700e-07,1.982702e-07,1.982703e-07,1.982704e-07,1.982706e-07,1.982707e-07,1.982708e-07,1.982710e-07,1.982711e-07,1.982712e-07,1.982714e-07,1.982715e-07,1.982716e-07,1.982718e-07,1.982719e-07,1.982721e-07,1.982722e-07,1.982723e-07,1.982725e-07,1.982726e-07,1.982727e-07,1.982729e-07,1.982730e-07,1.982731e-07,1.982733e-07,1.982734e-07,1.982735e-07,1.982737e-07,1.982738e-07,1.982739e-07,1.982741e-07,1.982742e-07,1.982744e-07,1.982745e-07,1.982746e-07,1.982748e-07,1.982749e-07,1.982750e-07,1.982752e-07,1.982753e-07,1.982754e-07,1.982756e-07,1.982757e-07,1.982758e-07,1.982760e-07,1.982761e-07,1.982762e-07,1.982764e-07,1.982765e-07,1.982767e-07,1.982768e-07,1.982769e-07,1.982771e-07,1.982772e-07,1.982773e-07,1.982775e-07,1.982776e-07,1.982777e-07,1.982779e-07,1.982780e-07,1.982781e-07,1.982783e-07,1.982784e-07,1.982786e-07,1.982787e-07,1.982788e-07,1.982790e-07,1.982791e-07,1.982792e-07,1.982794e-07,1.982795e-07,1.982796e-07,1.982798e-07,1.982799e-07,1.982800e-07,1.982802e-07,1.982803e-07,1.982804e-07,1.982806e-07,1.982807e-07,1.982809e-07,1.982810e-07,1.982811e-07,1.982813e-07,1.982814e-07,1.982815e-07,1.982817e-07,1.982818e-07,1.982819e-07,1.982821e-07,1.982822e-07,1.982823e-07,1.982825e-07,1.982826e-07,1.982827e-07,1.982829e-07,1.982830e-07,1.982832e-07,1.982833e-07,1.982834e-07,1.982836e-07,1.982837e-07,1.982838e-07,1.982840e-07,1.982841e-07,1.982842e-07,1.982844e-07,1.982845e-07,1.982846e-07,1.982848e-07,1.982849e-07,1.982850e-07,1.982852e-07,1.982853e-07,1.982854e-07,1.982856e-07,1.982857e-07,1.982859e-07,1.982860e-07,1.982861e-07,1.982863e-07,1.982864e-07,1.982865e-07,1.982867e-07,1.982868e-07,1.982869e-07,1.982871e-07,1.982872e-07,1.982873e-07,1.982875e-07,1.982876e-07,1.982877e-07,1.982879e-07,1.982880e-07,1.982882e-07,1.982883e-07,1.982884e-07,1.982886e-07,1.982887e-07,1.982888e-07,1.982890e-07,1.982891e-07,1.982892e-07,1.982894e-07,1.982895e-07,1.982896e-07,1.982898e-07,1.982899e-07,1.982900e-07,1.982902e-07,1.982903e-07,1.982905e-07,1.982906e-07,1.982907e-07,1.982909e-07,1.982910e-07,1.982911e-07,1.982913e-07,1.982914e-07,1.982915e-07,1.982917e-07,1.982918e-07,1.982919e-07,1.982921e-07,1.982922e-07,1.982923e-07,1.982925e-07,1.982926e-07,1.982928e-07,1.982929e-07,1.982930e-07,1.982932e-07,1.982933e-07,1.982934e-07,1.982936e-07,1.982937e-07,1.982938e-07,1.982940e-07,1.982941e-07,1.982942e-07,1.982944e-07,1.982945e-07,1.982946e-07,1.982948e-07,1.982949e-07,1.982950e-07,1.982952e-07,1.982953e-07,1.982955e-07,1.982956e-07,1.982957e-07,1.982959e-07,1.982960e-07,1.982961e-07,1.982963e-07,1.982964e-07,1.982965e-07,1.982967e-07,1.982968e-07,1.982969e-07,1.982971e-07,1.982972e-07,1.982973e-07,1.982975e-07,1.982976e-07,1.982978e-07,1.982979e-07,1.982980e-07,1.982982e-07,1.982983e-07,1.982984e-07,1.982986e-07,1.982987e-07,1.982988e-07,1.982990e-07,1.982991e-07,1.982992e-07,1.982994e-07,1.982995e-07,1.982996e-07,1.982998e-07,1.982999e-07,1.983000e-07,1.983002e-07,1.983003e-07,1.983005e-07,1.983006e-07,1.983007e-07,1.983009e-07,1.983010e-07,1.983011e-07,1.983013e-07,1.983014e-07,1.983015e-07,1.983017e-07,1.983018e-07,1.983019e-07,1.983021e-07,1.983022e-07,1.983023e-07,1.983025e-07,1.983026e-07,1.983027e-07,1.983029e-07,1.983030e-07,1.983032e-07,1.983033e-07,1.983034e-07,1.983036e-07,1.983037e-07,1.983038e-07,1.983040e-07,1.983041e-07,1.983042e-07,1.983044e-07,1.983045e-07,1.983046e-07,1.983048e-07,1.983049e-07,1.983050e-07,1.983052e-07,1.983053e-07,1.983054e-07,1.983056e-07,1.983057e-07,1.983059e-07,1.983060e-07,1.983061e-07,1.983063e-07,1.983064e-07,1.983065e-07,1.983067e-07,1.983068e-07,1.983069e-07,1.983071e-07,1.983072e-07,1.983073e-07,1.983075e-07,1.983076e-07,1.983077e-07,1.983079e-07,1.983080e-07,1.983081e-07,1.983083e-07,1.983084e-07,1.983086e-07,1.983087e-07,1.983088e-07,1.983090e-07,1.983091e-07,1.983092e-07,1.983094e-07,1.983095e-07,1.983096e-07,1.983098e-07,1.983099e-07,1.983100e-07,1.983102e-07,1.983103e-07,1.983104e-07,1.983106e-07,1.983107e-07,1.983108e-07,1.983110e-07,1.983111e-07,1.983113e-07,1.983114e-07,1.983115e-07,1.983117e-07,1.983118e-07,1.983119e-07,1.983121e-07,1.983122e-07,1.983123e-07,1.983125e-07,1.983126e-07,1.983127e-07,1.983129e-07,1.983130e-07,1.983131e-07,1.983133e-07,1.983134e-07,1.983135e-07,1.983137e-07,1.983138e-07,1.983140e-07,1.983141e-07,1.983142e-07,1.983144e-07,1.983145e-07,1.983146e-07,1.983148e-07,1.983149e-07,1.983150e-07,1.983152e-07,1.983153e-07,1.983154e-07,1.983156e-07,1.983157e-07,1.983158e-07,1.983160e-07,1.983161e-07,1.983162e-07,1.983164e-07,1.983165e-07,1.983166e-07,1.983168e-07,1.983169e-07,1.983171e-07,1.983172e-07,1.983173e-07,1.983175e-07,1.983176e-07,1.983177e-07,1.983179e-07,1.983180e-07,1.983181e-07,1.983183e-07,1.983184e-07,1.983185e-07,1.983187e-07,1.983188e-07,1.983189e-07,1.983191e-07,1.983192e-07,1.983193e-07,1.983195e-07,1.983196e-07,1.983198e-07,1.983199e-07,1.983200e-07,1.983202e-07,1.983203e-07,1.983204e-07,1.983206e-07,1.983207e-07,1.983208e-07,1.983210e-07,1.983211e-07,1.983212e-07,1.983214e-07,1.983215e-07,1.983216e-07,1.983218e-07,1.983219e-07,1.983220e-07,1.983222e-07,1.983223e-07,1.983224e-07,1.983226e-07,1.983227e-07,1.983229e-07,1.983230e-07,1.983231e-07,1.983233e-07,1.983234e-07,1.983235e-07,1.983237e-07,1.983238e-07,1.983239e-07,1.983241e-07,1.983242e-07,1.983243e-07,1.983245e-07,1.983246e-07,1.983247e-07,1.983249e-07,1.983250e-07,1.983251e-07,1.983253e-07,1.983254e-07,1.983255e-07,1.983257e-07,1.983258e-07,1.983260e-07,1.983261e-07,1.983262e-07,1.983264e-07,1.983265e-07,1.983266e-07,1.983268e-07,1.983269e-07,1.983270e-07,1.983272e-07,1.983273e-07,1.983274e-07,1.983276e-07,1.983277e-07,1.983278e-07,1.983280e-07,1.983281e-07,1.983282e-07,1.983284e-07,1.983285e-07,1.983286e-07,1.983288e-07,1.983289e-07,1.983291e-07,1.983292e-07,1.983293e-07,1.983295e-07,1.983296e-07,1.983297e-07,1.983299e-07,1.983300e-07,1.983301e-07,1.983303e-07,1.983304e-07,1.983305e-07,1.983307e-07,1.983308e-07,1.983309e-07,1.983311e-07,1.983312e-07,1.983313e-07,1.983315e-07,1.983316e-07,1.983317e-07,1.983319e-07,1.983320e-07,1.983322e-07,1.983323e-07,1.983324e-07,1.983326e-07,1.983327e-07,1.983328e-07,1.983330e-07,1.983331e-07,1.983332e-07,1.983334e-07,1.983335e-07,1.983336e-07,1.983338e-07,1.983339e-07,1.983340e-07,1.983342e-07,1.983343e-07,1.983344e-07,1.983346e-07,1.983347e-07,1.983348e-07,1.983350e-07,1.983351e-07,1.983352e-07,1.983354e-07,1.983355e-07,1.983357e-07,1.983358e-07,1.983359e-07,1.983361e-07,1.983362e-07,1.983363e-07,1.983365e-07,1.983366e-07,1.983367e-07,1.983369e-07,1.983370e-07,1.983371e-07,1.983373e-07,1.983374e-07,1.983375e-07,1.983377e-07,1.983378e-07,1.983379e-07,1.983381e-07,1.983382e-07,1.983383e-07,1.983385e-07,1.983386e-07,1.983387e-07,1.983389e-07,1.983390e-07,1.983392e-07,1.983393e-07,1.983394e-07,1.983396e-07,1.983397e-07,1.983398e-07,1.983400e-07,1.983401e-07,1.983402e-07,1.983404e-07,1.983405e-07,1.983406e-07,1.983408e-07,1.983409e-07,1.983410e-07,1.983412e-07,1.983413e-07,1.983414e-07,1.983416e-07,1.983417e-07,1.983418e-07,1.983420e-07,1.983421e-07,1.983422e-07,1.983424e-07,1.983425e-07,1.983427e-07,1.983428e-07,1.983429e-07,1.983431e-07,1.983432e-07,1.983433e-07,1.983435e-07,1.983436e-07,1.983437e-07,1.983439e-07,1.983440e-07,1.983441e-07,1.983443e-07,1.983444e-07,1.983445e-07,1.983447e-07,1.983448e-07,1.983449e-07,1.983451e-07,1.983452e-07,1.983453e-07,1.983455e-07,1.983456e-07,1.983457e-07,1.983459e-07,1.983460e-07,1.983462e-07,1.983463e-07,1.983464e-07,1.983466e-07,1.983467e-07,1.983468e-07,1.983470e-07,1.983471e-07,1.983472e-07,1.983474e-07,1.983475e-07,1.983476e-07,1.983478e-07,1.983479e-07,1.983480e-07,1.983482e-07,1.983483e-07,1.983484e-07,1.983486e-07,1.983487e-07,1.983488e-07,1.983490e-07,1.983491e-07,1.983492e-07,1.983494e-07,1.983495e-07,1.983496e-07,1.983498e-07,1.983499e-07,1.983501e-07,1.983502e-07,1.983503e-07,1.983505e-07,1.983506e-07,1.983507e-07,1.983509e-07,1.983510e-07,1.983511e-07,1.983513e-07,1.983514e-07,1.983515e-07,1.983517e-07,1.983518e-07,1.983519e-07,1.983521e-07,1.983522e-07,1.983523e-07,1.983525e-07,1.983526e-07,1.983527e-07,1.983529e-07,1.983530e-07,1.983531e-07,1.983533e-07,1.983534e-07,1.983535e-07,1.983537e-07,1.983538e-07,1.983540e-07,1.983541e-07,1.983542e-07,1.983544e-07,1.983545e-07,1.983546e-07,1.983548e-07,1.983549e-07,1.983550e-07,1.983552e-07,1.983553e-07,1.983554e-07,1.983556e-07,1.983557e-07,1.983558e-07,1.983560e-07,1.983561e-07,1.983562e-07,1.983564e-07,1.983565e-07,1.983566e-07,1.983568e-07,1.983569e-07,1.983570e-07,1.983572e-07,1.983573e-07,1.983574e-07,1.983576e-07,1.983577e-07,1.983579e-07,1.983580e-07,1.983581e-07,1.983583e-07,1.983584e-07,1.983585e-07,1.983587e-07,1.983588e-07,1.983589e-07,1.983591e-07,1.983592e-07,1.983593e-07,1.983595e-07,1.983596e-07,1.983597e-07,1.983599e-07,1.983600e-07,1.983601e-07,1.983603e-07,1.983604e-07,1.983605e-07,1.983607e-07,1.983608e-07,1.983609e-07,1.983611e-07,1.983612e-07,1.983613e-07,1.983615e-07,1.983616e-07,1.983617e-07,1.983619e-07,1.983620e-07,1.983622e-07,1.983623e-07,1.983624e-07,1.983626e-07,1.983627e-07,1.983628e-07,1.983630e-07,1.983631e-07,1.983632e-07,1.983634e-07,1.983635e-07,1.983636e-07,1.983638e-07,1.983639e-07,1.983640e-07,1.983642e-07,1.983643e-07,1.983644e-07,1.983646e-07,1.983647e-07,1.983648e-07,1.983650e-07,1.983651e-07,1.983652e-07,1.983654e-07,1.983655e-07,1.983656e-07,1.983658e-07,1.983659e-07,1.983660e-07,1.983662e-07,1.983663e-07,1.983664e-07,1.983666e-07,1.983667e-07,1.983669e-07,1.983670e-07,1.983671e-07,1.983673e-07,1.983674e-07,1.983675e-07,1.983677e-07,1.983678e-07,1.983679e-07,1.983681e-07,1.983682e-07,1.983683e-07,1.983685e-07,1.983686e-07,1.983687e-07,1.983689e-07,1.983690e-07,1.983691e-07,1.983693e-07,1.983694e-07,1.983695e-07,1.983697e-07,1.983698e-07,1.983699e-07,1.983701e-07,1.983702e-07,1.983703e-07,1.983705e-07,1.983706e-07,1.983707e-07,1.983709e-07,1.983710e-07,1.983711e-07,1.983713e-07,1.983714e-07,1.983716e-07,1.983717e-07,1.983718e-07,1.983720e-07,1.983721e-07,1.983722e-07,1.983724e-07,1.983725e-07,1.983726e-07,1.983728e-07,1.983729e-07,1.983730e-07,1.983732e-07,1.983733e-07,1.983734e-07,1.983736e-07,1.983737e-07,1.983738e-07,1.983740e-07,1.983741e-07,1.983742e-07,1.983744e-07,1.983745e-07,1.983746e-07,1.983748e-07,1.983749e-07,1.983750e-07,1.983752e-07,1.983753e-07,1.983754e-07,1.983756e-07,1.983757e-07,1.983758e-07,1.983760e-07,1.983761e-07,1.983762e-07,1.983764e-07,1.983765e-07,1.983767e-07,1.983768e-07,1.983769e-07,1.983771e-07,1.983772e-07,1.983773e-07,1.983775e-07,1.983776e-07,1.983777e-07,1.983779e-07,1.983780e-07,1.983781e-07,1.983783e-07,1.983784e-07,1.983785e-07,1.983787e-07,1.983788e-07,1.983789e-07,1.983791e-07,1.983792e-07,1.983793e-07,1.983795e-07,1.983796e-07,1.983797e-07,1.983799e-07,1.983800e-07,1.983801e-07,1.983803e-07,1.983804e-07,1.983805e-07,1.983807e-07,1.983808e-07,1.983809e-07,1.983811e-07,1.983812e-07,1.983813e-07,1.983815e-07,1.983816e-07,1.983818e-07,1.983819e-07,1.983820e-07,1.983822e-07,1.983823e-07,1.983824e-07,1.983826e-07,1.983827e-07,1.983828e-07,1.983830e-07,1.983831e-07,1.983832e-07,1.983834e-07,1.983835e-07,1.983836e-07,1.983838e-07,1.983839e-07,1.983840e-07,1.983842e-07,1.983843e-07,1.983844e-07,1.983846e-07,1.983847e-07,1.983848e-07,1.983850e-07,1.983851e-07,1.983852e-07,1.983854e-07,1.983855e-07,1.983856e-07,1.983858e-07,1.983859e-07,1.983860e-07,1.983862e-07,1.983863e-07,1.983864e-07,1.983866e-07,1.983867e-07,1.983868e-07,1.983870e-07,1.983871e-07,1.983872e-07,1.983874e-07,1.983875e-07,1.983877e-07,1.983878e-07,1.983879e-07,1.983881e-07,1.983882e-07,1.983883e-07,1.983885e-07,1.983886e-07,1.983887e-07,1.983889e-07,1.983890e-07,1.983891e-07,1.983893e-07,1.983894e-07,1.983895e-07,1.983897e-07,1.983898e-07,1.983899e-07,1.983901e-07,1.983902e-07,1.983903e-07,1.983905e-07,1.983906e-07,1.983907e-07,1.983909e-07,1.983910e-07,1.983911e-07,1.983913e-07,1.983914e-07,1.983915e-07,1.983917e-07,1.983918e-07,1.983919e-07,1.983921e-07,1.983922e-07,1.983923e-07,1.983925e-07,1.983926e-07,1.983927e-07,1.983929e-07,1.983930e-07,1.983931e-07,1.983933e-07,1.983934e-07,1.983935e-07,1.983937e-07,1.983938e-07,1.983940e-07,1.983941e-07,1.983942e-07,1.983944e-07,1.983945e-07,1.983946e-07,1.983948e-07,1.983949e-07,1.983950e-07,1.983952e-07,1.983953e-07,1.983954e-07,1.983956e-07,1.983957e-07,1.983958e-07,1.983960e-07,1.983961e-07,1.983962e-07,1.983964e-07,1.983965e-07,1.983966e-07,1.983968e-07,1.983969e-07,1.983970e-07,1.983972e-07,1.983973e-07,1.983974e-07,1.983976e-07,1.983977e-07,1.983978e-07,1.983980e-07,1.983981e-07,1.983982e-07,1.983984e-07,1.983985e-07,1.983986e-07,1.983988e-07,1.983989e-07,1.983990e-07,1.983992e-07,1.983993e-07,1.983994e-07,1.983996e-07,1.983997e-07,1.983998e-07,1.984000e-07,1.984001e-07,1.984002e-07,1.984004e-07,1.984005e-07,1.984006e-07,1.984008e-07,1.984009e-07,1.984010e-07,1.984012e-07,1.984013e-07,1.984015e-07,1.984016e-07,1.984017e-07,1.984019e-07,1.984020e-07,1.984021e-07,1.984023e-07,1.984024e-07,1.984025e-07,1.984027e-07,1.984028e-07,1.984029e-07,1.984031e-07,1.984032e-07,1.984033e-07,1.984035e-07,1.984036e-07,1.984037e-07,1.984039e-07,1.984040e-07,1.984041e-07,1.984043e-07,1.984044e-07,1.984045e-07,1.984047e-07,1.984048e-07,1.984049e-07,1.984051e-07,1.984052e-07,1.984053e-07,1.984055e-07,1.984056e-07,1.984057e-07,1.984059e-07,1.984060e-07,1.984061e-07,1.984063e-07,1.984064e-07,1.984065e-07,1.984067e-07,1.984068e-07,1.984069e-07,1.984071e-07,1.984072e-07,1.984073e-07,1.984075e-07,1.984076e-07,1.984077e-07,1.984079e-07,1.984080e-07,1.984081e-07,1.984083e-07,1.984084e-07,1.984085e-07,1.984087e-07,1.984088e-07,1.984089e-07,1.984091e-07,1.984092e-07,1.984093e-07,1.984095e-07,1.984096e-07,1.984098e-07,1.984099e-07,1.984100e-07,1.984102e-07,1.984103e-07,1.984104e-07,1.984106e-07,1.984107e-07,1.984108e-07,1.984110e-07,1.984111e-07,1.984112e-07,1.984114e-07,1.984115e-07,1.984116e-07,1.984118e-07,1.984119e-07,1.984120e-07,1.984122e-07,1.984123e-07,1.984124e-07,1.984126e-07,1.984127e-07,1.984128e-07,1.984130e-07,1.984131e-07,1.984132e-07,1.984134e-07,1.984135e-07,1.984136e-07,1.984138e-07,1.984139e-07,1.984140e-07,1.984142e-07,1.984143e-07,1.984144e-07,1.984146e-07,1.984147e-07,1.984148e-07,1.984150e-07,1.984151e-07,1.984152e-07,1.984154e-07,1.984155e-07,1.984156e-07,1.984158e-07,1.984159e-07,1.984160e-07,1.984162e-07,1.984163e-07,1.984164e-07,1.984166e-07,1.984167e-07,1.984168e-07,1.984170e-07,1.984171e-07,1.984172e-07,1.984174e-07,1.984175e-07,1.984176e-07,1.984178e-07,1.984179e-07,1.984180e-07,1.984182e-07,1.984183e-07,1.984184e-07,1.984186e-07,1.984187e-07,1.984188e-07,1.984190e-07,1.984191e-07,1.984192e-07,1.984194e-07,1.984195e-07,1.984196e-07,1.984198e-07,1.984199e-07,1.984200e-07,1.984202e-07,1.984203e-07,1.984205e-07,1.984206e-07,1.984207e-07,1.984209e-07,1.984210e-07,1.984211e-07,1.984213e-07,1.984214e-07,1.984215e-07,1.984217e-07,1.984218e-07,1.984219e-07,1.984221e-07,1.984222e-07,1.984223e-07,1.984225e-07,1.984226e-07,1.984227e-07,1.984229e-07,1.984230e-07,1.984231e-07,1.984233e-07,1.984234e-07,1.984235e-07,1.984237e-07,1.984238e-07,1.984239e-07,1.984241e-07,1.984242e-07,1.984243e-07,1.984245e-07,1.984246e-07,1.984247e-07,1.984249e-07,1.984250e-07,1.984251e-07,1.984253e-07,1.984254e-07,1.984255e-07,1.984257e-07,1.984258e-07,1.984259e-07,1.984261e-07,1.984262e-07,1.984263e-07,1.984265e-07,1.984266e-07,1.984267e-07,1.984269e-07,1.984270e-07,1.984271e-07,1.984273e-07,1.984274e-07,1.984275e-07,1.984277e-07,1.984278e-07,1.984279e-07,1.984281e-07,1.984282e-07,1.984283e-07,1.984285e-07,1.984286e-07,1.984287e-07,1.984289e-07,1.984290e-07,1.984291e-07,1.984293e-07,1.984294e-07,1.984295e-07,1.984297e-07,1.984298e-07,1.984299e-07,1.984301e-07,1.984302e-07,1.984303e-07,1.984305e-07,1.984306e-07,1.984307e-07,1.984309e-07,1.984310e-07,1.984311e-07,1.984313e-07,1.984314e-07,1.984315e-07,1.984317e-07,1.984318e-07,1.984319e-07,1.984321e-07,1.984322e-07,1.984323e-07,1.984325e-07,1.984326e-07,1.984327e-07,1.984329e-07,1.984330e-07,1.984331e-07,1.984333e-07,1.984334e-07,1.984335e-07,1.984337e-07,1.984338e-07,1.984339e-07,1.984341e-07,1.984342e-07,1.984343e-07,1.984345e-07,1.984346e-07,1.984347e-07,1.984349e-07,1.984350e-07,1.984351e-07,1.984353e-07,1.984354e-07,1.984355e-07,1.984357e-07,1.984358e-07,1.984359e-07,1.984361e-07,1.984362e-07,1.984363e-07,1.984365e-07,1.984366e-07,1.984368e-07,1.984369e-07,1.984370e-07,1.984372e-07,1.984373e-07,1.984374e-07,1.984376e-07,1.984377e-07,1.984378e-07,1.984380e-07,1.984381e-07,1.984382e-07,1.984384e-07,1.984385e-07,1.984386e-07,1.984388e-07,1.984389e-07,1.984390e-07,1.984392e-07,1.984393e-07,1.984394e-07,1.984396e-07,1.984397e-07,1.984398e-07,1.984400e-07,1.984401e-07,1.984402e-07,1.984404e-07,1.984405e-07,1.984406e-07,1.984408e-07,1.984409e-07,1.984410e-07,1.984412e-07,1.984413e-07,1.984414e-07,1.984416e-07,1.984417e-07,1.984418e-07,1.984420e-07,1.984421e-07,1.984422e-07,1.984424e-07,1.984425e-07,1.984426e-07,1.984428e-07,1.984429e-07,1.984430e-07,1.984432e-07,1.984433e-07,1.984434e-07,1.984436e-07,1.984437e-07,1.984438e-07,1.984440e-07,1.984441e-07,1.984442e-07,1.984444e-07,1.984445e-07,1.984446e-07,1.984448e-07,1.984449e-07,1.984450e-07,1.984452e-07,1.984453e-07,1.984454e-07,1.984456e-07,1.984457e-07,1.984458e-07,1.984460e-07,1.984461e-07,1.984462e-07,1.984464e-07,1.984465e-07,1.984466e-07,1.984468e-07,1.984469e-07,1.984470e-07,1.984472e-07,1.984473e-07,1.984474e-07,1.984476e-07,1.984477e-07,1.984478e-07,1.984480e-07,1.984481e-07,1.984482e-07,1.984484e-07,1.984485e-07,1.984486e-07,1.984488e-07,1.984489e-07,1.984490e-07,1.984492e-07,1.984493e-07,1.984494e-07,1.984496e-07,1.984497e-07,1.984498e-07,1.984500e-07,1.984501e-07,1.984502e-07,1.984504e-07,1.984505e-07,1.984506e-07,1.984508e-07,1.984509e-07,1.984510e-07,1.984512e-07,1.984513e-07,1.984514e-07,1.984516e-07,1.984517e-07,1.984518e-07,1.984520e-07,1.984521e-07,1.984522e-07,1.984524e-07,1.984525e-07,1.984526e-07,1.984528e-07,1.984529e-07,1.984530e-07,1.984532e-07,1.984533e-07,1.984534e-07,1.984536e-07,1.984537e-07,1.984538e-07,1.984540e-07,1.984541e-07,1.984542e-07,1.984544e-07,1.984545e-07,1.984546e-07,1.984548e-07,1.984549e-07,1.984550e-07,1.984552e-07,1.984553e-07,1.984554e-07,1.984556e-07,1.984557e-07,1.984558e-07,1.984560e-07,1.984561e-07,1.984562e-07,1.984564e-07,1.984565e-07,1.984566e-07,1.984568e-07,1.984569e-07,1.984570e-07,1.984572e-07,1.984573e-07,1.984574e-07,1.984576e-07,1.984577e-07,1.984578e-07,1.984580e-07,1.984581e-07,1.984582e-07,1.984584e-07,1.984585e-07,1.984586e-07,1.984588e-07,1.984589e-07,1.984590e-07,1.984592e-07,1.984593e-07,1.984594e-07,1.984596e-07,1.984597e-07,1.984598e-07,1.984600e-07,1.984601e-07,1.984602e-07,1.984604e-07,1.984605e-07,1.984606e-07,1.984608e-07,1.984609e-07,1.984610e-07,1.984612e-07,1.984613e-07,1.984614e-07,1.984616e-07,1.984617e-07,1.984618e-07,1.984620e-07,1.984621e-07,1.984622e-07,1.984624e-07,1.984625e-07,1.984626e-07,1.984628e-07,1.984629e-07,1.984630e-07,1.984632e-07,1.984633e-07,1.984634e-07,1.984636e-07,1.984637e-07,1.984638e-07,1.984640e-07,1.984641e-07,1.984642e-07,1.984644e-07,1.984645e-07,1.984646e-07,1.984648e-07,1.984649e-07,1.984650e-07,1.984652e-07,1.984653e-07,1.984654e-07,1.984656e-07,1.984657e-07,1.984658e-07,1.984660e-07,1.984661e-07,1.984662e-07,1.984664e-07,1.984665e-07,1.984666e-07,1.984668e-07,1.984669e-07,1.984670e-07,1.984672e-07,1.984673e-07,1.984674e-07,1.984675e-07,1.984677e-07,1.984678e-07,1.984679e-07,1.984681e-07,1.984682e-07,1.984683e-07,1.984685e-07,1.984686e-07,1.984687e-07,1.984689e-07,1.984690e-07,1.984691e-07,1.984693e-07,1.984694e-07,1.984695e-07,1.984697e-07,1.984698e-07,1.984699e-07,1.984701e-07,1.984702e-07,1.984703e-07,1.984705e-07,1.984706e-07,1.984707e-07,1.984709e-07,1.984710e-07,1.984711e-07,1.984713e-07,1.984714e-07,1.984715e-07,1.984717e-07,1.984718e-07,1.984719e-07,1.984721e-07,1.984722e-07,1.984723e-07,1.984725e-07,1.984726e-07,1.984727e-07,1.984729e-07,1.984730e-07,1.984731e-07,1.984733e-07,1.984734e-07,1.984735e-07,1.984737e-07,1.984738e-07,1.984739e-07,1.984741e-07,1.984742e-07,1.984743e-07,1.984745e-07,1.984746e-07,1.984747e-07,1.984749e-07,1.984750e-07,1.984751e-07,1.984753e-07,1.984754e-07,1.984755e-07,1.984757e-07,1.984758e-07,1.984759e-07,1.984761e-07,1.984762e-07,1.984763e-07,1.984765e-07,1.984766e-07,1.984767e-07,1.984769e-07,1.984770e-07,1.984771e-07,1.984773e-07,1.984774e-07,1.984775e-07,1.984777e-07,1.984778e-07,1.984779e-07,1.984781e-07,1.984782e-07,1.984783e-07,1.984785e-07,1.984786e-07,1.984787e-07,1.984789e-07,1.984790e-07,1.984791e-07,1.984793e-07,1.984794e-07,1.984795e-07,1.984797e-07,1.984798e-07,1.984799e-07,1.984801e-07,1.984802e-07,1.984803e-07,1.984805e-07,1.984806e-07,1.984807e-07,1.984809e-07,1.984810e-07,1.984811e-07,1.984813e-07,1.984814e-07,1.984815e-07,1.984817e-07,1.984818e-07,1.984819e-07,1.984821e-07,1.984822e-07,1.984823e-07,1.984825e-07,1.984826e-07,1.984827e-07,1.984829e-07,1.984830e-07,1.984831e-07,1.984833e-07,1.984834e-07,1.984835e-07,1.984837e-07,1.984838e-07,1.984839e-07,1.984840e-07,1.984842e-07,1.984843e-07,1.984844e-07,1.984846e-07,1.984847e-07,1.984848e-07,1.984850e-07,1.984851e-07,1.984852e-07,1.984854e-07,1.984855e-07,1.984856e-07,1.984858e-07,1.984859e-07,1.984860e-07,1.984862e-07,1.984863e-07,1.984864e-07,1.984866e-07,1.984867e-07,1.984868e-07,1.984870e-07,1.984871e-07,1.984872e-07,1.984874e-07,1.984875e-07,1.984876e-07,1.984878e-07,1.984879e-07,1.984880e-07,1.984882e-07,1.984883e-07,1.984884e-07,1.984886e-07,1.984887e-07,1.984888e-07,1.984890e-07,1.984891e-07,1.984892e-07,1.984894e-07,1.984895e-07,1.984896e-07,1.984898e-07,1.984899e-07,1.984900e-07,1.984902e-07,1.984903e-07,1.984904e-07,1.984906e-07,1.984907e-07,1.984908e-07,1.984910e-07,1.984911e-07,1.984912e-07,1.984914e-07,1.984915e-07,1.984916e-07,1.984918e-07,1.984919e-07,1.984920e-07,1.984922e-07,1.984923e-07,1.984924e-07,1.984926e-07,1.984927e-07,1.984928e-07,1.984930e-07,1.984931e-07,1.984932e-07,1.984934e-07,1.984935e-07,1.984936e-07,1.984938e-07,1.984939e-07,1.984940e-07,1.984942e-07,1.984943e-07,1.984944e-07,1.984945e-07,1.984947e-07,1.984948e-07,1.984949e-07,1.984951e-07,1.984952e-07,1.984953e-07,1.984955e-07,1.984956e-07,1.984957e-07,1.984959e-07,1.984960e-07,1.984961e-07,1.984963e-07,1.984964e-07,1.984965e-07,1.984967e-07,1.984968e-07,1.984969e-07,1.984971e-07,1.984972e-07,1.984973e-07,1.984975e-07,1.984976e-07,1.984977e-07,1.984979e-07,1.984980e-07,1.984981e-07,1.984983e-07,1.984984e-07,1.984985e-07,1.984987e-07,1.984988e-07,1.984989e-07,1.984991e-07,1.984992e-07,1.984993e-07,1.984995e-07,1.984996e-07,1.984997e-07,1.984999e-07,1.985000e-07,1.985001e-07,1.985003e-07,1.985004e-07,1.985005e-07,1.985007e-07,1.985008e-07,1.985009e-07,1.985011e-07,1.985012e-07,1.985013e-07,1.985015e-07,1.985016e-07,1.985017e-07,1.985019e-07,1.985020e-07,1.985021e-07,1.985023e-07,1.985024e-07,1.985025e-07,1.985026e-07,1.985028e-07,1.985029e-07,1.985030e-07,1.985032e-07,1.985033e-07,1.985034e-07,1.985036e-07,1.985037e-07,1.985038e-07,1.985040e-07,1.985041e-07,1.985042e-07,1.985044e-07,1.985045e-07,1.985046e-07,1.985048e-07,1.985049e-07,1.985050e-07,1.985052e-07,1.985053e-07,1.985054e-07,1.985056e-07,1.985057e-07,1.985058e-07,1.985060e-07,1.985061e-07,1.985062e-07,1.985064e-07,1.985065e-07,1.985066e-07,1.985068e-07,1.985069e-07,1.985070e-07,1.985072e-07,1.985073e-07,1.985074e-07,1.985076e-07,1.985077e-07,1.985078e-07,1.985080e-07,1.985081e-07,1.985082e-07,1.985084e-07,1.985085e-07,1.985086e-07,1.985088e-07,1.985089e-07,1.985090e-07,1.985092e-07,1.985093e-07,1.985094e-07,1.985096e-07,1.985097e-07,1.985098e-07,1.985099e-07,1.985101e-07,1.985102e-07,1.985103e-07,1.985105e-07,1.985106e-07,1.985107e-07,1.985109e-07,1.985110e-07,1.985111e-07,1.985113e-07,1.985114e-07,1.985115e-07,1.985117e-07,1.985118e-07,1.985119e-07,1.985121e-07,1.985122e-07,1.985123e-07,1.985125e-07,1.985126e-07,1.985127e-07,1.985129e-07,1.985130e-07,1.985131e-07,1.985133e-07,1.985134e-07,1.985135e-07,1.985137e-07,1.985138e-07,1.985139e-07,1.985141e-07,1.985142e-07,1.985143e-07,1.985145e-07,1.985146e-07,1.985147e-07,1.985149e-07,1.985150e-07,1.985151e-07,1.985153e-07,1.985154e-07,1.985155e-07,1.985157e-07,1.985158e-07,1.985159e-07,1.985161e-07,1.985162e-07,1.985163e-07,1.985164e-07,1.985166e-07,1.985167e-07,1.985168e-07,1.985170e-07,1.985171e-07,1.985172e-07,1.985174e-07,1.985175e-07,1.985176e-07,1.985178e-07,1.985179e-07,1.985180e-07,1.985182e-07,1.985183e-07,1.985184e-07,1.985186e-07,1.985187e-07,1.985188e-07,1.985190e-07,1.985191e-07,1.985192e-07,1.985194e-07,1.985195e-07,1.985196e-07,1.985198e-07,1.985199e-07,1.985200e-07,1.985202e-07,1.985203e-07,1.985204e-07,1.985206e-07,1.985207e-07,1.985208e-07,1.985210e-07,1.985211e-07,1.985212e-07,1.985214e-07,1.985215e-07,1.985216e-07,1.985218e-07,1.985219e-07,1.985220e-07,1.985221e-07,1.985223e-07,1.985224e-07,1.985225e-07,1.985227e-07,1.985228e-07,1.985229e-07,1.985231e-07,1.985232e-07,1.985233e-07,1.985235e-07,1.985236e-07,1.985237e-07,1.985239e-07,1.985240e-07,1.985241e-07,1.985243e-07,1.985244e-07,1.985245e-07,1.985247e-07,1.985248e-07,1.985249e-07,1.985251e-07,1.985252e-07,1.985253e-07,1.985255e-07,1.985256e-07,1.985257e-07,1.985259e-07,1.985260e-07,1.985261e-07,1.985263e-07,1.985264e-07,1.985265e-07,1.985267e-07,1.985268e-07,1.985269e-07,1.985271e-07,1.985272e-07,1.985273e-07,1.985274e-07,1.985276e-07,1.985277e-07,1.985278e-07,1.985280e-07,1.985281e-07,1.985282e-07,1.985284e-07,1.985285e-07,1.985286e-07,1.985288e-07,1.985289e-07,1.985290e-07,1.985292e-07,1.985293e-07,1.985294e-07,1.985296e-07,1.985297e-07,1.985298e-07,1.985300e-07,1.985301e-07,1.985302e-07,1.985304e-07,1.985305e-07,1.985306e-07,1.985308e-07,1.985309e-07,1.985310e-07,1.985312e-07,1.985313e-07,1.985314e-07,1.985316e-07,1.985317e-07,1.985318e-07,1.985320e-07,1.985321e-07,1.985322e-07,1.985323e-07,1.985325e-07,1.985326e-07,1.985327e-07,1.985329e-07,1.985330e-07,1.985331e-07,1.985333e-07,1.985334e-07,1.985335e-07,1.985337e-07,1.985338e-07,1.985339e-07,1.985341e-07,1.985342e-07,1.985343e-07,1.985345e-07,1.985346e-07,1.985347e-07,1.985349e-07,1.985350e-07,1.985351e-07,1.985353e-07,1.985354e-07,1.985355e-07,1.985357e-07,1.985358e-07,1.985359e-07,1.985361e-07,1.985362e-07,1.985363e-07,1.985365e-07,1.985366e-07,1.985367e-07,1.985369e-07,1.985370e-07,1.985371e-07,1.985372e-07,1.985374e-07,1.985375e-07,1.985376e-07,1.985378e-07,1.985379e-07,1.985380e-07,1.985382e-07,1.985383e-07,1.985384e-07,1.985386e-07,1.985387e-07,1.985388e-07,1.985390e-07,1.985391e-07,1.985392e-07,1.985394e-07,1.985395e-07,1.985396e-07,1.985398e-07,1.985399e-07,1.985400e-07,1.985402e-07,1.985403e-07,1.985404e-07,1.985406e-07,1.985407e-07,1.985408e-07,1.985410e-07,1.985411e-07,1.985412e-07,1.985414e-07,1.985415e-07,1.985416e-07,1.985417e-07,1.985419e-07,1.985420e-07,1.985421e-07,1.985423e-07,1.985424e-07,1.985425e-07,1.985427e-07,1.985428e-07,1.985429e-07,1.985431e-07,1.985432e-07,1.985433e-07,1.985435e-07,1.985436e-07,1.985437e-07,1.985439e-07,1.985440e-07,1.985441e-07,1.985443e-07,1.985444e-07,1.985445e-07,1.985447e-07,1.985448e-07,1.985449e-07,1.985451e-07,1.985452e-07,1.985453e-07,1.985455e-07,1.985456e-07,1.985457e-07,1.985458e-07,1.985460e-07,1.985461e-07,1.985462e-07,1.985464e-07,1.985465e-07,1.985466e-07,1.985468e-07,1.985469e-07,1.985470e-07,1.985472e-07,1.985473e-07,1.985474e-07,1.985476e-07,1.985477e-07,1.985478e-07,1.985480e-07,1.985481e-07,1.985482e-07,1.985484e-07,1.985485e-07,1.985486e-07,1.985488e-07,1.985489e-07,1.985490e-07,1.985492e-07,1.985493e-07,1.985494e-07,1.985496e-07,1.985497e-07,1.985498e-07,1.985499e-07,1.985501e-07,1.985502e-07,1.985503e-07,1.985505e-07,1.985506e-07,1.985507e-07,1.985509e-07,1.985510e-07,1.985511e-07,1.985513e-07,1.985514e-07,1.985515e-07,1.985517e-07,1.985518e-07,1.985519e-07,1.985521e-07,1.985522e-07,1.985523e-07,1.985525e-07,1.985526e-07,1.985527e-07,1.985529e-07,1.985530e-07,1.985531e-07,1.985533e-07,1.985534e-07,1.985535e-07,1.985537e-07,1.985538e-07,1.985539e-07,1.985540e-07,1.985542e-07,1.985543e-07,1.985544e-07,1.985546e-07,1.985547e-07,1.985548e-07,1.985550e-07,1.985551e-07,1.985552e-07,1.985554e-07,1.985555e-07,1.985556e-07,1.985558e-07,1.985559e-07,1.985560e-07,1.985562e-07,1.985563e-07,1.985564e-07,1.985566e-07,1.985567e-07,1.985568e-07,1.985570e-07,1.985571e-07,1.985572e-07,1.985574e-07,1.985575e-07,1.985576e-07,1.985577e-07,1.985579e-07,1.985580e-07,1.985581e-07,1.985583e-07,1.985584e-07,1.985585e-07,1.985587e-07,1.985588e-07,1.985589e-07,1.985591e-07,1.985592e-07,1.985593e-07,1.985595e-07,1.985596e-07,1.985597e-07,1.985599e-07,1.985600e-07,1.985601e-07,1.985603e-07,1.985604e-07,1.985605e-07,1.985607e-07,1.985608e-07,1.985609e-07,1.985611e-07,1.985612e-07,1.985613e-07,1.985614e-07,1.985616e-07,1.985617e-07,1.985618e-07,1.985620e-07,1.985621e-07,1.985622e-07,1.985624e-07,1.985625e-07,1.985626e-07,1.985628e-07,1.985629e-07,1.985630e-07,1.985632e-07,1.985633e-07,1.985634e-07,1.985636e-07,1.985637e-07,1.985638e-07,1.985640e-07,1.985641e-07,1.985642e-07,1.985644e-07,1.985645e-07,1.985646e-07,1.985647e-07,1.985649e-07,1.985650e-07,1.985651e-07,1.985653e-07,1.985654e-07,1.985655e-07,1.985657e-07,1.985658e-07,1.985659e-07,1.985661e-07,1.985662e-07,1.985663e-07,1.985665e-07,1.985666e-07,1.985667e-07,1.985669e-07,1.985670e-07,1.985671e-07,1.985673e-07,1.985674e-07,1.985675e-07,1.985677e-07,1.985678e-07,1.985679e-07,1.985680e-07,1.985682e-07,1.985683e-07,1.985684e-07,1.985686e-07,1.985687e-07,1.985688e-07,1.985690e-07,1.985691e-07,1.985692e-07,1.985694e-07,1.985695e-07,1.985696e-07,1.985698e-07,1.985699e-07,1.985700e-07,1.985702e-07,1.985703e-07,1.985704e-07,1.985706e-07,1.985707e-07,1.985708e-07,1.985710e-07,1.985711e-07,1.985712e-07,1.985713e-07,1.985715e-07,1.985716e-07,1.985717e-07,1.985719e-07,1.985720e-07,1.985721e-07,1.985723e-07,1.985724e-07,1.985725e-07,1.985727e-07,1.985728e-07,1.985729e-07,1.985731e-07,1.985732e-07,1.985733e-07,1.985735e-07,1.985736e-07,1.985737e-07,1.985739e-07,1.985740e-07,1.985741e-07,1.985743e-07,1.985744e-07,1.985745e-07,1.985746e-07,1.985748e-07,1.985749e-07,1.985750e-07,1.985752e-07,1.985753e-07,1.985754e-07,1.985756e-07,1.985757e-07,1.985758e-07,1.985760e-07,1.985761e-07,1.985762e-07,1.985764e-07,1.985765e-07,1.985766e-07,1.985768e-07,1.985769e-07,1.985770e-07,1.985772e-07,1.985773e-07,1.985774e-07,1.985776e-07,1.985777e-07,1.985778e-07,1.985779e-07,1.985781e-07,1.985782e-07,1.985783e-07,1.985785e-07,1.985786e-07,1.985787e-07,1.985789e-07,1.985790e-07,1.985791e-07,1.985793e-07,1.985794e-07,1.985795e-07,1.985797e-07,1.985798e-07,1.985799e-07,1.985801e-07,1.985802e-07,1.985803e-07,1.985805e-07,1.985806e-07,1.985807e-07,1.985808e-07,1.985810e-07,1.985811e-07,1.985812e-07,1.985814e-07,1.985815e-07,1.985816e-07,1.985818e-07,1.985819e-07,1.985820e-07,1.985822e-07,1.985823e-07,1.985824e-07,1.985826e-07,1.985827e-07,1.985828e-07,1.985830e-07,1.985831e-07,1.985832e-07,1.985834e-07,1.985835e-07,1.985836e-07,1.985837e-07,1.985839e-07,1.985840e-07,1.985841e-07,1.985843e-07,1.985844e-07,1.985845e-07,1.985847e-07,1.985848e-07,1.985849e-07,1.985851e-07,1.985852e-07,1.985853e-07,1.985855e-07,1.985856e-07,1.985857e-07,1.985859e-07,1.985860e-07,1.985861e-07,1.985863e-07,1.985864e-07,1.985865e-07,1.985866e-07,1.985868e-07,1.985869e-07,1.985870e-07,1.985872e-07,1.985873e-07,1.985874e-07,1.985876e-07,1.985877e-07,1.985878e-07,1.985880e-07,1.985881e-07,1.985882e-07,1.985884e-07,1.985885e-07,1.985886e-07,1.985888e-07,1.985889e-07,1.985890e-07,1.985892e-07,1.985893e-07,1.985894e-07,1.985895e-07,1.985897e-07,1.985898e-07,1.985899e-07,1.985901e-07,1.985902e-07,1.985903e-07,1.985905e-07,1.985906e-07,1.985907e-07,1.985909e-07,1.985910e-07,1.985911e-07,1.985913e-07,1.985914e-07,1.985915e-07,1.985917e-07,1.985918e-07,1.985919e-07,1.985921e-07,1.985922e-07,1.985923e-07,1.985924e-07,1.985926e-07,1.985927e-07,1.985928e-07,1.985930e-07,1.985931e-07,1.985932e-07,1.985934e-07,1.985935e-07,1.985936e-07,1.985938e-07,1.985939e-07,1.985940e-07,1.985942e-07,1.985943e-07,1.985944e-07,1.985946e-07,1.985947e-07,1.985948e-07,1.985950e-07,1.985951e-07,1.985952e-07,1.985953e-07,1.985955e-07,1.985956e-07,1.985957e-07,1.985959e-07,1.985960e-07,1.985961e-07,1.985963e-07,1.985964e-07,1.985965e-07,1.985967e-07,1.985968e-07,1.985969e-07,1.985971e-07,1.985972e-07,1.985973e-07,1.985975e-07,1.985976e-07,1.985977e-07,1.985978e-07,1.985980e-07,1.985981e-07,1.985982e-07,1.985984e-07,1.985985e-07,1.985986e-07,1.985988e-07,1.985989e-07,1.985990e-07,1.985992e-07,1.985993e-07,1.985994e-07,1.985996e-07,1.985997e-07,1.985998e-07,1.986000e-07,1.986001e-07,1.986002e-07,1.986003e-07,1.986005e-07,1.986006e-07,1.986007e-07,1.986009e-07,1.986010e-07,1.986011e-07,1.986013e-07,1.986014e-07,1.986015e-07,1.986017e-07,1.986018e-07,1.986019e-07,1.986021e-07,1.986022e-07,1.986023e-07,1.986025e-07,1.986026e-07,1.986027e-07,1.986029e-07,1.986030e-07,1.986031e-07,1.986032e-07,1.986034e-07,1.986035e-07,1.986036e-07,1.986038e-07,1.986039e-07,1.986040e-07,1.986042e-07,1.986043e-07,1.986044e-07,1.986046e-07,1.986047e-07,1.986048e-07,1.986050e-07,1.986051e-07,1.986052e-07,1.986054e-07,1.986055e-07,1.986056e-07,1.986057e-07,1.986059e-07,1.986060e-07,1.986061e-07,1.986063e-07,1.986064e-07,1.986065e-07,1.986067e-07,1.986068e-07,1.986069e-07,1.986071e-07,1.986072e-07,1.986073e-07,1.986075e-07,1.986076e-07,1.986077e-07,1.986079e-07,1.986080e-07,1.986081e-07,1.986082e-07,1.986084e-07,1.986085e-07,1.986086e-07,1.986088e-07,1.986089e-07,1.986090e-07,1.986092e-07,1.986093e-07,1.986094e-07,1.986096e-07,1.986097e-07,1.986098e-07,1.986100e-07,1.986101e-07,1.986102e-07,1.986104e-07,1.986105e-07,1.986106e-07,1.986107e-07,1.986109e-07,1.986110e-07,1.986111e-07,1.986113e-07,1.986114e-07,1.986115e-07,1.986117e-07,1.986118e-07,1.986119e-07,1.986121e-07,1.986122e-07,1.986123e-07,1.986125e-07,1.986126e-07,1.986127e-07,1.986128e-07,1.986130e-07,1.986131e-07,1.986132e-07,1.986134e-07,1.986135e-07,1.986136e-07,1.986138e-07,1.986139e-07,1.986140e-07,1.986142e-07,1.986143e-07,1.986144e-07,1.986146e-07,1.986147e-07,1.986148e-07,1.986150e-07,1.986151e-07,1.986152e-07,1.986153e-07,1.986155e-07,1.986156e-07,1.986157e-07,1.986159e-07,1.986160e-07,1.986161e-07,1.986163e-07,1.986164e-07,1.986165e-07,1.986167e-07,1.986168e-07,1.986169e-07,1.986171e-07,1.986172e-07,1.986173e-07,1.986175e-07,1.986176e-07,1.986177e-07,1.986178e-07,1.986180e-07,1.986181e-07,1.986182e-07,1.986184e-07,1.986185e-07,1.986186e-07,1.986188e-07,1.986189e-07,1.986190e-07,1.986192e-07,1.986193e-07,1.986194e-07,1.986196e-07,1.986197e-07,1.986198e-07,1.986199e-07,1.986201e-07,1.986202e-07,1.986203e-07,1.986205e-07,1.986206e-07,1.986207e-07,1.986209e-07,1.986210e-07,1.986211e-07,1.986213e-07,1.986214e-07,1.986215e-07,1.986217e-07,1.986218e-07,1.986219e-07,1.986221e-07,1.986222e-07,1.986223e-07,1.986224e-07,1.986226e-07,1.986227e-07,1.986228e-07,1.986230e-07,1.986231e-07,1.986232e-07,1.986234e-07,1.986235e-07,1.986236e-07,1.986238e-07,1.986239e-07,1.986240e-07,1.986242e-07,1.986243e-07,1.986244e-07,1.986245e-07,1.986247e-07,1.986248e-07,1.986249e-07,1.986251e-07,1.986252e-07,1.986253e-07,1.986255e-07,1.986256e-07,1.986257e-07,1.986259e-07,1.986260e-07,1.986261e-07,1.986263e-07,1.986264e-07,1.986265e-07,1.986267e-07,1.986268e-07,1.986269e-07,1.986270e-07,1.986272e-07,1.986273e-07,1.986274e-07,1.986276e-07,1.986277e-07,1.986278e-07,1.986280e-07,1.986281e-07,1.986282e-07,1.986284e-07,1.986285e-07,1.986286e-07,1.986288e-07,1.986289e-07,1.986290e-07,1.986291e-07,1.986293e-07,1.986294e-07,1.986295e-07,1.986297e-07,1.986298e-07,1.986299e-07,1.986301e-07,1.986302e-07,1.986303e-07,1.986305e-07,1.986306e-07,1.986307e-07,1.986309e-07,1.986310e-07,1.986311e-07,1.986312e-07,1.986314e-07,1.986315e-07,1.986316e-07,1.986318e-07,1.986319e-07,1.986320e-07,1.986322e-07,1.986323e-07,1.986324e-07,1.986326e-07,1.986327e-07,1.986328e-07,1.986330e-07,1.986331e-07,1.986332e-07,1.986333e-07,1.986335e-07,1.986336e-07,1.986337e-07,1.986339e-07,1.986340e-07,1.986341e-07,1.986343e-07,1.986344e-07,1.986345e-07,1.986347e-07,1.986348e-07,1.986349e-07,1.986351e-07,1.986352e-07,1.986353e-07,1.986354e-07,1.986356e-07,1.986357e-07,1.986358e-07,1.986360e-07,1.986361e-07,1.986362e-07,1.986364e-07,1.986365e-07,1.986366e-07,1.986368e-07,1.986369e-07,1.986370e-07,1.986372e-07,1.986373e-07,1.986374e-07,1.986375e-07,1.986377e-07,1.986378e-07,1.986379e-07,1.986381e-07,1.986382e-07,1.986383e-07,1.986385e-07,1.986386e-07,1.986387e-07,1.986389e-07,1.986390e-07,1.986391e-07,1.986393e-07,1.986394e-07,1.986395e-07,1.986396e-07,1.986398e-07,1.986399e-07,1.986400e-07,1.986402e-07,1.986403e-07,1.986404e-07,1.986406e-07,1.986407e-07,1.986408e-07,1.986410e-07,1.986411e-07,1.986412e-07,1.986414e-07,1.986415e-07,1.986416e-07,1.986417e-07,1.986419e-07,1.986420e-07,1.986421e-07,1.986423e-07,1.986424e-07,1.986425e-07,1.986427e-07,1.986428e-07,1.986429e-07,1.986431e-07,1.986432e-07,1.986433e-07,1.986435e-07,1.986436e-07,1.986437e-07,1.986438e-07,1.986440e-07,1.986441e-07,1.986442e-07,1.986444e-07,1.986445e-07,1.986446e-07,1.986448e-07,1.986449e-07,1.986450e-07,1.986452e-07,1.986453e-07,1.986454e-07,1.986456e-07,1.986457e-07,1.986458e-07,1.986459e-07,1.986461e-07,1.986462e-07,1.986463e-07,1.986465e-07,1.986466e-07,1.986467e-07,1.986469e-07,1.986470e-07,1.986471e-07,1.986473e-07,1.986474e-07,1.986475e-07,1.986476e-07,1.986478e-07,1.986479e-07,1.986480e-07,1.986482e-07,1.986483e-07,1.986484e-07,1.986486e-07,1.986487e-07,1.986488e-07,1.986490e-07,1.986491e-07,1.986492e-07,1.986494e-07,1.986495e-07,1.986496e-07,1.986497e-07,1.986499e-07,1.986500e-07,1.986501e-07,1.986503e-07,1.986504e-07,1.986505e-07,1.986507e-07,1.986508e-07,1.986509e-07,1.986511e-07,1.986512e-07,1.986513e-07,1.986515e-07,1.986516e-07,1.986517e-07,1.986518e-07,1.986520e-07,1.986521e-07,1.986522e-07,1.986524e-07,1.986525e-07,1.986526e-07,1.986528e-07,1.986529e-07,1.986530e-07,1.986532e-07,1.986533e-07,1.986534e-07,1.986535e-07,1.986537e-07,1.986538e-07,1.986539e-07,1.986541e-07,1.986542e-07,1.986543e-07,1.986545e-07,1.986546e-07,1.986547e-07,1.986549e-07,1.986550e-07,1.986551e-07,1.986553e-07,1.986554e-07,1.986555e-07,1.986556e-07,1.986558e-07,1.986559e-07,1.986560e-07,1.986562e-07,1.986563e-07,1.986564e-07,1.986566e-07,1.986567e-07,1.986568e-07,1.986570e-07,1.986571e-07,1.986572e-07,1.986573e-07,1.986575e-07,1.986576e-07,1.986577e-07,1.986579e-07,1.986580e-07,1.986581e-07,1.986583e-07,1.986584e-07,1.986585e-07,1.986587e-07,1.986588e-07,1.986589e-07,1.986591e-07,1.986592e-07,1.986593e-07,1.986594e-07,1.986596e-07,1.986597e-07,1.986598e-07,1.986600e-07,1.986601e-07,1.986602e-07,1.986604e-07,1.986605e-07,1.986606e-07,1.986608e-07,1.986609e-07,1.986610e-07,1.986611e-07,1.986613e-07,1.986614e-07,1.986615e-07,1.986617e-07,1.986618e-07,1.986619e-07,1.986621e-07,1.986622e-07,1.986623e-07,1.986625e-07,1.986626e-07,1.986627e-07,1.986629e-07,1.986630e-07,1.986631e-07,1.986632e-07,1.986634e-07,1.986635e-07,1.986636e-07,1.986638e-07,1.986639e-07,1.986640e-07,1.986642e-07,1.986643e-07,1.986644e-07,1.986646e-07,1.986647e-07,1.986648e-07,1.986649e-07,1.986651e-07,1.986652e-07,1.986653e-07,1.986655e-07,1.986656e-07,1.986657e-07,1.986659e-07,1.986660e-07,1.986661e-07,1.986663e-07,1.986664e-07,1.986665e-07,1.986666e-07,1.986668e-07,1.986669e-07,1.986670e-07,1.986672e-07,1.986673e-07,1.986674e-07,1.986676e-07,1.986677e-07,1.986678e-07,1.986680e-07,1.986681e-07,1.986682e-07,1.986683e-07,1.986685e-07,1.986686e-07,1.986687e-07,1.986689e-07,1.986690e-07,1.986691e-07,1.986693e-07,1.986694e-07,1.986695e-07,1.986697e-07,1.986698e-07,1.986699e-07,1.986701e-07,1.986702e-07,1.986703e-07,1.986704e-07,1.986706e-07,1.986707e-07,1.986708e-07,1.986710e-07,1.986711e-07,1.986712e-07,1.986714e-07,1.986715e-07,1.986716e-07,1.986718e-07,1.986719e-07,1.986720e-07,1.986721e-07,1.986723e-07,1.986724e-07,1.986725e-07,1.986727e-07,1.986728e-07,1.986729e-07,1.986731e-07,1.986732e-07,1.986733e-07,1.986735e-07,1.986736e-07,1.986737e-07,1.986738e-07,1.986740e-07,1.986741e-07,1.986742e-07,1.986744e-07,1.986745e-07,1.986746e-07,1.986748e-07,1.986749e-07,1.986750e-07,1.986752e-07,1.986753e-07,1.986754e-07,1.986755e-07,1.986757e-07,1.986758e-07,1.986759e-07,1.986761e-07,1.986762e-07,1.986763e-07,1.986765e-07,1.986766e-07,1.986767e-07,1.986769e-07,1.986770e-07,1.986771e-07,1.986772e-07,1.986774e-07,1.986775e-07,1.986776e-07,1.986778e-07,1.986779e-07,1.986780e-07,1.986782e-07,1.986783e-07,1.986784e-07,1.986786e-07,1.986787e-07,1.986788e-07,1.986789e-07,1.986791e-07,1.986792e-07,1.986793e-07,1.986795e-07,1.986796e-07,1.986797e-07,1.986799e-07,1.986800e-07,1.986801e-07,1.986803e-07,1.986804e-07,1.986805e-07,1.986806e-07,1.986808e-07,1.986809e-07,1.986810e-07,1.986812e-07,1.986813e-07,1.986814e-07,1.986816e-07,1.986817e-07,1.986818e-07,1.986820e-07,1.986821e-07,1.986822e-07,1.986823e-07,1.986825e-07,1.986826e-07,1.986827e-07,1.986829e-07,1.986830e-07,1.986831e-07,1.986833e-07,1.986834e-07,1.986835e-07,1.986837e-07,1.986838e-07,1.986839e-07,1.986840e-07,1.986842e-07,1.986843e-07,1.986844e-07,1.986846e-07,1.986847e-07,1.986848e-07,1.986850e-07,1.986851e-07,1.986852e-07,1.986854e-07,1.986855e-07,1.986856e-07,1.986857e-07,1.986859e-07,1.986860e-07,1.986861e-07,1.986863e-07,1.986864e-07,1.986865e-07,1.986867e-07,1.986868e-07,1.986869e-07,1.986871e-07,1.986872e-07,1.986873e-07,1.986874e-07,1.986876e-07,1.986877e-07,1.986878e-07,1.986880e-07,1.986881e-07,1.986882e-07,1.986884e-07,1.986885e-07,1.986886e-07,1.986888e-07,1.986889e-07,1.986890e-07,1.986891e-07,1.986893e-07,1.986894e-07,1.986895e-07,1.986897e-07,1.986898e-07,1.986899e-07,1.986901e-07,1.986902e-07,1.986903e-07,1.986904e-07,1.986906e-07,1.986907e-07,1.986908e-07,1.986910e-07,1.986911e-07,1.986912e-07,1.986914e-07,1.986915e-07,1.986916e-07,1.986918e-07,1.986919e-07,1.986920e-07,1.986921e-07,1.986923e-07,1.986924e-07,1.986925e-07,1.986927e-07,1.986928e-07,1.986929e-07,1.986931e-07,1.986932e-07,1.986933e-07,1.986935e-07,1.986936e-07,1.986937e-07,1.986938e-07,1.986940e-07,1.986941e-07,1.986942e-07,1.986944e-07,1.986945e-07,1.986946e-07,1.986948e-07,1.986949e-07,1.986950e-07,1.986952e-07,1.986953e-07,1.986954e-07,1.986955e-07,1.986957e-07,1.986958e-07,1.986959e-07,1.986961e-07,1.986962e-07,1.986963e-07,1.986965e-07,1.986966e-07,1.986967e-07,1.986968e-07,1.986970e-07,1.986971e-07,1.986972e-07,1.986974e-07,1.986975e-07,1.986976e-07,1.986978e-07,1.986979e-07,1.986980e-07,1.986982e-07,1.986983e-07,1.986984e-07,1.986985e-07,1.986987e-07,1.986988e-07,1.986989e-07,1.986991e-07,1.986992e-07,1.986993e-07,1.986995e-07,1.986996e-07,1.986997e-07,1.986999e-07,1.987000e-07,1.987001e-07,1.987002e-07,1.987004e-07,1.987005e-07,1.987006e-07,1.987008e-07,1.987009e-07,1.987010e-07,1.987012e-07,1.987013e-07,1.987014e-07,1.987015e-07,1.987017e-07,1.987018e-07,1.987019e-07,1.987021e-07,1.987022e-07,1.987023e-07,1.987025e-07,1.987026e-07,1.987027e-07,1.987029e-07,1.987030e-07,1.987031e-07,1.987032e-07,1.987034e-07,1.987035e-07,1.987036e-07,1.987038e-07,1.987039e-07,1.987040e-07,1.987042e-07,1.987043e-07,1.987044e-07,1.987046e-07,1.987047e-07,1.987048e-07,1.987049e-07,1.987051e-07,1.987052e-07,1.987053e-07,1.987055e-07,1.987056e-07,1.987057e-07,1.987059e-07,1.987060e-07,1.987061e-07,1.987062e-07,1.987064e-07,1.987065e-07,1.987066e-07,1.987068e-07,1.987069e-07,1.987070e-07,1.987072e-07,1.987073e-07,1.987074e-07,1.987076e-07,1.987077e-07,1.987078e-07,1.987079e-07,1.987081e-07,1.987082e-07,1.987083e-07,1.987085e-07,1.987086e-07,1.987087e-07,1.987089e-07,1.987090e-07,1.987091e-07,1.987092e-07,1.987094e-07,1.987095e-07,1.987096e-07,1.987098e-07,1.987099e-07,1.987100e-07,1.987102e-07,1.987103e-07,1.987104e-07,1.987106e-07,1.987107e-07,1.987108e-07,1.987109e-07,1.987111e-07,1.987112e-07,1.987113e-07,1.987115e-07,1.987116e-07,1.987117e-07,1.987119e-07,1.987120e-07,1.987121e-07,1.987122e-07,1.987124e-07,1.987125e-07,1.987126e-07,1.987128e-07,1.987129e-07,1.987130e-07,1.987132e-07,1.987133e-07,1.987134e-07,1.987136e-07,1.987137e-07,1.987138e-07,1.987139e-07,1.987141e-07,1.987142e-07,1.987143e-07,1.987145e-07,1.987146e-07,1.987147e-07,1.987149e-07,1.987150e-07,1.987151e-07,1.987152e-07,1.987154e-07,1.987155e-07,1.987156e-07,1.987158e-07,1.987159e-07,1.987160e-07,1.987162e-07,1.987163e-07,1.987164e-07,1.987165e-07,1.987167e-07,1.987168e-07,1.987169e-07,1.987171e-07,1.987172e-07,1.987173e-07,1.987175e-07,1.987176e-07,1.987177e-07,1.987179e-07,1.987180e-07,1.987181e-07,1.987182e-07,1.987184e-07,1.987185e-07,1.987186e-07,1.987188e-07,1.987189e-07,1.987190e-07,1.987192e-07,1.987193e-07,1.987194e-07,1.987195e-07,1.987197e-07,1.987198e-07,1.987199e-07,1.987201e-07,1.987202e-07,1.987203e-07,1.987205e-07,1.987206e-07,1.987207e-07,1.987209e-07,1.987210e-07,1.987211e-07,1.987212e-07,1.987214e-07,1.987215e-07,1.987216e-07,1.987218e-07,1.987219e-07,1.987220e-07,1.987222e-07,1.987223e-07,1.987224e-07,1.987225e-07,1.987227e-07,1.987228e-07,1.987229e-07,1.987231e-07,1.987232e-07,1.987233e-07,1.987235e-07,1.987236e-07,1.987237e-07,1.987238e-07,1.987240e-07,1.987241e-07,1.987242e-07,1.987244e-07,1.987245e-07,1.987246e-07,1.987248e-07,1.987249e-07,1.987250e-07,1.987251e-07,1.987253e-07,1.987254e-07,1.987255e-07,1.987257e-07,1.987258e-07,1.987259e-07,1.987261e-07,1.987262e-07,1.987263e-07,1.987265e-07,1.987266e-07,1.987267e-07,1.987268e-07,1.987270e-07,1.987271e-07,1.987272e-07,1.987274e-07,1.987275e-07,1.987276e-07,1.987278e-07,1.987279e-07,1.987280e-07,1.987281e-07,1.987283e-07,1.987284e-07,1.987285e-07,1.987287e-07,1.987288e-07,1.987289e-07,1.987291e-07,1.987292e-07,1.987293e-07,1.987294e-07,1.987296e-07,1.987297e-07,1.987298e-07,1.987300e-07,1.987301e-07,1.987302e-07,1.987304e-07,1.987305e-07,1.987306e-07,1.987307e-07,1.987309e-07,1.987310e-07,1.987311e-07,1.987313e-07,1.987314e-07,1.987315e-07,1.987317e-07,1.987318e-07,1.987319e-07,1.987321e-07,1.987322e-07,1.987323e-07,1.987324e-07,1.987326e-07,1.987327e-07,1.987328e-07,1.987330e-07,1.987331e-07,1.987332e-07,1.987334e-07,1.987335e-07,1.987336e-07,1.987337e-07,1.987339e-07,1.987340e-07,1.987341e-07,1.987343e-07,1.987344e-07,1.987345e-07,1.987347e-07,1.987348e-07,1.987349e-07,1.987350e-07,1.987352e-07,1.987353e-07,1.987354e-07,1.987356e-07,1.987357e-07,1.987358e-07,1.987360e-07,1.987361e-07,1.987362e-07,1.987363e-07,1.987365e-07,1.987366e-07,1.987367e-07,1.987369e-07,1.987370e-07,1.987371e-07,1.987373e-07,1.987374e-07,1.987375e-07,1.987376e-07,1.987378e-07,1.987379e-07,1.987380e-07,1.987382e-07,1.987383e-07,1.987384e-07,1.987386e-07,1.987387e-07,1.987388e-07,1.987389e-07,1.987391e-07,1.987392e-07,1.987393e-07,1.987395e-07,1.987396e-07,1.987397e-07,1.987399e-07,1.987400e-07,1.987401e-07,1.987403e-07,1.987404e-07,1.987405e-07,1.987406e-07,1.987408e-07,1.987409e-07,1.987410e-07,1.987412e-07,1.987413e-07,1.987414e-07,1.987416e-07,1.987417e-07,1.987418e-07,1.987419e-07,1.987421e-07,1.987422e-07,1.987423e-07,1.987425e-07,1.987426e-07,1.987427e-07,1.987429e-07,1.987430e-07,1.987431e-07,1.987432e-07,1.987434e-07,1.987435e-07,1.987436e-07,1.987438e-07,1.987439e-07,1.987440e-07,1.987442e-07,1.987443e-07,1.987444e-07,1.987445e-07,1.987447e-07,1.987448e-07,1.987449e-07,1.987451e-07,1.987452e-07,1.987453e-07,1.987455e-07,1.987456e-07,1.987457e-07,1.987458e-07,1.987460e-07,1.987461e-07,1.987462e-07,1.987464e-07,1.987465e-07,1.987466e-07,1.987468e-07,1.987469e-07,1.987470e-07,1.987471e-07,1.987473e-07,1.987474e-07,1.987475e-07,1.987477e-07,1.987478e-07,1.987479e-07,1.987481e-07,1.987482e-07,1.987483e-07,1.987484e-07,1.987486e-07,1.987487e-07,1.987488e-07,1.987490e-07,1.987491e-07,1.987492e-07,1.987494e-07,1.987495e-07,1.987496e-07,1.987497e-07,1.987499e-07,1.987500e-07,1.987501e-07,1.987503e-07,1.987504e-07,1.987505e-07,1.987507e-07,1.987508e-07,1.987509e-07,1.987510e-07,1.987512e-07,1.987513e-07,1.987514e-07,1.987516e-07,1.987517e-07,1.987518e-07,1.987520e-07,1.987521e-07,1.987522e-07,1.987523e-07,1.987525e-07,1.987526e-07,1.987527e-07,1.987529e-07,1.987530e-07,1.987531e-07,1.987533e-07,1.987534e-07,1.987535e-07,1.987536e-07,1.987538e-07,1.987539e-07,1.987540e-07,1.987542e-07,1.987543e-07,1.987544e-07,1.987546e-07,1.987547e-07,1.987548e-07,1.987549e-07,1.987551e-07,1.987552e-07,1.987553e-07,1.987555e-07,1.987556e-07,1.987557e-07,1.987559e-07,1.987560e-07,1.987561e-07,1.987562e-07,1.987564e-07,1.987565e-07,1.987566e-07,1.987568e-07,1.987569e-07,1.987570e-07,1.987572e-07,1.987573e-07,1.987574e-07,1.987575e-07,1.987577e-07,1.987578e-07,1.987579e-07,1.987581e-07,1.987582e-07,1.987583e-07,1.987584e-07,1.987586e-07,1.987587e-07,1.987588e-07,1.987590e-07,1.987591e-07,1.987592e-07,1.987594e-07,1.987595e-07,1.987596e-07,1.987597e-07,1.987599e-07,1.987600e-07,1.987601e-07,1.987603e-07,1.987604e-07,1.987605e-07,1.987607e-07,1.987608e-07,1.987609e-07,1.987610e-07,1.987612e-07,1.987613e-07,1.987614e-07,1.987616e-07,1.987617e-07,1.987618e-07,1.987620e-07,1.987621e-07,1.987622e-07,1.987623e-07,1.987625e-07,1.987626e-07,1.987627e-07,1.987629e-07,1.987630e-07,1.987631e-07,1.987633e-07,1.987634e-07,1.987635e-07,1.987636e-07,1.987638e-07,1.987639e-07,1.987640e-07,1.987642e-07,1.987643e-07,1.987644e-07,1.987646e-07,1.987647e-07,1.987648e-07,1.987649e-07,1.987651e-07,1.987652e-07,1.987653e-07,1.987655e-07,1.987656e-07,1.987657e-07,1.987659e-07,1.987660e-07,1.987661e-07,1.987662e-07,1.987664e-07,1.987665e-07,1.987666e-07,1.987668e-07,1.987669e-07,1.987670e-07,1.987671e-07,1.987673e-07,1.987674e-07,1.987675e-07,1.987677e-07,1.987678e-07,1.987679e-07,1.987681e-07,1.987682e-07,1.987683e-07,1.987684e-07,1.987686e-07,1.987687e-07,1.987688e-07,1.987690e-07,1.987691e-07,1.987692e-07,1.987694e-07,1.987695e-07,1.987696e-07,1.987697e-07,1.987699e-07,1.987700e-07,1.987701e-07,1.987703e-07,1.987704e-07,1.987705e-07,1.987707e-07,1.987708e-07,1.987709e-07,1.987710e-07,1.987712e-07,1.987713e-07,1.987714e-07,1.987716e-07,1.987717e-07,1.987718e-07,1.987719e-07,1.987721e-07,1.987722e-07,1.987723e-07,1.987725e-07,1.987726e-07,1.987727e-07,1.987729e-07,1.987730e-07,1.987731e-07,1.987732e-07,1.987734e-07,1.987735e-07,1.987736e-07,1.987738e-07,1.987739e-07,1.987740e-07,1.987742e-07,1.987743e-07,1.987744e-07,1.987745e-07,1.987747e-07,1.987748e-07,1.987749e-07,1.987751e-07,1.987752e-07,1.987753e-07,1.987755e-07,1.987756e-07,1.987757e-07,1.987758e-07,1.987760e-07,1.987761e-07,1.987762e-07,1.987764e-07,1.987765e-07,1.987766e-07,1.987767e-07,1.987769e-07,1.987770e-07,1.987771e-07,1.987773e-07,1.987774e-07,1.987775e-07,1.987777e-07,1.987778e-07,1.987779e-07,1.987780e-07,1.987782e-07,1.987783e-07,1.987784e-07,1.987786e-07,1.987787e-07,1.987788e-07,1.987790e-07,1.987791e-07,1.987792e-07,1.987793e-07,1.987795e-07,1.987796e-07,1.987797e-07,1.987799e-07,1.987800e-07,1.987801e-07,1.987803e-07,1.987804e-07,1.987805e-07,1.987806e-07,1.987808e-07,1.987809e-07,1.987810e-07,1.987812e-07,1.987813e-07,1.987814e-07,1.987815e-07,1.987817e-07,1.987818e-07,1.987819e-07,1.987821e-07,1.987822e-07,1.987823e-07,1.987825e-07,1.987826e-07,1.987827e-07,1.987828e-07,1.987830e-07,1.987831e-07,1.987832e-07,1.987834e-07,1.987835e-07,1.987836e-07,1.987838e-07,1.987839e-07,1.987840e-07,1.987841e-07,1.987843e-07,1.987844e-07,1.987845e-07,1.987847e-07,1.987848e-07,1.987849e-07,1.987850e-07,1.987852e-07,1.987853e-07,1.987854e-07,1.987856e-07,1.987857e-07,1.987858e-07,1.987860e-07,1.987861e-07,1.987862e-07,1.987863e-07,1.987865e-07,1.987866e-07,1.987867e-07,1.987869e-07,1.987870e-07,1.987871e-07,1.987872e-07,1.987874e-07,1.987875e-07,1.987876e-07,1.987878e-07,1.987879e-07,1.987880e-07,1.987882e-07,1.987883e-07,1.987884e-07,1.987885e-07,1.987887e-07,1.987888e-07,1.987889e-07,1.987891e-07,1.987892e-07,1.987893e-07,1.987895e-07,1.987896e-07,1.987897e-07,1.987898e-07,1.987900e-07,1.987901e-07,1.987902e-07,1.987904e-07,1.987905e-07,1.987906e-07,1.987907e-07,1.987909e-07,1.987910e-07,1.987911e-07,1.987913e-07,1.987914e-07,1.987915e-07,1.987917e-07,1.987918e-07,1.987919e-07,1.987920e-07,1.987922e-07,1.987923e-07,1.987924e-07,1.987926e-07,1.987927e-07,1.987928e-07,1.987929e-07,1.987931e-07,1.987932e-07,1.987933e-07,1.987935e-07,1.987936e-07,1.987937e-07,1.987939e-07,1.987940e-07,1.987941e-07,1.987942e-07,1.987944e-07,1.987945e-07,1.987946e-07,1.987948e-07,1.987949e-07,1.987950e-07,1.987952e-07,1.987953e-07,1.987954e-07,1.987955e-07,1.987957e-07,1.987958e-07,1.987959e-07,1.987961e-07,1.987962e-07,1.987963e-07,1.987964e-07,1.987966e-07,1.987967e-07,1.987968e-07,1.987970e-07,1.987971e-07,1.987972e-07,1.987974e-07,1.987975e-07,1.987976e-07,1.987977e-07,1.987979e-07,1.987980e-07,1.987981e-07,1.987983e-07,1.987984e-07,1.987985e-07,1.987986e-07,1.987988e-07,1.987989e-07,1.987990e-07,1.987992e-07,1.987993e-07,1.987994e-07,1.987996e-07,1.987997e-07,1.987998e-07,1.987999e-07,1.988001e-07,1.988002e-07,1.988003e-07,1.988005e-07,1.988006e-07,1.988007e-07,1.988008e-07,1.988010e-07,1.988011e-07,1.988012e-07,1.988014e-07,1.988015e-07,1.988016e-07,1.988018e-07,1.988019e-07,1.988020e-07,1.988021e-07,1.988023e-07,1.988024e-07,1.988025e-07,1.988027e-07,1.988028e-07,1.988029e-07,1.988030e-07,1.988032e-07,1.988033e-07,1.988034e-07,1.988036e-07,1.988037e-07,1.988038e-07,1.988040e-07,1.988041e-07,1.988042e-07,1.988043e-07,1.988045e-07,1.988046e-07,1.988047e-07,1.988049e-07,1.988050e-07,1.988051e-07,1.988052e-07,1.988054e-07,1.988055e-07,1.988056e-07,1.988058e-07,1.988059e-07,1.988060e-07,1.988062e-07,1.988063e-07,1.988064e-07,1.988065e-07,1.988067e-07,1.988068e-07,1.988069e-07,1.988071e-07,1.988072e-07,1.988073e-07,1.988074e-07,1.988076e-07,1.988077e-07,1.988078e-07,1.988080e-07,1.988081e-07,1.988082e-07,1.988084e-07,1.988085e-07,1.988086e-07,1.988087e-07,1.988089e-07,1.988090e-07,1.988091e-07,1.988093e-07,1.988094e-07,1.988095e-07,1.988096e-07,1.988098e-07,1.988099e-07,1.988100e-07,1.988102e-07,1.988103e-07,1.988104e-07,1.988105e-07,1.988107e-07,1.988108e-07,1.988109e-07,1.988111e-07,1.988112e-07,1.988113e-07,1.988115e-07,1.988116e-07,1.988117e-07,1.988118e-07,1.988120e-07,1.988121e-07,1.988122e-07,1.988124e-07,1.988125e-07,1.988126e-07,1.988127e-07,1.988129e-07,1.988130e-07,1.988131e-07,1.988133e-07,1.988134e-07,1.988135e-07,1.988137e-07,1.988138e-07,1.988139e-07,1.988140e-07,1.988142e-07,1.988143e-07,1.988144e-07,1.988146e-07,1.988147e-07,1.988148e-07,1.988149e-07,1.988151e-07,1.988152e-07,1.988153e-07,1.988155e-07,1.988156e-07,1.988157e-07,1.988159e-07,1.988160e-07,1.988161e-07,1.988162e-07,1.988164e-07,1.988165e-07,1.988166e-07,1.988168e-07,1.988169e-07,1.988170e-07,1.988171e-07,1.988173e-07,1.988174e-07,1.988175e-07,1.988177e-07,1.988178e-07,1.988179e-07,1.988180e-07,1.988182e-07,1.988183e-07,1.988184e-07,1.988186e-07,1.988187e-07,1.988188e-07,1.988190e-07,1.988191e-07,1.988192e-07,1.988193e-07,1.988195e-07,1.988196e-07,1.988197e-07,1.988199e-07,1.988200e-07,1.988201e-07,1.988202e-07,1.988204e-07,1.988205e-07,1.988206e-07,1.988208e-07,1.988209e-07,1.988210e-07,1.988211e-07,1.988213e-07,1.988214e-07,1.988215e-07,1.988217e-07,1.988218e-07,1.988219e-07,1.988221e-07,1.988222e-07,1.988223e-07,1.988224e-07,1.988226e-07,1.988227e-07,1.988228e-07,1.988230e-07,1.988231e-07,1.988232e-07,1.988233e-07,1.988235e-07,1.988236e-07,1.988237e-07,1.988239e-07,1.988240e-07,1.988241e-07,1.988242e-07,1.988244e-07,1.988245e-07,1.988246e-07,1.988248e-07,1.988249e-07,1.988250e-07,1.988252e-07,1.988253e-07,1.988254e-07,1.988255e-07,1.988257e-07,1.988258e-07,1.988259e-07,1.988261e-07,1.988262e-07,1.988263e-07,1.988264e-07,1.988266e-07,1.988267e-07,1.988268e-07,1.988270e-07,1.988271e-07,1.988272e-07,1.988273e-07,1.988275e-07,1.988276e-07,1.988277e-07,1.988279e-07,1.988280e-07,1.988281e-07,1.988283e-07,1.988284e-07,1.988285e-07,1.988286e-07,1.988288e-07,1.988289e-07,1.988290e-07,1.988292e-07,1.988293e-07,1.988294e-07,1.988295e-07,1.988297e-07,1.988298e-07,1.988299e-07,1.988301e-07,1.988302e-07,1.988303e-07,1.988304e-07,1.988306e-07,1.988307e-07,1.988308e-07,1.988310e-07,1.988311e-07,1.988312e-07,1.988314e-07,1.988315e-07,1.988316e-07,1.988317e-07,1.988319e-07,1.988320e-07,1.988321e-07,1.988323e-07,1.988324e-07,1.988325e-07,1.988326e-07,1.988328e-07,1.988329e-07,1.988330e-07,1.988332e-07,1.988333e-07,1.988334e-07,1.988335e-07,1.988337e-07,1.988338e-07,1.988339e-07,1.988341e-07,1.988342e-07,1.988343e-07,1.988344e-07,1.988346e-07,1.988347e-07,1.988348e-07,1.988350e-07,1.988351e-07,1.988352e-07,1.988354e-07,1.988355e-07,1.988356e-07,1.988357e-07,1.988359e-07,1.988360e-07,1.988361e-07,1.988363e-07,1.988364e-07,1.988365e-07,1.988366e-07,1.988368e-07,1.988369e-07,1.988370e-07,1.988372e-07,1.988373e-07,1.988374e-07,1.988375e-07,1.988377e-07,1.988378e-07,1.988379e-07,1.988381e-07,1.988382e-07,1.988383e-07,1.988384e-07,1.988386e-07,1.988387e-07,1.988388e-07,1.988390e-07,1.988391e-07,1.988392e-07,1.988394e-07,1.988395e-07,1.988396e-07,1.988397e-07,1.988399e-07,1.988400e-07,1.988401e-07,1.988403e-07,1.988404e-07,1.988405e-07,1.988406e-07,1.988408e-07,1.988409e-07,1.988410e-07,1.988412e-07,1.988413e-07,1.988414e-07,1.988415e-07,1.988417e-07,1.988418e-07,1.988419e-07,1.988421e-07,1.988422e-07,1.988423e-07,1.988424e-07,1.988426e-07,1.988427e-07,1.988428e-07,1.988430e-07,1.988431e-07,1.988432e-07,1.988433e-07,1.988435e-07,1.988436e-07,1.988437e-07,1.988439e-07,1.988440e-07,1.988441e-07,1.988443e-07,1.988444e-07,1.988445e-07,1.988446e-07,1.988448e-07,1.988449e-07,1.988450e-07,1.988452e-07,1.988453e-07,1.988454e-07,1.988455e-07,1.988457e-07,1.988458e-07,1.988459e-07,1.988461e-07,1.988462e-07,1.988463e-07,1.988464e-07,1.988466e-07,1.988467e-07,1.988468e-07,1.988470e-07,1.988471e-07,1.988472e-07,1.988473e-07,1.988475e-07,1.988476e-07,1.988477e-07,1.988479e-07,1.988480e-07,1.988481e-07,1.988482e-07,1.988484e-07,1.988485e-07,1.988486e-07,1.988488e-07,1.988489e-07,1.988490e-07,1.988492e-07,1.988493e-07,1.988494e-07,1.988495e-07,1.988497e-07,1.988498e-07,1.988499e-07,1.988501e-07,1.988502e-07,1.988503e-07,1.988504e-07,1.988506e-07,1.988507e-07,1.988508e-07,1.988510e-07,1.988511e-07,1.988512e-07,1.988513e-07,1.988515e-07,1.988516e-07,1.988517e-07,1.988519e-07,1.988520e-07,1.988521e-07,1.988522e-07,1.988524e-07,1.988525e-07,1.988526e-07,1.988528e-07,1.988529e-07,1.988530e-07,1.988531e-07,1.988533e-07,1.988534e-07,1.988535e-07,1.988537e-07,1.988538e-07,1.988539e-07,1.988540e-07,1.988542e-07,1.988543e-07,1.988544e-07,1.988546e-07,1.988547e-07,1.988548e-07,1.988549e-07,1.988551e-07,1.988552e-07,1.988553e-07,1.988555e-07,1.988556e-07,1.988557e-07,1.988559e-07,1.988560e-07,1.988561e-07,1.988562e-07,1.988564e-07,1.988565e-07,1.988566e-07,1.988568e-07,1.988569e-07,1.988570e-07,1.988571e-07,1.988573e-07,1.988574e-07,1.988575e-07,1.988577e-07,1.988578e-07,1.988579e-07,1.988580e-07,1.988582e-07,1.988583e-07,1.988584e-07,1.988586e-07,1.988587e-07,1.988588e-07,1.988589e-07,1.988591e-07,1.988592e-07,1.988593e-07,1.988595e-07,1.988596e-07,1.988597e-07,1.988598e-07,1.988600e-07,1.988601e-07,1.988602e-07,1.988604e-07,1.988605e-07,1.988606e-07,1.988607e-07,1.988609e-07,1.988610e-07,1.988611e-07,1.988613e-07,1.988614e-07,1.988615e-07,1.988616e-07,1.988618e-07,1.988619e-07,1.988620e-07,1.988622e-07,1.988623e-07,1.988624e-07,1.988625e-07,1.988627e-07,1.988628e-07,1.988629e-07,1.988631e-07,1.988632e-07,1.988633e-07,1.988634e-07,1.988636e-07,1.988637e-07,1.988638e-07,1.988640e-07,1.988641e-07,1.988642e-07,1.988643e-07,1.988645e-07,1.988646e-07,1.988647e-07,1.988649e-07,1.988650e-07,1.988651e-07,1.988653e-07,1.988654e-07,1.988655e-07,1.988656e-07,1.988658e-07,1.988659e-07,1.988660e-07,1.988662e-07,1.988663e-07,1.988664e-07,1.988665e-07,1.988667e-07,1.988668e-07,1.988669e-07,1.988671e-07,1.988672e-07,1.988673e-07,1.988674e-07,1.988676e-07,1.988677e-07,1.988678e-07,1.988680e-07,1.988681e-07,1.988682e-07,1.988683e-07,1.988685e-07,1.988686e-07,1.988687e-07,1.988689e-07,1.988690e-07,1.988691e-07,1.988692e-07,1.988694e-07,1.988695e-07,1.988696e-07,1.988698e-07,1.988699e-07,1.988700e-07,1.988701e-07,1.988703e-07,1.988704e-07,1.988705e-07,1.988707e-07,1.988708e-07,1.988709e-07,1.988710e-07,1.988712e-07,1.988713e-07,1.988714e-07,1.988716e-07,1.988717e-07,1.988718e-07,1.988719e-07,1.988721e-07,1.988722e-07,1.988723e-07,1.988725e-07,1.988726e-07,1.988727e-07,1.988728e-07,1.988730e-07,1.988731e-07,1.988732e-07,1.988734e-07,1.988735e-07,1.988736e-07,1.988737e-07,1.988739e-07,1.988740e-07,1.988741e-07,1.988743e-07,1.988744e-07,1.988745e-07,1.988746e-07,1.988748e-07,1.988749e-07,1.988750e-07,1.988752e-07,1.988753e-07,1.988754e-07,1.988755e-07,1.988757e-07,1.988758e-07,1.988759e-07,1.988761e-07,1.988762e-07,1.988763e-07,1.988764e-07,1.988766e-07,1.988767e-07,1.988768e-07,1.988770e-07,1.988771e-07,1.988772e-07,1.988773e-07,1.988775e-07,1.988776e-07,1.988777e-07,1.988779e-07,1.988780e-07,1.988781e-07,1.988782e-07,1.988784e-07,1.988785e-07,1.988786e-07,1.988788e-07,1.988789e-07,1.988790e-07,1.988791e-07,1.988793e-07,1.988794e-07,1.988795e-07,1.988797e-07,1.988798e-07,1.988799e-07,1.988800e-07,1.988802e-07,1.988803e-07,1.988804e-07,1.988806e-07,1.988807e-07,1.988808e-07,1.988809e-07,1.988811e-07,1.988812e-07,1.988813e-07,1.988815e-07,1.988816e-07,1.988817e-07,1.988818e-07,1.988820e-07,1.988821e-07,1.988822e-07,1.988824e-07,1.988825e-07,1.988826e-07,1.988827e-07,1.988829e-07,1.988830e-07,1.988831e-07,1.988833e-07,1.988834e-07,1.988835e-07,1.988836e-07,1.988838e-07,1.988839e-07,1.988840e-07,1.988842e-07,1.988843e-07,1.988844e-07,1.988845e-07,1.988847e-07,1.988848e-07,1.988849e-07,1.988851e-07,1.988852e-07,1.988853e-07,1.988854e-07,1.988856e-07,1.988857e-07,1.988858e-07,1.988860e-07,1.988861e-07,1.988862e-07,1.988863e-07,1.988865e-07,1.988866e-07,1.988867e-07,1.988869e-07,1.988870e-07,1.988871e-07,1.988872e-07,1.988874e-07,1.988875e-07,1.988876e-07,1.988878e-07,1.988879e-07,1.988880e-07,1.988881e-07,1.988883e-07,1.988884e-07,1.988885e-07,1.988887e-07,1.988888e-07,1.988889e-07,1.988890e-07,1.988892e-07,1.988893e-07,1.988894e-07,1.988896e-07,1.988897e-07,1.988898e-07,1.988899e-07,1.988901e-07,1.988902e-07,1.988903e-07,1.988905e-07,1.988906e-07,1.988907e-07,1.988908e-07,1.988910e-07,1.988911e-07,1.988912e-07,1.988914e-07,1.988915e-07,1.988916e-07,1.988917e-07,1.988919e-07,1.988920e-07,1.988921e-07,1.988922e-07,1.988924e-07,1.988925e-07,1.988926e-07,1.988928e-07,1.988929e-07,1.988930e-07,1.988931e-07,1.988933e-07,1.988934e-07,1.988935e-07,1.988937e-07,1.988938e-07,1.988939e-07,1.988940e-07,1.988942e-07,1.988943e-07,1.988944e-07,1.988946e-07,1.988947e-07,1.988948e-07,1.988949e-07,1.988951e-07,1.988952e-07,1.988953e-07,1.988955e-07,1.988956e-07,1.988957e-07,1.988958e-07,1.988960e-07,1.988961e-07,1.988962e-07,1.988964e-07,1.988965e-07,1.988966e-07,1.988967e-07,1.988969e-07,1.988970e-07,1.988971e-07,1.988973e-07,1.988974e-07,1.988975e-07,1.988976e-07,1.988978e-07,1.988979e-07,1.988980e-07,1.988982e-07,1.988983e-07,1.988984e-07,1.988985e-07,1.988987e-07,1.988988e-07,1.988989e-07,1.988991e-07,1.988992e-07,1.988993e-07,1.988994e-07,1.988996e-07,1.988997e-07,1.988998e-07,1.989000e-07,1.989001e-07,1.989002e-07,1.989003e-07,1.989005e-07,1.989006e-07,1.989007e-07,1.989009e-07,1.989010e-07,1.989011e-07,1.989012e-07,1.989014e-07,1.989015e-07,1.989016e-07,1.989017e-07,1.989019e-07,1.989020e-07,1.989021e-07,1.989023e-07,1.989024e-07,1.989025e-07,1.989026e-07,1.989028e-07,1.989029e-07,1.989030e-07,1.989032e-07,1.989033e-07,1.989034e-07,1.989035e-07,1.989037e-07,1.989038e-07,1.989039e-07,1.989041e-07,1.989042e-07,1.989043e-07,1.989044e-07,1.989046e-07,1.989047e-07,1.989048e-07,1.989050e-07,1.989051e-07,1.989052e-07,1.989053e-07,1.989055e-07,1.989056e-07,1.989057e-07,1.989059e-07,1.989060e-07,1.989061e-07,1.989062e-07,1.989064e-07,1.989065e-07,1.989066e-07,1.989068e-07,1.989069e-07,1.989070e-07,1.989071e-07,1.989073e-07,1.989074e-07,1.989075e-07,1.989076e-07,1.989078e-07,1.989079e-07,1.989080e-07,1.989082e-07,1.989083e-07,1.989084e-07,1.989085e-07,1.989087e-07,1.989088e-07,1.989089e-07,1.989091e-07,1.989092e-07,1.989093e-07,1.989094e-07,1.989096e-07,1.989097e-07,1.989098e-07,1.989100e-07,1.989101e-07,1.989102e-07,1.989103e-07,1.989105e-07,1.989106e-07,1.989107e-07,1.989109e-07,1.989110e-07,1.989111e-07,1.989112e-07,1.989114e-07,1.989115e-07,1.989116e-07,1.989118e-07,1.989119e-07,1.989120e-07,1.989121e-07,1.989123e-07,1.989124e-07,1.989125e-07,1.989126e-07,1.989128e-07,1.989129e-07,1.989130e-07,1.989132e-07,1.989133e-07,1.989134e-07,1.989135e-07,1.989137e-07,1.989138e-07,1.989139e-07,1.989141e-07,1.989142e-07,1.989143e-07,1.989144e-07,1.989146e-07,1.989147e-07,1.989148e-07,1.989150e-07,1.989151e-07,1.989152e-07,1.989153e-07,1.989155e-07,1.989156e-07,1.989157e-07,1.989159e-07,1.989160e-07,1.989161e-07,1.989162e-07,1.989164e-07,1.989165e-07,1.989166e-07,1.989168e-07,1.989169e-07,1.989170e-07,1.989171e-07,1.989173e-07,1.989174e-07,1.989175e-07,1.989176e-07,1.989178e-07,1.989179e-07,1.989180e-07,1.989182e-07,1.989183e-07,1.989184e-07,1.989185e-07,1.989187e-07,1.989188e-07,1.989189e-07,1.989191e-07,1.989192e-07,1.989193e-07,1.989194e-07,1.989196e-07,1.989197e-07,1.989198e-07,1.989200e-07,1.989201e-07,1.989202e-07,1.989203e-07,1.989205e-07,1.989206e-07,1.989207e-07,1.989209e-07,1.989210e-07,1.989211e-07,1.989212e-07,1.989214e-07,1.989215e-07,1.989216e-07,1.989217e-07,1.989219e-07,1.989220e-07,1.989221e-07,1.989223e-07,1.989224e-07,1.989225e-07,1.989226e-07,1.989228e-07,1.989229e-07,1.989230e-07,1.989232e-07,1.989233e-07,1.989234e-07,1.989235e-07,1.989237e-07,1.989238e-07,1.989239e-07,1.989241e-07,1.989242e-07,1.989243e-07,1.989244e-07,1.989246e-07,1.989247e-07,1.989248e-07,1.989250e-07,1.989251e-07,1.989252e-07,1.989253e-07,1.989255e-07,1.989256e-07,1.989257e-07,1.989258e-07,1.989260e-07,1.989261e-07,1.989262e-07,1.989264e-07,1.989265e-07,1.989266e-07,1.989267e-07,1.989269e-07,1.989270e-07,1.989271e-07,1.989273e-07,1.989274e-07,1.989275e-07,1.989276e-07,1.989278e-07,1.989279e-07,1.989280e-07,1.989282e-07,1.989283e-07,1.989284e-07,1.989285e-07,1.989287e-07,1.989288e-07,1.989289e-07,1.989290e-07,1.989292e-07,1.989293e-07,1.989294e-07,1.989296e-07,1.989297e-07,1.989298e-07,1.989299e-07,1.989301e-07,1.989302e-07,1.989303e-07,1.989305e-07,1.989306e-07,1.989307e-07,1.989308e-07,1.989310e-07,1.989311e-07,1.989312e-07,1.989314e-07,1.989315e-07,1.989316e-07,1.989317e-07,1.989319e-07,1.989320e-07,1.989321e-07,1.989322e-07,1.989324e-07,1.989325e-07,1.989326e-07,1.989328e-07,1.989329e-07,1.989330e-07,1.989331e-07,1.989333e-07,1.989334e-07,1.989335e-07,1.989337e-07,1.989338e-07,1.989339e-07,1.989340e-07,1.989342e-07,1.989343e-07,1.989344e-07,1.989346e-07,1.989347e-07,1.989348e-07,1.989349e-07,1.989351e-07,1.989352e-07,1.989353e-07,1.989354e-07,1.989356e-07,1.989357e-07,1.989358e-07,1.989360e-07,1.989361e-07,1.989362e-07,1.989363e-07,1.989365e-07,1.989366e-07,1.989367e-07,1.989369e-07,1.989370e-07,1.989371e-07,1.989372e-07,1.989374e-07,1.989375e-07,1.989376e-07,1.989377e-07,1.989379e-07,1.989380e-07,1.989381e-07,1.989383e-07,1.989384e-07,1.989385e-07,1.989386e-07,1.989388e-07,1.989389e-07,1.989390e-07,1.989392e-07,1.989393e-07,1.989394e-07,1.989395e-07,1.989397e-07,1.989398e-07,1.989399e-07,1.989401e-07,1.989402e-07,1.989403e-07,1.989404e-07,1.989406e-07,1.989407e-07,1.989408e-07,1.989409e-07,1.989411e-07,1.989412e-07,1.989413e-07,1.989415e-07,1.989416e-07,1.989417e-07,1.989418e-07,1.989420e-07,1.989421e-07,1.989422e-07,1.989424e-07,1.989425e-07,1.989426e-07,1.989427e-07,1.989429e-07,1.989430e-07,1.989431e-07,1.989432e-07,1.989434e-07,1.989435e-07,1.989436e-07,1.989438e-07,1.989439e-07,1.989440e-07,1.989441e-07,1.989443e-07,1.989444e-07,1.989445e-07,1.989447e-07,1.989448e-07,1.989449e-07,1.989450e-07,1.989452e-07,1.989453e-07,1.989454e-07,1.989455e-07,1.989457e-07,1.989458e-07,1.989459e-07,1.989461e-07,1.989462e-07,1.989463e-07,1.989464e-07,1.989466e-07,1.989467e-07,1.989468e-07,1.989470e-07,1.989471e-07,1.989472e-07,1.989473e-07,1.989475e-07,1.989476e-07,1.989477e-07,1.989479e-07,1.989480e-07,1.989481e-07,1.989482e-07,1.989484e-07,1.989485e-07,1.989486e-07,1.989487e-07,1.989489e-07,1.989490e-07,1.989491e-07,1.989493e-07,1.989494e-07,1.989495e-07,1.989496e-07,1.989498e-07,1.989499e-07,1.989500e-07,1.989502e-07,1.989503e-07,1.989504e-07,1.989505e-07,1.989507e-07,1.989508e-07,1.989509e-07,1.989510e-07,1.989512e-07,1.989513e-07,1.989514e-07,1.989516e-07,1.989517e-07,1.989518e-07,1.989519e-07,1.989521e-07,1.989522e-07,1.989523e-07,1.989525e-07,1.989526e-07,1.989527e-07,1.989528e-07,1.989530e-07,1.989531e-07,1.989532e-07,1.989533e-07,1.989535e-07,1.989536e-07,1.989537e-07,1.989539e-07,1.989540e-07,1.989541e-07,1.989542e-07,1.989544e-07,1.989545e-07,1.989546e-07,1.989547e-07,1.989549e-07,1.989550e-07,1.989551e-07,1.989553e-07,1.989554e-07,1.989555e-07,1.989556e-07,1.989558e-07,1.989559e-07,1.989560e-07,1.989562e-07,1.989563e-07,1.989564e-07,1.989565e-07,1.989567e-07,1.989568e-07,1.989569e-07,1.989570e-07,1.989572e-07,1.989573e-07,1.989574e-07,1.989576e-07,1.989577e-07,1.989578e-07,1.989579e-07,1.989581e-07,1.989582e-07,1.989583e-07,1.989585e-07,1.989586e-07,1.989587e-07,1.989588e-07,1.989590e-07,1.989591e-07,1.989592e-07,1.989593e-07,1.989595e-07,1.989596e-07,1.989597e-07,1.989599e-07,1.989600e-07,1.989601e-07,1.989602e-07,1.989604e-07,1.989605e-07,1.989606e-07,1.989608e-07,1.989609e-07,1.989610e-07,1.989611e-07,1.989613e-07,1.989614e-07,1.989615e-07,1.989616e-07,1.989618e-07,1.989619e-07,1.989620e-07,1.989622e-07,1.989623e-07,1.989624e-07,1.989625e-07,1.989627e-07,1.989628e-07,1.989629e-07,1.989630e-07,1.989632e-07,1.989633e-07,1.989634e-07,1.989636e-07,1.989637e-07,1.989638e-07,1.989639e-07,1.989641e-07,1.989642e-07,1.989643e-07,1.989645e-07,1.989646e-07,1.989647e-07,1.989648e-07,1.989650e-07,1.989651e-07,1.989652e-07,1.989653e-07,1.989655e-07,1.989656e-07,1.989657e-07,1.989659e-07,1.989660e-07,1.989661e-07,1.989662e-07,1.989664e-07,1.989665e-07,1.989666e-07,1.989668e-07,1.989669e-07,1.989670e-07,1.989671e-07,1.989673e-07,1.989674e-07,1.989675e-07,1.989676e-07,1.989678e-07,1.989679e-07,1.989680e-07,1.989682e-07,1.989683e-07,1.989684e-07,1.989685e-07,1.989687e-07,1.989688e-07,1.989689e-07,1.989690e-07,1.989692e-07,1.989693e-07,1.989694e-07,1.989696e-07,1.989697e-07,1.989698e-07,1.989699e-07,1.989701e-07,1.989702e-07,1.989703e-07,1.989705e-07,1.989706e-07,1.989707e-07,1.989708e-07,1.989710e-07,1.989711e-07,1.989712e-07,1.989713e-07,1.989715e-07,1.989716e-07,1.989717e-07,1.989719e-07,1.989720e-07,1.989721e-07,1.989722e-07,1.989724e-07,1.989725e-07,1.989726e-07,1.989727e-07,1.989729e-07,1.989730e-07,1.989731e-07,1.989733e-07,1.989734e-07,1.989735e-07,1.989736e-07,1.989738e-07,1.989739e-07,1.989740e-07,1.989741e-07,1.989743e-07,1.989744e-07,1.989745e-07,1.989747e-07,1.989748e-07,1.989749e-07,1.989750e-07,1.989752e-07,1.989753e-07,1.989754e-07,1.989756e-07,1.989757e-07,1.989758e-07,1.989759e-07,1.989761e-07,1.989762e-07,1.989763e-07,1.989764e-07,1.989766e-07,1.989767e-07,1.989768e-07,1.989770e-07,1.989771e-07,1.989772e-07,1.989773e-07,1.989775e-07,1.989776e-07,1.989777e-07,1.989778e-07,1.989780e-07,1.989781e-07,1.989782e-07,1.989784e-07,1.989785e-07,1.989786e-07,1.989787e-07,1.989789e-07,1.989790e-07,1.989791e-07,1.989792e-07,1.989794e-07,1.989795e-07,1.989796e-07,1.989798e-07,1.989799e-07,1.989800e-07,1.989801e-07,1.989803e-07,1.989804e-07,1.989805e-07,1.989807e-07,1.989808e-07,1.989809e-07,1.989810e-07,1.989812e-07,1.989813e-07,1.989814e-07,1.989815e-07,1.989817e-07,1.989818e-07,1.989819e-07,1.989821e-07,1.989822e-07,1.989823e-07,1.989824e-07,1.989826e-07,1.989827e-07,1.989828e-07,1.989829e-07,1.989831e-07,1.989832e-07,1.989833e-07,1.989835e-07,1.989836e-07,1.989837e-07,1.989838e-07,1.989840e-07,1.989841e-07,1.989842e-07,1.989843e-07,1.989845e-07,1.989846e-07,1.989847e-07,1.989849e-07,1.989850e-07,1.989851e-07,1.989852e-07,1.989854e-07,1.989855e-07,1.989856e-07,1.989857e-07,1.989859e-07,1.989860e-07,1.989861e-07,1.989863e-07,1.989864e-07,1.989865e-07,1.989866e-07,1.989868e-07,1.989869e-07,1.989870e-07,1.989871e-07,1.989873e-07,1.989874e-07,1.989875e-07,1.989877e-07,1.989878e-07,1.989879e-07,1.989880e-07,1.989882e-07,1.989883e-07,1.989884e-07,1.989886e-07,1.989887e-07,1.989888e-07,1.989889e-07,1.989891e-07,1.989892e-07,1.989893e-07,1.989894e-07,1.989896e-07,1.989897e-07,1.989898e-07,1.989900e-07,1.989901e-07,1.989902e-07,1.989903e-07,1.989905e-07,1.989906e-07,1.989907e-07,1.989908e-07,1.989910e-07,1.989911e-07,1.989912e-07,1.989914e-07,1.989915e-07,1.989916e-07,1.989917e-07,1.989919e-07,1.989920e-07,1.989921e-07,1.989922e-07,1.989924e-07,1.989925e-07,1.989926e-07,1.989928e-07,1.989929e-07,1.989930e-07,1.989931e-07,1.989933e-07,1.989934e-07,1.989935e-07,1.989936e-07,1.989938e-07,1.989939e-07,1.989940e-07,1.989942e-07,1.989943e-07,1.989944e-07,1.989945e-07,1.989947e-07,1.989948e-07,1.989949e-07,1.989950e-07,1.989952e-07,1.989953e-07,1.989954e-07,1.989956e-07,1.989957e-07,1.989958e-07,1.989959e-07,1.989961e-07,1.989962e-07,1.989963e-07,1.989964e-07,1.989966e-07,1.989967e-07,1.989968e-07,1.989970e-07,1.989971e-07,1.989972e-07,1.989973e-07,1.989975e-07,1.989976e-07,1.989977e-07,1.989978e-07,1.989980e-07,1.989981e-07,1.989982e-07,1.989984e-07,1.989985e-07,1.989986e-07,1.989987e-07,1.989989e-07,1.989990e-07,1.989991e-07,1.989992e-07,1.989994e-07,1.989995e-07,1.989996e-07,1.989998e-07,1.989999e-07,1.990000e-07,1.990001e-07,1.990003e-07,1.990004e-07,1.990005e-07,1.990006e-07,1.990008e-07,1.990009e-07,1.990010e-07,1.990012e-07,1.990013e-07,1.990014e-07,1.990015e-07,1.990017e-07,1.990018e-07,1.990019e-07,1.990020e-07,1.990022e-07,1.990023e-07,1.990024e-07,1.990026e-07,1.990027e-07,1.990028e-07,1.990029e-07,1.990031e-07,1.990032e-07,1.990033e-07,1.990034e-07,1.990036e-07,1.990037e-07,1.990038e-07,1.990040e-07,1.990041e-07,1.990042e-07,1.990043e-07,1.990045e-07,1.990046e-07,1.990047e-07,1.990048e-07,1.990050e-07,1.990051e-07,1.990052e-07,1.990054e-07,1.990055e-07,1.990056e-07,1.990057e-07,1.990059e-07,1.990060e-07,1.990061e-07,1.990062e-07,1.990064e-07,1.990065e-07,1.990066e-07,1.990067e-07,1.990069e-07,1.990070e-07,1.990071e-07,1.990073e-07,1.990074e-07,1.990075e-07,1.990076e-07,1.990078e-07,1.990079e-07,1.990080e-07,1.990081e-07,1.990083e-07,1.990084e-07,1.990085e-07,1.990087e-07,1.990088e-07,1.990089e-07,1.990090e-07,1.990092e-07,1.990093e-07,1.990094e-07,1.990095e-07,1.990097e-07,1.990098e-07,1.990099e-07,1.990101e-07,1.990102e-07,1.990103e-07,1.990104e-07,1.990106e-07,1.990107e-07,1.990108e-07,1.990109e-07,1.990111e-07,1.990112e-07,1.990113e-07,1.990115e-07,1.990116e-07,1.990117e-07,1.990118e-07,1.990120e-07,1.990121e-07,1.990122e-07,1.990123e-07,1.990125e-07,1.990126e-07,1.990127e-07,1.990129e-07,1.990130e-07,1.990131e-07,1.990132e-07,1.990134e-07,1.990135e-07,1.990136e-07,1.990137e-07,1.990139e-07,1.990140e-07,1.990141e-07,1.990143e-07,1.990144e-07,1.990145e-07,1.990146e-07,1.990148e-07,1.990149e-07,1.990150e-07,1.990151e-07,1.990153e-07,1.990154e-07,1.990155e-07,1.990156e-07,1.990158e-07,1.990159e-07,1.990160e-07,1.990162e-07,1.990163e-07,1.990164e-07,1.990165e-07,1.990167e-07,1.990168e-07,1.990169e-07,1.990170e-07,1.990172e-07,1.990173e-07,1.990174e-07,1.990176e-07,1.990177e-07,1.990178e-07,1.990179e-07,1.990181e-07,1.990182e-07,1.990183e-07,1.990184e-07,1.990186e-07,1.990187e-07,1.990188e-07,1.990190e-07,1.990191e-07,1.990192e-07,1.990193e-07,1.990195e-07,1.990196e-07,1.990197e-07,1.990198e-07,1.990200e-07,1.990201e-07,1.990202e-07,1.990203e-07,1.990205e-07,1.990206e-07,1.990207e-07,1.990209e-07,1.990210e-07,1.990211e-07,1.990212e-07,1.990214e-07,1.990215e-07,1.990216e-07,1.990217e-07,1.990219e-07,1.990220e-07,1.990221e-07,1.990223e-07,1.990224e-07,1.990225e-07,1.990226e-07,1.990228e-07,1.990229e-07,1.990230e-07,1.990231e-07,1.990233e-07,1.990234e-07,1.990235e-07,1.990237e-07,1.990238e-07,1.990239e-07,1.990240e-07,1.990242e-07,1.990243e-07,1.990244e-07,1.990245e-07,1.990247e-07,1.990248e-07,1.990249e-07,1.990250e-07,1.990252e-07,1.990253e-07,1.990254e-07,1.990256e-07,1.990257e-07,1.990258e-07,1.990259e-07,1.990261e-07,1.990262e-07,1.990263e-07,1.990264e-07,1.990266e-07,1.990267e-07,1.990268e-07,1.990270e-07,1.990271e-07,1.990272e-07,1.990273e-07,1.990275e-07,1.990276e-07,1.990277e-07,1.990278e-07,1.990280e-07,1.990281e-07,1.990282e-07,1.990283e-07,1.990285e-07,1.990286e-07,1.990287e-07,1.990289e-07,1.990290e-07,1.990291e-07,1.990292e-07,1.990294e-07,1.990295e-07,1.990296e-07,1.990297e-07,1.990299e-07,1.990300e-07,1.990301e-07,1.990303e-07,1.990304e-07,1.990305e-07,1.990306e-07,1.990308e-07,1.990309e-07,1.990310e-07,1.990311e-07,1.990313e-07,1.990314e-07,1.990315e-07,1.990316e-07,1.990318e-07,1.990319e-07,1.990320e-07,1.990322e-07,1.990323e-07,1.990324e-07,1.990325e-07,1.990327e-07,1.990328e-07,1.990329e-07,1.990330e-07,1.990332e-07,1.990333e-07,1.990334e-07,1.990336e-07,1.990337e-07,1.990338e-07,1.990339e-07,1.990341e-07,1.990342e-07,1.990343e-07,1.990344e-07,1.990346e-07,1.990347e-07,1.990348e-07,1.990349e-07,1.990351e-07,1.990352e-07,1.990353e-07,1.990355e-07,1.990356e-07,1.990357e-07,1.990358e-07,1.990360e-07,1.990361e-07,1.990362e-07,1.990363e-07,1.990365e-07,1.990366e-07,1.990367e-07,1.990368e-07,1.990370e-07,1.990371e-07,1.990372e-07,1.990374e-07,1.990375e-07,1.990376e-07,1.990377e-07,1.990379e-07,1.990380e-07,1.990381e-07,1.990382e-07,1.990384e-07,1.990385e-07,1.990386e-07,1.990388e-07,1.990389e-07,1.990390e-07,1.990391e-07,1.990393e-07,1.990394e-07,1.990395e-07,1.990396e-07,1.990398e-07,1.990399e-07,1.990400e-07,1.990401e-07,1.990403e-07,1.990404e-07,1.990405e-07,1.990407e-07,1.990408e-07,1.990409e-07,1.990410e-07,1.990412e-07,1.990413e-07,1.990414e-07,1.990415e-07,1.990417e-07,1.990418e-07,1.990419e-07,1.990420e-07,1.990422e-07,1.990423e-07,1.990424e-07,1.990426e-07,1.990427e-07,1.990428e-07,1.990429e-07,1.990431e-07,1.990432e-07,1.990433e-07,1.990434e-07,1.990436e-07,1.990437e-07,1.990438e-07,1.990440e-07,1.990441e-07,1.990442e-07,1.990443e-07,1.990445e-07,1.990446e-07,1.990447e-07,1.990448e-07,1.990450e-07,1.990451e-07,1.990452e-07,1.990453e-07,1.990455e-07,1.990456e-07,1.990457e-07,1.990459e-07,1.990460e-07,1.990461e-07,1.990462e-07,1.990464e-07,1.990465e-07,1.990466e-07,1.990467e-07,1.990469e-07,1.990470e-07,1.990471e-07,1.990472e-07,1.990474e-07,1.990475e-07,1.990476e-07,1.990478e-07,1.990479e-07,1.990480e-07,1.990481e-07,1.990483e-07,1.990484e-07,1.990485e-07,1.990486e-07,1.990488e-07,1.990489e-07,1.990490e-07,1.990491e-07,1.990493e-07,1.990494e-07,1.990495e-07,1.990497e-07,1.990498e-07,1.990499e-07,1.990500e-07,1.990502e-07,1.990503e-07,1.990504e-07,1.990505e-07,1.990507e-07,1.990508e-07,1.990509e-07,1.990510e-07,1.990512e-07,1.990513e-07,1.990514e-07,1.990516e-07,1.990517e-07,1.990518e-07,1.990519e-07,1.990521e-07,1.990522e-07,1.990523e-07,1.990524e-07,1.990526e-07,1.990527e-07,1.990528e-07,1.990529e-07,1.990531e-07,1.990532e-07,1.990533e-07,1.990535e-07,1.990536e-07,1.990537e-07,1.990538e-07,1.990540e-07,1.990541e-07,1.990542e-07,1.990543e-07,1.990545e-07,1.990546e-07,1.990547e-07,1.990548e-07,1.990550e-07,1.990551e-07,1.990552e-07,1.990554e-07,1.990555e-07,1.990556e-07,1.990557e-07,1.990559e-07,1.990560e-07,1.990561e-07,1.990562e-07,1.990564e-07,1.990565e-07,1.990566e-07,1.990567e-07,1.990569e-07,1.990570e-07,1.990571e-07,1.990573e-07,1.990574e-07,1.990575e-07,1.990576e-07,1.990578e-07,1.990579e-07,1.990580e-07,1.990581e-07,1.990583e-07,1.990584e-07,1.990585e-07,1.990586e-07,1.990588e-07,1.990589e-07,1.990590e-07,1.990592e-07,1.990593e-07,1.990594e-07,1.990595e-07,1.990597e-07,1.990598e-07,1.990599e-07,1.990600e-07,1.990602e-07,1.990603e-07,1.990604e-07,1.990605e-07,1.990607e-07,1.990608e-07,1.990609e-07,1.990611e-07,1.990612e-07,1.990613e-07,1.990614e-07,1.990616e-07,1.990617e-07,1.990618e-07,1.990619e-07,1.990621e-07,1.990622e-07,1.990623e-07,1.990624e-07,1.990626e-07,1.990627e-07,1.990628e-07,1.990630e-07,1.990631e-07,1.990632e-07,1.990633e-07,1.990635e-07,1.990636e-07,1.990637e-07,1.990638e-07,1.990640e-07,1.990641e-07,1.990642e-07,1.990643e-07,1.990645e-07,1.990646e-07,1.990647e-07,1.990648e-07,1.990650e-07,1.990651e-07,1.990652e-07,1.990654e-07,1.990655e-07,1.990656e-07,1.990657e-07,1.990659e-07,1.990660e-07,1.990661e-07,1.990662e-07,1.990664e-07,1.990665e-07,1.990666e-07,1.990667e-07,1.990669e-07,1.990670e-07,1.990671e-07,1.990673e-07,1.990674e-07,1.990675e-07,1.990676e-07,1.990678e-07,1.990679e-07,1.990680e-07,1.990681e-07,1.990683e-07,1.990684e-07,1.990685e-07,1.990686e-07,1.990688e-07,1.990689e-07,1.990690e-07,1.990691e-07,1.990693e-07,1.990694e-07,1.990695e-07,1.990697e-07,1.990698e-07,1.990699e-07,1.990700e-07,1.990702e-07,1.990703e-07,1.990704e-07,1.990705e-07,1.990707e-07,1.990708e-07,1.990709e-07,1.990710e-07,1.990712e-07,1.990713e-07,1.990714e-07,1.990716e-07,1.990717e-07,1.990718e-07,1.990719e-07,1.990721e-07,1.990722e-07,1.990723e-07,1.990724e-07,1.990726e-07,1.990727e-07,1.990728e-07,1.990729e-07,1.990731e-07,1.990732e-07,1.990733e-07,1.990734e-07,1.990736e-07,1.990737e-07,1.990738e-07,1.990740e-07,1.990741e-07,1.990742e-07,1.990743e-07,1.990745e-07,1.990746e-07,1.990747e-07,1.990748e-07,1.990750e-07,1.990751e-07,1.990752e-07,1.990753e-07,1.990755e-07,1.990756e-07,1.990757e-07,1.990759e-07,1.990760e-07,1.990761e-07,1.990762e-07,1.990764e-07,1.990765e-07,1.990766e-07,1.990767e-07,1.990769e-07,1.990770e-07,1.990771e-07,1.990772e-07,1.990774e-07,1.990775e-07,1.990776e-07,1.990777e-07,1.990779e-07,1.990780e-07,1.990781e-07,1.990783e-07,1.990784e-07,1.990785e-07,1.990786e-07,1.990788e-07,1.990789e-07,1.990790e-07,1.990791e-07,1.990793e-07,1.990794e-07,1.990795e-07,1.990796e-07,1.990798e-07,1.990799e-07,1.990800e-07,1.990801e-07,1.990803e-07,1.990804e-07,1.990805e-07,1.990807e-07,1.990808e-07,1.990809e-07,1.990810e-07,1.990812e-07,1.990813e-07,1.990814e-07,1.990815e-07,1.990817e-07,1.990818e-07,1.990819e-07,1.990820e-07,1.990822e-07,1.990823e-07,1.990824e-07,1.990826e-07,1.990827e-07,1.990828e-07,1.990829e-07,1.990831e-07,1.990832e-07,1.990833e-07,1.990834e-07,1.990836e-07,1.990837e-07,1.990838e-07,1.990839e-07,1.990841e-07,1.990842e-07,1.990843e-07,1.990844e-07,1.990846e-07,1.990847e-07,1.990848e-07,1.990850e-07,1.990851e-07,1.990852e-07,1.990853e-07,1.990855e-07,1.990856e-07,1.990857e-07,1.990858e-07,1.990860e-07,1.990861e-07,1.990862e-07,1.990863e-07,1.990865e-07,1.990866e-07,1.990867e-07,1.990868e-07,1.990870e-07,1.990871e-07,1.990872e-07,1.990874e-07,1.990875e-07,1.990876e-07,1.990877e-07,1.990879e-07,1.990880e-07,1.990881e-07,1.990882e-07,1.990884e-07,1.990885e-07,1.990886e-07,1.990887e-07,1.990889e-07,1.990890e-07,1.990891e-07,1.990892e-07,1.990894e-07,1.990895e-07,1.990896e-07,1.990898e-07,1.990899e-07,1.990900e-07,1.990901e-07,1.990903e-07,1.990904e-07,1.990905e-07,1.990906e-07,1.990908e-07,1.990909e-07,1.990910e-07,1.990911e-07,1.990913e-07,1.990914e-07,1.990915e-07,1.990916e-07,1.990918e-07,1.990919e-07,1.990920e-07,1.990921e-07,1.990923e-07,1.990924e-07,1.990925e-07,1.990927e-07,1.990928e-07,1.990929e-07,1.990930e-07,1.990932e-07,1.990933e-07,1.990934e-07,1.990935e-07,1.990937e-07,1.990938e-07,1.990939e-07,1.990940e-07,1.990942e-07,1.990943e-07,1.990944e-07,1.990945e-07,1.990947e-07,1.990948e-07,1.990949e-07,1.990951e-07,1.990952e-07,1.990953e-07,1.990954e-07,1.990956e-07,1.990957e-07,1.990958e-07,1.990959e-07,1.990961e-07,1.990962e-07,1.990963e-07,1.990964e-07,1.990966e-07,1.990967e-07,1.990968e-07,1.990969e-07,1.990971e-07,1.990972e-07,1.990973e-07,1.990975e-07,1.990976e-07,1.990977e-07,1.990978e-07,1.990980e-07,1.990981e-07,1.990982e-07,1.990983e-07,1.990985e-07,1.990986e-07,1.990987e-07,1.990988e-07,1.990990e-07,1.990991e-07,1.990992e-07,1.990993e-07,1.990995e-07,1.990996e-07,1.990997e-07,1.990998e-07,1.991000e-07,1.991001e-07,1.991002e-07,1.991004e-07,1.991005e-07,1.991006e-07,1.991007e-07,1.991009e-07,1.991010e-07,1.991011e-07,1.991012e-07,1.991014e-07,1.991015e-07,1.991016e-07,1.991017e-07,1.991019e-07,1.991020e-07,1.991021e-07,1.991022e-07,1.991024e-07,1.991025e-07,1.991026e-07,1.991027e-07,1.991029e-07,1.991030e-07,1.991031e-07,1.991033e-07,1.991034e-07,1.991035e-07,1.991036e-07,1.991038e-07,1.991039e-07,1.991040e-07,1.991041e-07,1.991043e-07,1.991044e-07,1.991045e-07,1.991046e-07,1.991048e-07,1.991049e-07,1.991050e-07,1.991051e-07,1.991053e-07,1.991054e-07,1.991055e-07,1.991056e-07,1.991058e-07,1.991059e-07,1.991060e-07,1.991062e-07,1.991063e-07,1.991064e-07,1.991065e-07,1.991067e-07,1.991068e-07,1.991069e-07,1.991070e-07,1.991072e-07,1.991073e-07,1.991074e-07,1.991075e-07,1.991077e-07,1.991078e-07,1.991079e-07,1.991080e-07,1.991082e-07,1.991083e-07,1.991084e-07,1.991085e-07,1.991087e-07,1.991088e-07,1.991089e-07,1.991091e-07,1.991092e-07,1.991093e-07,1.991094e-07,1.991096e-07,1.991097e-07,1.991098e-07,1.991099e-07,1.991101e-07,1.991102e-07,1.991103e-07,1.991104e-07,1.991106e-07,1.991107e-07,1.991108e-07,1.991109e-07,1.991111e-07,1.991112e-07,1.991113e-07,1.991114e-07,1.991116e-07,1.991117e-07,1.991118e-07,1.991120e-07,1.991121e-07,1.991122e-07,1.991123e-07,1.991125e-07,1.991126e-07,1.991127e-07,1.991128e-07,1.991130e-07,1.991131e-07,1.991132e-07,1.991133e-07,1.991135e-07,1.991136e-07,1.991137e-07,1.991138e-07,1.991140e-07,1.991141e-07,1.991142e-07,1.991143e-07,1.991145e-07,1.991146e-07,1.991147e-07,1.991149e-07,1.991150e-07,1.991151e-07,1.991152e-07,1.991154e-07,1.991155e-07,1.991156e-07,1.991157e-07,1.991159e-07,1.991160e-07,1.991161e-07,1.991162e-07,1.991164e-07,1.991165e-07,1.991166e-07,1.991167e-07,1.991169e-07,1.991170e-07,1.991171e-07,1.991172e-07,1.991174e-07,1.991175e-07,1.991176e-07,1.991177e-07,1.991179e-07,1.991180e-07,1.991181e-07,1.991183e-07,1.991184e-07,1.991185e-07,1.991186e-07,1.991188e-07,1.991189e-07,1.991190e-07,1.991191e-07,1.991193e-07,1.991194e-07,1.991195e-07,1.991196e-07,1.991198e-07,1.991199e-07,1.991200e-07,1.991201e-07,1.991203e-07,1.991204e-07,1.991205e-07,1.991206e-07,1.991208e-07,1.991209e-07,1.991210e-07,1.991211e-07,1.991213e-07,1.991214e-07,1.991215e-07,1.991217e-07,1.991218e-07,1.991219e-07,1.991220e-07,1.991222e-07,1.991223e-07,1.991224e-07,1.991225e-07,1.991227e-07,1.991228e-07,1.991229e-07,1.991230e-07,1.991232e-07,1.991233e-07,1.991234e-07,1.991235e-07,1.991237e-07,1.991238e-07,1.991239e-07,1.991240e-07,1.991242e-07,1.991243e-07,1.991244e-07,1.991245e-07,1.991247e-07,1.991248e-07,1.991249e-07,1.991251e-07,1.991252e-07,1.991253e-07,1.991254e-07,1.991256e-07,1.991257e-07,1.991258e-07,1.991259e-07,1.991261e-07,1.991262e-07,1.991263e-07,1.991264e-07,1.991266e-07,1.991267e-07,1.991268e-07,1.991269e-07,1.991271e-07,1.991272e-07,1.991273e-07,1.991274e-07,1.991276e-07,1.991277e-07,1.991278e-07,1.991279e-07,1.991281e-07,1.991282e-07,1.991283e-07,1.991285e-07,1.991286e-07,1.991287e-07,1.991288e-07,1.991290e-07,1.991291e-07,1.991292e-07,1.991293e-07,1.991295e-07,1.991296e-07,1.991297e-07,1.991298e-07,1.991300e-07,1.991301e-07,1.991302e-07,1.991303e-07,1.991305e-07,1.991306e-07,1.991307e-07,1.991308e-07,1.991310e-07,1.991311e-07,1.991312e-07,1.991313e-07,1.991315e-07,1.991316e-07,1.991317e-07,1.991318e-07,1.991320e-07,1.991321e-07,1.991322e-07,1.991324e-07,1.991325e-07,1.991326e-07,1.991327e-07,1.991329e-07,1.991330e-07,1.991331e-07,1.991332e-07,1.991334e-07,1.991335e-07,1.991336e-07,1.991337e-07,1.991339e-07,1.991340e-07,1.991341e-07,1.991342e-07,1.991344e-07,1.991345e-07,1.991346e-07,1.991347e-07,1.991349e-07,1.991350e-07,1.991351e-07,1.991352e-07,1.991354e-07,1.991355e-07,1.991356e-07,1.991357e-07,1.991359e-07,1.991360e-07,1.991361e-07,1.991363e-07,1.991364e-07,1.991365e-07,1.991366e-07,1.991368e-07,1.991369e-07,1.991370e-07,1.991371e-07,1.991373e-07,1.991374e-07,1.991375e-07,1.991376e-07,1.991378e-07,1.991379e-07,1.991380e-07,1.991381e-07,1.991383e-07,1.991384e-07,1.991385e-07,1.991386e-07,1.991388e-07,1.991389e-07,1.991390e-07,1.991391e-07,1.991393e-07,1.991394e-07,1.991395e-07,1.991396e-07,1.991398e-07,1.991399e-07,1.991400e-07,1.991401e-07,1.991403e-07,1.991404e-07,1.991405e-07,1.991407e-07,1.991408e-07,1.991409e-07,1.991410e-07,1.991412e-07,1.991413e-07,1.991414e-07,1.991415e-07,1.991417e-07,1.991418e-07,1.991419e-07,1.991420e-07,1.991422e-07,1.991423e-07,1.991424e-07,1.991425e-07,1.991427e-07,1.991428e-07,1.991429e-07,1.991430e-07,1.991432e-07,1.991433e-07,1.991434e-07,1.991435e-07,1.991437e-07,1.991438e-07,1.991439e-07,1.991440e-07,1.991442e-07,1.991443e-07,1.991444e-07,1.991445e-07,1.991447e-07,1.991448e-07,1.991449e-07,1.991451e-07,1.991452e-07,1.991453e-07,1.991454e-07,1.991456e-07,1.991457e-07,1.991458e-07,1.991459e-07,1.991461e-07,1.991462e-07,1.991463e-07,1.991464e-07,1.991466e-07,1.991467e-07,1.991468e-07,1.991469e-07,1.991471e-07,1.991472e-07,1.991473e-07,1.991474e-07,1.991476e-07,1.991477e-07,1.991478e-07,1.991479e-07,1.991481e-07,1.991482e-07,1.991483e-07,1.991484e-07,1.991486e-07,1.991487e-07,1.991488e-07,1.991489e-07,1.991491e-07,1.991492e-07,1.991493e-07,1.991495e-07,1.991496e-07,1.991497e-07,1.991498e-07,1.991500e-07,1.991501e-07,1.991502e-07,1.991503e-07,1.991505e-07,1.991506e-07,1.991507e-07,1.991508e-07,1.991510e-07,1.991511e-07,1.991512e-07,1.991513e-07,1.991515e-07,1.991516e-07,1.991517e-07,1.991518e-07,1.991520e-07,1.991521e-07,1.991522e-07,1.991523e-07,1.991525e-07,1.991526e-07,1.991527e-07,1.991528e-07,1.991530e-07,1.991531e-07,1.991532e-07,1.991533e-07,1.991535e-07,1.991536e-07,1.991537e-07,1.991538e-07,1.991540e-07,1.991541e-07,1.991542e-07,1.991543e-07,1.991545e-07,1.991546e-07,1.991547e-07,1.991549e-07,1.991550e-07,1.991551e-07,1.991552e-07,1.991554e-07,1.991555e-07,1.991556e-07,1.991557e-07,1.991559e-07,1.991560e-07,1.991561e-07,1.991562e-07,1.991564e-07,1.991565e-07,1.991566e-07,1.991567e-07,1.991569e-07,1.991570e-07,1.991571e-07,1.991572e-07,1.991574e-07,1.991575e-07,1.991576e-07,1.991577e-07,1.991579e-07,1.991580e-07,1.991581e-07,1.991582e-07,1.991584e-07,1.991585e-07,1.991586e-07,1.991587e-07,1.991589e-07,1.991590e-07,1.991591e-07,1.991592e-07,1.991594e-07,1.991595e-07,1.991596e-07,1.991597e-07,1.991599e-07,1.991600e-07,1.991601e-07,1.991602e-07,1.991604e-07,1.991605e-07,1.991606e-07,1.991608e-07,1.991609e-07,1.991610e-07,1.991611e-07,1.991613e-07,1.991614e-07,1.991615e-07,1.991616e-07,1.991618e-07,1.991619e-07,1.991620e-07,1.991621e-07,1.991623e-07,1.991624e-07,1.991625e-07,1.991626e-07,1.991628e-07,1.991629e-07,1.991630e-07,1.991631e-07,1.991633e-07,1.991634e-07,1.991635e-07,1.991636e-07,1.991638e-07,1.991639e-07,1.991640e-07,1.991641e-07,1.991643e-07,1.991644e-07,1.991645e-07,1.991646e-07,1.991648e-07,1.991649e-07,1.991650e-07,1.991651e-07,1.991653e-07,1.991654e-07,1.991655e-07,1.991656e-07,1.991658e-07,1.991659e-07,1.991660e-07,1.991661e-07,1.991663e-07,1.991664e-07,1.991665e-07,1.991666e-07,1.991668e-07,1.991669e-07,1.991670e-07,1.991672e-07,1.991673e-07,1.991674e-07,1.991675e-07,1.991677e-07,1.991678e-07,1.991679e-07,1.991680e-07,1.991682e-07,1.991683e-07,1.991684e-07,1.991685e-07,1.991687e-07,1.991688e-07,1.991689e-07,1.991690e-07,1.991692e-07,1.991693e-07,1.991694e-07,1.991695e-07,1.991697e-07,1.991698e-07,1.991699e-07,1.991700e-07,1.991702e-07,1.991703e-07,1.991704e-07,1.991705e-07,1.991707e-07,1.991708e-07,1.991709e-07,1.991710e-07,1.991712e-07,1.991713e-07,1.991714e-07,1.991715e-07,1.991717e-07,1.991718e-07,1.991719e-07,1.991720e-07,1.991722e-07,1.991723e-07,1.991724e-07,1.991725e-07,1.991727e-07,1.991728e-07,1.991729e-07,1.991730e-07,1.991732e-07,1.991733e-07,1.991734e-07,1.991735e-07,1.991737e-07,1.991738e-07,1.991739e-07,1.991740e-07,1.991742e-07,1.991743e-07,1.991744e-07,1.991745e-07,1.991747e-07,1.991748e-07,1.991749e-07,1.991751e-07,1.991752e-07,1.991753e-07,1.991754e-07,1.991756e-07,1.991757e-07,1.991758e-07,1.991759e-07,1.991761e-07,1.991762e-07,1.991763e-07,1.991764e-07,1.991766e-07,1.991767e-07,1.991768e-07,1.991769e-07,1.991771e-07,1.991772e-07,1.991773e-07,1.991774e-07,1.991776e-07,1.991777e-07,1.991778e-07,1.991779e-07,1.991781e-07,1.991782e-07,1.991783e-07,1.991784e-07,1.991786e-07,1.991787e-07,1.991788e-07,1.991789e-07,1.991791e-07,1.991792e-07,1.991793e-07,1.991794e-07,1.991796e-07,1.991797e-07,1.991798e-07,1.991799e-07,1.991801e-07,1.991802e-07,1.991803e-07,1.991804e-07,1.991806e-07,1.991807e-07,1.991808e-07,1.991809e-07,1.991811e-07,1.991812e-07,1.991813e-07,1.991814e-07,1.991816e-07,1.991817e-07,1.991818e-07,1.991819e-07,1.991821e-07,1.991822e-07,1.991823e-07,1.991824e-07,1.991826e-07,1.991827e-07,1.991828e-07,1.991829e-07,1.991831e-07,1.991832e-07,1.991833e-07,1.991834e-07,1.991836e-07,1.991837e-07,1.991838e-07,1.991839e-07,1.991841e-07,1.991842e-07,1.991843e-07,1.991844e-07,1.991846e-07,1.991847e-07,1.991848e-07,1.991849e-07,1.991851e-07,1.991852e-07,1.991853e-07,1.991855e-07,1.991856e-07,1.991857e-07,1.991858e-07,1.991860e-07,1.991861e-07,1.991862e-07,1.991863e-07,1.991865e-07,1.991866e-07,1.991867e-07,1.991868e-07,1.991870e-07,1.991871e-07,1.991872e-07,1.991873e-07,1.991875e-07,1.991876e-07,1.991877e-07,1.991878e-07,1.991880e-07,1.991881e-07,1.991882e-07,1.991883e-07,1.991885e-07,1.991886e-07,1.991887e-07,1.991888e-07,1.991890e-07,1.991891e-07,1.991892e-07,1.991893e-07,1.991895e-07,1.991896e-07,1.991897e-07,1.991898e-07,1.991900e-07,1.991901e-07,1.991902e-07,1.991903e-07,1.991905e-07,1.991906e-07,1.991907e-07,1.991908e-07,1.991910e-07,1.991911e-07,1.991912e-07,1.991913e-07,1.991915e-07,1.991916e-07,1.991917e-07,1.991918e-07,1.991920e-07,1.991921e-07,1.991922e-07,1.991923e-07,1.991925e-07,1.991926e-07,1.991927e-07,1.991928e-07,1.991930e-07,1.991931e-07,1.991932e-07,1.991933e-07,1.991935e-07,1.991936e-07,1.991937e-07,1.991938e-07,1.991940e-07,1.991941e-07,1.991942e-07,1.991943e-07,1.991945e-07,1.991946e-07,1.991947e-07,1.991948e-07,1.991950e-07,1.991951e-07,1.991952e-07,1.991953e-07,1.991955e-07,1.991956e-07,1.991957e-07,1.991958e-07,1.991960e-07,1.991961e-07,1.991962e-07,1.991963e-07,1.991965e-07,1.991966e-07,1.991967e-07,1.991968e-07,1.991970e-07,1.991971e-07,1.991972e-07,1.991973e-07,1.991975e-07,1.991976e-07,1.991977e-07,1.991978e-07,1.991980e-07,1.991981e-07,1.991982e-07,1.991983e-07,1.991985e-07,1.991986e-07,1.991987e-07,1.991988e-07,1.991990e-07,1.991991e-07,1.991992e-07,1.991993e-07,1.991995e-07,1.991996e-07,1.991997e-07,1.991998e-07,1.992000e-07,1.992001e-07,1.992002e-07,1.992003e-07,1.992005e-07,1.992006e-07,1.992007e-07,1.992008e-07,1.992010e-07,1.992011e-07,1.992012e-07,1.992013e-07,1.992015e-07,1.992016e-07,1.992017e-07,1.992018e-07,1.992020e-07,1.992021e-07,1.992022e-07,1.992023e-07,1.992025e-07,1.992026e-07,1.992027e-07,1.992028e-07,1.992030e-07,1.992031e-07,1.992032e-07,1.992033e-07,1.992035e-07,1.992036e-07,1.992037e-07,1.992038e-07,1.992040e-07,1.992041e-07,1.992042e-07,1.992043e-07,1.992045e-07,1.992046e-07,1.992047e-07,1.992048e-07,1.992050e-07,1.992051e-07,1.992052e-07,1.992053e-07,1.992055e-07,1.992056e-07,1.992057e-07,1.992058e-07,1.992060e-07,1.992061e-07,1.992062e-07,1.992063e-07,1.992065e-07,1.992066e-07,1.992067e-07,1.992068e-07,1.992070e-07,1.992071e-07,1.992072e-07,1.992073e-07,1.992075e-07,1.992076e-07,1.992077e-07,1.992078e-07,1.992080e-07,1.992081e-07,1.992082e-07,1.992083e-07,1.992085e-07,1.992086e-07,1.992087e-07,1.992088e-07,1.992090e-07,1.992091e-07,1.992092e-07,1.992093e-07,1.992095e-07,1.992096e-07,1.992097e-07,1.992098e-07,1.992100e-07,1.992101e-07,1.992102e-07,1.992103e-07,1.992105e-07,1.992106e-07,1.992107e-07,1.992108e-07,1.992110e-07,1.992111e-07,1.992112e-07,1.992113e-07,1.992115e-07,1.992116e-07,1.992117e-07,1.992118e-07,1.992120e-07,1.992121e-07,1.992122e-07,1.992123e-07,1.992125e-07,1.992126e-07,1.992127e-07,1.992128e-07,1.992130e-07,1.992131e-07,1.992132e-07,1.992133e-07,1.992135e-07,1.992136e-07,1.992137e-07,1.992138e-07,1.992140e-07,1.992141e-07,1.992142e-07,1.992143e-07,1.992145e-07,1.992146e-07,1.992147e-07,1.992148e-07,1.992150e-07,1.992151e-07,1.992152e-07,1.992153e-07,1.992155e-07,1.992156e-07,1.992157e-07,1.992158e-07,1.992160e-07,1.992161e-07,1.992162e-07,1.992163e-07,1.992165e-07,1.992166e-07,1.992167e-07,1.992168e-07,1.992170e-07,1.992171e-07,1.992172e-07,1.992173e-07,1.992175e-07,1.992176e-07,1.992177e-07,1.992178e-07,1.992180e-07,1.992181e-07,1.992182e-07,1.992183e-07,1.992185e-07,1.992186e-07,1.992187e-07,1.992188e-07,1.992190e-07,1.992191e-07,1.992192e-07,1.992193e-07,1.992195e-07,1.992196e-07,1.992197e-07,1.992198e-07,1.992200e-07,1.992201e-07,1.992202e-07,1.992203e-07,1.992205e-07,1.992206e-07,1.992207e-07,1.992208e-07,1.992210e-07,1.992211e-07,1.992212e-07,1.992213e-07,1.992215e-07,1.992216e-07,1.992217e-07,1.992218e-07,1.992220e-07,1.992221e-07,1.992222e-07,1.992223e-07,1.992225e-07,1.992226e-07,1.992227e-07,1.992228e-07,1.992230e-07,1.992231e-07,1.992232e-07,1.992233e-07,1.992235e-07,1.992236e-07,1.992237e-07,1.992238e-07,1.992240e-07,1.992241e-07,1.992242e-07,1.992243e-07,1.992245e-07,1.992246e-07,1.992247e-07,1.992248e-07,1.992250e-07,1.992251e-07,1.992252e-07,1.992253e-07,1.992255e-07,1.992256e-07,1.992257e-07,1.992258e-07,1.992260e-07,1.992261e-07,1.992262e-07,1.992263e-07,1.992265e-07,1.992266e-07,1.992267e-07,1.992268e-07,1.992270e-07,1.992271e-07,1.992272e-07,1.992273e-07,1.992275e-07,1.992276e-07,1.992277e-07,1.992278e-07,1.992280e-07,1.992281e-07,1.992282e-07,1.992283e-07,1.992285e-07,1.992286e-07,1.992287e-07,1.992288e-07,1.992290e-07,1.992291e-07,1.992292e-07,1.992293e-07,1.992295e-07,1.992296e-07,1.992297e-07,1.992298e-07,1.992300e-07,1.992301e-07,1.992302e-07,1.992303e-07,1.992305e-07,1.992306e-07,1.992307e-07,1.992308e-07,1.992310e-07,1.992311e-07,1.992312e-07,1.992313e-07,1.992314e-07,1.992316e-07,1.992317e-07,1.992318e-07,1.992319e-07,1.992321e-07,1.992322e-07,1.992323e-07,1.992324e-07,1.992326e-07,1.992327e-07,1.992328e-07,1.992329e-07,1.992331e-07,1.992332e-07,1.992333e-07,1.992334e-07,1.992336e-07,1.992337e-07,1.992338e-07,1.992339e-07,1.992341e-07,1.992342e-07,1.992343e-07,1.992344e-07,1.992346e-07,1.992347e-07,1.992348e-07,1.992349e-07,1.992351e-07,1.992352e-07,1.992353e-07,1.992354e-07,1.992356e-07,1.992357e-07,1.992358e-07,1.992359e-07,1.992361e-07,1.992362e-07,1.992363e-07,1.992364e-07,1.992366e-07,1.992367e-07,1.992368e-07,1.992369e-07,1.992371e-07,1.992372e-07,1.992373e-07,1.992374e-07,1.992376e-07,1.992377e-07,1.992378e-07,1.992379e-07,1.992381e-07,1.992382e-07,1.992383e-07,1.992384e-07,1.992386e-07,1.992387e-07,1.992388e-07,1.992389e-07,1.992391e-07,1.992392e-07,1.992393e-07,1.992394e-07,1.992396e-07,1.992397e-07,1.992398e-07,1.992399e-07,1.992401e-07,1.992402e-07,1.992403e-07,1.992404e-07,1.992406e-07,1.992407e-07,1.992408e-07,1.992409e-07,1.992411e-07,1.992412e-07,1.992413e-07,1.992414e-07,1.992416e-07,1.992417e-07,1.992418e-07,1.992419e-07,1.992420e-07,1.992422e-07,1.992423e-07,1.992424e-07,1.992425e-07,1.992427e-07,1.992428e-07,1.992429e-07,1.992430e-07,1.992432e-07,1.992433e-07,1.992434e-07,1.992435e-07,1.992437e-07,1.992438e-07,1.992439e-07,1.992440e-07,1.992442e-07,1.992443e-07,1.992444e-07,1.992445e-07,1.992447e-07,1.992448e-07,1.992449e-07,1.992450e-07,1.992452e-07,1.992453e-07,1.992454e-07,1.992455e-07,1.992457e-07,1.992458e-07,1.992459e-07,1.992460e-07,1.992462e-07,1.992463e-07,1.992464e-07,1.992465e-07,1.992467e-07,1.992468e-07,1.992469e-07,1.992470e-07,1.992472e-07,1.992473e-07,1.992474e-07,1.992475e-07,1.992477e-07,1.992478e-07,1.992479e-07,1.992480e-07,1.992482e-07,1.992483e-07,1.992484e-07,1.992485e-07,1.992487e-07,1.992488e-07,1.992489e-07,1.992490e-07,1.992492e-07,1.992493e-07,1.992494e-07,1.992495e-07,1.992496e-07,1.992498e-07,1.992499e-07,1.992500e-07,1.992501e-07,1.992503e-07,1.992504e-07,1.992505e-07,1.992506e-07,1.992508e-07,1.992509e-07,1.992510e-07,1.992511e-07,1.992513e-07,1.992514e-07,1.992515e-07,1.992516e-07,1.992518e-07,1.992519e-07,1.992520e-07,1.992521e-07,1.992523e-07,1.992524e-07,1.992525e-07,1.992526e-07,1.992528e-07,1.992529e-07,1.992530e-07,1.992531e-07,1.992533e-07,1.992534e-07,1.992535e-07,1.992536e-07,1.992538e-07,1.992539e-07,1.992540e-07,1.992541e-07,1.992543e-07,1.992544e-07,1.992545e-07,1.992546e-07,1.992548e-07,1.992549e-07,1.992550e-07,1.992551e-07,1.992553e-07,1.992554e-07,1.992555e-07,1.992556e-07,1.992558e-07,1.992559e-07,1.992560e-07,1.992561e-07,1.992562e-07,1.992564e-07,1.992565e-07,1.992566e-07,1.992567e-07,1.992569e-07,1.992570e-07,1.992571e-07,1.992572e-07,1.992574e-07,1.992575e-07,1.992576e-07,1.992577e-07,1.992579e-07,1.992580e-07,1.992581e-07,1.992582e-07,1.992584e-07,1.992585e-07,1.992586e-07,1.992587e-07,1.992589e-07,1.992590e-07,1.992591e-07,1.992592e-07,1.992594e-07,1.992595e-07,1.992596e-07,1.992597e-07,1.992599e-07,1.992600e-07,1.992601e-07,1.992602e-07,1.992604e-07,1.992605e-07,1.992606e-07,1.992607e-07,1.992609e-07,1.992610e-07,1.992611e-07,1.992612e-07,1.992614e-07,1.992615e-07,1.992616e-07,1.992617e-07,1.992619e-07,1.992620e-07,1.992621e-07,1.992622e-07,1.992623e-07,1.992625e-07,1.992626e-07,1.992627e-07,1.992628e-07,1.992630e-07,1.992631e-07,1.992632e-07,1.992633e-07,1.992635e-07,1.992636e-07,1.992637e-07,1.992638e-07,1.992640e-07,1.992641e-07,1.992642e-07,1.992643e-07,1.992645e-07,1.992646e-07,1.992647e-07,1.992648e-07,1.992650e-07,1.992651e-07,1.992652e-07,1.992653e-07,1.992655e-07,1.992656e-07,1.992657e-07,1.992658e-07,1.992660e-07,1.992661e-07,1.992662e-07,1.992663e-07,1.992665e-07,1.992666e-07,1.992667e-07,1.992668e-07,1.992670e-07,1.992671e-07,1.992672e-07,1.992673e-07,1.992674e-07,1.992676e-07,1.992677e-07,1.992678e-07,1.992679e-07,1.992681e-07,1.992682e-07,1.992683e-07,1.992684e-07,1.992686e-07,1.992687e-07,1.992688e-07,1.992689e-07,1.992691e-07,1.992692e-07,1.992693e-07,1.992694e-07,1.992696e-07,1.992697e-07,1.992698e-07,1.992699e-07,1.992701e-07,1.992702e-07,1.992703e-07,1.992704e-07,1.992706e-07,1.992707e-07,1.992708e-07,1.992709e-07,1.992711e-07,1.992712e-07,1.992713e-07,1.992714e-07,1.992716e-07,1.992717e-07,1.992718e-07,1.992719e-07,1.992720e-07,1.992722e-07,1.992723e-07,1.992724e-07,1.992725e-07,1.992727e-07,1.992728e-07,1.992729e-07,1.992730e-07,1.992732e-07,1.992733e-07,1.992734e-07,1.992735e-07,1.992737e-07,1.992738e-07,1.992739e-07,1.992740e-07,1.992742e-07,1.992743e-07,1.992744e-07,1.992745e-07,1.992747e-07,1.992748e-07,1.992749e-07,1.992750e-07,1.992752e-07,1.992753e-07,1.992754e-07,1.992755e-07,1.992757e-07,1.992758e-07,1.992759e-07,1.992760e-07,1.992762e-07,1.992763e-07,1.992764e-07,1.992765e-07,1.992766e-07,1.992768e-07,1.992769e-07,1.992770e-07,1.992771e-07,1.992773e-07,1.992774e-07,1.992775e-07,1.992776e-07,1.992778e-07,1.992779e-07,1.992780e-07,1.992781e-07,1.992783e-07,1.992784e-07,1.992785e-07,1.992786e-07,1.992788e-07,1.992789e-07,1.992790e-07,1.992791e-07,1.992793e-07,1.992794e-07,1.992795e-07,1.992796e-07,1.992798e-07,1.992799e-07,1.992800e-07,1.992801e-07,1.992803e-07,1.992804e-07,1.992805e-07,1.992806e-07,1.992807e-07,1.992809e-07,1.992810e-07,1.992811e-07,1.992812e-07,1.992814e-07,1.992815e-07,1.992816e-07,1.992817e-07,1.992819e-07,1.992820e-07,1.992821e-07,1.992822e-07,1.992824e-07,1.992825e-07,1.992826e-07,1.992827e-07,1.992829e-07,1.992830e-07,1.992831e-07,1.992832e-07,1.992834e-07,1.992835e-07,1.992836e-07,1.992837e-07,1.992839e-07,1.992840e-07,1.992841e-07,1.992842e-07,1.992844e-07,1.992845e-07,1.992846e-07,1.992847e-07,1.992848e-07,1.992850e-07,1.992851e-07,1.992852e-07,1.992853e-07,1.992855e-07,1.992856e-07,1.992857e-07,1.992858e-07,1.992860e-07,1.992861e-07,1.992862e-07,1.992863e-07,1.992865e-07,1.992866e-07,1.992867e-07,1.992868e-07,1.992870e-07,1.992871e-07,1.992872e-07,1.992873e-07,1.992875e-07,1.992876e-07,1.992877e-07,1.992878e-07,1.992880e-07,1.992881e-07,1.992882e-07,1.992883e-07,1.992884e-07,1.992886e-07,1.992887e-07,1.992888e-07,1.992889e-07,1.992891e-07,1.992892e-07,1.992893e-07,1.992894e-07,1.992896e-07,1.992897e-07,1.992898e-07,1.992899e-07,1.992901e-07,1.992902e-07,1.992903e-07,1.992904e-07,1.992906e-07,1.992907e-07,1.992908e-07,1.992909e-07,1.992911e-07,1.992912e-07,1.992913e-07,1.992914e-07,1.992916e-07,1.992917e-07,1.992918e-07,1.992919e-07,1.992920e-07,1.992922e-07,1.992923e-07,1.992924e-07,1.992925e-07,1.992927e-07,1.992928e-07,1.992929e-07,1.992930e-07,1.992932e-07,1.992933e-07,1.992934e-07,1.992935e-07,1.992937e-07,1.992938e-07,1.992939e-07,1.992940e-07,1.992942e-07,1.992943e-07,1.992944e-07,1.992945e-07,1.992947e-07,1.992948e-07,1.992949e-07,1.992950e-07,1.992952e-07,1.992953e-07,1.992954e-07,1.992955e-07,1.992956e-07,1.992958e-07,1.992959e-07,1.992960e-07,1.992961e-07,1.992963e-07,1.992964e-07,1.992965e-07,1.992966e-07,1.992968e-07,1.992969e-07,1.992970e-07,1.992971e-07,1.992973e-07,1.992974e-07,1.992975e-07,1.992976e-07,1.992978e-07,1.992979e-07,1.992980e-07,1.992981e-07,1.992983e-07,1.992984e-07,1.992985e-07,1.992986e-07,1.992987e-07,1.992989e-07,1.992990e-07,1.992991e-07,1.992992e-07,1.992994e-07,1.992995e-07,1.992996e-07,1.992997e-07,1.992999e-07,1.993000e-07,1.993001e-07,1.993002e-07,1.993004e-07,1.993005e-07,1.993006e-07,1.993007e-07,1.993009e-07,1.993010e-07,1.993011e-07,1.993012e-07,1.993014e-07,1.993015e-07,1.993016e-07,1.993017e-07,1.993018e-07,1.993020e-07,1.993021e-07,1.993022e-07,1.993023e-07,1.993025e-07,1.993026e-07,1.993027e-07,1.993028e-07,1.993030e-07,1.993031e-07,1.993032e-07,1.993033e-07,1.993035e-07,1.993036e-07,1.993037e-07,1.993038e-07,1.993040e-07,1.993041e-07,1.993042e-07,1.993043e-07,1.993045e-07,1.993046e-07,1.993047e-07,1.993048e-07,1.993049e-07,1.993051e-07,1.993052e-07,1.993053e-07,1.993054e-07,1.993056e-07,1.993057e-07,1.993058e-07,1.993059e-07,1.993061e-07,1.993062e-07,1.993063e-07,1.993064e-07,1.993066e-07,1.993067e-07,1.993068e-07,1.993069e-07,1.993071e-07,1.993072e-07,1.993073e-07,1.993074e-07,1.993076e-07,1.993077e-07,1.993078e-07,1.993079e-07,1.993080e-07,1.993082e-07,1.993083e-07,1.993084e-07,1.993085e-07,1.993087e-07,1.993088e-07,1.993089e-07,1.993090e-07,1.993092e-07,1.993093e-07,1.993094e-07,1.993095e-07,1.993097e-07,1.993098e-07,1.993099e-07,1.993100e-07,1.993102e-07,1.993103e-07,1.993104e-07,1.993105e-07,1.993106e-07,1.993108e-07,1.993109e-07,1.993110e-07,1.993111e-07,1.993113e-07,1.993114e-07,1.993115e-07,1.993116e-07,1.993118e-07,1.993119e-07,1.993120e-07,1.993121e-07,1.993123e-07,1.993124e-07,1.993125e-07,1.993126e-07,1.993128e-07,1.993129e-07,1.993130e-07,1.993131e-07,1.993133e-07,1.993134e-07,1.993135e-07,1.993136e-07,1.993137e-07,1.993139e-07,1.993140e-07,1.993141e-07,1.993142e-07,1.993144e-07,1.993145e-07,1.993146e-07,1.993147e-07,1.993149e-07,1.993150e-07,1.993151e-07,1.993152e-07,1.993154e-07,1.993155e-07,1.993156e-07,1.993157e-07,1.993159e-07,1.993160e-07,1.993161e-07,1.993162e-07,1.993163e-07,1.993165e-07,1.993166e-07,1.993167e-07,1.993168e-07,1.993170e-07,1.993171e-07,1.993172e-07,1.993173e-07,1.993175e-07,1.993176e-07,1.993177e-07,1.993178e-07,1.993180e-07,1.993181e-07,1.993182e-07,1.993183e-07,1.993185e-07,1.993186e-07,1.993187e-07,1.993188e-07,1.993189e-07,1.993191e-07,1.993192e-07,1.993193e-07,1.993194e-07,1.993196e-07,1.993197e-07,1.993198e-07,1.993199e-07,1.993201e-07,1.993202e-07,1.993203e-07,1.993204e-07,1.993206e-07,1.993207e-07,1.993208e-07,1.993209e-07,1.993211e-07,1.993212e-07,1.993213e-07,1.993214e-07,1.993215e-07,1.993217e-07,1.993218e-07,1.993219e-07,1.993220e-07,1.993222e-07,1.993223e-07,1.993224e-07,1.993225e-07,1.993227e-07,1.993228e-07,1.993229e-07,1.993230e-07,1.993232e-07,1.993233e-07,1.993234e-07,1.993235e-07,1.993237e-07,1.993238e-07,1.993239e-07,1.993240e-07,1.993241e-07,1.993243e-07,1.993244e-07,1.993245e-07,1.993246e-07,1.993248e-07,1.993249e-07,1.993250e-07,1.993251e-07,1.993253e-07,1.993254e-07,1.993255e-07,1.993256e-07,1.993258e-07,1.993259e-07,1.993260e-07,1.993261e-07,1.993263e-07,1.993264e-07,1.993265e-07,1.993266e-07,1.993267e-07,1.993269e-07,1.993270e-07,1.993271e-07,1.993272e-07,1.993274e-07,1.993275e-07,1.993276e-07,1.993277e-07,1.993279e-07,1.993280e-07,1.993281e-07,1.993282e-07,1.993284e-07,1.993285e-07,1.993286e-07,1.993287e-07,1.993289e-07,1.993290e-07,1.993291e-07,1.993292e-07,1.993293e-07,1.993295e-07,1.993296e-07,1.993297e-07,1.993298e-07,1.993300e-07,1.993301e-07,1.993302e-07,1.993303e-07,1.993305e-07,1.993306e-07,1.993307e-07,1.993308e-07,1.993310e-07,1.993311e-07,1.993312e-07,1.993313e-07,1.993314e-07,1.993316e-07,1.993317e-07,1.993318e-07,1.993319e-07,1.993321e-07,1.993322e-07,1.993323e-07,1.993324e-07,1.993326e-07,1.993327e-07,1.993328e-07,1.993329e-07,1.993331e-07,1.993332e-07,1.993333e-07,1.993334e-07,1.993336e-07,1.993337e-07,1.993338e-07,1.993339e-07,1.993340e-07,1.993342e-07,1.993343e-07,1.993344e-07,1.993345e-07,1.993347e-07,1.993348e-07,1.993349e-07,1.993350e-07,1.993352e-07,1.993353e-07,1.993354e-07,1.993355e-07,1.993357e-07,1.993358e-07,1.993359e-07,1.993360e-07,1.993361e-07,1.993363e-07,1.993364e-07,1.993365e-07,1.993366e-07,1.993368e-07,1.993369e-07,1.993370e-07,1.993371e-07,1.993373e-07,1.993374e-07,1.993375e-07,1.993376e-07,1.993378e-07,1.993379e-07,1.993380e-07,1.993381e-07,1.993382e-07,1.993384e-07,1.993385e-07,1.993386e-07,1.993387e-07,1.993389e-07,1.993390e-07,1.993391e-07,1.993392e-07,1.993394e-07,1.993395e-07,1.993396e-07,1.993397e-07,1.993399e-07,1.993400e-07,1.993401e-07,1.993402e-07,1.993404e-07,1.993405e-07,1.993406e-07,1.993407e-07,1.993408e-07,1.993410e-07,1.993411e-07,1.993412e-07,1.993413e-07,1.993415e-07,1.993416e-07,1.993417e-07,1.993418e-07,1.993420e-07,1.993421e-07,1.993422e-07,1.993423e-07,1.993425e-07,1.993426e-07,1.993427e-07,1.993428e-07,1.993429e-07,1.993431e-07,1.993432e-07,1.993433e-07,1.993434e-07,1.993436e-07,1.993437e-07,1.993438e-07,1.993439e-07,1.993441e-07,1.993442e-07,1.993443e-07,1.993444e-07,1.993446e-07,1.993447e-07,1.993448e-07,1.993449e-07,1.993450e-07,1.993452e-07,1.993453e-07,1.993454e-07,1.993455e-07,1.993457e-07,1.993458e-07,1.993459e-07,1.993460e-07,1.993462e-07,1.993463e-07,1.993464e-07,1.993465e-07,1.993467e-07,1.993468e-07,1.993469e-07,1.993470e-07,1.993471e-07,1.993473e-07,1.993474e-07,1.993475e-07,1.993476e-07,1.993478e-07,1.993479e-07,1.993480e-07,1.993481e-07,1.993483e-07,1.993484e-07,1.993485e-07,1.993486e-07,1.993488e-07,1.993489e-07,1.993490e-07,1.993491e-07,1.993492e-07,1.993494e-07,1.993495e-07,1.993496e-07,1.993497e-07,1.993499e-07,1.993500e-07,1.993501e-07,1.993502e-07,1.993504e-07,1.993505e-07,1.993506e-07,1.993507e-07,1.993509e-07,1.993510e-07,1.993511e-07,1.993512e-07,1.993513e-07,1.993515e-07,1.993516e-07,1.993517e-07,1.993518e-07,1.993520e-07,1.993521e-07,1.993522e-07,1.993523e-07,1.993525e-07,1.993526e-07,1.993527e-07,1.993528e-07,1.993530e-07,1.993531e-07,1.993532e-07,1.993533e-07,1.993534e-07,1.993536e-07,1.993537e-07,1.993538e-07,1.993539e-07,1.993541e-07,1.993542e-07,1.993543e-07,1.993544e-07,1.993546e-07,1.993547e-07,1.993548e-07,1.993549e-07,1.993551e-07,1.993552e-07,1.993553e-07,1.993554e-07,1.993555e-07,1.993557e-07,1.993558e-07,1.993559e-07,1.993560e-07,1.993562e-07,1.993563e-07,1.993564e-07,1.993565e-07,1.993567e-07,1.993568e-07,1.993569e-07,1.993570e-07,1.993571e-07,1.993573e-07,1.993574e-07,1.993575e-07,1.993576e-07,1.993578e-07,1.993579e-07,1.993580e-07,1.993581e-07,1.993583e-07,1.993584e-07,1.993585e-07,1.993586e-07,1.993588e-07,1.993589e-07,1.993590e-07,1.993591e-07,1.993592e-07,1.993594e-07,1.993595e-07,1.993596e-07,1.993597e-07,1.993599e-07,1.993600e-07,1.993601e-07,1.993602e-07,1.993604e-07,1.993605e-07,1.993606e-07,1.993607e-07,1.993609e-07,1.993610e-07,1.993611e-07,1.993612e-07,1.993613e-07,1.993615e-07,1.993616e-07,1.993617e-07,1.993618e-07,1.993620e-07,1.993621e-07,1.993622e-07,1.993623e-07,1.993625e-07,1.993626e-07,1.993627e-07,1.993628e-07,1.993629e-07,1.993631e-07,1.993632e-07,1.993633e-07,1.993634e-07,1.993636e-07,1.993637e-07,1.993638e-07,1.993639e-07,1.993641e-07,1.993642e-07,1.993643e-07,1.993644e-07,1.993646e-07,1.993647e-07,1.993648e-07,1.993649e-07,1.993650e-07,1.993652e-07,1.993653e-07,1.993654e-07,1.993655e-07,1.993657e-07,1.993658e-07,1.993659e-07,1.993660e-07,1.993662e-07,1.993663e-07,1.993664e-07,1.993665e-07,1.993666e-07,1.993668e-07,1.993669e-07,1.993670e-07,1.993671e-07,1.993673e-07,1.993674e-07,1.993675e-07,1.993676e-07,1.993678e-07,1.993679e-07,1.993680e-07,1.993681e-07,1.993683e-07,1.993684e-07,1.993685e-07,1.993686e-07,1.993687e-07,1.993689e-07,1.993690e-07,1.993691e-07,1.993692e-07,1.993694e-07,1.993695e-07,1.993696e-07,1.993697e-07,1.993699e-07,1.993700e-07,1.993701e-07,1.993702e-07,1.993703e-07,1.993705e-07,1.993706e-07,1.993707e-07,1.993708e-07,1.993710e-07,1.993711e-07,1.993712e-07,1.993713e-07,1.993715e-07,1.993716e-07,1.993717e-07,1.993718e-07,1.993719e-07,1.993721e-07,1.993722e-07,1.993723e-07,1.993724e-07,1.993726e-07,1.993727e-07,1.993728e-07,1.993729e-07,1.993731e-07,1.993732e-07,1.993733e-07,1.993734e-07,1.993736e-07,1.993737e-07,1.993738e-07,1.993739e-07,1.993740e-07,1.993742e-07,1.993743e-07,1.993744e-07,1.993745e-07,1.993747e-07,1.993748e-07,1.993749e-07,1.993750e-07,1.993752e-07,1.993753e-07,1.993754e-07,1.993755e-07,1.993756e-07,1.993758e-07,1.993759e-07,1.993760e-07,1.993761e-07,1.993763e-07,1.993764e-07,1.993765e-07,1.993766e-07,1.993768e-07,1.993769e-07,1.993770e-07,1.993771e-07,1.993772e-07,1.993774e-07,1.993775e-07,1.993776e-07,1.993777e-07,1.993779e-07,1.993780e-07,1.993781e-07,1.993782e-07,1.993784e-07,1.993785e-07,1.993786e-07,1.993787e-07,1.993789e-07,1.993790e-07,1.993791e-07,1.993792e-07,1.993793e-07,1.993795e-07,1.993796e-07,1.993797e-07,1.993798e-07,1.993800e-07,1.993801e-07,1.993802e-07,1.993803e-07,1.993805e-07,1.993806e-07,1.993807e-07,1.993808e-07,1.993809e-07,1.993811e-07,1.993812e-07,1.993813e-07,1.993814e-07,1.993816e-07,1.993817e-07,1.993818e-07,1.993819e-07,1.993821e-07,1.993822e-07,1.993823e-07,1.993824e-07,1.993825e-07,1.993827e-07,1.993828e-07,1.993829e-07,1.993830e-07,1.993832e-07,1.993833e-07,1.993834e-07,1.993835e-07,1.993837e-07,1.993838e-07,1.993839e-07,1.993840e-07,1.993841e-07,1.993843e-07,1.993844e-07,1.993845e-07,1.993846e-07,1.993848e-07,1.993849e-07,1.993850e-07,1.993851e-07,1.993853e-07,1.993854e-07,1.993855e-07,1.993856e-07,1.993857e-07,1.993859e-07,1.993860e-07,1.993861e-07,1.993862e-07,1.993864e-07,1.993865e-07,1.993866e-07,1.993867e-07,1.993869e-07,1.993870e-07,1.993871e-07,1.993872e-07,1.993873e-07,1.993875e-07,1.993876e-07,1.993877e-07,1.993878e-07,1.993880e-07,1.993881e-07,1.993882e-07,1.993883e-07,1.993885e-07,1.993886e-07,1.993887e-07,1.993888e-07,1.993889e-07,1.993891e-07,1.993892e-07,1.993893e-07,1.993894e-07,1.993896e-07,1.993897e-07,1.993898e-07,1.993899e-07,1.993901e-07,1.993902e-07,1.993903e-07,1.993904e-07,1.993905e-07,1.993907e-07,1.993908e-07,1.993909e-07,1.993910e-07,1.993912e-07,1.993913e-07,1.993914e-07,1.993915e-07,1.993917e-07,1.993918e-07,1.993919e-07,1.993920e-07,1.993921e-07,1.993923e-07,1.993924e-07,1.993925e-07,1.993926e-07,1.993928e-07,1.993929e-07,1.993930e-07,1.993931e-07,1.993933e-07,1.993934e-07,1.993935e-07,1.993936e-07,1.993937e-07,1.993939e-07,1.993940e-07,1.993941e-07,1.993942e-07,1.993944e-07,1.993945e-07,1.993946e-07,1.993947e-07,1.993949e-07,1.993950e-07,1.993951e-07,1.993952e-07,1.993953e-07,1.993955e-07,1.993956e-07,1.993957e-07,1.993958e-07,1.993960e-07,1.993961e-07,1.993962e-07,1.993963e-07,1.993965e-07,1.993966e-07,1.993967e-07,1.993968e-07,1.993969e-07,1.993971e-07,1.993972e-07,1.993973e-07,1.993974e-07,1.993976e-07,1.993977e-07,1.993978e-07,1.993979e-07,1.993981e-07,1.993982e-07,1.993983e-07,1.993984e-07,1.993985e-07,1.993987e-07,1.993988e-07,1.993989e-07,1.993990e-07,1.993992e-07,1.993993e-07,1.993994e-07,1.993995e-07,1.993997e-07,1.993998e-07,1.993999e-07,1.994000e-07,1.994001e-07,1.994003e-07,1.994004e-07,1.994005e-07,1.994006e-07,1.994008e-07,1.994009e-07,1.994010e-07,1.994011e-07,1.994013e-07,1.994014e-07,1.994015e-07,1.994016e-07,1.994017e-07,1.994019e-07,1.994020e-07,1.994021e-07,1.994022e-07,1.994024e-07,1.994025e-07,1.994026e-07,1.994027e-07,1.994028e-07,1.994030e-07,1.994031e-07,1.994032e-07,1.994033e-07,1.994035e-07,1.994036e-07,1.994037e-07,1.994038e-07,1.994040e-07,1.994041e-07,1.994042e-07,1.994043e-07,1.994044e-07,1.994046e-07,1.994047e-07,1.994048e-07,1.994049e-07,1.994051e-07,1.994052e-07,1.994053e-07,1.994054e-07,1.994056e-07,1.994057e-07,1.994058e-07,1.994059e-07,1.994060e-07,1.994062e-07,1.994063e-07,1.994064e-07,1.994065e-07,1.994067e-07,1.994068e-07,1.994069e-07,1.994070e-07,1.994072e-07,1.994073e-07,1.994074e-07,1.994075e-07,1.994076e-07,1.994078e-07,1.994079e-07,1.994080e-07,1.994081e-07,1.994083e-07,1.994084e-07,1.994085e-07,1.994086e-07,1.994087e-07,1.994089e-07,1.994090e-07,1.994091e-07,1.994092e-07,1.994094e-07,1.994095e-07,1.994096e-07,1.994097e-07,1.994099e-07,1.994100e-07,1.994101e-07,1.994102e-07,1.994103e-07,1.994105e-07,1.994106e-07,1.994107e-07,1.994108e-07,1.994110e-07,1.994111e-07,1.994112e-07,1.994113e-07,1.994115e-07,1.994116e-07,1.994117e-07,1.994118e-07,1.994119e-07,1.994121e-07,1.994122e-07,1.994123e-07,1.994124e-07,1.994126e-07,1.994127e-07,1.994128e-07,1.994129e-07,1.994130e-07,1.994132e-07,1.994133e-07,1.994134e-07,1.994135e-07,1.994137e-07,1.994138e-07,1.994139e-07,1.994140e-07,1.994142e-07,1.994143e-07,1.994144e-07,1.994145e-07,1.994146e-07,1.994148e-07,1.994149e-07,1.994150e-07,1.994151e-07,1.994153e-07,1.994154e-07,1.994155e-07,1.994156e-07,1.994158e-07,1.994159e-07,1.994160e-07,1.994161e-07,1.994162e-07,1.994164e-07,1.994165e-07,1.994166e-07,1.994167e-07,1.994169e-07,1.994170e-07,1.994171e-07,1.994172e-07,1.994173e-07,1.994175e-07,1.994176e-07,1.994177e-07,1.994178e-07,1.994180e-07,1.994181e-07,1.994182e-07,1.994183e-07,1.994185e-07,1.994186e-07,1.994187e-07,1.994188e-07,1.994189e-07,1.994191e-07,1.994192e-07,1.994193e-07,1.994194e-07,1.994196e-07,1.994197e-07,1.994198e-07,1.994199e-07,1.994200e-07,1.994202e-07,1.994203e-07,1.994204e-07,1.994205e-07,1.994207e-07,1.994208e-07,1.994209e-07,1.994210e-07,1.994212e-07,1.994213e-07,1.994214e-07,1.994215e-07,1.994216e-07,1.994218e-07,1.994219e-07,1.994220e-07,1.994221e-07,1.994223e-07,1.994224e-07,1.994225e-07,1.994226e-07,1.994227e-07,1.994229e-07,1.994230e-07,1.994231e-07,1.994232e-07,1.994234e-07,1.994235e-07,1.994236e-07,1.994237e-07,1.994239e-07,1.994240e-07,1.994241e-07,1.994242e-07,1.994243e-07,1.994245e-07,1.994246e-07,1.994247e-07,1.994248e-07,1.994250e-07,1.994251e-07,1.994252e-07,1.994253e-07,1.994254e-07,1.994256e-07,1.994257e-07,1.994258e-07,1.994259e-07,1.994261e-07,1.994262e-07,1.994263e-07,1.994264e-07,1.994266e-07,1.994267e-07,1.994268e-07,1.994269e-07,1.994270e-07,1.994272e-07,1.994273e-07,1.994274e-07,1.994275e-07,1.994277e-07,1.994278e-07,1.994279e-07,1.994280e-07,1.994281e-07,1.994283e-07,1.994284e-07,1.994285e-07,1.994286e-07,1.994288e-07,1.994289e-07,1.994290e-07,1.994291e-07,1.994293e-07,1.994294e-07,1.994295e-07,1.994296e-07,1.994297e-07,1.994299e-07,1.994300e-07,1.994301e-07,1.994302e-07,1.994304e-07,1.994305e-07,1.994306e-07,1.994307e-07,1.994308e-07,1.994310e-07,1.994311e-07,1.994312e-07,1.994313e-07,1.994315e-07,1.994316e-07,1.994317e-07,1.994318e-07,1.994320e-07,1.994321e-07,1.994322e-07,1.994323e-07,1.994324e-07,1.994326e-07,1.994327e-07,1.994328e-07,1.994329e-07,1.994331e-07,1.994332e-07,1.994333e-07,1.994334e-07,1.994335e-07,1.994337e-07,1.994338e-07,1.994339e-07,1.994340e-07,1.994342e-07,1.994343e-07,1.994344e-07,1.994345e-07,1.994346e-07,1.994348e-07,1.994349e-07,1.994350e-07,1.994351e-07,1.994353e-07,1.994354e-07,1.994355e-07,1.994356e-07,1.994358e-07,1.994359e-07,1.994360e-07,1.994361e-07,1.994362e-07,1.994364e-07,1.994365e-07,1.994366e-07,1.994367e-07,1.994369e-07,1.994370e-07,1.994371e-07,1.994372e-07,1.994373e-07,1.994375e-07,1.994376e-07,1.994377e-07,1.994378e-07,1.994380e-07,1.994381e-07,1.994382e-07,1.994383e-07,1.994384e-07,1.994386e-07,1.994387e-07,1.994388e-07,1.994389e-07,1.994391e-07,1.994392e-07,1.994393e-07,1.994394e-07,1.994396e-07,1.994397e-07,1.994398e-07,1.994399e-07,1.994400e-07,1.994402e-07,1.994403e-07,1.994404e-07,1.994405e-07,1.994407e-07,1.994408e-07,1.994409e-07,1.994410e-07,1.994411e-07,1.994413e-07,1.994414e-07,1.994415e-07,1.994416e-07,1.994418e-07,1.994419e-07,1.994420e-07,1.994421e-07,1.994422e-07,1.994424e-07,1.994425e-07,1.994426e-07,1.994427e-07,1.994429e-07,1.994430e-07,1.994431e-07,1.994432e-07,1.994434e-07,1.994435e-07,1.994436e-07,1.994437e-07,1.994438e-07,1.994440e-07,1.994441e-07,1.994442e-07,1.994443e-07,1.994445e-07,1.994446e-07,1.994447e-07,1.994448e-07,1.994449e-07,1.994451e-07,1.994452e-07,1.994453e-07,1.994454e-07,1.994456e-07,1.994457e-07,1.994458e-07,1.994459e-07,1.994460e-07,1.994462e-07,1.994463e-07,1.994464e-07,1.994465e-07,1.994467e-07,1.994468e-07,1.994469e-07,1.994470e-07,1.994471e-07,1.994473e-07,1.994474e-07,1.994475e-07,1.994476e-07,1.994478e-07,1.994479e-07,1.994480e-07,1.994481e-07,1.994482e-07,1.994484e-07,1.994485e-07,1.994486e-07,1.994487e-07,1.994489e-07,1.994490e-07,1.994491e-07,1.994492e-07,1.994494e-07,1.994495e-07,1.994496e-07,1.994497e-07,1.994498e-07,1.994500e-07,1.994501e-07,1.994502e-07,1.994503e-07,1.994505e-07,1.994506e-07,1.994507e-07,1.994508e-07,1.994509e-07,1.994511e-07,1.994512e-07,1.994513e-07,1.994514e-07,1.994516e-07,1.994517e-07,1.994518e-07,1.994519e-07,1.994520e-07,1.994522e-07,1.994523e-07,1.994524e-07,1.994525e-07,1.994527e-07,1.994528e-07,1.994529e-07,1.994530e-07,1.994531e-07,1.994533e-07,1.994534e-07,1.994535e-07,1.994536e-07,1.994538e-07,1.994539e-07,1.994540e-07,1.994541e-07,1.994542e-07,1.994544e-07,1.994545e-07,1.994546e-07,1.994547e-07,1.994549e-07,1.994550e-07,1.994551e-07,1.994552e-07,1.994554e-07,1.994555e-07,1.994556e-07,1.994557e-07,1.994558e-07,1.994560e-07,1.994561e-07,1.994562e-07,1.994563e-07,1.994565e-07,1.994566e-07,1.994567e-07,1.994568e-07,1.994569e-07,1.994571e-07,1.994572e-07,1.994573e-07,1.994574e-07,1.994576e-07,1.994577e-07,1.994578e-07,1.994579e-07,1.994580e-07,1.994582e-07,1.994583e-07,1.994584e-07,1.994585e-07,1.994587e-07,1.994588e-07,1.994589e-07,1.994590e-07,1.994591e-07,1.994593e-07,1.994594e-07,1.994595e-07,1.994596e-07,1.994598e-07,1.994599e-07,1.994600e-07,1.994601e-07,1.994602e-07,1.994604e-07,1.994605e-07,1.994606e-07,1.994607e-07,1.994609e-07,1.994610e-07,1.994611e-07,1.994612e-07,1.994613e-07,1.994615e-07,1.994616e-07,1.994617e-07,1.994618e-07,1.994620e-07,1.994621e-07,1.994622e-07,1.994623e-07,1.994624e-07,1.994626e-07,1.994627e-07,1.994628e-07,1.994629e-07,1.994631e-07,1.994632e-07,1.994633e-07,1.994634e-07,1.994635e-07,1.994637e-07,1.994638e-07,1.994639e-07,1.994640e-07,1.994642e-07,1.994643e-07,1.994644e-07,1.994645e-07,1.994646e-07,1.994648e-07,1.994649e-07,1.994650e-07,1.994651e-07,1.994653e-07,1.994654e-07,1.994655e-07,1.994656e-07,1.994657e-07,1.994659e-07,1.994660e-07,1.994661e-07,1.994662e-07,1.994664e-07,1.994665e-07,1.994666e-07,1.994667e-07,1.994669e-07,1.994670e-07,1.994671e-07,1.994672e-07,1.994673e-07,1.994675e-07,1.994676e-07,1.994677e-07,1.994678e-07,1.994680e-07,1.994681e-07,1.994682e-07,1.994683e-07,1.994684e-07,1.994686e-07,1.994687e-07,1.994688e-07,1.994689e-07,1.994691e-07,1.994692e-07,1.994693e-07,1.994694e-07,1.994695e-07,1.994697e-07,1.994698e-07,1.994699e-07,1.994700e-07,1.994702e-07,1.994703e-07,1.994704e-07,1.994705e-07,1.994706e-07,1.994708e-07,1.994709e-07,1.994710e-07,1.994711e-07,1.994713e-07,1.994714e-07,1.994715e-07,1.994716e-07,1.994717e-07,1.994719e-07,1.994720e-07,1.994721e-07,1.994722e-07,1.994724e-07,1.994725e-07,1.994726e-07,1.994727e-07,1.994728e-07,1.994730e-07,1.994731e-07,1.994732e-07,1.994733e-07,1.994735e-07,1.994736e-07,1.994737e-07,1.994738e-07,1.994739e-07,1.994741e-07,1.994742e-07,1.994743e-07,1.994744e-07,1.994746e-07,1.994747e-07,1.994748e-07,1.994749e-07,1.994750e-07,1.994752e-07,1.994753e-07,1.994754e-07,1.994755e-07,1.994757e-07,1.994758e-07,1.994759e-07,1.994760e-07,1.994761e-07,1.994763e-07,1.994764e-07,1.994765e-07,1.994766e-07,1.994768e-07,1.994769e-07,1.994770e-07,1.994771e-07,1.994772e-07,1.994774e-07,1.994775e-07,1.994776e-07,1.994777e-07,1.994778e-07,1.994780e-07,1.994781e-07,1.994782e-07,1.994783e-07,1.994785e-07,1.994786e-07,1.994787e-07,1.994788e-07,1.994789e-07,1.994791e-07,1.994792e-07,1.994793e-07,1.994794e-07,1.994796e-07,1.994797e-07,1.994798e-07,1.994799e-07,1.994800e-07,1.994802e-07,1.994803e-07,1.994804e-07,1.994805e-07,1.994807e-07,1.994808e-07,1.994809e-07,1.994810e-07,1.994811e-07,1.994813e-07,1.994814e-07,1.994815e-07,1.994816e-07,1.994818e-07,1.994819e-07,1.994820e-07,1.994821e-07,1.994822e-07,1.994824e-07,1.994825e-07,1.994826e-07,1.994827e-07,1.994829e-07,1.994830e-07,1.994831e-07,1.994832e-07,1.994833e-07,1.994835e-07,1.994836e-07,1.994837e-07,1.994838e-07,1.994840e-07,1.994841e-07,1.994842e-07,1.994843e-07,1.994844e-07,1.994846e-07,1.994847e-07,1.994848e-07,1.994849e-07,1.994851e-07,1.994852e-07,1.994853e-07,1.994854e-07,1.994855e-07,1.994857e-07,1.994858e-07,1.994859e-07,1.994860e-07,1.994862e-07,1.994863e-07,1.994864e-07,1.994865e-07,1.994866e-07,1.994868e-07,1.994869e-07,1.994870e-07,1.994871e-07,1.994873e-07,1.994874e-07,1.994875e-07,1.994876e-07,1.994877e-07,1.994879e-07,1.994880e-07,1.994881e-07,1.994882e-07,1.994884e-07,1.994885e-07,1.994886e-07,1.994887e-07,1.994888e-07,1.994890e-07,1.994891e-07,1.994892e-07,1.994893e-07,1.994894e-07,1.994896e-07,1.994897e-07,1.994898e-07,1.994899e-07,1.994901e-07,1.994902e-07,1.994903e-07,1.994904e-07,1.994905e-07,1.994907e-07,1.994908e-07,1.994909e-07,1.994910e-07,1.994912e-07,1.994913e-07,1.994914e-07,1.994915e-07,1.994916e-07,1.994918e-07,1.994919e-07,1.994920e-07,1.994921e-07,1.994923e-07,1.994924e-07,1.994925e-07,1.994926e-07,1.994927e-07,1.994929e-07,1.994930e-07,1.994931e-07,1.994932e-07,1.994934e-07,1.994935e-07,1.994936e-07,1.994937e-07,1.994938e-07,1.994940e-07,1.994941e-07,1.994942e-07,1.994943e-07,1.994945e-07,1.994946e-07,1.994947e-07,1.994948e-07,1.994949e-07,1.994951e-07,1.994952e-07,1.994953e-07,1.994954e-07,1.994955e-07,1.994957e-07,1.994958e-07,1.994959e-07,1.994960e-07,1.994962e-07,1.994963e-07,1.994964e-07,1.994965e-07,1.994966e-07,1.994968e-07,1.994969e-07,1.994970e-07,1.994971e-07,1.994973e-07,1.994974e-07,1.994975e-07,1.994976e-07,1.994977e-07,1.994979e-07,1.994980e-07,1.994981e-07,1.994982e-07,1.994984e-07,1.994985e-07,1.994986e-07,1.994987e-07,1.994988e-07,1.994990e-07,1.994991e-07,1.994992e-07,1.994993e-07,1.994995e-07,1.994996e-07,1.994997e-07,1.994998e-07,1.994999e-07,1.995001e-07,1.995002e-07,1.995003e-07,1.995004e-07,1.995005e-07,1.995007e-07,1.995008e-07,1.995009e-07,1.995010e-07,1.995012e-07,1.995013e-07,1.995014e-07,1.995015e-07,1.995016e-07,1.995018e-07,1.995019e-07,1.995020e-07,1.995021e-07,1.995023e-07,1.995024e-07,1.995025e-07,1.995026e-07,1.995027e-07,1.995029e-07,1.995030e-07,1.995031e-07,1.995032e-07,1.995034e-07,1.995035e-07,1.995036e-07,1.995037e-07,1.995038e-07,1.995040e-07,1.995041e-07,1.995042e-07,1.995043e-07,1.995044e-07,1.995046e-07,1.995047e-07,1.995048e-07,1.995049e-07,1.995051e-07,1.995052e-07,1.995053e-07,1.995054e-07,1.995055e-07,1.995057e-07,1.995058e-07,1.995059e-07,1.995060e-07,1.995062e-07,1.995063e-07,1.995064e-07,1.995065e-07,1.995066e-07,1.995068e-07,1.995069e-07,1.995070e-07,1.995071e-07,1.995073e-07,1.995074e-07,1.995075e-07,1.995076e-07,1.995077e-07,1.995079e-07,1.995080e-07,1.995081e-07,1.995082e-07,1.995083e-07,1.995085e-07,1.995086e-07,1.995087e-07,1.995088e-07,1.995090e-07,1.995091e-07,1.995092e-07,1.995093e-07,1.995094e-07,1.995096e-07,1.995097e-07,1.995098e-07,1.995099e-07,1.995101e-07,1.995102e-07,1.995103e-07,1.995104e-07,1.995105e-07,1.995107e-07,1.995108e-07,1.995109e-07,1.995110e-07,1.995112e-07,1.995113e-07,1.995114e-07,1.995115e-07,1.995116e-07,1.995118e-07,1.995119e-07,1.995120e-07,1.995121e-07,1.995122e-07,1.995124e-07,1.995125e-07,1.995126e-07,1.995127e-07,1.995129e-07,1.995130e-07,1.995131e-07,1.995132e-07,1.995133e-07,1.995135e-07,1.995136e-07,1.995137e-07,1.995138e-07,1.995140e-07,1.995141e-07,1.995142e-07,1.995143e-07,1.995144e-07,1.995146e-07,1.995147e-07,1.995148e-07,1.995149e-07,1.995150e-07,1.995152e-07,1.995153e-07,1.995154e-07,1.995155e-07,1.995157e-07,1.995158e-07,1.995159e-07,1.995160e-07,1.995161e-07,1.995163e-07,1.995164e-07,1.995165e-07,1.995166e-07,1.995168e-07,1.995169e-07,1.995170e-07,1.995171e-07,1.995172e-07,1.995174e-07,1.995175e-07,1.995176e-07,1.995177e-07,1.995178e-07,1.995180e-07,1.995181e-07,1.995182e-07,1.995183e-07,1.995185e-07,1.995186e-07,1.995187e-07,1.995188e-07,1.995189e-07,1.995191e-07,1.995192e-07,1.995193e-07,1.995194e-07,1.995196e-07,1.995197e-07,1.995198e-07,1.995199e-07,1.995200e-07,1.995202e-07,1.995203e-07,1.995204e-07,1.995205e-07,1.995206e-07,1.995208e-07,1.995209e-07,1.995210e-07,1.995211e-07,1.995213e-07,1.995214e-07,1.995215e-07,1.995216e-07,1.995217e-07,1.995219e-07,1.995220e-07,1.995221e-07,1.995222e-07,1.995224e-07,1.995225e-07,1.995226e-07,1.995227e-07,1.995228e-07,1.995230e-07,1.995231e-07,1.995232e-07,1.995233e-07,1.995234e-07,1.995236e-07,1.995237e-07,1.995238e-07,1.995239e-07,1.995241e-07,1.995242e-07,1.995243e-07,1.995244e-07,1.995245e-07,1.995247e-07,1.995248e-07,1.995249e-07,1.995250e-07,1.995252e-07,1.995253e-07,1.995254e-07,1.995255e-07,1.995256e-07,1.995258e-07,1.995259e-07,1.995260e-07,1.995261e-07,1.995262e-07,1.995264e-07,1.995265e-07,1.995266e-07,1.995267e-07,1.995269e-07,1.995270e-07,1.995271e-07,1.995272e-07,1.995273e-07,1.995275e-07,1.995276e-07,1.995277e-07,1.995278e-07,1.995279e-07,1.995281e-07,1.995282e-07,1.995283e-07,1.995284e-07,1.995286e-07,1.995287e-07,1.995288e-07,1.995289e-07,1.995290e-07,1.995292e-07,1.995293e-07,1.995294e-07,1.995295e-07,1.995297e-07,1.995298e-07,1.995299e-07,1.995300e-07,1.995301e-07,1.995303e-07,1.995304e-07,1.995305e-07,1.995306e-07,1.995307e-07,1.995309e-07,1.995310e-07,1.995311e-07,1.995312e-07,1.995314e-07,1.995315e-07,1.995316e-07,1.995317e-07,1.995318e-07,1.995320e-07,1.995321e-07,1.995322e-07,1.995323e-07,1.995324e-07,1.995326e-07,1.995327e-07,1.995328e-07,1.995329e-07,1.995331e-07,1.995332e-07,1.995333e-07,1.995334e-07,1.995335e-07,1.995337e-07,1.995338e-07,1.995339e-07,1.995340e-07,1.995342e-07,1.995343e-07,1.995344e-07,1.995345e-07,1.995346e-07,1.995348e-07,1.995349e-07,1.995350e-07,1.995351e-07,1.995352e-07,1.995354e-07,1.995355e-07,1.995356e-07,1.995357e-07,1.995359e-07,1.995360e-07,1.995361e-07,1.995362e-07,1.995363e-07,1.995365e-07,1.995366e-07,1.995367e-07,1.995368e-07,1.995369e-07,1.995371e-07,1.995372e-07,1.995373e-07,1.995374e-07,1.995376e-07,1.995377e-07,1.995378e-07,1.995379e-07,1.995380e-07,1.995382e-07,1.995383e-07,1.995384e-07,1.995385e-07,1.995386e-07,1.995388e-07,1.995389e-07,1.995390e-07,1.995391e-07,1.995393e-07,1.995394e-07,1.995395e-07,1.995396e-07,1.995397e-07,1.995399e-07,1.995400e-07,1.995401e-07,1.995402e-07,1.995403e-07,1.995405e-07,1.995406e-07,1.995407e-07,1.995408e-07,1.995410e-07,1.995411e-07,1.995412e-07,1.995413e-07,1.995414e-07,1.995416e-07,1.995417e-07,1.995418e-07,1.995419e-07,1.995421e-07,1.995422e-07,1.995423e-07,1.995424e-07,1.995425e-07,1.995427e-07,1.995428e-07,1.995429e-07,1.995430e-07,1.995431e-07,1.995433e-07,1.995434e-07,1.995435e-07,1.995436e-07,1.995438e-07,1.995439e-07,1.995440e-07,1.995441e-07,1.995442e-07,1.995444e-07,1.995445e-07,1.995446e-07,1.995447e-07,1.995448e-07,1.995450e-07,1.995451e-07,1.995452e-07,1.995453e-07,1.995455e-07,1.995456e-07,1.995457e-07,1.995458e-07,1.995459e-07,1.995461e-07,1.995462e-07,1.995463e-07,1.995464e-07,1.995465e-07,1.995467e-07,1.995468e-07,1.995469e-07,1.995470e-07,1.995472e-07,1.995473e-07,1.995474e-07,1.995475e-07,1.995476e-07,1.995478e-07,1.995479e-07,1.995480e-07,1.995481e-07,1.995482e-07,1.995484e-07,1.995485e-07,1.995486e-07,1.995487e-07,1.995489e-07,1.995490e-07,1.995491e-07,1.995492e-07,1.995493e-07,1.995495e-07,1.995496e-07,1.995497e-07,1.995498e-07,1.995499e-07,1.995501e-07,1.995502e-07,1.995503e-07,1.995504e-07,1.995506e-07,1.995507e-07,1.995508e-07,1.995509e-07,1.995510e-07,1.995512e-07,1.995513e-07,1.995514e-07,1.995515e-07,1.995516e-07,1.995518e-07,1.995519e-07,1.995520e-07,1.995521e-07,1.995523e-07,1.995524e-07,1.995525e-07,1.995526e-07,1.995527e-07,1.995529e-07,1.995530e-07,1.995531e-07,1.995532e-07,1.995533e-07,1.995535e-07,1.995536e-07,1.995537e-07,1.995538e-07,1.995540e-07,1.995541e-07,1.995542e-07,1.995543e-07,1.995544e-07,1.995546e-07,1.995547e-07,1.995548e-07,1.995549e-07,1.995550e-07,1.995552e-07,1.995553e-07,1.995554e-07,1.995555e-07,1.995556e-07,1.995558e-07,1.995559e-07,1.995560e-07,1.995561e-07,1.995563e-07,1.995564e-07,1.995565e-07,1.995566e-07,1.995567e-07,1.995569e-07,1.995570e-07,1.995571e-07,1.995572e-07,1.995573e-07,1.995575e-07,1.995576e-07,1.995577e-07,1.995578e-07,1.995580e-07,1.995581e-07,1.995582e-07,1.995583e-07,1.995584e-07,1.995586e-07,1.995587e-07,1.995588e-07,1.995589e-07,1.995590e-07,1.995592e-07,1.995593e-07,1.995594e-07,1.995595e-07,1.995597e-07,1.995598e-07,1.995599e-07,1.995600e-07,1.995601e-07,1.995603e-07,1.995604e-07,1.995605e-07,1.995606e-07,1.995607e-07,1.995609e-07,1.995610e-07,1.995611e-07,1.995612e-07,1.995614e-07,1.995615e-07,1.995616e-07,1.995617e-07,1.995618e-07,1.995620e-07,1.995621e-07,1.995622e-07,1.995623e-07,1.995624e-07,1.995626e-07,1.995627e-07,1.995628e-07,1.995629e-07,1.995630e-07,1.995632e-07,1.995633e-07,1.995634e-07,1.995635e-07,1.995637e-07,1.995638e-07,1.995639e-07,1.995640e-07,1.995641e-07,1.995643e-07,1.995644e-07,1.995645e-07,1.995646e-07,1.995647e-07,1.995649e-07,1.995650e-07,1.995651e-07,1.995652e-07,1.995654e-07,1.995655e-07,1.995656e-07,1.995657e-07,1.995658e-07,1.995660e-07,1.995661e-07,1.995662e-07,1.995663e-07,1.995664e-07,1.995666e-07,1.995667e-07,1.995668e-07,1.995669e-07,1.995671e-07,1.995672e-07,1.995673e-07,1.995674e-07,1.995675e-07,1.995677e-07,1.995678e-07,1.995679e-07,1.995680e-07,1.995681e-07,1.995683e-07,1.995684e-07,1.995685e-07,1.995686e-07,1.995687e-07,1.995689e-07,1.995690e-07,1.995691e-07,1.995692e-07,1.995694e-07,1.995695e-07,1.995696e-07,1.995697e-07,1.995698e-07,1.995700e-07,1.995701e-07,1.995702e-07,1.995703e-07,1.995704e-07,1.995706e-07,1.995707e-07,1.995708e-07,1.995709e-07,1.995711e-07,1.995712e-07,1.995713e-07,1.995714e-07,1.995715e-07,1.995717e-07,1.995718e-07,1.995719e-07,1.995720e-07,1.995721e-07,1.995723e-07,1.995724e-07,1.995725e-07,1.995726e-07,1.995727e-07,1.995729e-07,1.995730e-07,1.995731e-07,1.995732e-07,1.995734e-07,1.995735e-07,1.995736e-07,1.995737e-07,1.995738e-07,1.995740e-07,1.995741e-07,1.995742e-07,1.995743e-07,1.995744e-07,1.995746e-07,1.995747e-07,1.995748e-07,1.995749e-07,1.995750e-07,1.995752e-07,1.995753e-07,1.995754e-07,1.995755e-07,1.995757e-07,1.995758e-07,1.995759e-07,1.995760e-07,1.995761e-07,1.995763e-07,1.995764e-07,1.995765e-07,1.995766e-07,1.995767e-07,1.995769e-07,1.995770e-07,1.995771e-07,1.995772e-07,1.995774e-07,1.995775e-07,1.995776e-07,1.995777e-07,1.995778e-07,1.995780e-07,1.995781e-07,1.995782e-07,1.995783e-07,1.995784e-07,1.995786e-07,1.995787e-07,1.995788e-07,1.995789e-07,1.995790e-07,1.995792e-07,1.995793e-07,1.995794e-07,1.995795e-07,1.995797e-07,1.995798e-07,1.995799e-07,1.995800e-07,1.995801e-07,1.995803e-07,1.995804e-07,1.995805e-07,1.995806e-07,1.995807e-07,1.995809e-07,1.995810e-07,1.995811e-07,1.995812e-07,1.995813e-07,1.995815e-07,1.995816e-07,1.995817e-07,1.995818e-07,1.995820e-07,1.995821e-07,1.995822e-07,1.995823e-07,1.995824e-07,1.995826e-07,1.995827e-07,1.995828e-07,1.995829e-07,1.995830e-07,1.995832e-07,1.995833e-07,1.995834e-07,1.995835e-07,1.995836e-07,1.995838e-07,1.995839e-07,1.995840e-07,1.995841e-07,1.995843e-07,1.995844e-07,1.995845e-07,1.995846e-07,1.995847e-07,1.995849e-07,1.995850e-07,1.995851e-07,1.995852e-07,1.995853e-07,1.995855e-07,1.995856e-07,1.995857e-07,1.995858e-07,1.995859e-07,1.995861e-07,1.995862e-07,1.995863e-07,1.995864e-07,1.995866e-07,1.995867e-07,1.995868e-07,1.995869e-07,1.995870e-07,1.995872e-07,1.995873e-07,1.995874e-07,1.995875e-07,1.995876e-07,1.995878e-07,1.995879e-07,1.995880e-07,1.995881e-07,1.995882e-07,1.995884e-07,1.995885e-07,1.995886e-07,1.995887e-07,1.995889e-07,1.995890e-07,1.995891e-07,1.995892e-07,1.995893e-07,1.995895e-07,1.995896e-07,1.995897e-07,1.995898e-07,1.995899e-07,1.995901e-07,1.995902e-07,1.995903e-07,1.995904e-07,1.995905e-07,1.995907e-07,1.995908e-07,1.995909e-07,1.995910e-07,1.995912e-07,1.995913e-07,1.995914e-07,1.995915e-07,1.995916e-07,1.995918e-07,1.995919e-07,1.995920e-07,1.995921e-07,1.995922e-07,1.995924e-07,1.995925e-07,1.995926e-07,1.995927e-07,1.995928e-07,1.995930e-07,1.995931e-07,1.995932e-07,1.995933e-07,1.995935e-07,1.995936e-07,1.995937e-07,1.995938e-07,1.995939e-07,1.995941e-07,1.995942e-07,1.995943e-07,1.995944e-07,1.995945e-07,1.995947e-07,1.995948e-07,1.995949e-07,1.995950e-07,1.995951e-07,1.995953e-07,1.995954e-07,1.995955e-07,1.995956e-07,1.995957e-07,1.995959e-07,1.995960e-07,1.995961e-07,1.995962e-07,1.995964e-07,1.995965e-07,1.995966e-07,1.995967e-07,1.995968e-07,1.995970e-07,1.995971e-07,1.995972e-07,1.995973e-07,1.995974e-07,1.995976e-07,1.995977e-07,1.995978e-07,1.995979e-07,1.995980e-07,1.995982e-07,1.995983e-07,1.995984e-07,1.995985e-07,1.995987e-07,1.995988e-07,1.995989e-07,1.995990e-07,1.995991e-07,1.995993e-07,1.995994e-07,1.995995e-07,1.995996e-07,1.995997e-07,1.995999e-07,1.996000e-07,1.996001e-07,1.996002e-07,1.996003e-07,1.996005e-07,1.996006e-07,1.996007e-07,1.996008e-07,1.996009e-07,1.996011e-07,1.996012e-07,1.996013e-07,1.996014e-07,1.996016e-07,1.996017e-07,1.996018e-07,1.996019e-07,1.996020e-07,1.996022e-07,1.996023e-07,1.996024e-07,1.996025e-07,1.996026e-07,1.996028e-07,1.996029e-07,1.996030e-07,1.996031e-07,1.996032e-07,1.996034e-07,1.996035e-07,1.996036e-07,1.996037e-07,1.996038e-07,1.996040e-07,1.996041e-07,1.996042e-07,1.996043e-07,1.996045e-07,1.996046e-07,1.996047e-07,1.996048e-07,1.996049e-07,1.996051e-07,1.996052e-07,1.996053e-07,1.996054e-07,1.996055e-07,1.996057e-07,1.996058e-07,1.996059e-07,1.996060e-07,1.996061e-07,1.996063e-07,1.996064e-07,1.996065e-07,1.996066e-07,1.996067e-07,1.996069e-07,1.996070e-07,1.996071e-07,1.996072e-07,1.996074e-07,1.996075e-07,1.996076e-07,1.996077e-07,1.996078e-07,1.996080e-07,1.996081e-07,1.996082e-07,1.996083e-07,1.996084e-07,1.996086e-07,1.996087e-07,1.996088e-07,1.996089e-07,1.996090e-07,1.996092e-07,1.996093e-07,1.996094e-07,1.996095e-07,1.996096e-07,1.996098e-07,1.996099e-07,1.996100e-07,1.996101e-07,1.996103e-07,1.996104e-07,1.996105e-07,1.996106e-07,1.996107e-07,1.996109e-07,1.996110e-07,1.996111e-07,1.996112e-07,1.996113e-07,1.996115e-07,1.996116e-07,1.996117e-07,1.996118e-07,1.996119e-07,1.996121e-07,1.996122e-07,1.996123e-07,1.996124e-07,1.996125e-07,1.996127e-07,1.996128e-07,1.996129e-07,1.996130e-07,1.996132e-07,1.996133e-07,1.996134e-07,1.996135e-07,1.996136e-07,1.996138e-07,1.996139e-07,1.996140e-07,1.996141e-07,1.996142e-07,1.996144e-07,1.996145e-07,1.996146e-07,1.996147e-07,1.996148e-07,1.996150e-07,1.996151e-07,1.996152e-07,1.996153e-07,1.996154e-07,1.996156e-07,1.996157e-07,1.996158e-07,1.996159e-07,1.996160e-07,1.996162e-07,1.996163e-07,1.996164e-07,1.996165e-07,1.996167e-07,1.996168e-07,1.996169e-07,1.996170e-07,1.996171e-07,1.996173e-07,1.996174e-07,1.996175e-07,1.996176e-07,1.996177e-07,1.996179e-07,1.996180e-07,1.996181e-07,1.996182e-07,1.996183e-07,1.996185e-07,1.996186e-07,1.996187e-07,1.996188e-07,1.996189e-07,1.996191e-07,1.996192e-07,1.996193e-07,1.996194e-07,1.996195e-07,1.996197e-07,1.996198e-07,1.996199e-07,1.996200e-07,1.996202e-07,1.996203e-07,1.996204e-07,1.996205e-07,1.996206e-07,1.996208e-07,1.996209e-07,1.996210e-07,1.996211e-07,1.996212e-07,1.996214e-07,1.996215e-07,1.996216e-07,1.996217e-07,1.996218e-07,1.996220e-07,1.996221e-07,1.996222e-07,1.996223e-07,1.996224e-07,1.996226e-07,1.996227e-07,1.996228e-07,1.996229e-07,1.996230e-07,1.996232e-07,1.996233e-07,1.996234e-07,1.996235e-07,1.996237e-07,1.996238e-07,1.996239e-07,1.996240e-07,1.996241e-07,1.996243e-07,1.996244e-07,1.996245e-07,1.996246e-07,1.996247e-07,1.996249e-07,1.996250e-07,1.996251e-07,1.996252e-07,1.996253e-07,1.996255e-07,1.996256e-07,1.996257e-07,1.996258e-07,1.996259e-07,1.996261e-07,1.996262e-07,1.996263e-07,1.996264e-07,1.996265e-07,1.996267e-07,1.996268e-07,1.996269e-07,1.996270e-07,1.996271e-07,1.996273e-07,1.996274e-07,1.996275e-07,1.996276e-07,1.996278e-07,1.996279e-07,1.996280e-07,1.996281e-07,1.996282e-07,1.996284e-07,1.996285e-07,1.996286e-07,1.996287e-07,1.996288e-07,1.996290e-07,1.996291e-07,1.996292e-07,1.996293e-07,1.996294e-07,1.996296e-07,1.996297e-07,1.996298e-07,1.996299e-07,1.996300e-07,1.996302e-07,1.996303e-07,1.996304e-07,1.996305e-07,1.996306e-07,1.996308e-07,1.996309e-07,1.996310e-07,1.996311e-07,1.996312e-07,1.996314e-07,1.996315e-07,1.996316e-07,1.996317e-07,1.996319e-07,1.996320e-07,1.996321e-07,1.996322e-07,1.996323e-07,1.996325e-07,1.996326e-07,1.996327e-07,1.996328e-07,1.996329e-07,1.996331e-07,1.996332e-07,1.996333e-07,1.996334e-07,1.996335e-07,1.996337e-07,1.996338e-07,1.996339e-07,1.996340e-07,1.996341e-07,1.996343e-07,1.996344e-07,1.996345e-07,1.996346e-07,1.996347e-07,1.996349e-07,1.996350e-07,1.996351e-07,1.996352e-07,1.996353e-07,1.996355e-07,1.996356e-07,1.996357e-07,1.996358e-07,1.996360e-07,1.996361e-07,1.996362e-07,1.996363e-07,1.996364e-07,1.996366e-07,1.996367e-07,1.996368e-07,1.996369e-07,1.996370e-07,1.996372e-07,1.996373e-07,1.996374e-07,1.996375e-07,1.996376e-07,1.996378e-07,1.996379e-07,1.996380e-07,1.996381e-07,1.996382e-07,1.996384e-07,1.996385e-07,1.996386e-07,1.996387e-07,1.996388e-07,1.996390e-07,1.996391e-07,1.996392e-07,1.996393e-07,1.996394e-07,1.996396e-07,1.996397e-07,1.996398e-07,1.996399e-07,1.996400e-07,1.996402e-07,1.996403e-07,1.996404e-07,1.996405e-07,1.996407e-07,1.996408e-07,1.996409e-07,1.996410e-07,1.996411e-07,1.996413e-07,1.996414e-07,1.996415e-07,1.996416e-07,1.996417e-07,1.996419e-07,1.996420e-07,1.996421e-07,1.996422e-07,1.996423e-07,1.996425e-07,1.996426e-07,1.996427e-07,1.996428e-07,1.996429e-07,1.996431e-07,1.996432e-07,1.996433e-07,1.996434e-07,1.996435e-07,1.996437e-07,1.996438e-07,1.996439e-07,1.996440e-07,1.996441e-07,1.996443e-07,1.996444e-07,1.996445e-07,1.996446e-07,1.996447e-07,1.996449e-07,1.996450e-07,1.996451e-07,1.996452e-07,1.996453e-07,1.996455e-07,1.996456e-07,1.996457e-07,1.996458e-07,1.996459e-07,1.996461e-07,1.996462e-07,1.996463e-07,1.996464e-07,1.996466e-07,1.996467e-07,1.996468e-07,1.996469e-07,1.996470e-07,1.996472e-07,1.996473e-07,1.996474e-07,1.996475e-07,1.996476e-07,1.996478e-07,1.996479e-07,1.996480e-07,1.996481e-07,1.996482e-07,1.996484e-07,1.996485e-07,1.996486e-07,1.996487e-07,1.996488e-07,1.996490e-07,1.996491e-07,1.996492e-07,1.996493e-07,1.996494e-07,1.996496e-07,1.996497e-07,1.996498e-07,1.996499e-07,1.996500e-07,1.996502e-07,1.996503e-07,1.996504e-07,1.996505e-07,1.996506e-07,1.996508e-07,1.996509e-07,1.996510e-07,1.996511e-07,1.996512e-07,1.996514e-07,1.996515e-07,1.996516e-07,1.996517e-07,1.996518e-07,1.996520e-07,1.996521e-07,1.996522e-07,1.996523e-07,1.996525e-07,1.996526e-07,1.996527e-07,1.996528e-07,1.996529e-07,1.996531e-07,1.996532e-07,1.996533e-07,1.996534e-07,1.996535e-07,1.996537e-07,1.996538e-07,1.996539e-07,1.996540e-07,1.996541e-07,1.996543e-07,1.996544e-07,1.996545e-07,1.996546e-07,1.996547e-07,1.996549e-07,1.996550e-07,1.996551e-07,1.996552e-07,1.996553e-07,1.996555e-07,1.996556e-07,1.996557e-07,1.996558e-07,1.996559e-07,1.996561e-07,1.996562e-07,1.996563e-07,1.996564e-07,1.996565e-07,1.996567e-07,1.996568e-07,1.996569e-07,1.996570e-07,1.996571e-07,1.996573e-07,1.996574e-07,1.996575e-07,1.996576e-07,1.996577e-07,1.996579e-07,1.996580e-07,1.996581e-07,1.996582e-07,1.996583e-07,1.996585e-07,1.996586e-07,1.996587e-07,1.996588e-07,1.996589e-07,1.996591e-07,1.996592e-07,1.996593e-07,1.996594e-07,1.996595e-07,1.996597e-07,1.996598e-07,1.996599e-07,1.996600e-07,1.996602e-07,1.996603e-07,1.996604e-07,1.996605e-07,1.996606e-07,1.996608e-07,1.996609e-07,1.996610e-07,1.996611e-07,1.996612e-07,1.996614e-07,1.996615e-07,1.996616e-07,1.996617e-07,1.996618e-07,1.996620e-07,1.996621e-07,1.996622e-07,1.996623e-07,1.996624e-07,1.996626e-07,1.996627e-07,1.996628e-07,1.996629e-07,1.996630e-07,1.996632e-07,1.996633e-07,1.996634e-07,1.996635e-07,1.996636e-07,1.996638e-07,1.996639e-07,1.996640e-07,1.996641e-07,1.996642e-07,1.996644e-07,1.996645e-07,1.996646e-07,1.996647e-07,1.996648e-07,1.996650e-07,1.996651e-07,1.996652e-07,1.996653e-07,1.996654e-07,1.996656e-07,1.996657e-07,1.996658e-07,1.996659e-07,1.996660e-07,1.996662e-07,1.996663e-07,1.996664e-07,1.996665e-07,1.996666e-07,1.996668e-07,1.996669e-07,1.996670e-07,1.996671e-07,1.996672e-07,1.996674e-07,1.996675e-07,1.996676e-07,1.996677e-07,1.996678e-07,1.996680e-07,1.996681e-07,1.996682e-07,1.996683e-07,1.996684e-07,1.996686e-07,1.996687e-07,1.996688e-07,1.996689e-07,1.996690e-07,1.996692e-07,1.996693e-07,1.996694e-07,1.996695e-07,1.996696e-07,1.996698e-07,1.996699e-07,1.996700e-07,1.996701e-07,1.996702e-07,1.996704e-07,1.996705e-07,1.996706e-07,1.996707e-07,1.996709e-07,1.996710e-07,1.996711e-07,1.996712e-07,1.996713e-07,1.996715e-07,1.996716e-07,1.996717e-07,1.996718e-07,1.996719e-07,1.996721e-07,1.996722e-07,1.996723e-07,1.996724e-07,1.996725e-07,1.996727e-07,1.996728e-07,1.996729e-07,1.996730e-07,1.996731e-07,1.996733e-07,1.996734e-07,1.996735e-07,1.996736e-07,1.996737e-07,1.996739e-07,1.996740e-07,1.996741e-07,1.996742e-07,1.996743e-07,1.996745e-07,1.996746e-07,1.996747e-07,1.996748e-07,1.996749e-07,1.996751e-07,1.996752e-07,1.996753e-07,1.996754e-07,1.996755e-07,1.996757e-07,1.996758e-07,1.996759e-07,1.996760e-07,1.996761e-07,1.996763e-07,1.996764e-07,1.996765e-07,1.996766e-07,1.996767e-07,1.996769e-07,1.996770e-07,1.996771e-07,1.996772e-07,1.996773e-07,1.996775e-07,1.996776e-07,1.996777e-07,1.996778e-07,1.996779e-07,1.996781e-07,1.996782e-07,1.996783e-07,1.996784e-07,1.996785e-07,1.996787e-07,1.996788e-07,1.996789e-07,1.996790e-07,1.996791e-07,1.996793e-07,1.996794e-07,1.996795e-07,1.996796e-07,1.996797e-07,1.996799e-07,1.996800e-07,1.996801e-07,1.996802e-07,1.996803e-07,1.996805e-07,1.996806e-07,1.996807e-07,1.996808e-07,1.996809e-07,1.996811e-07,1.996812e-07,1.996813e-07,1.996814e-07,1.996815e-07,1.996817e-07,1.996818e-07,1.996819e-07,1.996820e-07,1.996821e-07,1.996823e-07,1.996824e-07,1.996825e-07,1.996826e-07,1.996827e-07,1.996829e-07,1.996830e-07,1.996831e-07,1.996832e-07,1.996833e-07,1.996835e-07,1.996836e-07,1.996837e-07,1.996838e-07,1.996839e-07,1.996841e-07,1.996842e-07,1.996843e-07,1.996844e-07,1.996845e-07,1.996847e-07,1.996848e-07,1.996849e-07,1.996850e-07,1.996851e-07,1.996853e-07,1.996854e-07,1.996855e-07,1.996856e-07,1.996857e-07,1.996859e-07,1.996860e-07,1.996861e-07,1.996862e-07,1.996863e-07,1.996865e-07,1.996866e-07,1.996867e-07,1.996868e-07,1.996869e-07,1.996871e-07,1.996872e-07,1.996873e-07,1.996874e-07,1.996875e-07,1.996877e-07,1.996878e-07,1.996879e-07,1.996880e-07,1.996881e-07,1.996883e-07,1.996884e-07,1.996885e-07,1.996886e-07,1.996887e-07,1.996889e-07,1.996890e-07,1.996891e-07,1.996892e-07,1.996893e-07,1.996895e-07,1.996896e-07,1.996897e-07,1.996898e-07,1.996899e-07,1.996901e-07,1.996902e-07,1.996903e-07,1.996904e-07,1.996905e-07,1.996907e-07,1.996908e-07,1.996909e-07,1.996910e-07,1.996911e-07,1.996913e-07,1.996914e-07,1.996915e-07,1.996916e-07,1.996917e-07,1.996919e-07,1.996920e-07,1.996921e-07,1.996922e-07,1.996923e-07,1.996925e-07,1.996926e-07,1.996927e-07,1.996928e-07,1.996929e-07,1.996931e-07,1.996932e-07,1.996933e-07,1.996934e-07,1.996935e-07,1.996937e-07,1.996938e-07,1.996939e-07,1.996940e-07,1.996941e-07,1.996943e-07,1.996944e-07,1.996945e-07,1.996946e-07,1.996947e-07,1.996949e-07,1.996950e-07,1.996951e-07,1.996952e-07,1.996953e-07,1.996955e-07,1.996956e-07,1.996957e-07,1.996958e-07,1.996959e-07,1.996961e-07,1.996962e-07,1.996963e-07,1.996964e-07,1.996965e-07,1.996967e-07,1.996968e-07,1.996969e-07,1.996970e-07,1.996971e-07,1.996973e-07,1.996974e-07,1.996975e-07,1.996976e-07,1.996977e-07,1.996979e-07,1.996980e-07,1.996981e-07,1.996982e-07,1.996983e-07,1.996985e-07,1.996986e-07,1.996987e-07,1.996988e-07,1.996989e-07,1.996991e-07,1.996992e-07,1.996993e-07,1.996994e-07,1.996995e-07,1.996997e-07,1.996998e-07,1.996999e-07,1.997000e-07,1.997001e-07,1.997003e-07,1.997004e-07,1.997005e-07,1.997006e-07,1.997007e-07,1.997009e-07,1.997010e-07,1.997011e-07,1.997012e-07,1.997013e-07,1.997015e-07,1.997016e-07,1.997017e-07,1.997018e-07,1.997019e-07,1.997021e-07,1.997022e-07,1.997023e-07,1.997024e-07,1.997025e-07,1.997027e-07,1.997028e-07,1.997029e-07,1.997030e-07,1.997031e-07,1.997032e-07,1.997034e-07,1.997035e-07,1.997036e-07,1.997037e-07,1.997038e-07,1.997040e-07,1.997041e-07,1.997042e-07,1.997043e-07,1.997044e-07,1.997046e-07,1.997047e-07,1.997048e-07,1.997049e-07,1.997050e-07,1.997052e-07,1.997053e-07,1.997054e-07,1.997055e-07,1.997056e-07,1.997058e-07,1.997059e-07,1.997060e-07,1.997061e-07,1.997062e-07,1.997064e-07,1.997065e-07,1.997066e-07,1.997067e-07,1.997068e-07,1.997070e-07,1.997071e-07,1.997072e-07,1.997073e-07,1.997074e-07,1.997076e-07,1.997077e-07,1.997078e-07,1.997079e-07,1.997080e-07,1.997082e-07,1.997083e-07,1.997084e-07,1.997085e-07,1.997086e-07,1.997088e-07,1.997089e-07,1.997090e-07,1.997091e-07,1.997092e-07,1.997094e-07,1.997095e-07,1.997096e-07,1.997097e-07,1.997098e-07,1.997100e-07,1.997101e-07,1.997102e-07,1.997103e-07,1.997104e-07,1.997106e-07,1.997107e-07,1.997108e-07,1.997109e-07,1.997110e-07,1.997112e-07,1.997113e-07,1.997114e-07,1.997115e-07,1.997116e-07,1.997118e-07,1.997119e-07,1.997120e-07,1.997121e-07,1.997122e-07,1.997124e-07,1.997125e-07,1.997126e-07,1.997127e-07,1.997128e-07,1.997130e-07,1.997131e-07,1.997132e-07,1.997133e-07,1.997134e-07,1.997136e-07,1.997137e-07,1.997138e-07,1.997139e-07,1.997140e-07,1.997141e-07,1.997143e-07,1.997144e-07,1.997145e-07,1.997146e-07,1.997147e-07,1.997149e-07,1.997150e-07,1.997151e-07,1.997152e-07,1.997153e-07,1.997155e-07,1.997156e-07,1.997157e-07,1.997158e-07,1.997159e-07,1.997161e-07,1.997162e-07,1.997163e-07,1.997164e-07,1.997165e-07,1.997167e-07,1.997168e-07,1.997169e-07,1.997170e-07,1.997171e-07,1.997173e-07,1.997174e-07,1.997175e-07,1.997176e-07,1.997177e-07,1.997179e-07,1.997180e-07,1.997181e-07,1.997182e-07,1.997183e-07,1.997185e-07,1.997186e-07,1.997187e-07,1.997188e-07,1.997189e-07,1.997191e-07,1.997192e-07,1.997193e-07,1.997194e-07,1.997195e-07,1.997197e-07,1.997198e-07,1.997199e-07,1.997200e-07,1.997201e-07,1.997203e-07,1.997204e-07,1.997205e-07,1.997206e-07,1.997207e-07,1.997209e-07,1.997210e-07,1.997211e-07,1.997212e-07,1.997213e-07,1.997214e-07,1.997216e-07,1.997217e-07,1.997218e-07,1.997219e-07,1.997220e-07,1.997222e-07,1.997223e-07,1.997224e-07,1.997225e-07,1.997226e-07,1.997228e-07,1.997229e-07,1.997230e-07,1.997231e-07,1.997232e-07,1.997234e-07,1.997235e-07,1.997236e-07,1.997237e-07,1.997238e-07,1.997240e-07,1.997241e-07,1.997242e-07,1.997243e-07,1.997244e-07,1.997246e-07,1.997247e-07,1.997248e-07,1.997249e-07,1.997250e-07,1.997252e-07,1.997253e-07,1.997254e-07,1.997255e-07,1.997256e-07,1.997258e-07,1.997259e-07,1.997260e-07,1.997261e-07,1.997262e-07,1.997264e-07,1.997265e-07,1.997266e-07,1.997267e-07,1.997268e-07,1.997270e-07,1.997271e-07,1.997272e-07,1.997273e-07,1.997274e-07,1.997276e-07,1.997277e-07,1.997278e-07,1.997279e-07,1.997280e-07,1.997281e-07,1.997283e-07,1.997284e-07,1.997285e-07,1.997286e-07,1.997287e-07,1.997289e-07,1.997290e-07,1.997291e-07,1.997292e-07,1.997293e-07,1.997295e-07,1.997296e-07,1.997297e-07,1.997298e-07,1.997299e-07,1.997301e-07,1.997302e-07,1.997303e-07,1.997304e-07,1.997305e-07,1.997307e-07,1.997308e-07,1.997309e-07,1.997310e-07,1.997311e-07,1.997313e-07,1.997314e-07,1.997315e-07,1.997316e-07,1.997317e-07,1.997319e-07,1.997320e-07,1.997321e-07,1.997322e-07,1.997323e-07,1.997325e-07,1.997326e-07,1.997327e-07,1.997328e-07,1.997329e-07,1.997330e-07,1.997332e-07,1.997333e-07,1.997334e-07,1.997335e-07,1.997336e-07,1.997338e-07,1.997339e-07,1.997340e-07,1.997341e-07,1.997342e-07,1.997344e-07,1.997345e-07,1.997346e-07,1.997347e-07,1.997348e-07,1.997350e-07,1.997351e-07,1.997352e-07,1.997353e-07,1.997354e-07,1.997356e-07,1.997357e-07,1.997358e-07,1.997359e-07,1.997360e-07,1.997362e-07,1.997363e-07,1.997364e-07,1.997365e-07,1.997366e-07,1.997368e-07,1.997369e-07,1.997370e-07,1.997371e-07,1.997372e-07,1.997374e-07,1.997375e-07,1.997376e-07,1.997377e-07,1.997378e-07,1.997379e-07,1.997381e-07,1.997382e-07,1.997383e-07,1.997384e-07,1.997385e-07,1.997387e-07,1.997388e-07,1.997389e-07,1.997390e-07,1.997391e-07,1.997393e-07,1.997394e-07,1.997395e-07,1.997396e-07,1.997397e-07,1.997399e-07,1.997400e-07,1.997401e-07,1.997402e-07,1.997403e-07,1.997405e-07,1.997406e-07,1.997407e-07,1.997408e-07,1.997409e-07,1.997411e-07,1.997412e-07,1.997413e-07,1.997414e-07,1.997415e-07,1.997417e-07,1.997418e-07,1.997419e-07,1.997420e-07,1.997421e-07,1.997422e-07,1.997424e-07,1.997425e-07,1.997426e-07,1.997427e-07,1.997428e-07,1.997430e-07,1.997431e-07,1.997432e-07,1.997433e-07,1.997434e-07,1.997436e-07,1.997437e-07,1.997438e-07,1.997439e-07,1.997440e-07,1.997442e-07,1.997443e-07,1.997444e-07,1.997445e-07,1.997446e-07,1.997448e-07,1.997449e-07,1.997450e-07,1.997451e-07,1.997452e-07,1.997454e-07,1.997455e-07,1.997456e-07,1.997457e-07,1.997458e-07,1.997460e-07,1.997461e-07,1.997462e-07,1.997463e-07,1.997464e-07,1.997465e-07,1.997467e-07,1.997468e-07,1.997469e-07,1.997470e-07,1.997471e-07,1.997473e-07,1.997474e-07,1.997475e-07,1.997476e-07,1.997477e-07,1.997479e-07,1.997480e-07,1.997481e-07,1.997482e-07,1.997483e-07,1.997485e-07,1.997486e-07,1.997487e-07,1.997488e-07,1.997489e-07,1.997491e-07,1.997492e-07,1.997493e-07,1.997494e-07,1.997495e-07,1.997497e-07,1.997498e-07,1.997499e-07,1.997500e-07,1.997501e-07,1.997502e-07,1.997504e-07,1.997505e-07,1.997506e-07,1.997507e-07,1.997508e-07,1.997510e-07,1.997511e-07,1.997512e-07,1.997513e-07,1.997514e-07,1.997516e-07,1.997517e-07,1.997518e-07,1.997519e-07,1.997520e-07,1.997522e-07,1.997523e-07,1.997524e-07,1.997525e-07,1.997526e-07,1.997528e-07,1.997529e-07,1.997530e-07,1.997531e-07,1.997532e-07,1.997534e-07,1.997535e-07,1.997536e-07,1.997537e-07,1.997538e-07,1.997539e-07,1.997541e-07,1.997542e-07,1.997543e-07,1.997544e-07,1.997545e-07,1.997547e-07,1.997548e-07,1.997549e-07,1.997550e-07,1.997551e-07,1.997553e-07,1.997554e-07,1.997555e-07,1.997556e-07,1.997557e-07,1.997559e-07,1.997560e-07,1.997561e-07,1.997562e-07,1.997563e-07,1.997565e-07,1.997566e-07,1.997567e-07,1.997568e-07,1.997569e-07,1.997571e-07,1.997572e-07,1.997573e-07,1.997574e-07,1.997575e-07,1.997576e-07,1.997578e-07,1.997579e-07,1.997580e-07,1.997581e-07,1.997582e-07,1.997584e-07,1.997585e-07,1.997586e-07,1.997587e-07,1.997588e-07,1.997590e-07,1.997591e-07,1.997592e-07,1.997593e-07,1.997594e-07,1.997596e-07,1.997597e-07,1.997598e-07,1.997599e-07,1.997600e-07,1.997602e-07,1.997603e-07,1.997604e-07,1.997605e-07,1.997606e-07,1.997607e-07,1.997609e-07,1.997610e-07,1.997611e-07,1.997612e-07,1.997613e-07,1.997615e-07,1.997616e-07,1.997617e-07,1.997618e-07,1.997619e-07,1.997621e-07,1.997622e-07,1.997623e-07,1.997624e-07,1.997625e-07,1.997627e-07,1.997628e-07,1.997629e-07,1.997630e-07,1.997631e-07,1.997633e-07,1.997634e-07,1.997635e-07,1.997636e-07,1.997637e-07,1.997638e-07,1.997640e-07,1.997641e-07,1.997642e-07,1.997643e-07,1.997644e-07,1.997646e-07,1.997647e-07,1.997648e-07,1.997649e-07,1.997650e-07,1.997652e-07,1.997653e-07,1.997654e-07,1.997655e-07,1.997656e-07,1.997658e-07,1.997659e-07,1.997660e-07,1.997661e-07,1.997662e-07,1.997664e-07,1.997665e-07,1.997666e-07,1.997667e-07,1.997668e-07,1.997669e-07,1.997671e-07,1.997672e-07,1.997673e-07,1.997674e-07,1.997675e-07,1.997677e-07,1.997678e-07,1.997679e-07,1.997680e-07,1.997681e-07,1.997683e-07,1.997684e-07,1.997685e-07,1.997686e-07,1.997687e-07,1.997689e-07,1.997690e-07,1.997691e-07,1.997692e-07,1.997693e-07,1.997694e-07,1.997696e-07,1.997697e-07,1.997698e-07,1.997699e-07,1.997700e-07,1.997702e-07,1.997703e-07,1.997704e-07,1.997705e-07,1.997706e-07,1.997708e-07,1.997709e-07,1.997710e-07,1.997711e-07,1.997712e-07,1.997714e-07,1.997715e-07,1.997716e-07,1.997717e-07,1.997718e-07,1.997720e-07,1.997721e-07,1.997722e-07,1.997723e-07,1.997724e-07,1.997725e-07,1.997727e-07,1.997728e-07,1.997729e-07,1.997730e-07,1.997731e-07,1.997733e-07,1.997734e-07,1.997735e-07,1.997736e-07,1.997737e-07,1.997739e-07,1.997740e-07,1.997741e-07,1.997742e-07,1.997743e-07,1.997745e-07,1.997746e-07,1.997747e-07,1.997748e-07,1.997749e-07,1.997750e-07,1.997752e-07,1.997753e-07,1.997754e-07,1.997755e-07,1.997756e-07,1.997758e-07,1.997759e-07,1.997760e-07,1.997761e-07,1.997762e-07,1.997764e-07,1.997765e-07,1.997766e-07,1.997767e-07,1.997768e-07,1.997770e-07,1.997771e-07,1.997772e-07,1.997773e-07,1.997774e-07,1.997775e-07,1.997777e-07,1.997778e-07,1.997779e-07,1.997780e-07,1.997781e-07,1.997783e-07,1.997784e-07,1.997785e-07,1.997786e-07,1.997787e-07,1.997789e-07,1.997790e-07,1.997791e-07,1.997792e-07,1.997793e-07,1.997795e-07,1.997796e-07,1.997797e-07,1.997798e-07,1.997799e-07,1.997800e-07,1.997802e-07,1.997803e-07,1.997804e-07,1.997805e-07,1.997806e-07,1.997808e-07,1.997809e-07,1.997810e-07,1.997811e-07,1.997812e-07,1.997814e-07,1.997815e-07,1.997816e-07,1.997817e-07,1.997818e-07,1.997820e-07,1.997821e-07,1.997822e-07,1.997823e-07,1.997824e-07,1.997825e-07,1.997827e-07,1.997828e-07,1.997829e-07,1.997830e-07,1.997831e-07,1.997833e-07,1.997834e-07,1.997835e-07,1.997836e-07,1.997837e-07,1.997839e-07,1.997840e-07,1.997841e-07,1.997842e-07,1.997843e-07,1.997845e-07,1.997846e-07,1.997847e-07,1.997848e-07,1.997849e-07,1.997850e-07,1.997852e-07,1.997853e-07,1.997854e-07,1.997855e-07,1.997856e-07,1.997858e-07,1.997859e-07,1.997860e-07,1.997861e-07,1.997862e-07,1.997864e-07,1.997865e-07,1.997866e-07,1.997867e-07,1.997868e-07,1.997870e-07,1.997871e-07,1.997872e-07,1.997873e-07,1.997874e-07,1.997875e-07,1.997877e-07,1.997878e-07,1.997879e-07,1.997880e-07,1.997881e-07,1.997883e-07,1.997884e-07,1.997885e-07,1.997886e-07,1.997887e-07,1.997889e-07,1.997890e-07,1.997891e-07,1.997892e-07,1.997893e-07,1.997895e-07,1.997896e-07,1.997897e-07,1.997898e-07,1.997899e-07,1.997900e-07,1.997902e-07,1.997903e-07,1.997904e-07,1.997905e-07,1.997906e-07,1.997908e-07,1.997909e-07,1.997910e-07,1.997911e-07,1.997912e-07,1.997914e-07,1.997915e-07,1.997916e-07,1.997917e-07,1.997918e-07,1.997919e-07,1.997921e-07,1.997922e-07,1.997923e-07,1.997924e-07,1.997925e-07,1.997927e-07,1.997928e-07,1.997929e-07,1.997930e-07,1.997931e-07,1.997933e-07,1.997934e-07,1.997935e-07,1.997936e-07,1.997937e-07,1.997939e-07,1.997940e-07,1.997941e-07,1.997942e-07,1.997943e-07,1.997944e-07,1.997946e-07,1.997947e-07,1.997948e-07,1.997949e-07,1.997950e-07,1.997952e-07,1.997953e-07,1.997954e-07,1.997955e-07,1.997956e-07,1.997958e-07,1.997959e-07,1.997960e-07,1.997961e-07,1.997962e-07,1.997963e-07,1.997965e-07,1.997966e-07,1.997967e-07,1.997968e-07,1.997969e-07,1.997971e-07,1.997972e-07,1.997973e-07,1.997974e-07,1.997975e-07,1.997977e-07,1.997978e-07,1.997979e-07,1.997980e-07,1.997981e-07,1.997982e-07,1.997984e-07,1.997985e-07,1.997986e-07,1.997987e-07,1.997988e-07,1.997990e-07,1.997991e-07,1.997992e-07,1.997993e-07,1.997994e-07,1.997996e-07,1.997997e-07,1.997998e-07,1.997999e-07,1.998000e-07,1.998002e-07,1.998003e-07,1.998004e-07,1.998005e-07,1.998006e-07,1.998007e-07,1.998009e-07,1.998010e-07,1.998011e-07,1.998012e-07,1.998013e-07,1.998015e-07,1.998016e-07,1.998017e-07,1.998018e-07,1.998019e-07,1.998021e-07,1.998022e-07,1.998023e-07,1.998024e-07,1.998025e-07,1.998026e-07,1.998028e-07,1.998029e-07,1.998030e-07,1.998031e-07,1.998032e-07,1.998034e-07,1.998035e-07,1.998036e-07,1.998037e-07,1.998038e-07,1.998040e-07,1.998041e-07,1.998042e-07,1.998043e-07,1.998044e-07,1.998045e-07,1.998047e-07,1.998048e-07,1.998049e-07,1.998050e-07,1.998051e-07,1.998053e-07,1.998054e-07,1.998055e-07,1.998056e-07,1.998057e-07,1.998059e-07,1.998060e-07,1.998061e-07,1.998062e-07,1.998063e-07,1.998064e-07,1.998066e-07,1.998067e-07,1.998068e-07,1.998069e-07,1.998070e-07,1.998072e-07,1.998073e-07,1.998074e-07,1.998075e-07,1.998076e-07,1.998078e-07,1.998079e-07,1.998080e-07,1.998081e-07,1.998082e-07,1.998083e-07,1.998085e-07,1.998086e-07,1.998087e-07,1.998088e-07,1.998089e-07,1.998091e-07,1.998092e-07,1.998093e-07,1.998094e-07,1.998095e-07,1.998097e-07,1.998098e-07,1.998099e-07,1.998100e-07,1.998101e-07,1.998102e-07,1.998104e-07,1.998105e-07,1.998106e-07,1.998107e-07,1.998108e-07,1.998110e-07,1.998111e-07,1.998112e-07,1.998113e-07,1.998114e-07,1.998116e-07,1.998117e-07,1.998118e-07,1.998119e-07,1.998120e-07,1.998121e-07,1.998123e-07,1.998124e-07,1.998125e-07,1.998126e-07,1.998127e-07,1.998129e-07,1.998130e-07,1.998131e-07,1.998132e-07,1.998133e-07,1.998135e-07,1.998136e-07,1.998137e-07,1.998138e-07,1.998139e-07,1.998140e-07,1.998142e-07,1.998143e-07,1.998144e-07,1.998145e-07,1.998146e-07,1.998148e-07,1.998149e-07,1.998150e-07,1.998151e-07,1.998152e-07,1.998154e-07,1.998155e-07,1.998156e-07,1.998157e-07,1.998158e-07,1.998159e-07,1.998161e-07,1.998162e-07,1.998163e-07,1.998164e-07,1.998165e-07,1.998167e-07,1.998168e-07,1.998169e-07,1.998170e-07,1.998171e-07,1.998173e-07,1.998174e-07,1.998175e-07,1.998176e-07,1.998177e-07,1.998178e-07,1.998180e-07,1.998181e-07,1.998182e-07,1.998183e-07,1.998184e-07,1.998186e-07,1.998187e-07,1.998188e-07,1.998189e-07,1.998190e-07,1.998192e-07,1.998193e-07,1.998194e-07,1.998195e-07,1.998196e-07,1.998197e-07,1.998199e-07,1.998200e-07,1.998201e-07,1.998202e-07,1.998203e-07,1.998205e-07,1.998206e-07,1.998207e-07,1.998208e-07,1.998209e-07,1.998210e-07,1.998212e-07,1.998213e-07,1.998214e-07,1.998215e-07,1.998216e-07,1.998218e-07,1.998219e-07,1.998220e-07,1.998221e-07,1.998222e-07,1.998224e-07,1.998225e-07,1.998226e-07,1.998227e-07,1.998228e-07,1.998229e-07,1.998231e-07,1.998232e-07,1.998233e-07,1.998234e-07,1.998235e-07,1.998237e-07,1.998238e-07,1.998239e-07,1.998240e-07,1.998241e-07,1.998243e-07,1.998244e-07,1.998245e-07,1.998246e-07,1.998247e-07,1.998248e-07,1.998250e-07,1.998251e-07,1.998252e-07,1.998253e-07,1.998254e-07,1.998256e-07,1.998257e-07,1.998258e-07,1.998259e-07,1.998260e-07,1.998261e-07,1.998263e-07,1.998264e-07,1.998265e-07,1.998266e-07,1.998267e-07,1.998269e-07,1.998270e-07,1.998271e-07,1.998272e-07,1.998273e-07,1.998275e-07,1.998276e-07,1.998277e-07,1.998278e-07,1.998279e-07,1.998280e-07,1.998282e-07,1.998283e-07,1.998284e-07,1.998285e-07,1.998286e-07,1.998288e-07,1.998289e-07,1.998290e-07,1.998291e-07,1.998292e-07,1.998294e-07,1.998295e-07,1.998296e-07,1.998297e-07,1.998298e-07,1.998299e-07,1.998301e-07,1.998302e-07,1.998303e-07,1.998304e-07,1.998305e-07,1.998307e-07,1.998308e-07,1.998309e-07,1.998310e-07,1.998311e-07,1.998312e-07,1.998314e-07,1.998315e-07,1.998316e-07,1.998317e-07,1.998318e-07,1.998320e-07,1.998321e-07,1.998322e-07,1.998323e-07,1.998324e-07,1.998326e-07,1.998327e-07,1.998328e-07,1.998329e-07,1.998330e-07,1.998331e-07,1.998333e-07,1.998334e-07,1.998335e-07,1.998336e-07,1.998337e-07,1.998339e-07,1.998340e-07,1.998341e-07,1.998342e-07,1.998343e-07,1.998344e-07,1.998346e-07,1.998347e-07,1.998348e-07,1.998349e-07,1.998350e-07,1.998352e-07,1.998353e-07,1.998354e-07,1.998355e-07,1.998356e-07,1.998358e-07,1.998359e-07,1.998360e-07,1.998361e-07,1.998362e-07,1.998363e-07,1.998365e-07,1.998366e-07,1.998367e-07,1.998368e-07,1.998369e-07,1.998371e-07,1.998372e-07,1.998373e-07,1.998374e-07,1.998375e-07,1.998376e-07,1.998378e-07,1.998379e-07,1.998380e-07,1.998381e-07,1.998382e-07,1.998384e-07,1.998385e-07,1.998386e-07,1.998387e-07,1.998388e-07,1.998389e-07,1.998391e-07,1.998392e-07,1.998393e-07,1.998394e-07,1.998395e-07,1.998397e-07,1.998398e-07,1.998399e-07,1.998400e-07,1.998401e-07,1.998403e-07,1.998404e-07,1.998405e-07,1.998406e-07,1.998407e-07,1.998408e-07,1.998410e-07,1.998411e-07,1.998412e-07,1.998413e-07,1.998414e-07,1.998416e-07,1.998417e-07,1.998418e-07,1.998419e-07,1.998420e-07,1.998421e-07,1.998423e-07,1.998424e-07,1.998425e-07,1.998426e-07,1.998427e-07,1.998429e-07,1.998430e-07,1.998431e-07,1.998432e-07,1.998433e-07,1.998434e-07,1.998436e-07,1.998437e-07,1.998438e-07,1.998439e-07,1.998440e-07,1.998442e-07,1.998443e-07,1.998444e-07,1.998445e-07,1.998446e-07,1.998448e-07,1.998449e-07,1.998450e-07,1.998451e-07,1.998452e-07,1.998453e-07,1.998455e-07,1.998456e-07,1.998457e-07,1.998458e-07,1.998459e-07,1.998461e-07,1.998462e-07,1.998463e-07,1.998464e-07,1.998465e-07,1.998466e-07,1.998468e-07,1.998469e-07,1.998470e-07,1.998471e-07,1.998472e-07,1.998474e-07,1.998475e-07,1.998476e-07,1.998477e-07,1.998478e-07,1.998479e-07,1.998481e-07,1.998482e-07,1.998483e-07,1.998484e-07,1.998485e-07,1.998487e-07,1.998488e-07,1.998489e-07,1.998490e-07,1.998491e-07,1.998493e-07,1.998494e-07,1.998495e-07,1.998496e-07,1.998497e-07,1.998498e-07,1.998500e-07,1.998501e-07,1.998502e-07,1.998503e-07,1.998504e-07,1.998506e-07,1.998507e-07,1.998508e-07,1.998509e-07,1.998510e-07,1.998511e-07,1.998513e-07,1.998514e-07,1.998515e-07,1.998516e-07,1.998517e-07,1.998519e-07,1.998520e-07,1.998521e-07,1.998522e-07,1.998523e-07,1.998524e-07,1.998526e-07,1.998527e-07,1.998528e-07,1.998529e-07,1.998530e-07,1.998532e-07,1.998533e-07,1.998534e-07,1.998535e-07,1.998536e-07,1.998537e-07,1.998539e-07,1.998540e-07,1.998541e-07,1.998542e-07,1.998543e-07,1.998545e-07,1.998546e-07,1.998547e-07,1.998548e-07,1.998549e-07,1.998550e-07,1.998552e-07,1.998553e-07,1.998554e-07,1.998555e-07,1.998556e-07,1.998558e-07,1.998559e-07,1.998560e-07,1.998561e-07,1.998562e-07,1.998563e-07,1.998565e-07,1.998566e-07,1.998567e-07,1.998568e-07,1.998569e-07,1.998571e-07,1.998572e-07,1.998573e-07,1.998574e-07,1.998575e-07,1.998577e-07,1.998578e-07,1.998579e-07,1.998580e-07,1.998581e-07,1.998582e-07,1.998584e-07,1.998585e-07,1.998586e-07,1.998587e-07,1.998588e-07,1.998590e-07,1.998591e-07,1.998592e-07,1.998593e-07,1.998594e-07,1.998595e-07,1.998597e-07,1.998598e-07,1.998599e-07,1.998600e-07,1.998601e-07,1.998603e-07,1.998604e-07,1.998605e-07,1.998606e-07,1.998607e-07,1.998608e-07,1.998610e-07,1.998611e-07,1.998612e-07,1.998613e-07,1.998614e-07,1.998616e-07,1.998617e-07,1.998618e-07,1.998619e-07,1.998620e-07,1.998621e-07,1.998623e-07,1.998624e-07,1.998625e-07,1.998626e-07,1.998627e-07,1.998629e-07,1.998630e-07,1.998631e-07,1.998632e-07,1.998633e-07,1.998634e-07,1.998636e-07,1.998637e-07,1.998638e-07,1.998639e-07,1.998640e-07,1.998642e-07,1.998643e-07,1.998644e-07,1.998645e-07,1.998646e-07,1.998647e-07,1.998649e-07,1.998650e-07,1.998651e-07,1.998652e-07,1.998653e-07,1.998655e-07,1.998656e-07,1.998657e-07,1.998658e-07,1.998659e-07,1.998660e-07,1.998662e-07,1.998663e-07,1.998664e-07,1.998665e-07,1.998666e-07,1.998668e-07,1.998669e-07,1.998670e-07,1.998671e-07,1.998672e-07,1.998673e-07,1.998675e-07,1.998676e-07,1.998677e-07,1.998678e-07,1.998679e-07,1.998681e-07,1.998682e-07,1.998683e-07,1.998684e-07,1.998685e-07,1.998686e-07,1.998688e-07,1.998689e-07,1.998690e-07,1.998691e-07,1.998692e-07,1.998694e-07,1.998695e-07,1.998696e-07,1.998697e-07,1.998698e-07,1.998699e-07,1.998701e-07,1.998702e-07,1.998703e-07,1.998704e-07,1.998705e-07,1.998707e-07,1.998708e-07,1.998709e-07,1.998710e-07,1.998711e-07,1.998712e-07,1.998714e-07,1.998715e-07,1.998716e-07,1.998717e-07,1.998718e-07,1.998720e-07,1.998721e-07,1.998722e-07,1.998723e-07,1.998724e-07,1.998725e-07,1.998727e-07,1.998728e-07,1.998729e-07,1.998730e-07,1.998731e-07,1.998733e-07,1.998734e-07,1.998735e-07,1.998736e-07,1.998737e-07,1.998738e-07,1.998740e-07,1.998741e-07,1.998742e-07,1.998743e-07,1.998744e-07,1.998745e-07,1.998747e-07,1.998748e-07,1.998749e-07,1.998750e-07,1.998751e-07,1.998753e-07,1.998754e-07,1.998755e-07,1.998756e-07,1.998757e-07,1.998758e-07,1.998760e-07,1.998761e-07,1.998762e-07,1.998763e-07,1.998764e-07,1.998766e-07,1.998767e-07,1.998768e-07,1.998769e-07,1.998770e-07,1.998771e-07,1.998773e-07,1.998774e-07,1.998775e-07,1.998776e-07,1.998777e-07,1.998779e-07,1.998780e-07,1.998781e-07,1.998782e-07,1.998783e-07,1.998784e-07,1.998786e-07,1.998787e-07,1.998788e-07,1.998789e-07,1.998790e-07,1.998792e-07,1.998793e-07,1.998794e-07,1.998795e-07,1.998796e-07,1.998797e-07,1.998799e-07,1.998800e-07,1.998801e-07,1.998802e-07,1.998803e-07,1.998805e-07,1.998806e-07,1.998807e-07,1.998808e-07,1.998809e-07,1.998810e-07,1.998812e-07,1.998813e-07,1.998814e-07,1.998815e-07,1.998816e-07,1.998818e-07,1.998819e-07,1.998820e-07,1.998821e-07,1.998822e-07,1.998823e-07,1.998825e-07,1.998826e-07,1.998827e-07,1.998828e-07,1.998829e-07,1.998830e-07,1.998832e-07,1.998833e-07,1.998834e-07,1.998835e-07,1.998836e-07,1.998838e-07,1.998839e-07,1.998840e-07,1.998841e-07,1.998842e-07,1.998843e-07,1.998845e-07,1.998846e-07,1.998847e-07,1.998848e-07,1.998849e-07,1.998851e-07,1.998852e-07,1.998853e-07,1.998854e-07,1.998855e-07,1.998856e-07,1.998858e-07,1.998859e-07,1.998860e-07,1.998861e-07,1.998862e-07,1.998864e-07,1.998865e-07,1.998866e-07,1.998867e-07,1.998868e-07,1.998869e-07,1.998871e-07,1.998872e-07,1.998873e-07,1.998874e-07,1.998875e-07,1.998877e-07,1.998878e-07,1.998879e-07,1.998880e-07,1.998881e-07,1.998882e-07,1.998884e-07,1.998885e-07,1.998886e-07,1.998887e-07,1.998888e-07,1.998889e-07,1.998891e-07,1.998892e-07,1.998893e-07,1.998894e-07,1.998895e-07,1.998897e-07,1.998898e-07,1.998899e-07,1.998900e-07,1.998901e-07,1.998902e-07,1.998904e-07,1.998905e-07,1.998906e-07,1.998907e-07,1.998908e-07,1.998910e-07,1.998911e-07,1.998912e-07,1.998913e-07,1.998914e-07,1.998915e-07,1.998917e-07,1.998918e-07,1.998919e-07,1.998920e-07,1.998921e-07,1.998923e-07,1.998924e-07,1.998925e-07,1.998926e-07,1.998927e-07,1.998928e-07,1.998930e-07,1.998931e-07,1.998932e-07,1.998933e-07,1.998934e-07,1.998935e-07,1.998937e-07,1.998938e-07,1.998939e-07,1.998940e-07,1.998941e-07,1.998943e-07,1.998944e-07,1.998945e-07,1.998946e-07,1.998947e-07,1.998948e-07,1.998950e-07,1.998951e-07,1.998952e-07,1.998953e-07,1.998954e-07,1.998956e-07,1.998957e-07,1.998958e-07,1.998959e-07,1.998960e-07,1.998961e-07,1.998963e-07,1.998964e-07,1.998965e-07,1.998966e-07,1.998967e-07,1.998968e-07,1.998970e-07,1.998971e-07,1.998972e-07,1.998973e-07,1.998974e-07,1.998976e-07,1.998977e-07,1.998978e-07,1.998979e-07,1.998980e-07,1.998981e-07,1.998983e-07,1.998984e-07,1.998985e-07,1.998986e-07,1.998987e-07,1.998989e-07,1.998990e-07,1.998991e-07,1.998992e-07,1.998993e-07,1.998994e-07,1.998996e-07,1.998997e-07,1.998998e-07,1.998999e-07,1.999000e-07,1.999001e-07,1.999003e-07,1.999004e-07,1.999005e-07,1.999006e-07,1.999007e-07,1.999009e-07,1.999010e-07,1.999011e-07,1.999012e-07,1.999013e-07,1.999014e-07,1.999016e-07,1.999017e-07,1.999018e-07,1.999019e-07,1.999020e-07,1.999022e-07,1.999023e-07,1.999024e-07,1.999025e-07,1.999026e-07,1.999027e-07,1.999029e-07,1.999030e-07,1.999031e-07,1.999032e-07,1.999033e-07,1.999034e-07,1.999036e-07,1.999037e-07,1.999038e-07,1.999039e-07,1.999040e-07,1.999042e-07,1.999043e-07,1.999044e-07,1.999045e-07,1.999046e-07,1.999047e-07,1.999049e-07,1.999050e-07,1.999051e-07,1.999052e-07,1.999053e-07,1.999054e-07,1.999056e-07,1.999057e-07,1.999058e-07,1.999059e-07,1.999060e-07,1.999062e-07,1.999063e-07,1.999064e-07,1.999065e-07,1.999066e-07,1.999067e-07,1.999069e-07,1.999070e-07,1.999071e-07,1.999072e-07,1.999073e-07,1.999075e-07,1.999076e-07,1.999077e-07,1.999078e-07,1.999079e-07,1.999080e-07,1.999082e-07,1.999083e-07,1.999084e-07,1.999085e-07,1.999086e-07,1.999087e-07,1.999089e-07,1.999090e-07,1.999091e-07,1.999092e-07,1.999093e-07,1.999095e-07,1.999096e-07,1.999097e-07,1.999098e-07,1.999099e-07,1.999100e-07,1.999102e-07,1.999103e-07,1.999104e-07,1.999105e-07,1.999106e-07,1.999107e-07,1.999109e-07,1.999110e-07,1.999111e-07,1.999112e-07,1.999113e-07,1.999115e-07,1.999116e-07,1.999117e-07,1.999118e-07,1.999119e-07,1.999120e-07,1.999122e-07,1.999123e-07,1.999124e-07,1.999125e-07,1.999126e-07,1.999127e-07,1.999129e-07,1.999130e-07,1.999131e-07,1.999132e-07,1.999133e-07,1.999135e-07,1.999136e-07,1.999137e-07,1.999138e-07,1.999139e-07,1.999140e-07,1.999142e-07,1.999143e-07,1.999144e-07,1.999145e-07,1.999146e-07,1.999148e-07,1.999149e-07,1.999150e-07,1.999151e-07,1.999152e-07,1.999153e-07,1.999155e-07,1.999156e-07,1.999157e-07,1.999158e-07,1.999159e-07,1.999160e-07,1.999162e-07,1.999163e-07,1.999164e-07,1.999165e-07,1.999166e-07,1.999168e-07,1.999169e-07,1.999170e-07,1.999171e-07,1.999172e-07,1.999173e-07,1.999175e-07,1.999176e-07,1.999177e-07,1.999178e-07,1.999179e-07,1.999180e-07,1.999182e-07,1.999183e-07,1.999184e-07,1.999185e-07,1.999186e-07,1.999188e-07,1.999189e-07,1.999190e-07,1.999191e-07,1.999192e-07,1.999193e-07,1.999195e-07,1.999196e-07,1.999197e-07,1.999198e-07,1.999199e-07,1.999200e-07,1.999202e-07,1.999203e-07,1.999204e-07,1.999205e-07,1.999206e-07,1.999208e-07,1.999209e-07,1.999210e-07,1.999211e-07,1.999212e-07,1.999213e-07,1.999215e-07,1.999216e-07,1.999217e-07,1.999218e-07,1.999219e-07,1.999220e-07,1.999222e-07,1.999223e-07,1.999224e-07,1.999225e-07,1.999226e-07,1.999228e-07,1.999229e-07,1.999230e-07,1.999231e-07,1.999232e-07,1.999233e-07,1.999235e-07,1.999236e-07,1.999237e-07,1.999238e-07,1.999239e-07,1.999240e-07,1.999242e-07,1.999243e-07,1.999244e-07,1.999245e-07,1.999246e-07,1.999247e-07,1.999249e-07,1.999250e-07,1.999251e-07,1.999252e-07,1.999253e-07,1.999255e-07,1.999256e-07,1.999257e-07,1.999258e-07,1.999259e-07,1.999260e-07,1.999262e-07,1.999263e-07,1.999264e-07,1.999265e-07,1.999266e-07,1.999267e-07,1.999269e-07,1.999270e-07,1.999271e-07,1.999272e-07,1.999273e-07,1.999275e-07,1.999276e-07,1.999277e-07,1.999278e-07,1.999279e-07,1.999280e-07,1.999282e-07,1.999283e-07,1.999284e-07,1.999285e-07,1.999286e-07,1.999287e-07,1.999289e-07,1.999290e-07,1.999291e-07,1.999292e-07,1.999293e-07,1.999295e-07,1.999296e-07,1.999297e-07,1.999298e-07,1.999299e-07,1.999300e-07,1.999302e-07,1.999303e-07,1.999304e-07,1.999305e-07,1.999306e-07,1.999307e-07,1.999309e-07,1.999310e-07,1.999311e-07,1.999312e-07,1.999313e-07,1.999315e-07,1.999316e-07,1.999317e-07,1.999318e-07,1.999319e-07,1.999320e-07,1.999322e-07,1.999323e-07,1.999324e-07,1.999325e-07,1.999326e-07,1.999327e-07,1.999329e-07,1.999330e-07,1.999331e-07,1.999332e-07,1.999333e-07,1.999334e-07,1.999336e-07,1.999337e-07,1.999338e-07,1.999339e-07,1.999340e-07,1.999342e-07,1.999343e-07,1.999344e-07,1.999345e-07,1.999346e-07,1.999347e-07,1.999349e-07,1.999350e-07,1.999351e-07,1.999352e-07,1.999353e-07,1.999354e-07,1.999356e-07,1.999357e-07,1.999358e-07,1.999359e-07,1.999360e-07,1.999362e-07,1.999363e-07,1.999364e-07,1.999365e-07,1.999366e-07,1.999367e-07,1.999369e-07,1.999370e-07,1.999371e-07,1.999372e-07,1.999373e-07,1.999374e-07,1.999376e-07,1.999377e-07,1.999378e-07,1.999379e-07,1.999380e-07,1.999381e-07,1.999383e-07,1.999384e-07,1.999385e-07,1.999386e-07,1.999387e-07,1.999389e-07,1.999390e-07,1.999391e-07,1.999392e-07,1.999393e-07,1.999394e-07,1.999396e-07,1.999397e-07,1.999398e-07,1.999399e-07,1.999400e-07,1.999401e-07,1.999403e-07,1.999404e-07,1.999405e-07,1.999406e-07,1.999407e-07,1.999408e-07,1.999410e-07,1.999411e-07,1.999412e-07,1.999413e-07,1.999414e-07,1.999416e-07,1.999417e-07,1.999418e-07,1.999419e-07,1.999420e-07,1.999421e-07,1.999423e-07,1.999424e-07,1.999425e-07,1.999426e-07,1.999427e-07,1.999428e-07,1.999430e-07,1.999431e-07,1.999432e-07,1.999433e-07,1.999434e-07,1.999435e-07,1.999437e-07,1.999438e-07,1.999439e-07,1.999440e-07,1.999441e-07,1.999443e-07,1.999444e-07,1.999445e-07,1.999446e-07,1.999447e-07,1.999448e-07,1.999450e-07,1.999451e-07,1.999452e-07,1.999453e-07,1.999454e-07,1.999455e-07,1.999457e-07,1.999458e-07,1.999459e-07,1.999460e-07,1.999461e-07,1.999462e-07,1.999464e-07,1.999465e-07,1.999466e-07,1.999467e-07,1.999468e-07,1.999470e-07,1.999471e-07,1.999472e-07,1.999473e-07,1.999474e-07,1.999475e-07,1.999477e-07,1.999478e-07,1.999479e-07,1.999480e-07,1.999481e-07,1.999482e-07,1.999484e-07,1.999485e-07,1.999486e-07,1.999487e-07,1.999488e-07,1.999489e-07,1.999491e-07,1.999492e-07,1.999493e-07,1.999494e-07,1.999495e-07,1.999497e-07,1.999498e-07,1.999499e-07,1.999500e-07,1.999501e-07,1.999502e-07,1.999504e-07,1.999505e-07,1.999506e-07,1.999507e-07,1.999508e-07,1.999509e-07,1.999511e-07,1.999512e-07,1.999513e-07,1.999514e-07,1.999515e-07,1.999516e-07,1.999518e-07,1.999519e-07,1.999520e-07,1.999521e-07,1.999522e-07,1.999524e-07,1.999525e-07,1.999526e-07,1.999527e-07,1.999528e-07,1.999529e-07,1.999531e-07,1.999532e-07,1.999533e-07,1.999534e-07,1.999535e-07,1.999536e-07,1.999538e-07,1.999539e-07,1.999540e-07,1.999541e-07,1.999542e-07,1.999543e-07,1.999545e-07,1.999546e-07,1.999547e-07,1.999548e-07,1.999549e-07,1.999550e-07,1.999552e-07,1.999553e-07,1.999554e-07,1.999555e-07,1.999556e-07,1.999558e-07,1.999559e-07,1.999560e-07,1.999561e-07,1.999562e-07,1.999563e-07,1.999565e-07,1.999566e-07,1.999567e-07,1.999568e-07,1.999569e-07,1.999570e-07,1.999572e-07,1.999573e-07,1.999574e-07,1.999575e-07,1.999576e-07,1.999577e-07,1.999579e-07,1.999580e-07,1.999581e-07,1.999582e-07,1.999583e-07,1.999584e-07,1.999586e-07,1.999587e-07,1.999588e-07,1.999589e-07,1.999590e-07,1.999592e-07,1.999593e-07,1.999594e-07,1.999595e-07,1.999596e-07,1.999597e-07,1.999599e-07,1.999600e-07,1.999601e-07,1.999602e-07,1.999603e-07,1.999604e-07,1.999606e-07,1.999607e-07,1.999608e-07,1.999609e-07,1.999610e-07,1.999611e-07,1.999613e-07,1.999614e-07,1.999615e-07,1.999616e-07,1.999617e-07,1.999618e-07,1.999620e-07,1.999621e-07,1.999622e-07,1.999623e-07,1.999624e-07,1.999626e-07,1.999627e-07,1.999628e-07,1.999629e-07,1.999630e-07,1.999631e-07,1.999633e-07,1.999634e-07,1.999635e-07,1.999636e-07,1.999637e-07,1.999638e-07,1.999640e-07,1.999641e-07,1.999642e-07,1.999643e-07,1.999644e-07,1.999645e-07,1.999647e-07,1.999648e-07,1.999649e-07,1.999650e-07,1.999651e-07,1.999652e-07,1.999654e-07,1.999655e-07,1.999656e-07,1.999657e-07,1.999658e-07,1.999660e-07,1.999661e-07,1.999662e-07,1.999663e-07,1.999664e-07,1.999665e-07,1.999667e-07,1.999668e-07,1.999669e-07,1.999670e-07,1.999671e-07,1.999672e-07,1.999674e-07,1.999675e-07,1.999676e-07,1.999677e-07,1.999678e-07,1.999679e-07,1.999681e-07,1.999682e-07,1.999683e-07,1.999684e-07,1.999685e-07,1.999686e-07,1.999688e-07,1.999689e-07,1.999690e-07,1.999691e-07,1.999692e-07,1.999693e-07,1.999695e-07,1.999696e-07,1.999697e-07,1.999698e-07,1.999699e-07,1.999701e-07,1.999702e-07,1.999703e-07,1.999704e-07,1.999705e-07,1.999706e-07,1.999708e-07,1.999709e-07,1.999710e-07,1.999711e-07,1.999712e-07,1.999713e-07,1.999715e-07,1.999716e-07,1.999717e-07,1.999718e-07,1.999719e-07,1.999720e-07,1.999722e-07,1.999723e-07,1.999724e-07,1.999725e-07,1.999726e-07,1.999727e-07,1.999729e-07,1.999730e-07,1.999731e-07,1.999732e-07,1.999733e-07,1.999734e-07,1.999736e-07,1.999737e-07,1.999738e-07,1.999739e-07,1.999740e-07,1.999742e-07,1.999743e-07,1.999744e-07,1.999745e-07,1.999746e-07,1.999747e-07,1.999749e-07,1.999750e-07,1.999751e-07,1.999752e-07,1.999753e-07,1.999754e-07,1.999756e-07,1.999757e-07,1.999758e-07,1.999759e-07,1.999760e-07,1.999761e-07,1.999763e-07,1.999764e-07,1.999765e-07,1.999766e-07,1.999767e-07,1.999768e-07,1.999770e-07,1.999771e-07,1.999772e-07,1.999773e-07,1.999774e-07,1.999775e-07,1.999777e-07,1.999778e-07,1.999779e-07,1.999780e-07,1.999781e-07,1.999782e-07,1.999784e-07,1.999785e-07,1.999786e-07,1.999787e-07,1.999788e-07,1.999790e-07,1.999791e-07,1.999792e-07,1.999793e-07,1.999794e-07,1.999795e-07,1.999797e-07,1.999798e-07,1.999799e-07,1.999800e-07,1.999801e-07,1.999802e-07,1.999804e-07,1.999805e-07,1.999806e-07,1.999807e-07,1.999808e-07,1.999809e-07,1.999811e-07,1.999812e-07,1.999813e-07,1.999814e-07,1.999815e-07,1.999816e-07,1.999818e-07,1.999819e-07,1.999820e-07,1.999821e-07,1.999822e-07,1.999823e-07,1.999825e-07,1.999826e-07,1.999827e-07,1.999828e-07,1.999829e-07,1.999830e-07,1.999832e-07,1.999833e-07,1.999834e-07,1.999835e-07,1.999836e-07,1.999837e-07,1.999839e-07,1.999840e-07,1.999841e-07,1.999842e-07,1.999843e-07,1.999845e-07,1.999846e-07,1.999847e-07,1.999848e-07,1.999849e-07,1.999850e-07,1.999852e-07,1.999853e-07,1.999854e-07,1.999855e-07,1.999856e-07,1.999857e-07,1.999859e-07,1.999860e-07,1.999861e-07,1.999862e-07,1.999863e-07,1.999864e-07,1.999866e-07,1.999867e-07,1.999868e-07,1.999869e-07,1.999870e-07,1.999871e-07,1.999873e-07,1.999874e-07,1.999875e-07,1.999876e-07,1.999877e-07,1.999878e-07,1.999880e-07,1.999881e-07,1.999882e-07,1.999883e-07,1.999884e-07,1.999885e-07,1.999887e-07,1.999888e-07,1.999889e-07,1.999890e-07,1.999891e-07,1.999892e-07,1.999894e-07,1.999895e-07,1.999896e-07,1.999897e-07,1.999898e-07,1.999899e-07,1.999901e-07,1.999902e-07,1.999903e-07,1.999904e-07,1.999905e-07,1.999906e-07,1.999908e-07,1.999909e-07,1.999910e-07,1.999911e-07,1.999912e-07,1.999914e-07,1.999915e-07,1.999916e-07,1.999917e-07,1.999918e-07,1.999919e-07,1.999921e-07,1.999922e-07,1.999923e-07,1.999924e-07,1.999925e-07,1.999926e-07,1.999928e-07,1.999929e-07,1.999930e-07,1.999931e-07,1.999932e-07,1.999933e-07,1.999935e-07,1.999936e-07,1.999937e-07,1.999938e-07,1.999939e-07,1.999940e-07,1.999942e-07,1.999943e-07,1.999944e-07,1.999945e-07,1.999946e-07,1.999947e-07,1.999949e-07,1.999950e-07,1.999951e-07,1.999952e-07,1.999953e-07,1.999954e-07,1.999956e-07,1.999957e-07,1.999958e-07,1.999959e-07,1.999960e-07,1.999961e-07,1.999963e-07,1.999964e-07,1.999965e-07,1.999966e-07,1.999967e-07,1.999968e-07,1.999970e-07,1.999971e-07,1.999972e-07,1.999973e-07,1.999974e-07,1.999975e-07,1.999977e-07,1.999978e-07,1.999979e-07,1.999980e-07,1.999981e-07,1.999982e-07,1.999984e-07,1.999985e-07,1.999986e-07,1.999987e-07,1.999988e-07,1.999989e-07,1.999991e-07,1.999992e-07,1.999993e-07,1.999994e-07,1.999995e-07,1.999996e-07,1.999998e-07,1.999999e-07,2.000000e-07 PRINTFOOTER=false
