Netlist to Test the Xyce Voltage Controlled Current Source Model, multiplier version
******************************************************************************
*	Based on the original vccs.cir test, but current is 10x larger.
*
* This is modified from vccs_m, to use the expression library.  This means that
* behind the scenes, Xyce will convert this to a Bsource.  So, this test 
* effectively tests is (1) the Bsrc multiplier works and (2) if the internal 
* conversion from Gsource to Bsource works correctly.
*
* This test has been modified from vccs_nl1_m.cir to place the G-source inside 
* a subcircuit.   There is a multiplier on the subcircuit, that is subsequently
* applied to the G-source.
*
* This case is linear, but the use of expressions allows for nonlinear G-sources.
****************************************************************************** 
VIN 1 0 DC 12V
Xtest 3 0 2 0 gsrcSub m=10

.subckt gsrcSub A B C D M=1
G A B cur='v(C,D)*0.02' M='M'
.ends

R1 1 2 300
R2 2 0 900
R3 3 0 200
R4 3 0 200
.DC VIN 1 12 1
.PRINT DC V(1) V(2) V(3) 
* NOTE: XYCE DOES NOT CURRENTLY SUPPORT TRANSFER FUNCTION ANALYSIS 
* THIS PORTION HAS BEEN COMMENTED OUT UNTIL TF IS SUPPORTED
*.TF V(3) V
.END
