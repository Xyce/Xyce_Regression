Test for bug 797 SON.  Direct sensitivity baseline.
********************************************************************************

.param cap=1e-6
.param res=1e3

V1 1 0 0.0 sin (0.0 1.0 200 0.0 0.0 0.0 )
R1 1 2 {res}
C1 2 0 {V(5)}

B2 5 0 V={cap+0.01*(time)}
R2 5 0 

.tran 1.0e-6 0.5e-2

.print tran V(1) V(2) 
.print TRANADJOINT 

.options timeint method=gear  debuglevel=-100 conststep=0  
.options device debuglevel=-100

.SENS objfunc={V(2)} param=R1:R
.options SENSITIVITY direct=0 adjoint=1  diagnosticfile=0  stdoutput=0 

.end

