A test of .OPTIONS MEASURE MEASFAIL=1  
* That option value takes precedence over the DEFAULT_VAL qualifier
* on the .MEASURE lines.  It also takes precedence over 
* .OPTIONS MEASURE DEFAULT_VAL=<val>.
*
* This test uses new TRIG-TARG mode,  so it tests the
* TrigTarg classes.  See gitlab-ex issue 303 for more details.
*******************************************************************
VS2  2  0  SIN(0 -1.0 1KHz 0 0.9)
R2  2  0  100

.TRAN 0  1ms
.OPTIONS OUTPUT INITIAL_INTERVAL=0.00001
.PRINT TRAN FORMAT=NOINDEX V(2)
.OPTIONS MEASURE DEFAULT_VAL=-100
.OPTIONS MEASURE MEASFAIL=1

*TRIG/TARG
.measure tran trigTargAtFail TRIG AT=2e-3 TARG V(2)=0.5 DEFAULT_VAL=2

* for testing convenience do not make separate .mt0 files
* for each TRAN_CONT measure
.OPTIONS MEASURE USE_CONT_FILES=0
.measure tran_cont trigTargContAtFail TRIG AT=2e-3 TARG V(2)=0.5 DEFAULT_VAL=2

.END
