*** Simple amplifier sensitivity test for transient adjoints
*
* Taken from Spice OPUS website: http://fides.fe.uni-lj.si/spice/opt001.html
vcc 1 0 dc 12V
i1 2 0 sin(100uA 600uA 1e6 )

r1 1 3 5k
r2 2 3 20k

q1 3 2 0 2n3510

.model 2n3510 npn
+ bf=100 br=1.35e-4 xtb=1.5 is=8.35e-14 eg=1.11 cjc=9.63e-12
+ cje=9.47e-12 rb=16.7 rc=1.66 vaf=90 tf=1e-10 tr=1.27e-4
+ cjs=1e-15 vjs=0.8 mjs=0.5 var=100 ise=4.77e-11 isc=1e-16
+ ikf=0.18 ikr=1000 irb=1 rbm=0 vtf=1000

.SENS param=R1:R
+objfunc={V(3)} 

.options SENSITIVITY direct=1 adjoint=0  diagnosticfile=0 STDOUTPUT=0 debuglevel=-100 

.options timeint method=gear debuglevel=-100 
*maxord=1 

.tran 2ns 1us
.print tran v(3)
.print sens 

.end
