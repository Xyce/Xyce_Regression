UA555 Timer Circuit
********************************************************************************
* Tier No.: 2
* Directory/Circuit Name:SANDLER21/sandler21.cir
* Description:  UA555 timer circuit netlist developed by Steve Sandler to 
*       compare the validity of simulations using 3 different circuit
*       simulation tools.  The results were compared to measured data.
* Input: V2=V(6)
* Output: V(1), V(4), V(6)
* Analysis:
********************************************************************************
*
.SUBCKT UA555  32 30 19 23 33 1  21 
*              TR O  R  F  TH D  V  
*
Q4 25 2 3 QP
Q5 0 6 3 QP
Q6 6 6 8 QP
R1 9 21 4.7K
R2 3 21 830
R3 8 21 4.7K
Q7 2 33 5 QN
Q8 2 5 17 QN
Q9 6 4 17 QN
Q10 6 23 4 QN
Q11 12 20 10 QP
R4 10 21 1K
Q12 22 11 12 QP
Q13 14 13 12 QP
Q14 0 32 11 QP
Q15 14 18 13 QP
R5 14 0 100K
R6 22 0 100K
R7 17 0 10K
Q16 1 15 0 QN
Q17 15 19 31 QP
R8 18 23 5K
R9 18 0 5K
R10 21 23 5K
Q18 27 20 21 QP
Q19 20 20 21 QP
R11 20 31 5K
D1 31 24 DA
Q20 24 25 0 QN
Q21 25 22 0 QN
Q22 27 24 0 QN
R12 25 27 4.7K
R13 21 29 6.8K
Q23 21 29 28 QN
Q24 29 27 16 QN
Q25 30 26 0 QN
Q26 21 28 30 QN
D2 30 29 DA
R14 16 15 100
R15 16 26 220
R16 16 0 4.7K
R17 28 30 3.9K
Q3 2 2 9 QP
*
.MODEL DA D (RS=40 IS=1.0E-14 CJO=1PF)
.MODEL QP PNP (BF=20 BR=0.02 RC=4 RB=25 IS=1.0E-14 VAF=50 NE=2
+ CJE=12.4P VJE=1.1 MJE=.5 CJC=4.02P VJC=.3 MJC=.3 TF=229P TR=159N)
.MODEL QN NPN (IS=5.07F NF=1 BF=100 VAF=161 IKF=30M ISE=3.9P NE=2       
+ BR=4 NR=1 VAR=16 IKR=45M RE=1.03 RB=4.12 RC=.412 XTB=1.5      
+ CJE=12.4P VJE=1.1 MJE=.5 CJC=4.02P VJC=.3 MJC=.3 TF=229P TR=959P)
.ENDS
**********************************************************************************
*
.param RVAL={76K+i(c2)}
* MAIN CIRCUIT
C1 1 0 2140P
R2 3 1 {RVAL}
C2 5 0 .01U
X2 6 4 3 5 1 1 3 UA555
V2 6 0 PULSE(0 15 0U .1U .1U 900U 1M)
V1 3 0 15
*
.TRAN 1U 5M
.PRINT TRAN V(4)  V(1)  V(6)
*ALIAS  V(4)=OUT V(1)=RAMP V(6)=TRIGGER
.END

