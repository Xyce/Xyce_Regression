*******************************************************
* Test of AC output with FILE= and FORMAT= qualifiers.
* This netlist has a .OP statement so that the .TD.csv
* file is also made.  See SON Bug 701 for more
* details.
*
* Trivial high-pass filter (V-C-R) circuit, just do
* an AC sweep and watch the output.
*
*****************************************************
R1 b 0 2
C1 a b 1u
V1 a 0 DC 0V AC 1

* Generate the time-domain output with a fallback
* .PRINT AC_IC line
.print AC FILE=ac_foo_csv FORMAT=CSV vr(b) vi(b)

.OP
.ac dec 5 100Hz 10e6

.end

