Bug 1358:  test for quoted expressions. (regression)

.param resistance = '2.0'

VT1 4 0 0V
R1  4 0 'resistance*5.0' 

.DC VT1 -0.2 0.5 0.01  
.print DC v(4) '(abs(I(VT1)))' '(V(4)**2.0)' I(VT1) 

.END

