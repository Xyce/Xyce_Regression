Regression test to show transient adjoint sensitivities for second order Gear time integration.
********************************************************************************

.param cap=1e-6
.param res=1e3

V1 1 0 0.0 sin (0.0 1.0 200 0.0 0.0 0.0 )
R1 1 2 {res}
C1 2 0 {cap}

.tran 1.0e-6 0.5e-2

*comp   {V(2)}  offset=0.7
*comp d{V(2)}/d(R1:R)_Adj offset=0.0004
*comp d{V(2)}/d(C1:C)_Adj offset=400000

.print tran V(1) V(2) 
.print TRANADJOINT 
* this is here to fool xyce verify.
.print sens

.options timeint method=gear  debuglevel=-100 conststep=0  reltol=1.0e-6 abstol=1e-6
.options device debuglevel=-100

.SENS objfunc={V(2)} param=R1:R,C1:C
.options SENSITIVITY direct=0 adjoint=1  diagnosticfile=0  stdoutput=0 
+ adjointTimePoints=0.1e-2, 0.2e-2, 0.3e-2, 0.4e-2, 0.5e-2

.end

