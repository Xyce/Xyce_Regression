* A test of whether DC mode for .MEASURE statements works with I, P and W
* 
* This bug covers:
*   1) the case of one variable in the .DC line, 
*      without a .STEP statement.
*
*   2) the use of a FROM and TO statement, where the FROM
*      value is less than TO value.
*
* See SON Bug 886 for more details.
*******************************************************************************
*

vsrc1   1a 0 1
rload1a 1a 1b 0.1
rload1b 1b 0 1

.DC vsrc1 1 5 1
* Note: vsrc1:DCV0 is the syntax for printing the DC value of vsrc1,
* at it is swept. 
.print dc vsrc1:DCV0 I(Rload1a) P(Rload1a) W(Rload1a) N(VSRC1_BRANCH)

* tests
.measure dc maxI max I(Rload1a)
.measure dc maxIFT max I(Rload1a) FROM=2 TO=4
.measure dc maxP max P(Rload1a)
.measure dc maxW max W(Rload1a)
.measure dc maxN max N(VSRC1_BRANCH)

.END

