Power test for MOSFET Level 2
*
VDS 4 0  5V
VGS  1   0  pulse (0 1 1ns 1ns 1ns 1us 5us)
VMOND 4 3 0V
VMONS 0 2 0V
VMONG 1 1a 0
VMONB 0 6 0

M1 3 1a 2 6 CD4012_NMOS L=5u W=175u
.MODEL cd4012_nmos NMOS (LEVEL = 2) 

.options timeint method=gear
.options nonlin-tran rhstol=1.0e-8
.tran 1ns 20us

* test that P(M1) and W(M1) are equal to the formula (Id*Vds + Ig*Vgs)
* and also equal to the combined power dissipation of the two
* source VDS and VGS.
.PRINT TRAN PRECISION=10 
+ P(M1) W(M1) {ID(M1)*V(4) + IG(M1)*V(1)} {-1*(P(VDS)+P(VGS))}
+ ID(M1) IG(M1) IS(M1) IB(M1) I(VDS) I(VGS) V(4) V(1) 

.END
