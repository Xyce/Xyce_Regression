Test for solution dependent resistor.

Vcontrol cntl 0 2.0
Rcontrol cntl 0 1.0

.param scalar=2.0

V1 1 0 2.0
R1 1 2 1.0
R2 2 0 R={1.0+scalar*V(cntl)}

.DC V1 2 2 1
.Print dc V(1) V(2) R2:R V(cntl) 
+ {1.0+scalar*V(cntl)}
+ {ddx(1.0+scalar*V(cntl),v(cntl))}
+ {1.0/(1.0+scalar*V(cntl))}
+ {ddx(1.0/(1.0+scalar*V(cntl)),v(cntl))}
+ I(V1)
+ {V(2)/(1.0+scalar*V(cntl))}
+ {ddx(V(2)/(1.0+scalar*V(cntl)),v(cntl))}

