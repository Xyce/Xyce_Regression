Lowpass filter from https://www.electronics-tutorials.ws/filter/filter_2.html
* this is identical to the lowpass.cir sensitivity test, except that I am intentionally 
* excluding v1:acmag.  The purpose of this circuit is to provide a "gold" standard for
* the lowpass_forceDeviceFD test.

* device parameters:
.param rval=4.7k
.param cval=47n
.param vinval=10.0

* Circuit:
v1 1 0 ac {vinval}
r1 1 2 {rval}
c1 2 0 {cval}

.ac dec 10 1 10k

* Output vp() in degrees
.OPTIONS OUTPUT PHASE_OUTPUT_RADIANS=true

.print ac 
+ vm(1) vp(1) vm(2) vp(2)   

.print sens 

.sens objvars=2 param=r1:r,c1:c
.options sensitivity direct=1 adjoint=1  stdoutput=1  

.options device debuglevel=-100

.end 
