*Trivial sweep of diode to produce I/V curve
* This netlist is intended to test the PSPICE-compatible model of 
* temperature-dependent diode breakdown voltage, as defined by the 
* parameters TBV1 and TBV2.  Until 6 May 2010, this feature did not work,
* and this netlist would fail when compared to the gold standard provided
* here.  The failure between pre-fix and post-fix code is evidenced by a 
* mere 1.09% integrated error, but it is definitely significant.  

.tran 0 1 0 100m
.step TEMP list -55 25 72 

*.print tran V(1) V(2) {-I(VIN)} TEMP
*.print tran format=probe  V(1) V(2) {-I(VIN)} TEMP
.print tran V(2) TEMP

* NOTE:  DO not loosen this tolerance, it needs to be this tight to catch
* the regression!
*COMP V(2) reltol=0.005

*We start the pulse pretty high, because we're really only interested in
* seeing where the breakdown is, and if we don't do this, the places where
* breakdown isn't happening make it look like the simulation is better than
* it is (i.e. they artificially reduce the integrated error).
VIN 1 0 pulse ( 7.5 10 1m 1 1 3 6)
R1  1 2 1k
DZR 0 2 DZR  
.MODEL DZR D( level=2
+         IS = 1E-14
+         RS = 0
+          N = 1
+         TT = 0
+        CJO = 1P
+         VJ = 1
+          M = .5
+         EG = 1.11
+        XTI = 3
+         KF = 0
+         AF = 1
+         FC = .5
+         BV = 7.255;7.25 yields vout=5V @25C;6.9504;Vref determines Vout
+        IBV = .001
+ tbv1 = 0.00013
+ tbv2 = -5e-8
+        
+ )
