*Xyce netlist for testing H-sources syntaxes

.TRAN 0 1000ns
.PRINT TRAN FORMAT=PROBE V(N390192) V(N390144) I(V_V8) I(R_R15) 
*+ V(N390344) V(N390288)

R_R12         0 N390186  1 
R_R13         0 N390144  1
V_V7         N390192 0  SIN(0V 1 1e6 0 0 0)
X_H1    N390192 N390186 N390144 0 SCHEMATIC1_H1 

.subckt SCHEMATIC1_H1 1 2 3 4  
H_H1         3 4 VH_H1 2
VH_H1         1 2 0V
.ends SCHEMATIC1_H1

* test POLY form of the H-source
R_R14        0 N390338  1
V_V8         N390338 0  SIN (0V 2V 1e6 0 0 0)
R_R15        0 N390388  1

H_H2 N390388 0 POLY(1) V_V8 0 2

* test POLY Form of H-Source.  This is commented out since
* the gold and translated Xyce netlists do not give the same
* results for this sub-circuit version of the POLY H-Source
* produced by the OrCAD Capture UI.
*V_V8         N390344 0  SIN(0 2 1e6 0 0 0)
*R_R14         0 N390338  1 
*R_R15         0 N390288  1 TC=0,0 
*X_H2    N390344 N390338 N390288 0 SCHEMATIC1_H2

*.subckt SCHEMATIC1_H2 1 2 3 4  
*H_H2         3 4 POLY(1) VH_H2 2
*VH_H2         1 2 0
*.ends SCHEMATIC1_H2

.END