* Test the BINSIZ parameter for the ENOB, SFDR and SNDR
* measure types for .MEASURE FFT for a .TRAN analysis.
*
* See git issue 256 for more details
******************************************************

.TRAN 0 1
.OPTIONS FFT FFT_ACCURATE=1 FFTOUT=1

V7 7 0 SIN(0 2 1)
V8 8 0 SIN(0 1 2)
V9 9 0 SIN(0 2 4)
R7 7 10 1
R8 8 10 1
R9 9 10 1
R10 10 0 1

.FFT V(10) NP=16 WINDOW=HANN FREQ=4

.MEASURE FFT SFDR_BINSIZDEFAULT SFDR V(10) MINFREQ=2
.MEASURE FFT SFDR_BINSIZ0 SFDR V(10) BINSIZ=0 MINFREQ=2
.MEASURE FFT SFDR_BINSIZ1 SFDR V(10) BINSIZ=1 MINFREQ=2
.MEASURE FFT SFDR_BINSIZ2 SFDR V(10) BINSIZ=2 MINFREQ=2

.MEASURE FFT SNDR_BINSIZDEFAULT SNDR V(10)
.MEASURE FFT SNDR_BINSIZ0 SNDR V(10) BINSIZ=0
.MEASURE FFT SNDR_BINSIZ1 SNDR V(10) BINSIZ=1
.MEASURE FFT SNDR_BINSIZ2 SNDR V(10) BINSIZ=2

.MEASURE FFT ENOB_BINSIZDEFAULT ENOB V(10)
.MEASURE FFT ENOB_BINSIZ0 ENOB V(10) BINSIZ=0
.MEASURE FFT ENOB_BINSIZ1 ENOB V(10) BINSIZ=1
.MEASURE FFT ENOB_BINSIZ2 ENOB V(10) BINSIZ=2

.PRINT TRAN  V(10)
.END
