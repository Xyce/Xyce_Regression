Testing the use of .param in objective functions

.DC V1 1 1 1
.param res=1
V1 1 0 1
R1 1 2 1
R2 2 0 0.5

.print sens
.SENS objfunc={res*I(V1)} param=R1:R

.end
