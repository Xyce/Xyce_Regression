HB test of print output format
*
* Because we use VP and IP here, it is pretty essential that there be nontrivial
* power in frequencies other than the fundamental -- using a sinusoidal
* input source and only linear devices would have what is essentially
* roundoff error in all frequencies other than the fundamental.   This
* leads to platform-dependent failure when comparing the VP signal.
*
* Thus, we're driving this with a roughly square wave and making the 
* circuit slightly non-linear.
* 
*

R1 1 0 1k
C1 1 0 1p
D1 2 1 D1N3940
.MODEL D1N3940 D (IS=4e-10 RS=.105 N=1.48 TT=8e-7 CJO=1.95E-11 VJ=.4 M=.38 EG=1.36 XTI=-8 KF=0 AF=1 FC=.9 BV=600 IBV=1e-4)
*            low high td tr  tf  pulsewidth    period
v1 2 0 pulse 1V 2V  0 1e-5 1e-5 {1/1e4/2-1e-5 } {1/1e4}

.hb 1e4

* The .PRINT HB FILE=hbfile line should produce the output file hbfile.HB.FD.prn, after the fix
* for SON Bug 701.
.print HB file=hbfile vr(1) {vr(1)} vi(1) {vi(1)} vm(1) {vm(1)} vp(1) {vp(1)} vdb(1) {vdb(1)} ir(v1) {ir(v1)} ii(v1) {ii(v1)} im(v1) {im(v1)} ip(v1) {ip(v1)} idb(v1) {idb(v1)}

* An attempt to overwrite the netlist with an explicit .PRINT HB_TD line
* should produce the file printFilename.cir.HB.TD.prn
.print HB_TD file=printFilename.cir vr(1) {vr(1)} vi(1) {vi(1)} vm(1) {vm(1)} vp(1) {vp(1)} vdb(1) {vdb(1)} ir(v1) {ir(v1)} ii(v1) {ii(v1)} im(v1) {im(v1)} ip(v1) {ip(v1)} idb(v1) {idb(v1)}

* An attempt to write to a file that ends in .cir with an explicit
* .PRINT HB_IC line should produce the file hbfileic.cir.hb_ic.prn
.print HB_IC file=hbfileic.cir vr(1) {vr(1)} vi(1) {vi(1)} vm(1) {vm(1)} vp(1) {vp(1)} vdb(1) {vdb(1)} ir(v1) {ir(v1)} ii(v1) {ii(v1)} im(v1) {im(v1)} ip(v1) {ip(v1)} idb(v1) {idb(v1)}

.options hbint numfreq=50

* Output vp() and ip() in degrees
.OPTIONS OUTPUT PHASE_OUTPUT_RADIANS=true

.end
