* Transient sensitivity example, pulse source, analytical version
.param cap=0.1u
.param res=1K

c1 1 0 cap
c2 2 0 cap
R1 1 3 res
R2 1 2 res

Vin 3 0 PULSE(0V 1V 0S 10US 10US 100US 220US)

* Transient commands
.tran 0 1.5ms 
.options timeint reltol=1e-6 abstol=1e-6

.print tran v(1) v(2) v(3)

* Sensitivity commands
.print sens 
.SENS objfunc={V(2)} param=Vin:v1,Vin:v2,Vin:td,Vin:tr,Vin:tf,Vin:pw,Vin:per
.options SENSITIVITY direct=1 adjoint=0  forceanalytic=true
.end

