Static Latch
*
* ERK.  4/16/2021.  This circuit runs fine with embedded sampling, but fails with PCE.
*
* It previous seg faulted, but I added an error trap to the Xyce source to prevent that.   
* It segfaulted when it attempted to do gmin stepping after straight Newton failed.
* There are one or more functions in the PCEBuilder that need to be implemented to 
* properly support GMIN stepping.
*
***   resistors
rcc2 6 8 3.33k
ree2 9 0 200
***   transistors
q1 6 8 4 npn1
q2 8 4 9 npn1
***   models
.model npn1 npn(
+ bf={agauss(50,20,1)}
+ br=0.2 rb=81 rc=100 re=6.1 
+ cjs={agauss(0.3pf,0.03pf,1)}
+ tf=0.36ns
+tr=10ns 
+ cje={agauss(0.13pf, 0.013pf, 1)}
+ cjc={agauss(0.1pf,0.01pf,1)}
+ is=1e-16 ne=1 nc=1.082 vje=0.84v
+vjc=1.1v mje=0.36 mjc=0.76 vaf=50v eg=1.1)
***   sources
vcc 6 0 5v
vref 3 0 2.5v
vrset 1 0 pulse(0v 3v 1ns 1ns 1ns 10ns 40ns)
vset 7 0 pulse(0v 3v 20ns 1ns 1ns 10ns 40ns)
***   subcircuits
.subckt eclg2 1 2 3 4 5 6
**  resistors
rs 6 11 619
rc2 11 10 900
re4 12 0 200
re6 5 0 6k
**  transistors
q1 9 1 8 npn1
q2 9 2 8 npn1
q3 11 3 8 npn1
q4 8 4 12 npn1
q5 10 10 9 npn1
q6 6 9 5 npn1
.ends eclg2
x1 1 2 3 4 5 6 eclg2
x2 5 7 3 4 2 6 eclg2
***   control cards
*.tran 1ns 75ns
.tran 1ns 40ns
.print tran v(1) v(7) v(5) v(2)

.PCE
+ useExpr=true

.options PCES outputs={v(5)},{v(2)} 
+ projection_pce=true
* As the number of samples will be small, don't output the mean, variance, std dev from the original samples.
* Just output the PCE statistics:
+ sparse_grid=true

.options device debuglevel=-100

.end
