Basic function test of delay device
VIN 1 0 PULSE(0 5 0 10N 10N 20N 40N)
R0 1 0 1

VIN_delayed 4 0 PULSE(0 5 .1N 10N 10N 20N 40N)
R2 4 0 1

YDELAY delay1 2 0 1 0 TD=.1N
R1 2 0 1

.TRAN 0.25N 50N
*comp {V(4)-V(2)} offset=1e-14
.PRINT TRAN V(1) V(2) V(4) {V(4)-V(2)}
*.PRINT TRAN V(1) V(2)
.END
