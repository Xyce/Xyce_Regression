Netlist to Test out the period "." separator for device instance parameters
*
* this netlist must be run with either -hspice-ext all, or -hspice-ext separator
*
R1 1 0 1K 
V1 1 0 5V
.DC V1 1V 1V 1V
.PRINT DC V(1) R1.R  {R1.R}
.END
