*****************************************************************
* This netlist tests the -noise_names_file command line option.
*
* This netlist should produce entries in that file for all of
* the R, Q and M devices in the netlist.  There should be no
* entries for the V, L or C devices, since they don't have
* noise sources.  
* 
* The BSIMCMG device (M1) was chosen because it has duplicate
* noise source names.  So, the test verifies that each of
* those duplicate entries only appears once in the noise 
* names file.
*
* The EKV MOSFET has some bad characters, like ( and ), in the
* noise type string in the source code auto-generated by the ADMS 
* parser.  So, this tests that those characters are removed in 
* the noise type name that output by -noise_names_file
*****************************************************************

* BJT noise test circuit
V2 N001 0 15
V1 N003 0 0 AC 1
Q1 N002 N005 N006 0 2N2222
R3 N001 N002 1K
R5 N006 0 100
R1 N001 N005 75K
R2 N005 0 10K
C1 N005 N004 .1u
C2 N006 0 10u
R4 OUT 0 100K
C3 OUT N002 1u
R6 N004 N003 1K

.model 2N2222 NPN(IS=1E-14 VAF=100
+   BF=200 IKF=0.3 XTB=1.5 BR=3
+   CJC=8E-12 CJE=25E-12 TR=100E-9 TF=400E-12
+   ITF=1 VTF=2 XTF=3 RB=10 RC=.3 RE=.2  KF=5.0E-16  AF=1.0
+ )

********************************************
* BSIMCMG has duplicate noise-source names
********************************************
.include "modelcard.nmos_xyce"
vds 1 0 dc 1v
vgs gate 0 dc 0.5v ac 1
vbs bulk 0 dc 0v

lbias 1 drain 1m
cload drain 2 1m
rload 2 0 1
M1 drain gate 0 bulk nmos1 TFIN=15n L=30n NFIN=10 NRS=1 NRD=1

**************************************************
* EKV has "bad characters" in its noise type name
* autogenerated by the ADMS parser.  See SON Bug
* 926 for more details.
**************************************************
.include "150nm.mod"
M2 D G S B NMOS150 W=150e-9 L=150e-9  NF=1

Vg G Ga DC .5v AC 1
Vgprobe 0 Ga 0
Vd 1 Da DC 1v
Ldrain 1 D 1m
Cdrain D 0 1m
*Rdrain 2 0 1
Vdprobe 0 Da 0
Vs S Sa DC 0v
Vsprobe 0 Sa 0
Vb B Ba DC 0v
Vbprobe 0 Ba 0

.noise V(out) V1 dec 10 1e3 1e5 1
.PRINT NOISE ONOISE INOISE 
 
.end

