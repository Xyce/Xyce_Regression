
V1   1   0   1
r   1   2   {rval}
r2  2   3   {rval2}

* Select low, nom, or high for the library.  The values of V(2) and V(3)are:
*       V(2)   V(3)
* low   0.9   0.7
* nom   0.85  0.55
* high  0.8   0.4

.lib exclude
.erroneous dot line to be excluded in pass one
erroneous device to be excluded in pass two
.endl exclude

.lib rvals.lib nom

.tran 1ps 1ns
.print tran V(2) V(3)

.end
