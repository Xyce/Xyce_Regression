LOAD TEST CIRCUIT
*
V1 3 0 -15
V2 2 0 15
V3 4 0 10
R2 15 8 63.4K
R3 4 7 3.65K
R4 7 11 2.53K
R5 11 0 3.83K
Q1 15 7 9 QN2222
R6 9 8 26.7K
Q2 15 11 5 QN2222
R7 5 8 8.66K
R8 8 6 8.45K
R9 6 0 1K
V4 13 0 
R10 13 16 10K
R11 16 0 2.53K
D2 16 15 DN4148
R12 12 15 100K
D3 13 12 DN4148
X1 15 4 8 3 2 UA741
.DC V4 5 55 .05
.PRINT DC  V(13) V(6) V(8) 

*V(6)=VOUT V(13)=VIN V(8)=ILIMIT
*
************************************
* SUBCIRCUIT AND MODEL DEFINITIONS *
************************************
*
.MODEL QN2222 NPN (IS=15.2F NF=1 BF=105 VAF=98.5 IKF=.5
+ ISE=8.2P NE=2 BR=4 NR=1 VAR=20 IKR=.225 RE=.373 RB=1.49
+ RC=.149 XTB=1.5 CJE=35.5P CJC=12.2P TF=500P TR=85N)
*
.MODEL DN4148 D(RS=.8 CJO=4PF IS=7E-09 N=2 VJ=.6V    
+ TT=6E-09 M=.45 BV=100V)
*
.SUBCKT UA741 2    3  6   7   4
*             - IN + OUT VCC VEE
RP 4 7 10K
RXX 4 0 10MEG
*
IBP 3 0 80NA
RIP 3 0 10MEG
CIP 3 0 1.4PF
IBN 2 0 100NA
RIN 2 0 10MEG
CIN 2 0 1.4PF
VOFST 2 10 1MV
RID 10 3 200K
EA 11 0 10 3 1
R1 11 12 5K
R2 12 13 50K
C1 12 0 13PF
GA 0 14 0 13 2700
C2 13 14 2.7PF
RO 14 0 75
L 14 6 30UHY
RL 14 6 1000
CL 6 0 3PF
.ENDS UA741

.END 

