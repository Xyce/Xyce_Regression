* 51 stage Ring-Osc.

vin in out 2 pulse 2 0 0.1n 5n 1 1 1
*vdd dd 0 dc 0 pulse 0 2 0 1n 1 1 1
vdd dd 0 2
vss ss 0 dc 0
ve  sub  0 dc 0

xinv1 dd ss sub in out25 inv25
xinv2 dd ss sub out25 out50 inv25
xinv5 dd ss sub out50 out inv1
xinv11 dd ss sub out buf inv1
cout  buf ss 1pF

xdum ss dum

.tran 0.2n 1n
*.print tran format=tecplot V(in) V(out)
.print tran V(in) V(out)

************************************
* **** Start Homotopy Setup ****
************************************
.options nonlin nlstrategy=0 searchmethod=0
+ maxstep=50 maxsearchstep=20 continuation=1

.options loca stepper=0 stepcontrol=1
+ conparam=vdd
+ initialvalue=0.0 minvalue=-1.0 maxvalue=2.0
+ initialstepsize=0.05 minstepsize=0.01 maxstepsize=2.0 aggressiveness=1.0
+ maxsteps=5000 maxnliters=200
**********************************
* **** End Homotopy Setup ****
**********************************

.options device debuglevel=-10
.options timeint debuglevel=-10
.options linsol type=aztecoo AZ_kspace=100

.include nmos_3_2.mod
.include pmos_3_2.mod
.include lib.h
.end


