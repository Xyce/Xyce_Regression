* Transient sensitivity example, sine source, finite difference
.param cap=0.1u
.param res=1K

.param v0=0
.param va=1
.param f=100k 
.param td=-2.5u
.param theta=0.0
.param phase=-90.0

c1 1 0 cap
c2 2 0 cap
R1 1 3 res
R2 1 2 res

Vin 3 0 SIN({V0} {VA} {F} {TD} {THETA} {PHASE} )

* Transient commands
.tran 0 10us uic
.options timeint reltol=1e-6 abstol=1e-6

.print tran v(1) v(2) v(3)

* Sensitivity commands
.print sens
.SENS objfunc={V(2)} param=v0,va,f,td,theta,phase

.options SENSITIVITY direct=1 adjoint=0 forcefd=true
.end

