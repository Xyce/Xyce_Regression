4049 Circuit

X2 3 8 2 0 CD4049UB
V1 2 0 5
C1 8 5 1.088N
R1 3 5 46.5K
R2 1 5 98.6K
X1 1 3 2 0 CD4049UB

*
* NOOP used to forego the operating point
* This circuit does not perform as an oscillator if an operating point
* calculation is done --- the transient solution simply has to start from
* an all-0 initial condition.
*
.tran .05U 500U NOOP

* Xyce option needed when default is changed to 1 (Backward Euler).
* Also serves as useful test of non-default method.

*.options timeint method=2 abstol=1.0e-7 reltol=1.0e-6
.options timeint method=7 newlte=1 reltol=0.5e-3 
*.options timeint method=7 erroption=1 delmax=4e-7 

* speed comparison for above different options:
* with trap and erroption=1, 1255 steps
* with trap and new LTE, 419 steps 

*COMP V(8) reltol=0.02
.print tran precision=10 width=19 {V(8)+4} {v(5)+4} {V(1)+4} {V(3)+4}

* Subcircuit and Model Definitions
.SUBCKT CD4049UB 1  2   3   4
*HEX BUFFER    IN OUT VCC VSS
M1 2 1 3 3 CD4049P
M2 2 1 4 4 CD4049N
.MODEL CD4049P PMOS (LEVEL=1 VTO=-2.9 KP=2M GAMMA=3.97U
+ PHI=.75 LAMBDA=1.87M RD=28.2 RS=45.2 IS=31.2F PB=.8 MJ=.46
+ CBD=148P CBS=177P CGSO=218N CGDO=182N CGBO=299N)
.MODEL CD4049N NMOS (LEVEL=1 VTO=2.1 KP=5M GAMMA=3.97U
+ PHI=.75 LAMBDA=1.87M RD=4.2 RS=4.2 IS=31.2F PB=.8 MJ=.46
+ CBD=105P CBS=127P CGSO=156N CGDO=130N CGBO=214N)
.ENDS

.END

