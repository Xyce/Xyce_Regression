* Xyce netlist, with two identical Resistor-Diode-Resistor circuits

.OPTIONS DEVICE TNOM=25 TEMP=25

*Analysis directives and print statement
.TRAN  0.1ms 1ms
.PRINT TRAN FORMAT=PROBE V(N01192) V(N011460) V(N07223)
+ V(N07602) V(N075620) V(N07662)

R1         N01192 N011460  R=1000
V1         N01192 0  SIN(0 1 1KHz 0 0 0)
R2         N07223 0  R=1k
D1         N011460 N07223 D1N3940

R3         N07602 N075620  R=1000
R4         N07662 0  R=1k
D2         N075620 N07662 D1N3940
V2         N07602 0 SIN(0 1 1KHz 0 0 0)

* Diode model from the Diode Clipper example in the
* Xyce Users' Guide
.MODEL D1N3940 D(
+ LEVEL=2
+ IS = 4E-10
+ RS = .105
+ N = 1.48
+ TT = 8E-7
+ CJO = 1.95E-11
+ VJ = .4
+ M = .38
+ EG = 1.36
+ XTI = -8
+ KF = 0
+ AF = 1
+ FC = .9
+ BV = 600
+ IBV = 1E-4)

.END
