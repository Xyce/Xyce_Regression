* Test AC mode support for the FIND-WHEN and WHEN measures.
* To be conservative, there are subtests for each
* valid operator (V, VR, VI, VP, VM and VDB) for
* each measure type.
*
* See SON Bug 1270 for more details.
*****************************************************

* trivial high-pass filter (V-C-R) circuit

R2 c 0 1
R1 b c 1
C1 a b 1u
V1 a 0 DC 0V AC 1

.print AC vr(b) vi(b) vm(b) vp(b) vdb(b)
+ vr(b) vi(b) vm(b) vp(b) vdb(b)
.ac dec 5 100Hz 1e6

* WHEN
.MEASURE AC whenvmb0.5 WHEN vm(b)= 0.5
.MEASURE AC whenvrb0.5 WHEN vr(b)= 0.5
.MEASURE AC whenvib0.1 WHEN vi(b)= 0.1
.MEASURE AC whenvbp50 WHEN vp(b)= 50

* FIND-WHEN
.MEASURE AC findvmcwhenvmb0.5 find vm(c) when vm(b)= 0.5
.MEASURE AC findvrcwhenvrb0.5 find vr(c) when vr(b)= 0.5
.MEASURE AC findvicwhenvib0.1 find vi(c) when vi(b)= 0.1
.MEASURE AC findvpcwhenvpb50 find vp(c) when vp(b)= 50.0

.END
