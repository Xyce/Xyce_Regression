CMOS INVERTER  - test of .FOUR with transient sensitivities
*
M1 2 1 0 0 NMOS W = 20U L = 5U
M2 2 1 3 3 PMOS W = 40U L = 5U
VDD 3 0 5
VIN 1 0 SIN 2.5 2.5 20MEG
.MODEL NMOS NMOS LEVEL = 3 CGDO = .2N CGSO = .2N CGBO = 2N
.MODEL PMOS PMOS LEVEL = 3 CGDO = .2N CGSO = .2N CGBO = 2N

.sens objfunc={V(2)}  param=M1:L,M2:L
.print sens
.options sensitivity direct=1 adjoint=0

.TRAN 1N 100N

.FOUR 20MEG V(2) V(1) V(3)
.FOUR 40MEG V(3) V(2)
*
* do every sensitivity, along with a (redundant) signal.  Check the redudant ones match.
.FOUR 20MEG v(3) sens 
.FOUR 40MEG v(2) sens

.PRINT TRAN V(2) V(1)
.END
