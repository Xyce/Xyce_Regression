TEST OF A 1-BIT ADDER WITH SWITCHES
*
* Will add comments to this netlist at a later time. Regina Schells 6/1
*
* MAIN CIRCUIT 
* 
X1 1 2 3 9 13 99 ONEBIT
RINA 1 0 1K
RINB 2 0 1K
RCIN 3 0 1K
RBIT0 9 0 1K
RCOUT 13 0 1K
VCC 99 0 5
VINA 1 0 PULSE(0 3 0 10N 10N 10N 50N)
VINB 2 0 PULSE(0 3 0 10N 10N 20N 100N)
VCIN 3 0 PULSE(0 3 100N 10N 10N 100N 200N)
.TRAN 0.5N 200N
.PRINT TRAN V(1) V(2) V(3) V(9) V(13)
.OPTIONS TIMEINT ABSTOL=1.0E-3 RELTOL=1.0E-3
*
.MODEL SW VSWITCH (RON=1 ROFF=1MEG VON=2.51 VOFF=2.5)
*
.SUBCKT ONEBIT 1 2 3 4 5 6
* TERMINALS: A B CIN OUT COUT VCC
X1 1 2 7 6 XOR
X2 1 2 8 6 AND
X3 7 3 4 6 XOR
X4 3 7 9 6 AND
X5 8 9 5 6 OR
*
.SUBCKT OR 1 2 3 4
* TERMINALS A B OUT VCC
RL 3 0 1K
S1 3 4 1 0 SW
S2 3 4 2 0 SW
.ENDS OR
*
.SUBCKT AND 1 2 3 4
* TERMINALS A B OUT VCC
RL 3 0 1K
S1 4 5 1 0 SW
S2 5 3 2 0 SW
.ENDS AND
*
.SUBCKT XOR 1 2 3 4
* TERMINALS A B OUT VCC
RL 3 0 1K
S1 4 3 1 2 SW
S2 4 3 2 1 SW
.ENDS XOR
*
.ENDS ONEBIT
*
.END   
