* **********************************************************
* Test non-default value (0) for .OPTIONS FFT FFT_ACCURATE,
* which then uses interpolation to get the waveform values
* at the requested sample times.  Also test that the WINDOW
* qualifier defaults to RECT.
*
************************************************************
.TRAN 0 1
.OPTIONS FFT FFT_ACCURATE=0 FFTOUT=1

V1 1 0 SIN(0 500 1)
V3 3 0 SIN(0 200 2)
R1 1 2 1
R2 2 0 1
R3 3 2 1

.FFT V(2) NP=8 WINDOW=HANN FORMAT=UNORM
.PRINT TRAN V(1) V(2) V(3)

.END
