* Test to make sure that the "override" type of raw file 
* does not include adjoint information, as it is not supported.
*
* The correct behavior is for this circuit to run successfully via :
*
*     Xyce -r xyce.raw
*
* The resulting file, xyce.raw should be identical to the raw file 
* produced by an equivalent netlist that lacks .SENS commands.
*

V1 1 0 PWL 0 0 1 1
R1 1 2 1
R2 2 0 1
M1 2 1 0 0 PMOS
.model PMOS PMOS (W=1.5u L=1u)

.TRAN 0 1

.OPTIONS OUTPUT initial_interval=0.1 

.options timeint breakpoints=0.25,0.5,0.75

.PRINT TRAN R1:R R2:R V(1) V(2)

.end

