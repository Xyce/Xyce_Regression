A neuron cable example
*
* A copy of the rallpack1 test, modified to use a user-defined equation 
* to specify the leak current rather than using the passive membrane model
*


.param length = 0.1e-2 ; [m]
.param radius = 0.5e-6  ; [m]
.param memC = 1.0e-2  ; [F/m^2] ok
.param restV = -0.065 ; [V]
.param Rm = 4.0 ; [ohms m^2]
.param memG = {1.0/Rm}    
.param Ra = 1.0 ; [ohms m]


.model pcParams neuron level=6 
+ ionchannelmodel = UD 
+ indvars = { {Ipas} }
+ indfequs = { { memG * (V -  restV) } }
+ indqequs = { {0} }
+ cMem = {memC}
+ gMem = {memG}
+ vRest = {restV}

*
* Using the above neuron model
*

* This is a standard current pulse to start an activation
*          pulse( initial_value pulse_value delay_time rise_time fall_time pulse_width period)
Iin 0 a PULSE( 0 1.0e-10 1.0e-12 0.0 0.0 1.0e10 1.0e10)

* the parameters R (intra-cellular resistivity Ohm/cm), A= radius (cm), L = length (cm)
* can be specified in the .model statement or as part of the instance.  Instance level
* parameters override model level ones.  N = number of segments.

* intra cellular resistivity, rl,  is typically 1-3 kOhm mm.  Resistance along the long axis (longitudinal resistance Rl = rl L / (pi a^2)
* 1 kOhm mm = 1000 Ohm mm = 100 Ohm cm 

yneuron neuron1  a b pcParams 
* R=1.0e2 A=1.0e-4 L=0.4 
+ R = {Ra}
+ A = {radius}
+ L = {length}
+ N = 1000

.tran 0 0.25

.options output initial_interval=5.0e-5
.options timeint method=7 newlte=1 newbpstepping=1 reltol=1e-3
.print tran 
*+ i(iin) 
+ V(a) 
*+ n(y%neuron%neuron1_V1) 
+ V(b)



.end


