*Sample netlist for BSIM6
*Inverter Transient

.options timeint method=gear debuglevel=-100
.options device temp=25 debuglevel=-100

*.hdl "bsim6.va"
.include "modelcard_xyce.nmos"
.include "modelcard_xyce.pmos"

* --- Voltage Sources ---
vdd   supply  0 dc 1.0
VIN1 vi 0 PWL(0S 0V  7.0e-8 0V 0.1us 1.0V )

* --- Inverter Subcircuit ---
.subckt inverter vin vout vdd gnd
Mp1 vout vin vdd gnd pmos W=10u L=10u 
Mn1 vout vin gnd gnd nmos W=10u L=10u 
.ends

* --- Inverter ---
Xinv1  vi vo supply 0 inverter

* --- Transient Analysis ---
.tran 2ns 1us

.print tran v(vi) v(vo) {ddt(v(vo))} 

.SENS objfunc={V(VO)}
+ param=
+ XINV1:MP1:W,
+ XINV1:MP1:L,
+ XINV1:MN1:W,
+ XINV1:MN1:L

.options SENSITIVITY STDOUTPUT=1 DIAGNOSTICFILE=0 adjoint=0 direct=1  
.print sens 

.end

