TRAN test of print output format
*
* Trivial resistor circuit, just do a transient and watch the output
*

R1 1 0 10
V1 1 0 sin (0 1 1 0 0)

.OPTIONS OUTPUT INITIAL_INTERVAL=0.01

.print TRAN FORMAT=NOINDEX v(1) I(v1)
.tran 0 1

.end
