* Xyce netlist for testing Spectre V-Sources.  Note that
* the device "names" in the Spectre netlist are (for example)
* R5 and V5.  However, the Spectre instance lines are of the 
* form:
*
*   R5 (net3 V6) resistor r=1K
*   V5 (net3 0) vsource dc=1 type=dc
*
* So, on a Spectre instance line, it is the "resistor" and "vsource" 
* keywords that identify the devices as Resistors or Voltage Sources.
* So, the xdm translation will turn those devices into RR5 and VV5 
* in the translated Xyce netlist.  For this reason, the device names 
* in this "Gold" Xyce netlist are (for example) RR5 and VV5, to match
* what the device names will be in the xdm-translated Xyce netlist.

*Analysis directives: 
.TRAN  0 1ms 0
.PRINT TRAN V(V2) V(V4) V(V6) V(V8) V(V10) V(V12)

**********************************************************
*AC Source syntaxes
**********************************************************
* SIN source, no DC offset.  1V amplitude.  Freq. of 1KHz
RR1        net7 V2  1k 
RR2        0 V2 2K 
VV1        net7 0 SIN(0 1 1KHz 0 0 0)

* SIN source, With DC Offset of 1V
RR9        net9 V10  1k 
RR10       0 V10 2K 
VV9        net9 0 SIN(1 1 1KHz 0 0 0)

* Pulse source.  Xyce parameters within pulse( ) spec are:
* V1 (initial value), V2 (pulse value), TD (delay time),
* TR (rise time), TF (fall time), PW (pulse width) and PER (period)
VV11 net11 0 pulse(1 10 50e-6 50e-6 70e-6 200e-6 400e-6) 
RR12 V12 0 R=1K
RR11 net11 V12 R=1K

* Exp source.  Xyce parameters within exp() spec are:
* V1 (initial amplitude), V2 (amplitude), TD1 (rise delay time),
* TAU1 (rise time constant), TD2 (fall delay time) and
* TAU2 (fall time constant)
RR7        net1 V8  1k 
RR8        0 V8   2K 
VV7        net1 0  exp(0 1 100e-6 20e-6 600e-6 40e-6)

****************************************************
* DC source syntaxes
****************************************************
RR3        net5 V4  1k 
RR4        0 V4 2K 
VV3        net5 0  5

RR5        net3 V6  1k 
RR6        0 V6 2K 
VV5        net3 0  1

.END

