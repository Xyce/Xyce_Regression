* Transient sensitivity example, PWL source, analytical version, device-level specification
.param cap=1u
.param res=1K

c1 1 0 cap
c2 2 0 cap
R1 1 3 res
R2 1 2 res

Vin 3 0 PWL(0 0 1ms 1 2ms -1 3ms -0.5 4ms 0.25 5ms 0.75 6ms 0.0  )

* Transient commands
.tran 0 10ms 
.options timeint reltol=1e-6 abstol=1e-6

.print tran v(2)

* Sensitivity commands
.print sens 
.sens objfunc={v(2)} sensdevicename=vin
.options sensitivity direct=1 adjoint=0
.end

