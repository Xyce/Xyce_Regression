Test circuit for AC output through expressions

* It is important to have a signal with significant harmonics throught
* the HB spectrum.  Using a sin source here leads to most solution magnitudes
* being *very* small (roundoff error) and therefore the phase is effectively
* a random number, leading to cross-platform compare failures.  
* Using a PULSE source instead makes the phase meaningful.
* Here, the period is 1e-4, and the PW parameter is half of that minus the
* rise and fall times
*             TL TH TD TR TF PW          PER
v1 a 0 PULSE( 1V 5V 0  5n 5n {.5e-4-10n} 1e-4) AC 1
R1 a b 1
R2 b 0 2
C1 a b 1u

* Output vp() in degrees
.OPTIONS OUTPUT PHASE_OUTPUT_RADIANS=true

.hb 1e4
.print hb V(A) V(B) V(A,B) VR(A,B) VI(A,B) VM(A,B) VDB(A,B) VP(A,B)
.end
