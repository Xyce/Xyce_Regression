* This .LIN analysis was used to generate the input files for
* the ylin-5port-yparam.cir test.  However, it is not run as
* part of any regression test.

* RC ladder circuit
* Note that all ports (P devices) must use a common
* Reference Node, which is 0 here.
P1 2   0  port=1  z0=50
P2 5   0  port=2  z0=50
P3 6   0  port=3  Z0=50
P4 7   0  port=4  Z0=50
P5 12  0  port=5  Z0=50

C1 2 0 1e-2
Rgs 1 2 0.02

.subckt RCBlock IN OUT GND
R1 IN OUT 20
C1 IN OUT 1p
Cg1 OUT GND 1p
.ends

X1 2 3 0 RCBlock
X2 3 4 0 RCBlock
X3 4 5 0 RCBlock
X4 5 6 0 RCBlock
X5 6 7 0 RCBlock
X6 7 8 0 RCBlock
X7 8 9 0 RCBlock
X8 9 10 0 RCBlock
X9 10 11 0 RCBlock
X10 11 12 0 RCBlock

.AC LIN 11 0 10e4
.LIN LINTYPE=Y FILE=ylin-5port-yparam.cir.y5p format=touchstone2 precision=12
.LIN LINTYPE=Y FILE=ylin-5port-yparam.cir-ts1.y5p format=touchstone precision=12

.END
