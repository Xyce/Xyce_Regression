* Sensitivity of collector current to amplifier component
* This circuit was found  on page 298 of the book, 
* "PSPICE and MATLAB for Electronics: An Integrated Approach" by John Okyere Attia.  
*
* The relevant pages are excerpted in google books, and includes a printout of the 
* PSPICE output.
*

.global_param VCCvalue=10V
.global_param Mval=6


VCC 4 0 DC {VCCvalue}
RB1 4 1 40k
RB2 1 0 10k
RE 2 0 1K
RC 5 3 6K
VM 4 5 DC 0; monitor collector current
XQ1 3 1 2 npnSub m={Mval}

.subckt npnSub A B C 
Q1 A B C Q2N2222 
.ends

.model Q2N2222 NPN(BF=100 IS=3.295e-14 VA=200)

.DC VCCvalue 1 10 0.2
.print dc v(4) I(VM)
.print sens v(4)

.SENS param=RB1:R,RB2:R,RE:R,RC:R,VM:DCV0,
+ Q2N2222:bf,
+ Q2N2222:is,
+ Q2N2222:nf,
+ Q2N2222:tnom,
+ Q2N2222:vaf
+objfunc={I(VM)} 

.options SENSITIVITY direct=1 adjoint=0  difference=forward  diagnosticfile=0 STDOUTPUT=0 debuglevel=-100 REUSEFACTORS=0

