*****************************************************************
* A test of .OPTIONS MEASURE MEASFAIL for successful measures.
* This tests .OPTIONS MEASURE MEASFAIL=1 for successful measures.
*
* See gitlab issue 221 for more details.
*****************************************************************

VS1  1  0  SIN(0 1.0 1KHZ 0 0.9)
VS2  2  0  SIN(0 -1.0 1KHz 0 0.9)
R1  1  0  100
R2  2  0  100

.OPTIONS MEASURE MEASFAIL=1

.TRAN 0  1ms
.PRINT TRAN FORMAT=NOINDEX V(1) V(2)

.measure tran avgVal avg V(1)

.measure tran derivValWhen deriv V(1) WHEN V(1)=0.5
.measure tran derivValAt deriv V(1) AT=5e-04

.measure tran dutyVal duty V(1)

.measure tran eqnVal EQN {V(1)+10}

.measure tran errorVal ERROR v(1) FILE=issue_221_comp_file.prn
+ COMP_FUNCTION=L1NORM INDEPVARCOL=1 DEPVARCOL=2

.measure tran whenVal WHEN V(1)=0.5
.measure tran findWhenVal FIND V(2) WHEN V(1)=0.5

.measure tran fourfail FOUR V(1) AT=1e6 TD=2e-3

.measure tran freqVal FREQ v(1) ON=0.75 OFF=0.25

.measure tran integVal integ V(1)

.measure tran maxVal max V(1)
.measure tran minVal min V(1)

.measure tran ppVal pp V(1)
.measure tran rmsVal rms V(1)

.measure tran trigTargVal TRIG v(1)=0.1 TARG v(1)=0.99

.END
