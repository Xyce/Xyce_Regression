* 51 stage Ring-Osc.

vin in out 2 pulse 2 0 0.1n 5n 1 1 1
vdd dd 0 2.0
*dc 0 pulse 0 2 0 1n 1 1 1
vss ss 0 dc 0
ve  sub  0 dc 0

xinv1 dd ss sub in out25 inv25 
xinv2 dd ss sub out25 out50 inv25
xinv5 dd ss sub out50 out inv1
xinv11 dd ss sub out buf inv1
cout  buf ss 1pF

xdum ss dum

.options timeint reltol=1e-4
*.option itl1=500 gmin=1e-15 itl4=10 
*.tran 0.2n 50n

*.tran 1n 10n
*COMP TIME zerotol=1e-14
*.print tran v(dd) v(in) v(out) 
.dc vin 0 2 0.5
.print dc v(dd) v(in) v(out) 
.options diagnostic 


*
* NMOS model
*
* bsimsoi3.2 model card
.model  n1 nmos  level = 10 
+mobmod  = 1    capmod  = 2    shmod   = 1 
+soimod  = 1    igcmod  = 0	igbmod  = 0
+dtoxcv  = 0   llc     = 0   lwc     = 0    lwlc    = 0
+wlc = 0          wwc = 0               wwlc    = 0  tsi = 9e-008 
+tox = 5e-009   toxref = 5e-009     tbox = 5e-007   tnom  = 25
+rbody = 1	rbsh = 0	rsh = 0    rhalo = 1e+015
+wint = 0	lint = 0	wth0 = 0	ll = 0
+wl = 0		lln  = 1	wln = 1		lw = 0
+ww = 0		lwn  = 1	wwn = 1		lwl = 0 
+wwl = 0	ln = 2e-006	xpart = 1	xj = 1e-007
+k1b = 0	k2b = 0		dk2b = 0	vbsa = 0.10         
+aigc = 1  bigc = 1  cigc = 1  aigsd = 1 
+bigsd = 1    cigsd = 1  nigc = 1   poxedge = 1  pigcd = 1 
+vth0 = 0.5	k1 = 0.1	k1w1 = 0 
+k1w2 = 0	k2 = 0		k3 = -2		k3b = 0             
+kb1 = 1	w0 = 0          nlx = 0                          
+nch = 8e+017	nsub = 5e+015        
+ngate = 2e+020 dvt0 = 1        dvt1 = 0.15	dvt2 = 0             
+dvt0w = 0	dvt1w  = 2000000 dvt2w = 0	eta0    = 0.5           
+etab    = 0               dsub    = 0.35            voff    = -0.15           nfactor = 0.4           
+cdsc    = 0.005           cdscb   = -0.01           cdscd   = 0               cit     = 0             
+u0 = 0.05	ua = 0		ub = 1.2e-018        uc      = 0             
+prwg = 0               prwb = 0               wr      = 1               rdsw    = 100           
+a0 = 0		ags = 0       a1      = 0               a2      = 0.99       
+b0      = 0               b1      = 0               vsat    = 80000           keta    = 0             
+ketas   = 0               dwg     = 0               dwb     = 0               dwbc    = 0             
+pclm    = 1               pdiblc1 = 0.15            pdiblc2 = 0               pdiblcb = 0             
+drout   = 0.4             pvag    = 0               delta   = 0.001           alpha0  = 8e-009        
+beta0   = 0               beta1   = 0               beta2   = 0.05            fbjtii  = 0             
+vdsatii0= 0.8             tii     = -0.2         lii     = 5e-008          esatii  = 1e+008        
+sii0    = 0.5             sii1    = 0               sii2    = 0               siid    = 0             
+agidl   = 2e-009          bgidl   = 2e+009          ngidl   = 0.5             ebg     = 1.2           
+vgb1    = 300             vgb2    = 17           
+voxh    = 5               deltavox= 0.005         
+ntox    = 1               ntun    = 3.6             ndiode  = 1               nrecf0  = 1.8           
+nrecr0  = 1               isbjt   = 3e-007          isdif   = 3e-008          isrec   = 0.0005        
+istun   = 1e-008          vrec0   = 0.05            vtun0   = 5               nbjt    = 1             
+lbjt0   = 2e-007          vabjt   = 10              aely    = 0               ahli    = 1e-015        
+vevb    = 0.075           vecb    = 0.026         
+cjswg  = 5e-010	mjswg = 0.5	pbswg = 0.8	tt = 5e-010        
+ldif0   = 0.001           cgeo    = 0               cgso    = 6.5e-010        cgdo    = 6e-010      
+dlc     = 0               dwc     = 0               dlcb    = 0               dlbg    = 0             
+fbody   = 1               clc     = 1e-007          cle     = 0.6             cf      = 0             
+csdmin  = 2.5e-005        asd     = 0.5             csdesw  = 0               vsdfb   = -0.8          
+vsdth   = -0.3            delvt   = 0               acde    = 0               moin    = 15            
+ckappa  = 0.6             cgdl    = 0               cgsl    = 0               ndif    = -1            
+rth0    = 0.09            cth0    = 1e-005    
+tpbswg = 0  
+tcjswg  = 0.0005
+kt1 = -0.2	kt1l = 8e-009          kt2 = -0.06         ute = -1.5        
+ua1 = 3e-010	ub1 = -3e-018      uc1 = -6.0e-011       prt = 10         
+at = 65000	ntrecf  = 0.1	ntrecr = -1              xbjt    = 1e-020      
+xdif    = 1.6             xrec    = 0.8             xtun    = 6
*+fnoimod = 1 tnoimod = 1   tnoia = 1  tnoib = 2.5   rnoia = 0.577 rnoib = 0.37
*+ntnoi = 1.0	em = 41000000  af = 1	ef = 1      kf = 0
*+noif = 1.0	
+rgateMod = 2 rshg = 0.1 xrcrg1 = 12 xrcrG2 = 1


*
* PMOS model
*
* bsimsoi3.2 model card
.model  p1 pmos  level = 10 
+mobmod  = 1    capmod  = 2    shmod   = 1 
+soimod  = 1    igcmod  = 0	igbmod  = 0
+dtoxcv  = 0	llc     = 0   lwc     = 0    lwlc    = 0
+wlc = 0	wwc = 0               wwlc    = 0  tsi = 9e-008 
+tox = 5e-009   toxref = 5e-009     tbox = 5e-007   tnom  = 25
+rbody = 1	rbsh = 0	rsh = 0    rhalo = 1e+015
+wint = 0	lint = 0	wth0 = 0	ll = 0
+wl = 0		lln  = 1	wln = 1		lw = 0
+ww = 0		lwn  = 1	wwn = 1		lwl = 0 
+wwl = 0	ln = 2e-006	xpart = 1	xj = 1e-007
+k1b = 0	k2b = 0		dk2b = 0	vbsa = 0.10         
+aigc = 1  bigc = 1  cigc = 1  aigsd = 1 
+bigsd = 1    cigsd = 1  nigc = 1   poxedge = 1  pigcd = 1 
+vth0 = -0.5	k1 = 0.1	k1w1 = 0 
+k1w2 = 0	k2 = 0		k3 = -2		k3b = 0             
+kb1 = 1	w0 = 0          nlx = 0           
+nch = 8e+017	nsub = 5e+015        
+ngate = 2e+020 dvt0 = 1        dvt1 = 0.15	dvt2 = 0             
+dvt0w = 0	dvt1w  = 2000000 dvt2w = 0	eta0    = 0.5           
+etab    = 0               dsub    = 0.35            voff    = -0.15           nfactor = 0.4           
+cdsc    = 0.005           cdscb   = -0.01           cdscd   = 0               cit     = 0             
+u0 = 0.05	ua = 0		ub = 1.2e-018        uc      = 0             
+prwg = 0               prwb = 0               wr      = 1               rdsw    = 100           
+a0 = 0		ags = 0       a1      = 0               a2      = 0.99       
+b0      = 0               b1      = 0               vsat    = 80000           keta    = 0             
+ketas   = 0               dwg     = 0               dwb     = 0               dwbc    = 0             
+pclm    = 1               pdiblc1 = 0.15            pdiblc2 = 0               pdiblcb = 0             
+drout   = 0.4             pvag    = 0               delta   = 0.001           alpha0  = 8e-009        
+beta0   = 0               beta1   = 0               beta2   = 0.05            fbjtii  = 0             
+vdsatii0= 0.8             tii     = -0.2         lii     = 5e-008          esatii  = 1e+008        
+sii0    = 0.5             sii1    = 0               sii2    = 0               siid    = 0             
+agidl   = 2e-009          bgidl   = 2e+009          ngidl   = 0.5             ebg     = 1.2           
+vgb1    = 300             vgb2    = 17           
+voxh    = 5               deltavox= 0.005         
+ntox    = 1               ntun    = 3.6             ndiode  = 1               nrecf0  = 1.8           
+nrecr0  = 1               isbjt   = 3e-007          isdif   = 3e-008          isrec   = 0.0005        
+istun   = 1e-008          vrec0   = 0.05            vtun0   = 5               nbjt    = 1             
+lbjt0   = 2e-007          vabjt   = 10              aely    = 0               ahli    = 1e-015        
+vevb    = 0.075           vecb    = 0.026         
+cjswg  = 5e-010	mjswg = 0.5	pbswg = 0.8	tt = 5e-010        
+ldif0   = 0.001           cgeo    = 0               cgso    = 6.5e-010        cgdo    = 6e-010      
+dlc     = 0               dwc     = 0               dlcb    = 0               dlbg    = 0             
+fbody   = 1               clc     = 1e-007          cle     = 0.6             cf      = 0             
+csdmin  = 2.5e-005        asd     = 0.5             csdesw  = 0               vsdfb   = -0.8          
+vsdth   = -0.3            delvt   = 0               acde    = 0               moin    = 15            
+ckappa  = 0.6             cgdl    = 0               cgsl    = 0               ndif    = -1            
+rth0    = 0.09            cth0    = 1e-005    
+tpbswg = 0  
+tcjswg  = 0.0005
+kt1 = -0.2	kt1l = 8e-009          kt2 = -0.06         ute = -1.5        
+ua1 = 3e-010	ub1 = -3e-018      uc1 = -6.0e-011       prt = 10         
+at = 65000	ntrecf  = 0.1	ntrecr = -1              xbjt    = 1e-020      
+xdif    = 1.6             xrec    = 0.8             xtun    = 6
*+fnoimod = 1 tnoimod = 1   tnoia = 1  tnoib = 2.5   rnoia = 0.577 rnoib = 0.37
*+ntnoi = 1.0	em = 41000000  af = 1	ef = 1      kf = 0
*+noif = 1.0	
+rgateMod = 2 rshg = 0.1 xrcrg1 = 12 xrcrG2 = 1

*
* subcircuits that build up gates
*

.subckt dum ss
mn1 ss ss ss ss ss n1 w=4u l=0.15u debug=1 AS=6p AD=6p PS=7u PD=7u
.ends dum

* XOR2
.subckt xnor2 dd ss sub A B out
mn1  T1  A   C1  sub  n1  w=4u  l=0.15u  AS=6p AD=6p PS=7u PD=7u
mn2  C1  B   ss  sub  n1  w=4u  l=0.15u   AS=6p AD=6p PS=7u PD=7u
mn3  out A   C2  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mn4  out B   C2  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mn5  C2  T1  ss  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mp1  T1  A   dd  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
mp2  T1  B   dd  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
mp3  out A   C3  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
mp4  C3  B   dd  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
mp5  out T1  dd  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
.ends xnor2

.subckt nor2 dd ss sub A B out
mn1  out A   ss  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mn2  out B   ss  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mp1  out A   C1  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
mp2  C1  B   dd  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
.ends nor2

.subckt nand2 dd ss sub A B out
mn1  out A   C1  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mn2  C1  B   ss  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mp1  out A   dd  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
mp2  out B   dd  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
.ends nand2

.subckt nor3 dd ss sub A B C out
mn1  out A   ss  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mn2  out B   ss  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mn3  out C   ss  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mp1  out A   C1  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
mp2  C1  B   C2  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
mp3  C2  C   dd  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
.ends nor3

.subckt nand3 dd ss sub A B C out
mn1  out A   C1  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mn2  C1  B   C2  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mn3  C2  C   ss  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mp1  out A   dd  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
mp2  out B   dd  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
mp3  out C   dd  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
.ends nand3

.subckt nor4 dd ss sub A B C D out
mn1  out A   ss  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mn2  out B   ss  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mn3  out C   ss  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mn4  out C   ss  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mp1  out A   C1  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
mp2  C1  B   C2  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
mp3  C2  C   C3  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
mp4  C3  C   dd  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
.ends nor4

.subckt nand4 dd ss sub A B C D out
mn1  out A   C1  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mn2  C1  B   C2  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mn3  C2  C   C3  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mn4  C3  C   ss  sub  n1  w=4u  l=0.15u AS=6p AD=6p PS=7u PD=7u
mp1  out A   dd  sub  p1  w=10u l=0.15u AS=15p AD=15p PS=13u PD=13u
mp2  out B   dd  sub  p1  w=10u l=0.15u AS=15p AD=15p PS=13u PD=13u
mp3  out C   dd  sub  p1  w=10u l=0.15u AS=15p AD=15p PS=13u PD=13u
mp4  out C   dd  sub  p1  w=10u l=0.15u AS=15p AD=15p PS=13u PD=13u
.ends nand4

.subckt inv1 dd ss sub in out
mn1  out in  ss  sub  n1  w=4u  l=0.15u  AS=6p AD=6p PS=7u PD=7u
mp1  out in  dd  sub  p1  w=10u l=0.15u  AS=15p AD=15p PS=13u PD=13u
.ends inv1

.subckt inv5 dd ss sub in out
xinv1 dd ss sub in 1 inv1
xinv2 dd ss sub 1  2 inv1
xinv3 dd ss sub 2  3 inv1
xinv4 dd ss sub 3  4 inv1
xinv5 dd ss sub 4 out inv1
.ends inv5

.subckt inv25 dd ss sub in out
xinv1 dd ss sub in 1 inv5
xinv2 dd ss sub 1  2 inv5
xinv3 dd ss sub 2  3 inv5
xinv4 dd ss sub 3  4 inv5
xinv5 dd ss sub 4 out inv5
.ends inv25

.subckt inv125 dd ss sub in out
xinv1 dd ss sub in 1 inv25
xinv2 dd ss sub 1  2 inv25
xinv3 dd ss sub 2  3 inv25
xinv4 dd ss sub 3  4 inv25
xinv5 dd ss sub 4 out inv25
.ends inv125

.subckt inv625 dd ss sub in out
xinv1 dd ss sub in 1 inv125
xinv2 dd ss sub 1  2 inv125
xinv3 dd ss sub 2  3 inv125
xinv4 dd ss sub 3  4 inv125
xinv5 dd ss sub 4 out inv125
.ends inv625


.end
