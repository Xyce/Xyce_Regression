A simple test case of a resistor with zero resistance

* test case when resistance is given a zero
V1 a 0 5V
R1 a b 0
R2 b 0 1K

.DC V1 0 5V 1V
.PRINT dc V(a) I(R1) I(R2)

.END
