Transmission Line Test Circuit
*
.OPTIONS TIMEINT ABSTOL=1e-04 RELTOL=1e-02 

* Slow pulse to drive 10K lump dual microstrip or simple transfer load
VSLOW 1 22 DC 0 EXP(0v 10v 3ms 10ms 200ms 10ms)
RS 1 11 50

* Enable xtstcir for 10K lump dual microstrip transmission line
* Or enable RT, RB, & RG for simple transfer load
xtstcir 11 22 33 44 microstrip
* RT 11 33 50
* RB 22 44 50
* RG 22 0 1u

* Terminator
RL 33 44 10K

**************************************************************
.subckt microstrip 1 2 3 4 
xcouple1 1 2 3 4 l3dsub1
.ends microstrip
***********************************
*** subcircuit: l3dsc1
*** Parasitic Model: microstrip
*** Only one segment
***
.subckt l3dsc1 1 3 2 4 
C01 1 0 4.540e-12
RG01 1 0 7.816e+03
L1 1 5 3.718e-08
R1 5 2 4.300e-01
C1 2 0 4.540e-12
RG1 2 0 7.816e+03
C02 3 0 4.540e-12
RG02 3 0 7.816e+03
L2 3 6 3.668e-08
R2 6 4 4.184e-01
C2 4 0 4.540e-12
RG2 4 0 7.816e+03
CM012 1 3 5.288e-13
KM12 L1 L2 2.229e-01
CM12 2 4 5.288e-13
.ends l3dsc1
***********************************
*** subcircuit: l3dsub1
*** Parasitic Model: microstrip
*** All segments
***
.subckt l3dsub1 1 2 41 42 
X1 1 2 3 4 l3dsc1
X2 3 4 5 6 l3dsc1
X3 5 6 7 8 l3dsc1
X4 7 8 9 10 l3dsc1
X5 9 10 11 12 l3dsc1
X6 11 12 13 14 l3dsc1
X7 13 14 15 16 l3dsc1
X8 15 16 17 18 l3dsc1
X9 17 18 19 20 l3dsc1
X10 19 20 21 22 l3dsc1
X11 21 22 23 24 l3dsc1
X12 23 24 25 26 l3dsc1
X13 25 26 27 28 l3dsc1
X14 27 28 29 30 l3dsc1
X15 29 30 31 32 l3dsc1
X16 31 32 33 34 l3dsc1
X17 33 34 35 36 l3dsc1
X18 35 36 37 38 l3dsc1
X19 37 38 39 40 l3dsc1
X20 39 40 41 42 l3dsc1
.ends l3dsub1

* Isolated High Speed Circuit
*
* High Speed source
* VFAST 8 0 DC 0 SIN(5v 10v 400MEGhz 1ms) NO CHANCE, Too expensive
*VFAST 8 0 DC 0 SIN(5v 10v 400Khz 1ms 0)
*VFAST 8 0 DC 0 SIN(5v 10v 4Khz 1ms 0)
*RFSS 8 9 0.5

* High Speed RLC load
*LFS  8 9 3n
*RFSP 9 0 1K
*CFS  9 0 680p

.tran 100us 300ms 

*COMP v(1) reltol=0.02 abstol=2e-6
*COMP v(11) reltol=0.02 abstol=1e-6
*COMP v(22) reltol=0.02 abstol=1e-6
*COMP v(33) reltol=0.02 abstol=1e-6
*COMP v(44) reltol=0.02 abstol=1e-6

.print  tran v(1) v(11) v(22) v(33) v(44)

.END
