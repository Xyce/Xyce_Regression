VBIC MODEL EXERCISER

**********  Solver Settings **********************************************************
.options device debuglevel=-1000 
.options timeint debuglevel=-1000 

********* Include Settings ************************************************************

*------------NPN Gummel curve generator-----------------*
VC       coll         0         0V
VB       basel        0         0V
RB       baseh        basel     1.0
VE       emit         0         0V
Qtest    coll        baseh     emit  dtn2   q2n2222B

rxth1 dtn1  0 1e9
rxth2 dtn2  0 1.0

* VBIC model 
.model q2n2222 npn
+ level=10 AFN=1 AJC=-0.5 AJE=-0.5 AJS=-0.5 ART=1000 
+ AVC1=0 AVC2=0 TAVC=0 BFN=1 CBCO=2.5e-14 CBEO=6e-14 CCSO=0 
+ CJC=3.63e-13 CJCP=0 CJE=1.07e-012 CJEP=0 CTH=5e-9
+ DEAR=-9.976E-005 DTEMP=-6.15 EA=1.529 EAIC=1.418 EAIE=1.533 
+ EAIS=1.529 EANC=1.625 EANE=1.932 EANS=1.529 EAP=1.12 EBBE=0 FC=0.9 
+ IBCI=1.0e-11 IBCIP=1.0e-11 IBCN=1.0E-11 IBCNP=1.0e-11 IBEI=1.64E-024 
+ IBEIP=0.6e-11 IBEN=6.0E-017 IBENP=0.6e-11 IKF=2.40168e-08 IKP=0
+ IKR=0.005 IS=3.99127e-26 ISMIN=1E-034 ISP=0 ISPMIN=0 ISRR=0.9247
+ ITF=0 KFN=0 MC=0.35 ME=0.33 MS=0.33 NCI=1.0 NCIP=1 NCN=1.0 
+ NCNP=2 NEI=1.155 NEN=2.20 NF=0.949660 NFP=1.0 NKF=0.122164 NR=1.012
+ PC=0.96 PE=3.18 PS=0.75 QBM=0 QTF=0 RBI=0.1 RBP=0.1 RBPMIN=0 
+ RBX=0.1 RCX=0.1 RE=0.2 RS=1E+06 RTH=1.0 TD=8.56E-13 TF=1.14e-11 
+ TNBBE=0 TNF=-0.0001 TNOM=20.85 TR=1.14e-11 TVBBE1=0.586e-3 
+ TVBBE2=0 VBBE=7.7 IBBE=1E-004 NBBE=1.0 VEF=0 VER=0 VRT=0 VTF=0
+ WBE=1 WSP=1 XII=5.758 XIKF=-2.572 XIN=1.903 XIS=3.834 XISR=0.7797 
+ XRBI=0 XRBP=0 XRBX=0 XRCX=0.0 XRE=0 XRS=0 XTF=0 HRCF=0
+ QCO=0 XRCI=0 RCI=0.1 VO=0 GAMM=0 XVO=1.0


* VBIC model generated by sgp2vbic.pl from q2n2222 level 1 BJT model (
.model q2n2222B npn
+ LEVEL=10  rcx=0.001 rci=0.001 rbx=0.001 rbi=0 re=0.001 rb=0.001 rc=0.001
+ is=3.295e-14 nf=1 nr=1 fc=0.5 cje=0 pe=0.75 me=0.33 cjc=0 cjep=0 pc=0.75
+ mc=0.33 cjcp=0 ps=0.75 ms=0.001 ibei=3.295e-16 nei=1 iben=0 nen=1.5
+ ibci=3.295e-14 nci=1 ibcn=0 ncn=2 vef=134.605947186551 ver=6485118644.83438
+ ikf=1e-11 nkf=0.2
+ ikr=0 tf=0 xtf=0 vtf=0 itf=0 tr=0 td=0 ea=1.11 eaie=1.11 eaic=1.11
+ eane=1.11 eanc=1.11 xis=3 xii=3 xin=3 kfn=0 afn=1 tnom=27

*.SENS param=
*+ q2n2222b:is,
*+ q2n2222b:ikf,
*+ q2n2222b:nkf,
*+ q2n2222b:nf
*+objfunc={(log10(abs(I(VC)))-(16.363*(abs(V(emit)))-23.41))}

.DC VE 0 -1.4 -1.0e-2
*.rol VE 0 -1.0 -1.0e-2
.PRINT DC FORMAT = tecplot {abs(V(emit))} {abs(I(VC))}  {abs(I(VB))}  

*.PRINT DC FORMAT = tecplot V(emit) {(log10(abs(I(VC)))-(16.363*(abs(V(emit)))-23.41))}

*.PRINT SENS FORMAT = noindex  {abs(V(emit))}

*.PRINT SENS FORMAT = tecplot {abs(V(emit))}

.end




