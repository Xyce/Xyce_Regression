* Test FIND measure type for .MEASURE FFT for a .TRAN
* analysis.  Test covers voltage-difference operators
* and lead currents.
*
* See SON Bugs 1280 and 1327 for more details.
******************************************************

.TRAN 0 1
.OPTIONS FFT FFT_ACCURATE=1 FFTOUT=1

V1 1 0 1
R1 1 2 1
R2 2 0 1

V3 3 0 SIN(0 1 1)
R3 3 0 1

* test with multiple .FFT lines.  Use UNORM format, because
* the FFT coeffs are returned in unnormalized format.
.FFT V(1) NP=8 WINDOW=HANN FORMAT=UNORM
.FFT V(1,2) NP=8 WINDOW=HARRIS FORMAT=UNORM
.FFT I(R3) NP=8 WINDOW=HARRIS FORMAT=UNORM

.MEASURE FFT FINDV1AT0 FIND V(1) AT=0
.MEASURE FFT FINDVR1AT0 FIND VR(1) AT=0
.MEASURE FFT FINDVI1AT0 FIND VI(1) AT=0
.MEASURE FFT FINDVM1AT0 FIND VM(1) AT=0
.MEASURE FFT FINDVP1AT0 FIND VP(1) AT=0
.MEASURE FFT FINDVDB1AT0 FIND VDB(1) AT=0

.MEASURE FFT FINDV1AT1 FIND v(1) AT=1.0
.MEASURE FFT FINDVR1AT1 FIND vr(1) AT=1.0
.MEASURE FFT FINDVI1AT1 FIND vi(1) AT=1.0
.MEASURE FFT FINDVM1AT1 FIND vm(1) AT=1.0
.MEASURE FFT FINDVP1AT1 FIND vp(1) AT=1.0
.MEASURE FFT FINDVDB1AT1 FIND vdb(1) AT=1.0

.MEASURE FFT FINDV1AT2 FIND V(1) AT=2.0
.MEASURE FFT FINDVR1AT2 FIND VR(1) AT=2.0
.MEASURE FFT FINDVI1AT2 FIND VI(1) AT=2.0
.MEASURE FFT FINDVM1AT2 FIND VM(1) AT=2.0
.MEASURE FFT FINDVP1AT2 FIND VP(1) AT=2.0
.MEASURE FFT FINDVDB1AT2 FIND VDB(1) AT=2.0

.MEASURE FFT FINDV1AT3 FIND V(1) AT=3.0
.MEASURE FFT FINDVR1AT3 FIND VR(1) AT=3.0
.MEASURE FFT FINDVI1AT3 FIND VI(1) AT=3.0
.MEASURE FFT FINDVM1AT3 FIND VM(1) AT=3.0
.MEASURE FFT FINDVP1AT3 FIND VP(1) AT=3.0
.MEASURE FFT FINDVDB1AT3 FIND VDB(1) AT=3.0

* Test with voltage difference syntax
.MEASURE FFT FINDV12 find VM(1,2) at=1.0

* lead current
.MEASURE FFT FINDI3 FIND I(R3) AT=1.0
.MEASURE FFT FINDDIR3 FIND Ir(R3) AT=1.0
.MEASURE FFT FINDII3 FIND ii(R3) AT=1.0
.MEASURE FFT FINDIM3 FIND IM(R3) AT=1.0
.MEASURE FFT FINDIP3 FIND IP(R3) AT=1.0
.MEASURE FFT FINDIDB3 FIND Idb(R3) AT=1.0

* Test rounding
.MEASURE FFT FINDVR1ROUND1 FIND VR(1) AT=1.25
.MEASURE FFT FINDVI1ROUND2a FIND VI(1) AT=1.75
.MEASURE FFT FINDVM1ROUND2b FIND VM(1) AT=2.4
.MEASURE FFT FINDVP1ROUND3 FIND VP(1) AT=2.9
.MEASURE FFT FINDVDB1ROUND0 FIND VDB(1) AT=0.3

.PRINT TRAN V(1) V(2) V(3)
.END
