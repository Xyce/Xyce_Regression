* This netlist is equivalent to Step 1 for the AllMeasures.cir
* netlist. It has V1:VA=600.

.TRAN 0 1
.PRINT TRAN V(1) V(2) V(3)

V1 1 0 SIN(0 600 1)
V3 3 0 SIN(0 200 2)
R1 1 2 1
R2 2 0 1
R3 3 2 1

.FFT V(2) NP=16 WINDOW=HANN FORMAT=UNORM


.MEASURE FFT ENOB ENOB V(2)
.MEASURE FFT SFDR SFDR V(2)
.MEASURE FFT SNDR SNDR V(2)
.MEASURE FFT THD THD V(2)

.MEASURE FFT FINDV2AT1 FIND v(2) AT=1.0
.MEASURE FFT FINDVR2AT1 FIND vr(2) AT=1.0
.MEASURE FFT FINDVI2AT1 FIND vi(2) AT=1.0
.MEASURE FFT FINDVM2AT1 FIND vm(2) AT=1.0
.MEASURE FFT FINDVP2AT1 FIND vp(2) AT=1.0
.MEASURE FFT FINDVDB2AT1 FIND vdb(2) AT=1.0

.END
