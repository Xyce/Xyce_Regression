*Sample netlist for BSIM-MG
*Drain current symmetry


.options device temp=25

* --- Voltage Sources ---
vdrain drain 0 dc 0
esource source 0 drain 0 -1
vgate gate  0 dc -1.0
vbulk bulk 0 dc 0


* --- Transistor ---
M1 drain gate source bulk pmos1 TFIN=15n L=30n NFIN=10 NRS=1 NRD=1

* --- DC Analysis ---
.dc vdrain -0.1 0.1 0.001 vgate 0.0 -1.0 -0.2
.print dc v(drain) v(gate) {-I(vdrain)}
.print sens v(drain) v(gate)

.sens param=pmos1:toxp,pmos1:vsat objfunc={I(vdrain)}
.options sensitivity direct=1 adjoint=0


******** BSIM-MG 105 Sample Modelcard for PMOS ********

** The BSIM-MG sample modelcard below was not extracted/obtained
** from/based on any real technologies. It should not be used for any
** other purposes except for benchmarking the implementation of BSIM-MG
** against BSIM Team's standard results

.model pmos1 pmos LEVEL=110
+ BULKMOD = 1
+ CAPMOD = 0
+ COREMOD = 0
+ CGEOMOD = 0
+ DEVTYPE = 0
+ GEOMOD = 0
+ GIDLMOD = 1
+ IGBMOD = 0
+ IGCMOD = 1
+ IIMOD = 0
+ NGATE  = 0
+ NQSMOD = 0
+ RDSMOD = 0
+ RGATEMOD = 0
+ RGEOMOD = 0
+ NSEG = 5
+ SDTERM = 0
+ SHMOD = 0
+ AGIDL = 2E-12
+ AGISL = 2E-12
+ AIGC = 0.007
+ AIGD = 0.006
+ AIGS = 0.006
+ AT  = 0.0008234
+ BG0SUB  = 1.17
+ BGIDL = 1.50E+08
+ BGISL = 1.50E+08
+ BIGC = 0.0015
+ BIGD = 0.001944
+ BIGS = 0.001944
+ CDSC = 0.003469
+ CDSCD = 0.001486
+ CFD = 0.2e-10
+ CFS = 0.2e-10
+ CGBL  = 0
+ CGBO  = 0
+ CGDL  = 0
+ CGDO = 1E-10
+ CGSL  = 0
+ CGSO = 1E-10
+ CIGC = 1
+ CIGD = 1
+ CIGS = 1
+ CIT = 0
+ CKAPPAD  = 0.6
+ CKAPPAS  = 0.6
+ CTH0  = 1.243E-06
+ DELTAVSAT  = 11.56
+ DELTAW  = 0
+ DELTAWCV  = -1.00E-08
+ DLBIN  = 0
+ DLC  = -9.2E-09
+ DLCIGD = 5.00E-09
+ DLCIGS = 5.00E-09
+ DROUT = 4.97
+ DSUB = 0.5
+ DVT0 = 0.05006
+ DVT1 = 0.4
+ DVTSHIFT = 0
+ EASUB  = 4.05
+ EGIDL = 1.142
+ EGISL = 1.142
+ EOT  = 2.10E-09
+ EOTACC  = 3.00E-10
+ EOTBOX  = 1.40E-07
+ EPSROX  = 3.9
+ EPSRSP  = 3.9
+ EPSRSUB  = 11.9
+ ETA0  = 0.03952
+ ETAMOB = 4
+ ETAQM  = 0.54
+ EU = 0.05
+ FPITCH  = 4.00E-08
+ HFIN  = 3.00E-08
+ IGT  = 3.5
+ K1RSCE = 0
+ KSATIV = 1.592
+ KT1 = 0.08387
+ KT1L = 0
+ L  = 2.50E-08
+ LINT  = -2.5E-09
+ LPE0 = 0
+ LCDSCD = 0
+ LCDSCDR = 0
+ LRDSW = 1.3
+ LVSAT = 1441
+ MEXP = 2.491
+ NBODY  = 1E+22
+ NC0SUB  = 2.86E+25
+ NI0SUB  = 1.1E+16
+ NIGC = 0.5
+ NSD  = 2E+26
+ PCLM = 0.01
+ PCLMCV = 0.013
+ PCLMG = 1
+ PCLMGCV = 0
+ PDIBL1 = 800
+ PDIBL2 = 0.005704
+ PHIG  = 4.678
+ PHIN = 0.05
+ POXEDGE = 1.152
+ PQM  = 0.66
+ PRT  = 0.002477
+ PRWG  = 0
+ PTWG  = 6.322
+ PTWGT  = 0.0015
+ PVAG = 200
+ QM0  = 2.183E-12
+ QMFACTOR  = 0
+ RDSW  = 190.6
+ RDSWMIN  = 0
+ RDWMIN  = 0
+ RSHD  = 0
+ RSHS  = 0
+ RSWMIN  = 0
+ RTH0  = 0.15
+ TBGASUB = 0.000473
+ TBGBSUB = 636
+ TFIN  = 1.40E-08
+ TGIDL  = -0.01
+ TMEXP  = 0
+ TNOM = 25
+ TOXP  = 2.1E-09
+ TOXG  = 2.1E-09
+ U0 = 0.02935
+ UA = 1.133
+ UA1 = 0.00134
+ UCS = 0.2672
+ UCSTE = 0
+ UD = 0.0105
+ UD1 = 0
+ UP = 0
+ UTE = 0
+ UTL = 0.001
+ VSAT = 48390
+ VSAT1 = 48390
+ VSATCV = 48390
+ WR  = 1
+ WTH0  = 2.60E-07
+ XL  = 0

.end
