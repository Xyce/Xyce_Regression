*******************************************************************************
* This netlist is equivalent to Step 0 for the RiseFallCrossTest.cir netlist.
* It has VS1:VA=1
*
*******************************************************************************
*
** use a damped sinusoid
VS  1  0  SIN(0 1.0 1KHZ 0 2.0)
VP  2  0  PULSE( 0 100 0.2ms 0.2ms 0.2ms 1ms 2ms )

R1  1  0  100
R2  2  0  100

.TRAN 0  10ms
.PRINT TRAN FORMAT=NOINDEX V(1) V(2)

* test RISE, FALL and CROSS qualifiers
.measure tran Rise4 min V(1) RISE=4
.measure tran Fall3 min V(1) FALL=3
.measure tran Cross8 min V(1) CROSS=8

* this test should return -1 since the RISE, FALl and CROSS 
* values are too high
.measure tran returnNegOneRise min V(1) RISE=12
.measure tran returnNegOneFall min V(1) FALL=11
.measure tran returnNegOneCross min V(1) CROSS=20

.measure tran v2Rise4 min V(2) RISE=4

.END

