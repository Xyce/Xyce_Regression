N-Channel MESFET Circuit
*
VDS 2 0 2V
VGS 3 0 pulse (-1 1 1ns 1ns 1ns 1us 2us)
VSS 4 0 0
Z1 2 3 4 MESMOD AREA=1.4
.MODEL MESMOD NMF
+ LEVEL=1 BETA=1.4E-3
+ RD=46 RS=46 VTO=-1.3 LAMBDA=0.03 ALPHA=3 CGS=1uf CGD=1uf

.options timeint method=trap
.options nonlin-tran rhstol=1.0e-7

.tran 1ns 10us 
.PRINT TRAN PRECISION=10 
+ P(Z1) W(Z1) {ID(Z1)*V(2) + IG(Z1)*V(3)} {-1*(P(VDS)+P(VGS))}
+ ID(Z1) IG(Z1) IS(Z1) I(VDS) I(VGS) V(2) V(3) 

.END

