* Unit test of Power Grid Branch Device, in I=YV format

* Vary the voltage at bus 1 to check if the answers match theory,
* given on pg.250-254 of Kundar. Ammeter is defined so that power
* flows from bus 1 into the branch between buses 1 and 2
V1R bus1R ammBus1R 1V
V1I bus1I ammBus1I 0V
Vamm1R 0 ammBus1R 0V
Vamm1I 0 ammBus1I 0V

* Have bus 2 be the slack bus. Ammeter is defined so that power 
* flows from branch between buses 1 and 2 into bus 2, so as to match
* equations in Kundar.
V2R bus2R ammBus2R 1V
V2I bus2I ammBus2I 0V
Vamm2R ammBus2R 0 0V
Vamm2I ammBus2I 0 0V

* simple reactance-only branch has closed form solution for power flow
YPowerGridBranch pg1 bus1R bus2R bus1I bus2I AT=IV R=0.0 X=2.0 B=0.0

.DC V1I -0.5 1.0 0.5 V1R -0.5 1.0 0.5
.PRINT DC width=10 precision=6 V(bus1R) V(bus1I)
+ {V(bus1R)*I(Vamm1R)+V(bus1I)*I(Vamm1I)}
+ {V(bus1I)*I(Vamm1R)-V(bus1R)*I(Vamm1I)}
+ {V(bus2R)*I(Vamm2R)+V(bus2I)*I(Vamm2I)}
+ {V(bus2I)*I(Vamm2R)-V(bus2R)*I(Vamm2I)}
 
.end
