MMSZ5229BT1 Zener Subcircuit using Pspice level 2 diode at elevated temperature
********************************************************************************
VIN 20 0 DC 1V
VMON 20 10 0
*
X1 10 0 MMSZ5229
.OPTIONS DEVICE TEMP=35
*
.OPTIONS DEVICE GMIN=1.0E-15
*
.SUBCKT MMSZ5229 1 2 
D1 1 2  DFOR 
D2 4 1  DLEAKLO 
D4 2 4  DLEAKHI 
D3 2 3  DBLOCK 
IC 1 3 83.27758 
RC 1 3 0.0311172 RTEMP
*
.MODEL DFOR D  ( LEVEL=2  ISR=3.4E-11  NR=2.00  IKF=0 
+ IS = 0.27E-14  N = 1.05  BV = 75  IBV = 0.001  RS = 0.14 
+ CJO = 2.682354E-10  VJ = 0.5259017  M = 0.3225012  FC = 0.5
+ TT = 150E-09  EG = 1.11  XTI = 4 )
*
.MODEL DLEAKLO D (
+ IS = 9.354E-11  N = 6.156  XTI = 50.11872  EG = 0.1  RS = 0 )
.MODEL DLEAKHI D (
+ IS = 2.49E-05  N = 7.691304  XTI = 90.78205  EG = 0.1  RS = 1 )
.MODEL DBLOCK D ( 
+ IS = 1.45E-12  N = 2.987045  RS = 0.05324657  XTI = 0.1  EG = 0.1  CJO = 0 )
.MODEL RTEMP R (
+ TC1 = -0.00233213  TC2 = 2.3137E-06 )
.ENDS
*
.DC VIN 0.2 1.001 0.016 
*.DC VIN 0.1 1.001 0.018 
*.DC VIN -0.5 -5.51 -0.07
*.DC VIN -0.5 -4.01 -0.1
*.DC VIN -3.76 -4.77 -0.02
.PRINT DC  V(20) I(VMON)
*
.END

