CD4020B PMOS Test Circuit - Level 1 Mosfet with temp effects

VD 1 0 DC 0
VG 3 0 DC 0
VS 4 0 DC 0
VID 1 2 DC 0

.options device TEMP=15
*.options device TEMP=27
*.options device TEMP=66

M1 2 3 4 4 CD4020 W=80u L=6.3u 

.MODEL CD4020 PMOS (  LEVEL=1  TNOM=15 TEMPMODEL=QUADRATIC
+  UO=466.5  VTO=-1.45 TOX=1.1E-07 KP=2.3e-5
+  NSUB=1.379E+16 LD=0 NSS=1E10
+  RSH=0  RS=0  RD=10  IS =1E-14 
+  LAMBDA=0.3
+  CGDO=1PF CGSO=1PF CGBO=1PF CBD=1PF CBS=1PF 
+  ALPHANINT=1.3e-11  ALPHANOXT=0   )

.MODEL CD4020 PMOS (  LEVEL=1  TNOM=27 TEMPMODEL=QUADRATIC
+  UO=566.5  VTO=-1.40 TOX=1.1E-07 KP=2.3e-5
+  NSUB=1.379E+15 LD=0 NSS=1E10
+  RSH=0  RS=0  RD=1  IS =1E-14 
+  LAMBDA=0.3
+  CGDO=1PF CGSO=1PF CGBO=1PF CBD=1PF CBS=1PF 
+  ALPHANINT=1.3e-11  ALPHANOXT=0   )

.MODEL CD4020 PMOS (  LEVEL=1  TNOM=66 TEMPMODEL=QUADRATIC
+  UO=666.5  VTO=-1.55 TOX=1.1E-07 KP=2.3e-5
+  NSUB=1.379E+14 LD=0 NSS=1E10
+  RSH=0  RS=0  RD=0  IS =1E-14 
+  LAMBDA=0.3
+  CGDO=1PF CGSO=1PF CGBO=1PF CBD=1PF CBS=1PF 
+  ALPHANINT=1.3e-11  ALPHANOXT=0   )

.DC VD 0 -1.0 -0.1v VG -1.6 -2.01 -0.1v
*.DC VD 0 -8.0 -1.0v VG -2.0 -5.01 -0.5v

.PRINT DC V(1) V(3) I(VID)
.END
*
