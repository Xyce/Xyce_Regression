**********************************************************
* Test M=0 error condition for the multiplicity factor (M)
* for Resistor, Thermal Resistor, Inductor and Capacitor
* devices.  M must be non-negative.
*
*
*
* See SON Bug 834 for more details.
**********************************************************

* Test with and without a model card for Level 1 Resistor.
V1  1   0 1
R1  1  1a 1.25 M=0
R1a 1a  0 1 M=0
.MODEL R1amodel R R=4 LEVEL=1

* Test Level 2 Resistor
V2  2   0  1
R2a 2  2a  1.68e-4
R2  2a  0 copperConstant L=0.1 a=1e-5 M=0
* model card
.include copper.constant

* Inductor
I3 3 0 PULSE(0 5V 0 1MS 1MS 10MS 25MS) 
L3 3a 0 L=10mH M=0
R3 3 3a 0.001 

* Capacitor
* C value missing from instance line.
c4 4  0 C=1uf IC=1 M=0 
r4 4 4a 1K 
v4 4a 0 0V 

* analysis and print statements.
.DC V1 1 1 1
.PRINT DC V(1a) V(2a) V(3a) V(4a)

.END
