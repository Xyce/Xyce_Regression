**********************************************************
* Netlist tests that DC output in TOUCHSTONE or TOUCHSTONE2
* formats default to STD format (.prn file with an Index column)
*
*********************************************************

V1 1 0 1
R1 1 0 1

.DC V1 1 5 1
.PRINT DC FORMAT=TOUCHSTONE V(1)
.PRINT DC FILE=dc-touchstone-defaults-to-prn.cir.ts2 FORMAT=TOUCHSTONE2 V(1)

.END

