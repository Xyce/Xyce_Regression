****************************************************
* Test Touchstone1 output using a 1-Port S-Parameter
* analysis.  This also verifies DATAFORMAT=MA and
* DATAFORMAT=DB for a number-of-ports not equal to 2.
*
* It also verifies that specifying SPARCALC=1 on a
* .LIN line is okay.
*
* There is no .PRINT AC line.  So, there should
* not be any .AC output.
****************************************************

* RC ladder circuit
* Note that all ports (P devices) must use a common
* Reference Node, which is 0 here.
P1 1  0  port=1  z0=50

C1 2 0 1e-2
Rgs 1 2 0.02

.subckt RCBlock IN OUT GND
R1 IN OUT 20
C1 IN OUT 1p
Cg1 OUT GND 1p
.ends

X1 2 3 0 RCBlock
X2 3 4 0 RCBlock
X3 4 5 0 RCBlock
X4 5 6 0 RCBlock
X5 6 7 0 RCBlock
X6 7 8 0 RCBlock
X7 8 9 0 RCBlock
X8 9 10 0 RCBlock
X9 10 11 0 RCBlock
X10 11 12 0 RCBlock

.AC DEC 10 10  1e5

.LIN FORMAT=TOUCHSTONE SPARCALC=1
.LIN FORMAT=TOUCHSTONE DATAFORMAT=MA FILE=sparams-ts1-1port.cir.ma.s1p
.LIN FORMAT=TOUCHSTONE DATAFORMAT=DB FILE=sparams-ts1-1port.cir.db.s1p

.END
