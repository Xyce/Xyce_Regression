dup-subcircuit.cir
* this circuit demonstrates a parser error, in which 2 sources of the same
* name are specified, and not trapped.


.subckt rNodes a b 
R1 a b 1
R1 b 0 1
.ends

V1 22 0 4
V2 1 0 5

.dc V1 7 7 1
.print dc V(1) V(22)

XvNodes 1 22 rNodes

.end
