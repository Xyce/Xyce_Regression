TEST A1_DUP of subcircuit regression tests
* **********************************************************************
* A simple pair of MOSFET level 3 inverters
* The inverters are constructed from dissimilar mosfets, just for testing 
* purposes
*
* Test A1 puts the two inverters of test A0 into separate subcircuits.
* No parameters are used, and separate versions of global model statements
* are kept.
*
*Note added by ERK on 10/22/09:
* This test is identical to subckt_a1.cir, except that the SUBCKT definitions
* now all have some node duplications in the definition, per bug 1665.  It
* should produce the same answer.
*
* Author:   $Author$
* Revision: $Revision$
* Date:     $Date$
*
* **********************************************************************

.subckt INV1 IN OUT VDD GND VDD
MN1 OUT IN GND GND CD4012_NMOS L=5u W=175u
MP1 OUT IN VDD VDD CD4012_PMOS L=5u W=270u
.ends

.subckt INV2 IN OUT VDD GND OUT
MN1a OUT IN GND GND CD4012_NMOS1 L=5u W=175u
MP1a OUT IN VDD VDD CD4012_PMOS1 L=5u W=270u
.ends

Xinv1 IN MID VDD 0 VDD INV1
Xinv2 MID OUT VDD 0 OUT INV2
VDDdev 	VDD	0	5V
RIN	IN	1	1K
VIN1  1	0  5V PULSE (5V 0V 1.5us 5ns 5ns 1.5us 3.01us)
R1    OUT  0  10K  
C2    OUT  0  0.1p

.tran 20ns 30us
.print tran PRECISION=10 WIDTH=19 v(out) v(in) v(1)


***** original mosfets
.MODEL cd4012_nmos NMOS (
+ LEVEL = 3 UO = 190   VTO = 1.679   TOX = 6E-08   NSUB = 8.601E+15
+ NSS = 0   RS = 13.21   RD = 11.59   RSH = 0   IS = 1E-14
+ VMAX = 4.206E+04 NFS=1E10  GAMMA=0.37 PHI=0.65 
+ XJ = 7.1E-06   LD = 8.6E-07   DELTA = 0   THETA = 0.0021   ETA = 0.057   KAPPA = 0.15
+ KP = 2.161E-05  L=5u W=175u
+ CBD=0.1P CBS=0.1P PB=0.81 CGSO=2P CGBO=4P CGDO=2P CJ=2E-4 MJ=0.5 CJSW=1E-9
+ MJSW=0.5 JS=1E-8 TPG=0 KF=1E-25 AF=1 FC=0.5 TNOM=27)
.MODEL cd4012_pmos PMOS (
+ LEVEL = 3  UO = 310  VTO = -1.6  TOX = 6E-08  NSUB = 5.701E+15
+ NSS = 0    VMAX = 5.374E+04   RS = 5.359   RD = 93.66   RSH = 0   IS = 1E-14
+ XJ = 7.9E-06   LD = 3E-08   DELTA = 0   THETA = 0.0278   ETA = 0.535   KAPPA = 0.643
+ KP = 1.711E-05 L=5u W=270u GAMMA=0.37 PHI=0.65 NFS=1E10
+ CBD=0.1P CBS=0.1P PB=0.81 CGSO=2P CGBO=4P CGDO=2P CJ=2E-4 MJ=0.5 CJSW=1E-9
+ MJSW=0.5 JS=1E-8 TPG=0 KF=1E-25 AF=1 FC=0.5 TNOM=27)
******slightly modified mosfets (changed VTO of both)
.MODEL cd4012_nmos1 NMOS (
+ LEVEL = 3 UO = 190   VTO = 1.0   TOX = 6E-08   NSUB = 8.601E+15
+ NSS = 0   RS = 13.21   RD = 11.59   RSH = 0   IS = 1E-14
+ VMAX = 4.206E+04 NFS=1E10  GAMMA=0.37 PHI=0.65 
+ XJ = 7.1E-06   LD = 8.6E-07   DELTA = 0   THETA = 0.0021   ETA = 0.057   KAPPA = 0.15
+ KP = 2.161E-05  L=5u W=175u
+ CBD=0.1P CBS=0.1P PB=0.81 CGSO=2P CGBO=4P CGDO=2P CJ=2E-4 MJ=0.5 CJSW=1E-9
+ MJSW=0.5 JS=1E-8 TPG=0 KF=1E-25 AF=1 FC=0.5 TNOM=27)
.MODEL cd4012_pmos1 PMOS (
+ LEVEL = 3  UO = 310  VTO = -1.0  TOX = 6E-08  NSUB = 5.701E+15
+ NSS = 0    VMAX = 5.374E+04   RS = 5.359   RD = 93.66   RSH = 0   IS = 1E-14
+ XJ = 7.9E-06   LD = 3E-08   DELTA = 0   THETA = 0.0278   ETA = 0.535   KAPPA = 0.643
+ KP = 1.711E-05 L=5u W=270u GAMMA=0.37 PHI=0.65 NFS=1E10
+ CBD=0.1P CBS=0.1P PB=0.81 CGSO=2P CGBO=4P CGDO=2P CJ=2E-4 MJ=0.5 CJSW=1E-9
+ MJSW=0.5 JS=1E-8 TPG=0 KF=1E-25 AF=1 FC=0.5 TNOM=27)
.end
