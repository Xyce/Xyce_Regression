* Test .FFT and .MEASURE FFT for lead currents for
* multiterminal devices.  They should work for all
* measures but FIND-AT.
*
* See SON Bugs 1280 and 1332 for more details.
****************************************************

.OPTIONS FFT FFT_ACCURATE=1 FFTOUT=1
.options nonlin-tran rhstol=1.0e-7

.tran 1ns 1us
.PRINT TRAN IB(Q1) IC(Q1) IE(Q1) ID(J1) IG(J1) IS(J1)

.FFT IB(Q1) NP=64 WINDOW=HAMM
.FFT IC(Q1) NP=64 WINDOW=HAMM
.FFT IE(Q1) NP=64 WINDOW=HAMM

.FFT ID(J1) NP=64 WINDOW=HAMM
.FFT IG(J1) NP=64 WINDOW=HAMM
.FFT IS(J1) NP=64 WINDOW=HAMM

.MEASURE FFT THDIB THD IB(Q1)
.MEASURE FFT SNDRIB SNDR IB(Q1)
.MEASURE FFT ENOBIB ENOB IB(Q1)
.MEASURE FFT SNRIB SNR IB(Q1)
.MEASURE FFT SFDRIB SFDR IB(Q1)

.MEASURE FFT THDIC THD IC(Q1)
.MEASURE FFT SNDRIC SNDR IC(Q1)
.MEASURE FFT ENOBIC ENOB IC(Q1)
.MEASURE FFT SNRIC SNR IC(Q1)
.MEASURE FFT SFDRIC SFDR IC(Q1)

.MEASURE FFT THDIE THD IE(Q1)
.MEASURE FFT SNDRIE SNDR IE(Q1)
.MEASURE FFT ENOBIE ENOB IE(Q1)
.MEASURE FFT SNRIE SNR IE(Q1)
.MEASURE FFT SFDRIE SFDR IE(Q1)

.MEASURE FFT THDID THD ID(J1)
.MEASURE FFT SNDRID SNDR ID(J1)
.MEASURE FFT ENOBID ENOB ID(J1)
.MEASURE FFT SNRID SNR ID(J1)
.MEASURE FFT SFDRID SFDR ID(J1)

.MEASURE FFT THDIG THD IG(J1)
.MEASURE FFT SNDRIG SNDR IG(J1)
.MEASURE FFT ENOBIG ENOB IG(J1)
.MEASURE FFT SNRIG SNR IG(J1)
.MEASURE FFT SFDRIG SFDR IG(J1)

.MEASURE FFT THDIS THD IS(J1)
.MEASURE FFT SNDRIS SNDR IS(J1)
.MEASURE FFT ENOBIS ENOB IS(J1)
.MEASURE FFT SNRIS SNR IS(J1)
.MEASURE FFT SFDRIS SFDR IS(J1)

* bjt
vie 0 1b 0
vic 0 3b 5
vib 0 2b pulse(0 1 50ns 400s 50ns 1us)
q1 3b 2b 1b qjunk

.model qjunk npn
+bf=130 br=1 is=3e-14
+tf=1e-8 vjs=0.68 ne=1.6 nc=2.0 rb=450
+cje=1uf cjc=1uf cjs=1uf ikf=0.002 ikr=0.002 vaf=50 var=50
+nf=1.0 ise=0 nr=1 isc=0 irb=0 rbm=450 re=0 rc=0 vje=0.75
+mje=0.33 xtf=0 vtf=100 itf=0 ptf=0 vjc=0.75 mjs=0 xtb=0
+eg=1.11 xti=3 kf=0 af=1 fc=0.5 tnom=27

*Drain curves
Vds2 1 0 5V
Vgs2 2 0 pulse (0 1 10ns 80ns 10ns 1us)
J1 1 2 0 SA2109
*
.MODEL SA2109 NJF
+ LEVEL=2
+ BETA= 0.0003790
+ VTO = -3.760
+ PB = 0.650
+ LAMBDA = 0.01240
+ DELTA = 0.370;
+ THETA = 0.01120;
+ RD = 0.0
+ RS = 104.5
+ FC = 0.5
+ IS = 1.393E-10
+ AF = 1.0
+ KF = 0.05
+ CGS= 1uf
+ CGD= 1uf
*

.end
