Test of multiple print lines
* This tests that multiple .print TRAN lines to the default file are the
* same as a single .print TRAN line with all arguments aggregated.
* It further tests that a second pair of print lines to a different file
* also aggregate the output list.
* both outputs should be compared to the output of the associated _baseline
* netlist.
*
* This differs from test 2 because it uses continuation, and therefore produces
* an extra output file of continuation data, called "netlist.HOMOTOPY.prn" in
* this case.  This extra output file should also have its lines of data
* built up from the combined variable lists of the two print lines.

R1 1 0 10
V1 1 0 sin (0 10 10MEG 0 0)

.print TRAN v(1)
.print TRAN I(v1)
.print HOMOTOPY v(1)
.print HOMOTOPY I(v1)

.tran 1ns 10ns
.options nonlin maxstep=200 continuation=gmin reltol=1.0e-2 abstol=1.0e-6 rhstol=1.0e-4

.options loca stepper=natural predictor=constant stepcontrol=adaptive

.end
