Test for bug 1190 SON, for mutual inductors.
*
* This is re-purposed from the bug 28 SON test.
*
* The point of this test, like all tests in this directory, is to
* prove that a complex device, which has a "processParams" functions,
* can have a device parameter depend on a .param, which in turn 
* depends on a .global_param, which in turn is modified during
* the calculation via .STEP.
*
* This is possible now, with the new expression library, as it does 
* not treat .param as constants.  
*
* This circuit is the "baseline" in that it doesn't use .param to set the scalefac.
*

.global_param winding1=10
.global_param winding2=100
.global_param scalefac=1
.subckt transformer node1 node6
Llead4 node1 0 {winding1}
Llead5 node5 node6 {winding2*scalefac}
Llead6 node6 node7 {winding2*scalefac}
Ktrans2 Llead4 Llead5 Llead6 1.0 nlcore

.model nlcore CORE c=0.001

rload3  node5 0 100
rpathtg2 node7 0 1
.ends

Vinput node1 0 sin(0 14 120 0 0)
X1 node1 node6 transformer
rload4  node6 0 100

.tran 0 10m 
.print tran v(node1) v(node6)
.step scalefac list 0.5 .75 1
.end

