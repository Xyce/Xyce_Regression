* test of coupled inductor parameters on the .PRINT line
V1 1 0 SIN(0 1 1KHz)
R1 1 0 1
R2 2 0 1

* mutual inductor definition
L1 1 0 1e-3
L2 2 0 2mH
K1 L1 L2 0.75

.TRAN 0 1ms 
.PRINT TRAN V(1) V(2) L1:L {L1:L}

.END 

