Local Variation test
*
V1 1 0 1.0

.param c=2
.param myvar=c+rand()


r1 1 2 myvar
r2 2 0 1.0

.dc V1 1 1 1
.print dc precision=12 width=21 v(1) v(2) 

.sampling useExpr=true

.options samples numsamples=10 seed=1923635719
+ outputs={v(1)+0.2}
+ sample_type=lhs
+ stdoutput=false

.result {r1:R}

.END

