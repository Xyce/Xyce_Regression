*************************************************
* Test of various invalid combinations of FREQ,
* FMIN and FMAX values on .FFT lines.
*
*************************************************
.TRAN 0 1

V1 1 0 1
R1 1 2 1
R2 2 3 1
R3 3 4 1
R4 4 5 1
R5 5 6 1
R6 6 0 1

.PRINT TRAN V(1)

.FFT V(1) FREQ=0
.FFT V(2) NP=16 FREQ=9 ; max frequency in FFT is 8
.FFT V(3) NP=16 FMIN=9
.FFT V(4) FMAX=1 ; This implicitly has FREQ=1
.FFT V(5) FREQ=2 FMAX=0
.FFT V(6) FMIN=5 FMAX=4

.END
