***************************************************************
* Test for P() and W() for devices that do not implement
* those calculations for .AC.
*
* The goal of this test is to ensure that Xyce exits gracefully
* with a reasonable error message, instead of printing "all
* zeros" for those devices.  See SON Bug 855 for more details.
*
***************************************************************

* AC ANALYSIS: RESISTOR DIVIDER, AMP, AND LP FILTER
*
* RESISTOR DIVIDER
V1  1 0 DC 5.0 AC  1.0
R1  1 2 100K
R2  2 0 100K
*
* AMP AND LP FILTER
EAMP  3 0 2 0 1
RLP1  3 4 100
CLP1  4 0 1.59NF

I3 3 0 DC 5.0 AC 1.0
R3 3 0 100K

* It is important to test the case of the .OP statement coming
* before the .AC statement.
.OP
.AC DEC 5 100 1MEG

* I() is not supported for the R, I and C devices, amongst others
* for .AC analyses.
.PRINT AC I(V1) I(I3) I(R1) II(CLP1) IP(R2) IM(RLP1) IDB(R3)

.END

