1D PDE Diode test circuit 
*
* This is a very simple test of the 1-D PDE diode device
* in Xyce.  DC sweep.  Full Newton only, serves as a baseline for the
* corresponding 2-level test.
*
* Creator: Eric Keiter
* Date   : 2/25/2019
*
R 1 2 1000.0
V1 2 0 -0.21
V2 3 0  0.0

YPDE d1 1 3 DIODE na=1.0e15 nd=1.0e15  tecplotlevel=0 gnuplotlevel=0
+ graded=0 l=5.0e-4 wj=0.1e-3 nx=101  area=1.0 
+ mobmodel=carr
+ useOldNi=true

.MODEL DIODE  ZOD 
.DC V1 0.0 -0.21 -0.01
*.options NONLIN maxstep=50 maxsearchstep=3 searchmethod=1 abstol=1.0e-17 nox=0 debuglevel=-100
.options device debuglevel=-100 
.options timeint debuglevel=-100   

.print DC v(2) {v(1)+0.1} {I(V1)+1.0e-9} {I(V2)-1.0e-9}
.END
