********************************************************
* Test error messsage when .DATA line has an freq
* entry that is not > 0
*
* See SON Bug 1146 for more details.
********************************************************

.global_param mag=1
.global_param phase=0.1

* Trivial high-pass filter (V-C-R) circuit.
R1 b 0 2
C1 a b 1u
V1 a 0 AC {mag} {phase}

.DATA table
+  mag  phase   freq
+  1.0   0.1   1.0e0
+  2.0   0.2   1.0e1
+  3.0   0.3   1.0e2
+  4.0   0.4   1.0e3
+  5.0   0.5   1.0e4
+  6.0   0.6   1.0e5
+  1.0   0.1   0.0e0
.enddata

.print AC vm(b)
*.ac dec 5 100 1e6
.ac data=table

.end
