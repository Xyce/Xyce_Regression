************************************************
* Test .DATA and its use with .MEASURE and 
* -remeasure for .TRAN.
*
* See SON Bug 1160 for more details.
************************************************
VT1 4 0 PWL 0 0 1 1
R1  4 5 10
R2  5 0 5

.data test
+ r1   r2  
+ 1.0000e+00  4.0000e+00 
+ 2.0000e+00  2.0000e+00 
.enddata

.STEP data=test
.TRAN 0 1
.OPTIONS OUTPUT INITIAL_INTERVAL=0.1
.print TRAN {R1:R} {R2:R} V(4) V(5)
.MEASURE TRAN MAXV5 MAX V(5)

.END

