* Test DC mode support for AVG Measures. This bug covers:
*
*   1) The case of one variable (vsrc1) on the .DC line,
*      with one variable (vsrc2) in the .STEP statement.
*
*   2) The DC values of the swept variable (vsrc1) are
*      monotonically decreasing.
*
* See SON Bug 1270 for more details.
****************************************************************

vsrc1   1a 0 1
rload1a 1a 1b 0.1
rload1b 1b 0 1

vsrc2   2a 0 1
rload2a 2a 2b 0.1
rload2b 2b 1b 0.1

* Reverse the step order on vsrc1 (from the test in MEASURE_DC)
* to make sure that both increasing and decreasing sequences of
* values are tested.
.DC vsrc1 5 1 -1
.STEP VSRC2 1 4 3

* Note: vsrc1:DCV0 is the syntax for printing the DC value of vsrc1,
* at it is swept.
.print dc vsrc1:DCV0 vsrc2:DCV0 v(1a) v(2a) v(1b) v(2b)

* WHEN
.MEASURE DC whenv1b3 WHEN v(1b)=3
.MEASURE DC whenExp1 when v(1b)={v(2b)+0.1}
.MEASURE DC whenExp2 when {v(1b)-0.1}=v(2b)

* FIND-WHEN
.MEASURE DC findv2bwhenv1b3 find v(2b) when v(1b)=3

* Signifies end of test. .sh file looks for a measure named lastMeasure.
* This is needed for compatibility for testing with a verbose build, which
* is often used by the Xyce developers.
.measure dc lastMeasure max v(1b)

.end
