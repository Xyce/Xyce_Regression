*******************************************************************************
* This netlist is equivalent to Step 3 for the MinTest.cir netlist.
* It has VS1:VA=2 and VS3:V0=-0.5
*
*******************************************************************************
*
* a few sources of different types
VS1  1  0  SIN(0 2 1KHz 0 0)
VP  2  0  PULSE( 0 100 0.2ms 0.2ms 0.2ms 1ms 2ms )
VS3  3  0  SIN(-0.5 1.0 1KHZ 0 500)
VS4  4  0  SIN(0.5 -1.0 1KHZ 0 500)

R1  1  0  100
R2  2  0  100
R3  3  0  100
R4  4  0  100

.TRAN 0  3ms
.PRINT TRAN FORMAT=NOINDEX V(1) V(2) V(3) V(4)

* plain test
.measure tran minSine min V(1)
.measure tran min2 MIN v(2)

* add TO-FROM modifiers
.measure tran minHalfSine min V(1) from=0 to=0.5e-3

* mix in TDs before and after FROM value.
.measure tran sine10 min V(1) FROM=0 TO=0.25e-3 TD=0.1e-3
.measure tran sine15 min V(1) FROM=0.00015 TO=0.25e-3 TD=0.1e-3
.measure tran sine20 min V(1) FROM=0.0002 TO=0.25e-3 TD=0.1e-3

* these tests should return -1 and -100
.measure tran returnNegOne min V(1) FROM=0.2e-3 TO=0.25e-3 TD=0.5e-3
.measure tran returnNeg100 min V(1) FROM=0.2e-3 TO=0.25e-3 TD=0.5e-3 default_val=-100

* add tests for rise/fall/cross.  VS2 and VS3 have a DC offset
* and are damped sinusoids
.measure tran minv3fall2 min v(3) fall=2
.measure tran minv4rise1 min v(4) rise=1
.measure tran minv3cross3 min v(3) cross=3

* test LAST for rise/fall/cross
.measure tran minv3falllast min v(3) fall=last
.measure tran minv4riselast min v(4) rise=last
.measure tran minv3crosslast min v(3) cross=last
.measure tran minv4crosslast min v(4) cross=last

*test RFC_LEVEL keyword
.measure tran minv1Rise1RFClevel50 min V(1) RFC_LEVEL=0.5 RISE=1
.measure tran minv1Fall1RFClevel50 min V(1) RFC_LEVEL=0.5 FALL=1
.measure tran minv1Cross1RFClevel50 min V(1) RFC_LEVEL=0.5 CROSS=1 

*test Failed measures for rise/fall/cross
.measure tran minv3fallfail min v(3) fall=10
.measure tran minv4risefail min v(4) rise=10
.measure tran minv3crossfail min v(3) cross=10

.END

