test errors for measure types that are not supported for DC_CONT
**********************************************************************
* Only the DERIV-AT, DERIV-WHEN, FIND-AT, FIND-WHEN, WHEN,
* TRIG and TARG  measure types are supported for DC_CONT
* mode for .MEASURE.  This tests the error messages from the
* other valid types, that aren't supported for DC_CONT.
*
* The netlist and .DC print/analysis statements in this netlist
* don't really matter.
*
*******************************************************************
vsrc1   1a 0 1
rload1a 1a 1b 0.1
rload1b 1b 0 1
.DC vsrc1 1 5 1

* Note: vsrc1:DCV0 is the syntax for printing the DC value of vsrc1,
* at it is swept.
.print dc vsrc1:DCV0 v(1a) v(1b)

* These measure types are not supported for DC_CONT mode. The exact syntax
* of each measure line doesn't matter.  Just that it has dc as the
* second word.
.measure dc_cont avgVal avg V(1)
.measure dc_cont dutyVal duty V(1)
.measure dc_cont eqnVal EQN {V(1)+10}
.measure dc_cont err1Val ERR1 v(1a) v(1b)
.measure dc_cont err2Val ERR2 v(1a) v(1b)
.measure dc_cont errorVal ERROR v(1b) file=bogo.prn comp_function=infnorm indepvarcol=2 depvarcol=3
.measure dc_cont fourfail FOUR V(1) AT=1e6 TD=2e-3
.measure dc_cont freqVal FREQ v(1) ON=0.75 OFF=0.25
.measure dc_cont integVal integ V(1)
.measure dc_cont offVal off_time V(1) OFF=0
.measure dc_cont onVal on_time V(1) ON=0
.measure dc_cont maxVal max V(1)
.measure dc_cont minVal min V(1)
.measure dc_cont ppVal pp V(1)
.measure dc_cont rmsVal rms V(1)

.END
