* test the TABLE form of the G-Source

*COMP v(node1) OFFSET=.0
*COMP v(node2) OFFSET=3.0

.TRAN 0 1us
.PRINT TRAN V(node1) V(node2)
R1         node2 0  1
G1         node2 0 TABLE V(node1,0) = (-1,-3) (1,3)
V1         node1 0 SIN(0V 0.75V 1e6 0 0 0)
