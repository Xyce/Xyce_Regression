* Test AC mode support for the AC_CONT version of
* DERIV-AT and DERIV-WHEN measures.
*
* See SON Bugs 1274, 1304 and 1313 for more details
*****************************************************

* Used to adjust reference frequency from 1Hz to 10Hz
.PARAM scaleFactor=10

V1 a 0 DC 0V AC 1

* 7th order Chebychev LPF with 2dB of passband ripple.
* This is not a realistic passbad ripple level, but is
* useful for this test.
RS a b 1
C1 b 0 {2.865/scaleFactor}
L2 b c {0.912/scaleFactor}
C3 c 0 {3.8774/scaleFactor}
L4 c d {0.9537/scaleFactor}
C5 d 0 {3.8774/scaleFactor}
L6 d e {0.912/scaleFactor}
C7 e 0 {2.8650/scaleFactor}

* The magnitude at DC is RL/(RL + RS)
RL e 0 1.0

.ac dec 20 1e-2 10
.print AC vm(a) vm(b) vm(c) vm(d) vm(e)
+ derivCrossContTest2 derivCrossContTest3 derivCrossContTest4
+ derivCrossNeg2 derivCrossContNeg2 derivCrossNeg6 derivCrossContNeg6

* The non-continuous version should return the first crossing.
* The continuous version should return all crossings.
.MEASURE AC derivCrossTest1 DERIV vm(d) WHEN vm(e)=0.45
.MEASURE AC_CONT derivCrossContTest1 DERIVATIVE vm(d) WHEN vm(e)=0.45

* Non-continuous version should return first crossing.
* Continuous version should return all crossings, starting
* with the first one.
.MEASURE AC derivCrossTest2 DERIV vm(d) WHEN vm(e)=0.45 CROSS=1
.MEASURE AC_CONT derivCrossContTest2 DERIV vm(d) WHEN vm(e)=0.45 CROSS=1

* Non-continuous version should return second crossing.
* Continuous version should return all crossings, starting
* with the second one.
.MEASURE AC derivCrossTest3 DERIV vm(d) WHEN vm(e)=0.45 CROSS=2
.MEASURE AC_CONT derivCrossContTest3 DERIV vm(d) WHEN vm(e)=0.45 CROSS=2

* These should both return the last crossing
.MEASURE AC derivCrossTest4 DERIV vm(d)  WHEN VM(e)=0.45 CROSS=LAST
.MEASURE AC_CONT derivCrossContTest4 DERIV vm(d) WHEN VM(e)=0.45 CROSS=LAST

* DERIV-AT measures
* These should give the same answer
.MEASURE AC atTest DERIV VM(e) AT=2
.MEASURE AC_CONT atContTest DERIV VM(e) AT=2

*****************************************************
* test RISE and FAll qualifiers for DERIV-WHEN
.MEASURE AC_CONT derivRiseContTest1 DERIV VM(d) WHEN VM(e)=0.45 RISE=1
.MEASURE AC_CONT derivRiseContTest2 DERIV VM(d) WHEN VM(e)=0.45 RISE=2
.MEASURE AC_CONT derivRiseContTest3 DERIV VM(d) WHEN VM(e)=0.45 RISE=LAST

.MEASURE AC_CONT derivFallContTest1 DERIV VM(d) WHEN VM(e)=0.45 FALL=1
.MEASURE AC_CONT derivFallContTest2 DERIV VM(d) WHEN VM(e)=0.45 FALL=2
.MEASURE AC_CONT derivFallContTest3 DERIV VM(d) WHEN VM(e)=0.45 FALL=LAST

************************************************************************
* Use of FROM-TO.  Only the rise, fall or cross values within the
* FROM-TO windows should be returned, starting at the requested value.
* For CROSS=LAST, only the last one within the FROM-TO window is returned
.MEASURE AC_CONT derivCross1ContFrom DERIV VM(d) WHEN VM(e)=0.45 CROSS=1 FROM=0.5
.MEASURE AC_CONT derivCross2ContFrom DERIV VM(d) WHEN VM(e)=0.45 CROSS=2 FROM=0.5
.MEASURE AC_CONT derivCrossContTo DERIV VM(d) WHEN VM(e)=0.45 CROSS=1 TO=1
.MEASURE AC_CONT derivRiseContTo DERIV VM(d) WHEN VM(e)=0.45 RISE=1 TO=1
.MEASURE AC_CONT derivFallContFrom DERIV VM(d) WHEN VM(e)=0.45 FALL=1 FROM=0.5
.MEASURE AC_CONT derivCrossContToLast DERIV VM(d) WHEN VM(e)=0.45 CROSS=LAST TO=1

*********************************************************
* Test negative values
.MEASURE AC derivCrossNeg2 DERIV VM(d) WHEN VM(e)=0.45 CROSS=-2
.MEASURE AC derivCrossNeg3 DERIV VM(d) WHEN VM(e)=0.45 CROSS=-3
.MEASURE AC derivCrossNeg6 DERIV VM(d) WHEN VM(e)=0.45 CROSS=-6
.MEASURE AC_CONT derivCrossContNeg1 DERIV VM(d) WHEN VM(e)=0.45 CROSS=-1
.MEASURE AC_CONT derivCrossContNeg2 DERIV VM(d) WHEN VM(e)=0.45 CROSS=-2
.MEASURE AC_CONT derivCrossContNeg3 DERIV VM(d) WHEN VM(e)=0.45 CROSS=-3
.MEASURE AC_CONT derivCrossContNeg6 DERIV VM(d) WHEN VM(e)=0.45 CROSS=-6

.MEASURE AC derivRiseNeg2 DERIV VM(d) WHEN VM(e)=0.45 RISE=-2
.MEASURE AC derivRiseNeg3 DERIV VM(d) WHEN VM(e)=0.45 RISE=-3
.MEASURE AC_CONT derivRiseContNeg1 DERIV VM(d) WHEN VM(e)=0.45 RISE=-1
.MEASURE AC_CONT derivRiseContNeg2 DERIV VM(d) WHEN VM(e)=0.45 RISE=-2
.MEASURE AC_CONT derivRiseContNeg3 DERIV VM(d) WHEN VM(e)=0.45 RISE=-3

.MEASURE AC derivFallNeg2 DERIV VM(d) WHEN VM(e)=0.45 FALL=-2
.MEASURE AC derivFallNeg4 DERIV VM(d) WHEN VM(e)=0.45 FALL=-4
.MEASURE AC_CONT derivFallContNeg1 DERIV VM(d) WHEN VM(e)=0.45 FALL=-1
.MEASURE AC_CONT derivFallContNeg2 DERIV VM(d) WHEN VM(e)=0.45 FALL=-2
.MEASURE AC_CONT derivFallContNeg4 DERIV VM(d) WHEN VM(e)=0.45 FALL=-4

*************************************************
* test failed measures
.MEASURE AC_CONT derivCrossContFail1 DERIV VM(b) WHEN VM(e)=1
.MEASURE AC_CONT atContFail DERIV VM(b) at=200
.MEASURE AC_CONT derivCrossContFail2 DERIV VM(b) WHEN VM(e)=0.45 CROSS=6
.MEASURE AC_CONT derivRiseContFail DERIV VM(b) WHEN VM(e)=0.45 RISE=4
.MEASURE AC_CONT derivFallContFail DERIV VM(b) WHEN VM(e)=0.45 FALL=4

.END
