* DC simulation for xyce
.options device temp=27
.subckt mysub c_x b_x e_x s_x
e_c c_v 0 c_x 0 -1
v_c c_v c 0
f_c c_x 0 v_c   1
e_b b_v 0 b_x 0 -1
v_b b_v b 0
f_b b_x 0 v_b   1
e_e e_v 0 e_x 0 -1
v_e e_v e 0
f_e e_x 0 v_e   1
e_s s_v 0 s_x 0 -1
v_s s_v s 0
f_s s_x 0 v_s   1
q1 c b e s mymodel
+ sw_et=0
.model mymodel pnp level=12
+ IS=1e-16
+ IBEI=1e-18
+ IBEN=5e-15
+ IBCI=2e-17
+ IBCN=5e-15
+ ISP=1e-15
+ RCX=10
+ RCI=60
+ RBX=10
+ RBI=40
+ RE=2
+ RS=20
+ RBP=40
+ VEF=10
+ VER=4
+ IKF=2e-3
+ ITF=8e-2
+ XTF=20
+ IKR=2e-4
+ IKP=2e-4
+ CJE=1e-13
+ CJC=2e-14
+ CJEP=1e-13
+ CJCP=4e-13
+ VO=2
+ GAMM=2e-11
+ HRCF=2
+ QCO=1e-12
+ AVC1=2
+ AVC2=15
+ TF=10e-12
+ TR=100e-12
+ TD=1.0e-20
+ RTH=300
+ GMIN=0.0
.ends
v_c c 0 -0.05
v_b b 0 1.00
v_e e 0 0
v_s s 0 0
x1 c b e s mysub
.dc v_c 0.00 5.00 0.05
.step v_b list 0.70 0.75 0.80 0.85 0.90 0.95 1.00
.print dc V(c) V(b)
+ i(v_c)
+ i(v_b)
+ i(v_s)
.end
