************************************************
* Test .DATA and its use with .MEASURE and 
* -remeasure for .DC.
*
* See SON Bug 1160 for more details.
************************************************

VT1 4 0 10V
R1  4 5 10
R2  5 0 5

.data test
+ r1   r2  
+ 8.0000e+00  4.0000e+00 
+ 9.0000e+00  4.0000e+00 
+ 1.0000e+01  4.0000e+00 
+ 1.1000e+01  4.0000e+00 
+ 1.2000e+01  4.0000e+00 
+ 8.0000e+00  5.0000e+00 
+ 9.0000e+00  5.0000e+00 
+ 1.0000e+01  5.0000e+00 
+ 1.1000e+01  5.0000e+00 
+ 1.2000e+01  5.0000e+00 
+ 8.0000e+00  6.0000e+00 
+ 9.0000e+00  6.0000e+00 
+ 1.0000e+01  6.0000e+00 
+ 1.1000e+01  6.0000e+00 
+ 1.2000e+01  6.0000e+00 
.enddata

.DC data=test

.print DC {R1:R} {R2:R} V(4) V(5)
.MEASURE DC MAXV4 MAX V(5)

.END

