***********************************************************************
* DC remeasure assumes that the remeasured .prn file has an 
* Index column.  It should produce a fatal netlist error if 
* there isn't one.
*
* See SON Bug 885 for more details.
***********************************************************************

vsrc1   1a 0 1
rload1a 1a 1b 0.1
rload1b 1b 0 1

.DC vsrc1 1 5 1
.PRINT DC FORMAT=NOINDEX v(1b)

* MAX measure
.measure dc maxv1b  max v(1b)

.end

