A test of re-measure of .CSD formatted output file
*******************************************************************************
* The data portion of a .CSD file (made by Xyce) is formatted as follows.
* The #N line is followed by a list of the data column headers.
* The subsequent #C line has the time value and the number of data points.  
* It is followed by a list of values (0.00000000e+00:1) that may span multiple 
* lines.  The :1 says this is the value for the first data column.
* 
* #N
* 'V(1)' 'V(2)' 'V(3)' 'V(4)' 'V(5)'
* #C 0.00000000e+00 5
* 0.00000000e+00:1   -5.00000000e-01:2   5.00000000e-01:3   0.00000000e+00:4
* 0.00000000e+00:5   
* #C 1.00000000e-05 5
* 6.27773973e-02:1   -4.37569034e-01:2   4.37569034e-01:3   1.25554795e-01:4
* -1.25554795e-01:5   
*
* So, it is important to use a CSD file where the data values span at 
* least two lines
*
* collection of SIN sources
VS1  1  0  SIN(0 1.0 1KHZ 0 0)
VS2  2  0  SIN(-0.5 1.0 1KHZ 0 500)
VS3  3  0  SIN(0.5 -1.0 1KHZ 0 500)
VS4  4  0  SIN(0 2.0 1KHZ 0 0)
VS5  5  0  SIN(0 -2.0 1KHZ 0 0)

R1  1  0  100
R2  2  0  100
R3  3  0  100
R4  4  0  100
R5  5  0  100

.TRAN 0  3ms
.PRINT TRAN FORMAT=PROBE V(1) V(2) V(3) V(4) V(5)

* check re-measure for the first and last data column on the first line
* after each #C, and also for the value on the second line after each #C.
* This should be sufficient.
.measure tran minSineOne min V(1) 
.measure tran minSinFour min V(4)
.measure tran minSinFive min V(5)

* also test that a measure of V(1) works for all measure types, 
* with a reasonable set of syntaxes.  FOUR will be tested
* separately.

* AVG
.measure tran avgVal avg V(1)

*DERIV
.measure tran derivValWhen deriv V(1) WHEN V(1)=0.5
.measure tran derivValAt deriv V(1) AT=5e-04

* DUTY
.measure tran dutyVal duty V(1)

*EQN
.measure tran eqnVal EQN {V(1)+10}

* FIND WHEN
.measure tran whenVal WHEN V(1)=0.5
.measure tran findWhenVal FIND V(2) WHEN V(1)=0.5

*FREQ
.measure tran freqVal FREQ v(1) ON=0.75 OFF=0.25

* INTEG
.measure tran integVal integ V(1)

* MAX
.measure tran maxVal max V(1)

* OFF_TIME
.measure tran offVal off_time V(1) OFF=0

* ON_TIME
.measure tran onVal on_time V(1) ON=0

* PP
.measure tran ppVal pp V(1) 

* RMS
.measure tran rmsVal rms V(1)

*TRIG/TARG (RiseFallDelay)
.measure tran trigTargVal TRIG v(1)=0.1 TARG v(1)=0.99
.measure tran trigTargAt TRIG AT=1e-3 TARG V(4)=1

.END

