module main;
initial $ADCtest;
endmodule
