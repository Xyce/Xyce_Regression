Testing .MEASURE lines that are mismatched with the Analysis Types
*********************************************************************
* This tests the error messages that should occur if a TRAN, TRAN_CONT,
* NOISE, NOISE_CONT, FFT, DC or DC_CONT mode measure is requested for a netlist
* that is doing a .AC analysis.
*
* See SON Bugs 889, 1274 and 1280 for more details.
*
*
*********************************************************************

* Trivial high-pass filter (V-C-R) circuit
R1 b 0 2
C1 a b 1u
V1 a 0 DC 0V AC 1

.print AC v(b) 

.ac dec 5 100Hz 10e6

* Test what happens when a TRAN, TRAN_CONT, DC, DC_CONT, FFT, NOISE or NOISE_CONT
* measure is requested for a .AC netlist
.MEASURE DC dcmax max v(b)
.MEASURE DC_CONT dc_cont_when when vm(b)=0.5
.MEASURE TRAN tranmax max v(b)
.MEASURE TRAN_CONT tran_cont_find find vi(b) when vm(b)=0.5
.MEASURE NOISE noisemax max v(b)
.MEASURE NOISE_CONT noise_cont_find find vi(b) when vm(b)=0.5
.MEASURE FFT THD THD v(b)

.END

