* Test DC mode support for TRIG-TARG Measures
*
* This bug covers:
*   1) the case of one variable in the .DC line,
*      without a .STEP statement. where the swept
*      variable is increasing.
*
*   2) An ascending sweep variable.
*****************************************************

.DC V1 1 10 1
.PRINT DC V(1) V(2) V(3)

V1 1 0 1
R1 1 0 1

B2 2 0 V={(V(1)-2.5)*(V(1)-2.5)*(V(1)-7.5)*(V(1)-7.5)/4}
R2 2 3 1
R3 3 0 1

.MEASURE DC TRIGTARGAT TRIG AT=2.5 TARG AT=7.5
.MEASURE DC TRIGTARGAT1 TRIG AT=2.5 TARG V(2)=5 CROSS=1
.MEASURE DC TRIGTARGAT2 TRIG V(2)=5 CROSS=1 TARG AT=7.5

.MEASURE DC TRIGTARG1 TRIG V(2)=3 CROSS=1 TARG V(2)=7 CROSS=1 
.MEASURE DC TRIGTARG2 TRIG V(2)=3 CROSS=1 TARG V(2)=7 CROSS=2
.MEASURE DC TRIGTARG3 TRIG V(2)=3 CROSS=2 TARG V(2)=7 CROSS=1

* Variables for TRIG and TARG, with and without expressions
.MEASURE DC TRIGTARGVAR TRIG V(2)=V(1) CROSS=1 TARG V(2)=V(1) CROSS=2
.MEASURE DC TRIGTARGVAREXP TRIG {V(2)}={V(1)} CROSS=1 TARG {V(2)}={V(1)} CROSS=2

.END
