* 2-port example. Input uses a default Option line, with just a #
* character on it.  In that case:
*
*   1) the [Network Data] is assumed to S-parameter data in MA format.
*
*   2) the default frequency multiplier is GHz.
*
*   3) No Z0 information is given by the [Reference] line, so a default of
*      50 ohms is assumed for each port.
*
* Note that this netlist does not have the R2 load resistor in it.
* This is because that resistance is already included in the
* S-parameter model used by YLIN_MOD1.

.model diod d

.options hbint numfreq=10 tahb=0
.hb 1e5
.print hb v(1) v(2) i(v1)

v1 1 0  sin  0 5 1e5
YLIN YLIN1 1 0 2 0 YLIN_MOD1
.MODEL YLIN_MOD1 LIN TSTONEFILE=ylin-2port-defaultOptions.cir.s2p
d1  2 0 diod

.end
