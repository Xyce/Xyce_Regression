* Transient sensitivity example, sine source, analytical sensitivity
.param cap=0.1u
.param res=1K

c1 1 0 cap
c2 2 0 cap
R1 1 3 res
R2 1 2 res

Vin 3 0 SIN(0 1 100K -2.5U 0.0 -90.0

* Transient commands
.tran 0 10us uic
.options timeint reltol=1e-6 abstol=1e-6

.print tran v(1) v(2) v(3)

* Sensitivity commands
.print sens 
.SENS objfunc={V(2)} param=Vin:V0,Vin:VA,Vin:FREQ,Vin:TD,Vin:THETA,Vin:PHASE

.options SENSITIVITY direct=1 adjoint=0 forceanalytic=true
.end

