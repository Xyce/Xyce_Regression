Mx  Drain Gate Source Back-gate(substrate) Body  Tx  W  L (body ommitted for FB)
* Modified by Darsen Lu 03/11/2009

* Modified also by Eric R. Keiter 04/30/2010 to use the SOI model version 3.2.
* To get it to work I had to increase the L instance parameter somewhat.

.include ./nmos3p2.mod
.include ./pmos3p2.mod
.option TEMP=27C

Vpower VD 0 1.5
Vgnd VS 0 0

Vgate   Gate   VS PULSE(0v 1.5v 100ps 50ps 50ps 200ps 500ps)

MN0 VS Gate Out VS N1 W=10u L=0.35u
MP0 VD Gate Out VS P1 W=20u L=0.35u

.tran 0.01n 600ps
.print tran v(gate) v(out)
.END
