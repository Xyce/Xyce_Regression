* Test DC mode support for TRIG-TARG measures
*
* This bug covers:
*   1) The case of two variables on the .DC line.  (Note:
*      since there is no .STEP statement, the output is treated
*      like one STEP.)
*
*   2) Have one sweep variable (vsrc1) be monotonically decreasing,
*      while the other (vsrc2) is monotonically increasing
*
* See gitlab-ex issue 289 for more details.
**************************************************************

vsrc1   1a 0 1
rload1a 1a 1b 0.1
rload1b 1b 0 1

vsrc2   2a 0 5
rload2a 2a 2b 0.1
rload2b 2b 1b 0.1

.DC vsrc1 5 1 -1 vsrc2 2 5 3

* Note: vsrc1:DCV0 is the syntax for printing the DC value of vsrc1,
* as it is swept.
.print dc vsrc1:DCV0 vsrc2:DCV0 v(1a) v(2a) v(1b) v(2b)

* This measure should TRIG in the first sweep of vsrc1 and TARG in
* the second sweep of vsrc1.
.MEASURE DC trigtarg1 TRIG V(1b)=3 CROSS=1 TARG V(1b)=3 CROSS=2

* This measure should not find a TRIG and TARG in the second sweep
* of vsrc1.
.MEASURE DC trigtarg2 TRIG V(1b)=3 RISE=1 TARG V(1b)=4 CROSS=1

.end
