* Test AC mode support for the DERIV / DERIVATIVE measure.
* To be conservative, there are subtests for each
* valid operator (V, VR, VI, VP, VM and VDB) for
* each measure type.  Expressions are also tested.
* One current operator (IM) is tested for a branch current.
*
* See SON Bug 1282 for more details.
*****************************************************

* Trivial high-pass filter (V-C-R) circuit
R1 b 0 2
C1 a b 1m
V1 a 0 DC 0V AC 1

.print AC vr(b) vi(b) vm(b) vp(b) vdb(b) im(v1)
.ac dec 5 1Hz 1e3

* AT syntaxes
.MEASURE AC DERIVVMBAT100 DERIV VM(b) AT=100
.MEASURE AC DERIVVMBAT50 DERIVATIVE VM(b) AT=50

.MEASURE AC DERIVVRBAT50 DERIV VR(b) AT=50
.MEASURE AC DERIVVIBAT50 DERIV VI(b) AT=50
.MEASURE AC DERIVVPBAT50 DERIV VP(b) AT=50
.MEASURE AC DERIVVDBBAT50 DERIV VDB(b) AT=50

* Test AT value at start of sweep
.MEASURE AC DERIVVMBAT1 DERIV VM(b) AT=1

* WHEN syntaxes
.MEASURE AC DERIVWHENVMB0.5 DERIV VM(b) WHEN VM(b)=0.5

* Expressions in WHEN clause
.MEASURE AC derivExp1 DERIV VM(b) when vr(b)=vi(b)
.MEASURE AC derivExp2 DERIV VM(b) when {vm(b)+0.1}=0.5
.MEASURE AC derivExp3 DERIV VM(b) when vm(b)={0.3+0.2}
.MEASURE AC derivExp4 DERIV VM(b) when vr(b)={vi(b)+0.3}

* Expression in DERIV clause
.MEASURE AC derivExp5 DERIV {VR(b)+VI(b)} when vm(b)=0.5

* branch current
.MEASURE AC derivimv1at50 deriv im(v1) AT=50

* Tests should return -1 or -100
.measure ac derivRetNeg1 deriv v(b) AT=1e4
.measure ac derivReturnNeg100 deriv vm(b) when vm(b)=2 DEFAULT_VAL=-100

.end
