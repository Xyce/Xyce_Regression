* Transient sensitivity example, SFFM source, FD derivatives
.param cap=0.1u
.param res=1K

.param v0=0.0
.param va=1.0
.param fc=1meg
.param mdi=2.0
.param fs=250k

c1 1 0 cap
c2 2 0 cap
R1 1 3 res
R2 1 2 res

Vin 3 0 SFFM({v0} {va} {fc} {MDI} {fs})

* Transient commands
.tran 0 10us 
.options timeint reltol=1e-6 abstol=1e-6

.print tran v(1) v(2) v(3)

* Sensitivity commands
.print sens 
.SENS objfunc={V(2)} param=V0,VA,FC,MDI,FS
.options SENSITIVITY direct=1 adjoint=0 forcefd=true
.end

