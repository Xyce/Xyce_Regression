* Test the use of .STEP with .FFT when interpolation (fft_accurate=0)
* is used to get the waveform value at the requested sample points.
*
* See SON Bug 1327 for more details.
*********************************************************************

.STEP V1:VA 500 600 100

.TRAN 0 1
.OPTIONS FFT FFT_ACCURATE=0 FFTOUT=1

V1 1 0 SIN(0 500 1)
V3 3 0 SIN(0 200 2)
R1 1 2 1
R2 2 0 1
R3 3 2 1

.FFT V(2) NP=16 WINDOW=HANN FORMAT=UNORM
.PRINT TRAN V(1) V(2) V(3)

.END
