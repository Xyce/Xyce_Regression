A neuron cable example
*
* This is a simple test of simulating a neuron cable
* via the cable equation (6.29 in Theorteical Neuroscience,
* by P. Dayan and L. Abbot)
*
* in this case there will be no ion channel currents, so
* the cable is entirely passive
*

* units for model parameters
* cMem = F/cm^2
* gMem = S/cm^2
* vRest = V
* eNa = V
* gNa = S/cm^2
* eK = V
* gK = S/cm^2
* r  = ohms cm
*
* NOTE: length scale is immaterial as long as it's always a consistent unit
* parameters from Dayan's book pg 173, 157, 155
* cMem  = 1.0 uF/cm^2   =>  1.0e-6 F/cm^2
* gMem  = 0.003 mS/mm^2 =>  0.000003 S/mm^2  => 0.0003 S/cm^2
* vRest = -17 mV        => -0.017 V
*
* cMem  = 10 nF/mm^2    =>  1.0e-8 F/mm^2    => 1.0e-6 F/cm^2 
* r     = 1 kOhm mm     =>  1000 Ohm mm      => 100 Ohm cm 

*.param length = 0.1 ; [cm]
*.param radius = 0.5e-4  ; [cm]
*.param memC = 1.0e-6  ; [uF/cm^2]
*.param restV = -0.065 ; [V]
*.param Rm = 4.0e4 ; [40000 ohms cm^2]
*.param memG = {1.0/Rm}    ; TODO - make sure that's what Rm is for
*.param Ra = 100.0 ; [ohms cm]

.param length = 0.1e-2 ; [m]
.param radius = 0.5e-6  ; [m]
.param memC = 1.0e-2  ; [F/m^2] ok
.param restV = -0.065 ; [V]
.param Rm = 4.0 ; [ohms m^2]
.param memG = {1.0/Rm}    ; TODO - make sure that's what Rm is for
.param Ra = 1.0 ; [ohms m]


.model pcParams neuron level=6
*+ cmem=1.0e-6   gmem=0.0003  vrest=-0.017 n=100
*+  R=1.0e2 A=1.0e-4 L=0.4 
+ cMem = {memC}
+ gMem = {memG}
+ vRest = {restV}

*
* Using the above neuron model
*

* This is a standard current pulse to start an activation
*          pulse( initial_value pulse_value delay_time rise_time fall_time pulse_width period)
Iin 0 a PULSE( 0 1.0e-10 1.0e-12 0.0 0.0 1.0e10 1.0e10)

* the parameters R (intra-cellular resistivity Ohm/cm), A= radius (cm), L = length (cm)
* can be specified in the .model statement or as part of the instance.  Instance level
* parameters override model level ones.  N = number of segments.

* intra cellular resistivity, rl,  is typically 1-3 kOhm mm.  Resistance along the long axis (longitudinal resistance Rl = rl L / (pi a^2)
* 1 kOhm mm = 1000 Ohm mm = 100 Ohm cm 

yneuron neuron1  a b pcParams 
* R=1.0e2 A=1.0e-4 L=0.4 
+ R = {Ra}
+ A = {radius}
+ L = {length}
+ N = 1000

.tran 0 0.25

.options output initial_interval=5.0e-5
.options timeint method=7 newlte=1 newbpstepping=1 reltol=1e-3
.options linsol type=klu
.print tran 
*+ i(iin) 
+ V(a) 
*+ n(y%neuron%neuron1_V1) 
+ V(b)
   



.end


