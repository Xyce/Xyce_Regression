* Unit test of Power Grid Branch Transformer, in I=YV format 

*********************************************
* Bus 1 is the slack bus.  Ammeter          *
* is wired so that current flows into Bus 1 *
*********************************************
V1R Bus1R ammBus1R 1V
V1I Bus1I ammBus1I 0V
Vamm1R 0 ammBus1R 0V
Vamm1I 0 ammBus1I 0V

*********************************************
* Transformer Definition                    *
*********************************************
YPowerGridTransformer pg1_2 bus1R bus2R bus1I bus2I AT=IV R=0.05 X=0.2 TR=0.978

*********************************************
* Load Definitions                          *
*********************************************
XLoad2 bus2R bus2I CPL PARAMS: P=0.9 Q=0.1

*********************************************
* Simulation Control and Output Statements  *
*********************************************
.DC V1R 1 1 1
.PRINT DC width=10 precision=6
+ V(bus1R) V(bus1I) V(bus2R) V(bus2I) 
+ {V(bus1R)*I(Vamm1R)+V(bus1I)*I(Vamm1I)}
+ {V(bus1I)*I(Vamm1R)-V(bus1R)*I(Vamm1I)}
+ {V(bus2R)*I(Xload2:VammR)+V(bus2I)*I(Xload2:VammI)}
+ {V(bus2I)*I(Xload2:VammR)-V(bus2R)*I(Xload2:VammI)}

**************************************************************
* Subcircuit defintion of a constant power load for I=YV form*
**************************************************************
.SUBCKT CPL RNode INode PARAMS: P=0.5 Q=0.0 CurrLim=1000

* Ammeter at load is defined so that power flows into the load from the bus
VammR ammR 0 0V
VammI ammI 0 0V
BloadR RNode ammR I={limit((P*V(RNode)+Q*V(INode))/(V(RNode)*V(RNode)+V(INode)*V(INode)),
+ -CurrLim,CurrLim)}
BloadI INode ammI  I={limit((P*V(INode)-Q*V(RNode))/(V(RNode)*V(RNode)+V(INode)*V(INode)),
+ -CurrLim,CurrLim)}

.ENDS

.end
