Test Circuit for the Arcsine and Arccosine Functions
*******************************************************************************
* Tier No.:     1			
* Directory/Circuit Name: ABM_ACOS_ASIN/acos_asin.cir
* Description:  Test of analog behavioral modeling arcsine and arccosine 
*	functions.								
* Input: V1								
* Output: V(1), V(2), V(3)					
* Analysis:						
*	The netlist contains an independent voltage source, V1 or V(1),  that is swept from
*	-0.99V to 0.99V in 0.01V steps.  Two nonlinear dependent voltage sources are 	
*	used to define the functions as follows:				
*		V(2)=B2=ASIN(V(1)) = inverse sine of V(1)		
*		V(3)=B3=ACOS(V(1)) = inverse cosine of V(1)	
*	A DC analysis is performed and the output recorded is voltages defined by the
*	arccosine and arcsine functions.					
*									
*	This table is a set of hand calculations for the functions of ACOS and ASIN of X
*	          X	       ACOS(X)		        ASIN(X) 		
*		-1.0		3.14			-1.570	
*		-0.5		2.09			-0.524
*		 0.0		1.57		  	 0.000	
*		 0.5		1.05			 0.524
*		 1.0		0.00			 1.570
*******************************************************************************
V1  1  0  0
R1  1  0  1
B2  2  0  V = {ASIN(V(1))}
R2  2  0  1
B3  3  0  V = {ACOS(V(1))}
R3  3  0  1
.DC V1 -0.99 0.99 0.01
.PRINT DC V(1) V(2) V(3) 
.END
