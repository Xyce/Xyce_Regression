* The contents of this netlist doesn't really matter
V1 1 0 1
R1 1 0 1
.DC V1 1 2 1
.PRINT DC V(1)
.END
