Resistor Circuit Netlist - top level

VIN1 1 0 DC 0V
VIN2 2 0 DC 0V

YEXT y1 1 2 externcode=xyce netlist=capInner.cir

.print tran v(1) 
.tran 0 1ms

.options nonlin maxstep=10 nox=1
.options timeint reltol=1e-6 abstol=1e-6
*
.END
