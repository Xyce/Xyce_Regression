DTEMP Test circuit for P-Channel JFET 
***********************************
*Drain curves
vds 1 0 0
vgs 2 0 0
*
vidmon 1 1a 0
vigmon 2 2a 0
vismon 0 3 0
*
.dc vgs 0 1.5 0.5 vds -15 0 1
.print dc v(1) v(2) i(vidmon)
.step tempParam list 15 25 35
*
.param tempParam=10
ztest 1a 2a 3 sa2108 temp={tempParam}
*
.model sa2108 pmf
+ level=1 beta= 0.000278
+ vto = -2.10
+ pb = 0.265
+ lambda = 0.0055
+ b = 0.590;
+ rd = 302.5
+ rs = 0.0
+ fc = 0.5
+ is = 1.393e-10
+ af = 1.0
+ kf = 0.05
+ cgs= 0
+ cgd= 0
*
.end

