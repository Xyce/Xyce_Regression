* Test FOUR measure with .STEP.  Also test PRECISION qualifier for
* FOUR measure.

* Jfet Transient Sine wave 6 volt input signal to output 

Vdd   Vdd     0       DC 20
*                          SIN(Voffset Vamplitude Frequency)
*                          ---------------------------------
V1    Vin     0       DC 0 SIN(0       6        1e6)
Rload Vout    0       1Meg
Xamp1 Vin Vdd 0 Vout  amp2n3819
*
*     STEP STOP
*     TIME TIME
*     ---- ---
.TRAN 1e-8 1e-6 

.STEP V1:freq 1e6 2e6 1e6 

.PRINT TRAN V(Vin) V(Vout)

.MEASURE TRAN fourVP FOUR V(Vout) AT=1e6 PRECISION=7
.MEASURE TRAN LASTMEASURE MAX V(Vout) PRECISION=7

* Amplifier subcircuit

.subckt amp2n3819 Vin Vdd Vss Vout
Rd  Vdd     Vout           1462
J1  Vout    Vin    Nsource J2N3819
Rs  Nsource Vss            188
Rg  Vin     Vss            1Meg
*
.model J2N3819 NJF(Beta=1.304m Rd=1 Rs=1 Lambda=2.25m Vto=-3
+ Is=33.57f Cgd=1.6p Pb=1 Fc=.5 Cgs=2.414p Kf=9.882E-18 Af=1)
*
.ENDS

.END

 
