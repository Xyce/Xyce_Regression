Regression test for simple normal distribution sampling

Isrc 1 0 AC 1 0 sin(0 1 1e+5 0 0)
R1 1 0 1e3
C1 1 0 2e-6

.print ac v(1)
.ac dec 10 1 1e5

.EMBEDDEDSAMPLING 
+ param=R1
+ type=normal
+ means=1K
+ std_deviations=0.2K

.options EMBEDDEDSAMPLES numsamples=10

.end

