simple RC

.options nonlin continuation=1

.options loca stepper=natural predictor=constant stepcontrol=1 conparam=GSTEPPING
+ initialvalue=4 minvalue=-4 maxvalue=4 initialstepsize=-2 minstepsize=1e-6 maxstepsize=1e12
+ aggressiveness=0.01 residualconductance=1e-10 maxsteps=200 maxnliters=20 voltagelist=DOFS

.tran   0    50e-5

.print tran  v(1) v(2)   v(3)

v1 1 0 1

r1 1 2 1k
c1 2 3 2u

c2 3 0 1u

r2 3 5 1k
.end
