****************************************************************
* A simple test of a fourier transform using I(), P(), W() and
* expressions when I() is not on the .PRINT TRAN line.
* The Fourier transform of I(R1) should be a tone with magnitude
* 2 at 1 HZ.  The Fourier transform of P(R1) and W(R1) should 
* have tones at DC and 2 HZ with magnitude of 2.  Etc.
*
*
****************************************************************
V1 1 0 SIN(0 2 1)
R1 1 0 1

V2 2 0 SIN(0 1 2)
R2 2 0 1

V3 3 0 SIN(0 1 3)
R3 3 0 1

V4 4 0 SIN(0 2 3)
R4 4 0 1

V5 5 0 SIN(0 1 4)
R5 5 0 1

V6 6 0 SIN(0 2 4)
R6 6 0 1

V7 7 0 SIN(0 1 5)
R7 7 0 1

V8 8 0 SIN(0 2 5)
R8 8 0 1

.TRAN 10ms 1 
.PRINT TRAN V(1) I(V1)
.OPTIONS OUTPUT INITIAL_INTERVAL=0.01

* These lines test that .FOUR works even if the I(), P()
* or W() is not on the .PRINT TRAN line.  See SON Bug 703.
.four 1 I(R1) P(R1) W(R1)
.four 2 I(R2) P(R2) W(R2)

* Make sure that multiple lead current requests can be 
* parsed out of an expression.
.four 3 {I(R4) - I(R3)}
.four 4 {P(R6) - P(R5)}
.four 5 {W(R8) - W(R7)}

* used to make sure that lead current requests work if they
* come from a combo of .PRINT TRAN, .FOUR and .MEASURE lines
.MEASURE TRAN MAXIV1 max I(V1) 
.MEASURE TRAN MAXIV2 max I(V2)

.end
