test of table, without "file" suffix.  Also, using data file that is not in order.

b1 1 0 v={table("sinewaveOutOfOrder.dat")}
r1 1 0 500
.tran 1us 10us

*COMP V(1) OFFSET=6
.print tran v(1)

.end
