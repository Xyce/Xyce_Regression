NOISE test of -r output format with .OP
*
V1  1 0 DC 5.0 AC  1.0   
R1  1 0 100K

* For testing SON Bug 1026, the .NOISE statement
* precedes the .OP statement.
.NOISE  V(1) V1  DEC  5 100 100K 1
.OP
.PRINT NOISE INOISE ONOISE

.END

