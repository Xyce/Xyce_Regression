*******************************************************************
* This netlist is used, along with the netlist hb-files.cir,
* to test SON Bugs 941 and 1011.  This netlist:
*
*  1) should produce the same .HB.FD.prn file as the 
*     netlist hb-files.cir.
*
*  2) should NOT produce the hb-files-fd.startup.prn and 
*     hb-files-fd.hb_ic.prn output files since .PRINT HB_FD 
*     no longer produces "fallback" print lines, as of Xyce 6.10.
*
*   3) should not produce the hb-files-fd.HB.TD.prn file, per
*      the fix for SON Bug 1011
*
* The netlist hb-files.cir should produce all four output files. 
*   
*******************************************************************

* Qucs 0.0.19  /users/russo/src/qucs/examples/xyce/hb-test.sch
D1 Node3 0 DMOD_D1 AREA=1.0 Temp=26.85
.MODEL DMOD_D1 D (LEVEL = 2 Is=1e-15 N=1 Cj0=0 M=0.5 Vj=0.7 Fc=0.5 Rs=0 Tt=0 Ikf=0 Kf=0 Af=1 Bv=0.7 Ibv=0.001 Xti=3 Eg=1.11 Tbv1=0 Trs1=0 Tnom=26.85 )

R1 Node1 _net0  100
R2 _net1 Node3  100
VPr2 _net0 _net1 DC 0 AC 0
EPr1 Pr1 0 Node3 0 1.0
V1 Node1 0 DC 0 SIN(0 4 1MEG 0 0) AC 4

.options hbint numfreq=17 STARTUPPERIODS=2 saveicdata=1

.HB 1MEG

.PRINT HB_FD I(VPr2) v(Node3) v(Pr1) 

.END
