* This test will use an absolute path to a file in
* subdirectory two levels down.

.DC V1 1 5 1
.PRINT DC V(1) V(2)

V1 1 0 1
R1 1 2 1

* The absolute path for the file on this line will be
* filled in by the .sh file.
.INC

.END
