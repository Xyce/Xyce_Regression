* The bug this is intended to test, bug 204, was one in which any netlist
* with a ".DC" analysis line, which lacked a 3rd parameter to indicate the step
* size, would fail by going into an infinite loop.
*
* This circuit tests it by having such a .DC statement.  This is the
* "diode" circuit from the test suite, but with the .DC analysis statement
* changed to set up the bug.  Xyce should take this in stride now.

VIN 1 0 DC 5V
R1 1 2 2K
D1 3 0 DMOD
VMON 2 3 0
.MODEL DMOD D (IS=100FA)
.DC VIN 5 5
.PRINT DC V(1) I(VMON) V(3)
*
.END
