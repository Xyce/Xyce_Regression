* Test NOISE mode support for the INTEG measure. It was deemed sufficient
* to mostly just test with the VR and VI operators.  Expressions
* are also tested. One current operator (IM) is tested for a branch
* current.
*
* See SON Bug 1301 for more details.
********************************************************************

* RESISTOR DIVIDER
V1  1 0 DC 5.0 AC  1.0
R1  1 2 100K
R2  2 0 100K
*
* AMP AND LP FILTER
EAMP  3 0 2 0 1
RLP1  3 4 100
CLP1  4 0 1.59NF

.NOISE  V(4)  V1  DEC  5 1 1e3 1
.PRINT NOISE VR(4) VI(4) IM(EAMP) integvr4 INOISE ONOISE

* RMS
.MEASURE NOISE integvr4 INTEG vr(4)
.meas    noise integralvi4 integral vi(4)

* Use expression
.MEASURE NOISE integvr4Exp integ {1+vr(4)}

* add FROM-TO
.MEASURE NOISE integvr4FromTo integ vr(4) FROM=1e1 TO=1e2

* branch current
.MEASURE NOISE integimeamp integ IM(EAMP)

* FROM=TO value yields a value of 0, by definition
* for INTEG measure.
.MEASURE NOISE integvm4FromTo1Pt integ vm(4) FROM=1e2 TO=1e2

* Tests should return -1 or -100, since the FROM-T0 window
* has various problems.
.measure noise integReturnNegOne integ v(4) FROM=1e4 TO=1e5
.measure noise integReturnNeg100 integ vr(4) FROM=1e3 TO=1e0 DEFAULT_VAL=-100

.END
