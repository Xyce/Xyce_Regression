N-Channel Mosfet Circuit
**************************************************************
*
* Full Newton version of the nmos1.cir circuit.
*
VDD 5 0 DC 5V
R1 5 1 47MEG
R2 1 0 22MEG
RD 5 4 2.2K
RS 2 0 500
VMON 4 3 0
YPDE NMOSB 3 2 1 4 NFET sgplotLevel=0 tecplotLevel=0
+ mobmodel=carr
+ nx=81 l=1.0e-3
+ ny=41 w=5.0e-4
+ node = { name  =   source,     gate,   drain,     sub
+          start =      0.0,   3.0e-4,  8.0e-4,     0.0
+            end =   2.0e-4,   7.0e-4,  1.0e-3,  1.0e-3
+           side =      top,      top,     top,  bottom
+       material =   neutral, neutral, neutral, neutral
+ oxideBndryFlag =         0,       0,       0,       0}
*
.MODEL NFET ZOD level=2

* Nonlinear solver params:
.options NONLIN maxstep=40 maxsearchstep=2 searchmethod=0 nox=0 debuglevel=-100

* Time integration params:
.options DEVICE debuglevel=-100 

* Linear solver params:
.options LINSOL type=klu

*.DC VDD 0 5 0.5 
.DC VDD 0 3 0.5 
*.print DC I(VMON) V(3,2) V(1,2)
.print DC V(5) {abs(I(VMON))}
.END

