****************************************************
* This test uses SPARCALC=0 on the .LIN line.
* So it should do an AC analysis rather than an
* S-Parameter analysis.
****************************************************

* RC ladder circuit
P1 1  0  port=1  z0=50 AC 1

C1 2 0 1e-2
Rgs 1 2 0.02

.subckt RCBlock IN OUT GND
R1 IN OUT 20
C1 IN OUT 1p
Cg1 OUT GND 1p
.ends

X1 2 3 0 RCBlock
X2 3 4 0 RCBlock
X3 4 5 0 RCBlock
X4 5 6 0 RCBlock
X5 6 7 0 RCBlock
X6 7 8 0 RCBlock
X7 8 9 0 RCBlock
X8 9 10 0 RCBlock
X9 10 11 0 RCBlock
X10 11 12 0 RCBlock

.AC DEC 10 10  1e5
.PRINT AC VM(1) VM(2)
.LIN SPARCALC=0

.END
