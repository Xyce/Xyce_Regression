*******************************************************************************
* This netlist is equivalent to Step 2 for the FindWhenTest.cir netlist.
* It has VS1:VA=1 and VS4:V0=-0.5
*
*******************************************************************************
*
* a few sources of different types
VS1  1  0  SIN(0 1.0 1KHZ 0 0)
VP2  2  0  PULSE( 0 100 0.2ms 0.2ms 0.2ms 1ms 2ms )
VS3  3  0  SIN(0 -1.0 1KHZ 0 0)
VS4  4  0  SIN(-0.5 1.0 1KHZ 0 0.5)
VS5  5  0  SIN(0.5 -1.0 1KHZ 0 0.5)


R1  1  0  100
R2  2  0  100
R3  3  0  100
R4  4  0  100
R5  5  0  100

.TRAN 0  5ms 0 1.0e-5
.PRINT TRAN FORMAT=NOINDEX V(1) V(2) V(3) V(4) V(5)

* WHEN measures
.measure tran hit1_75 when v(1)=0.75 MINVAL=0.02
.measure tran hit2_75 when v(1)=0.75 MINVAL=0.08 RISE=2
.measure tran riseLast_minus75 when v(1)=-0.75 RISE=LAST
.measure tran riseLast_75 when v(1)=0.75 RISE=LAST
.measure tran hit1_75_ft when v(1)=0.75 FROM=0.002 TO=0.006
.measure tran hit1_75_td when v(1)=0.75 TD=0.004

.measure tran cross1_90 WHEN V(1)=0.9 cross=1
.measure tran cross4_90 WHEN V(1)=0.9 CROSS=4
.measure tran cross4_90_wtd WHEN V(1)=0.9 Cross=4 TD=0.001
.measure tran crossLast_90 WHEN V(1)=0.9 CROSS=LAST

.measure tran fall1_80 WHEN V(1)=0.8 fall=1
.measure tran fall4_80 WHEN V(1)=0.8 FALL=4
.measure tran fall4_80_wtd WHEN V(1)=0.8 Fall=4 TD=0.001
.measure tran fallLast_80 WHEN V(1)=0.8 fall=LAST

* FIND-WHEN measures
.measure tran find3hit1_75 find v(3) when v(1)=0.75 MINVAL=0.02
.measure tran find3rise2_75 FIND v(3) When v(1)=0.75 RISE=2
.measure tran find3riseLast_minus75 find v(3) when v(1)=-0.75 RISE=LAST
.measure tran riseFindWhenLast_75 find v(3) when v(1)=0.75 RISE=LAST
.measure tran find3hit1_75_ft find v(3) when v(1)=0.75 FROM=0.002 TO=0.006
.measure tran find3hit1_75_td find v(3) when v(1)=0.75 TD=0.004

.measure tran find3cross1_90 find v(3) WHEN V(1)=0.9 cross=1
.measure tran find3cross4_90 find v(3) WHEN V(1)=0.9 CROSS=4
.measure tran find3cross4_90_wtd find v(3) WHEN V(1)=0.9 Cross=4 TD=0.001
.measure tran find3crossLast_90 find v(3) WHEN V(1)=0.9 CROSS=LAST

.measure tran find3fall1_80 find v(3) WHEN V(1)=0.8 fall=1
.measure tran find3fall4_80 find v(3) WHEN V(1)=0.8 FALL=4
.measure tran find3fall4_80_wtd find v(3) WHEN V(1)=0.8 Fall=4 TD=0.001
.measure tran find3fallLast_80 find v(3) WHEN V(1)=0.8 fall=LAST

* add tests for rise/fall/cross.  VS4 and VS5 have a DC offset
* and are damped sinusoids
.measure tran v4fall2 when v(4)=0.25 fall=2
.measure tran v5rise1 when v(5)=0.25 rise=1
.measure tran v4cross2 when v(4)=0.25 cross=2

* test LAST for rise/fall/cross
.measure tran v4falllast when v(4)=0.25 fall=last
.measure tran v5riselast when v(5)=0.25 rise=last
.measure tran v4crosslast when v(4)=0.25 cross=last
.measure tran findv1_v4falllast find v(1) when v(4)=0.25 fall=last
.measure tran findv1_v5riselast find v(1) when v(5)=0.25 rise=last
.measure tran findv1_v4crosslast find v(1) when v(4)=0.25 cross=last

* test RFC_LEVEL keyword
.measure tran v4Rise2RFClevel20 when v(4)=0.1 RFC_LEVEL=0.2 RISE=2
.measure tran v4Fall2RFClevel20 when v(4)=0.1 RFC_LEVEL=0.2 FALL=2
.measure tran v4Cross2RFClevel20 when v(4)=0.1 RFC_LEVEL=0.2 CROSS=2

*test Failed measures for rise/fall/cross
.measure tran v4fallfail when v(4)=0 fall=250
.measure tran v5risefail when v(5)=0 rise=250
.measure tran v4crossfail when v(4)=0 cross=250

.END

