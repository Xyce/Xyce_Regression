A neuron cable example
*
* This is a simple test of simulating a neuron cable
* via the cable equation (6.29 in Theorteical Neuroscience,
* by P. Dayan and L. Abbot)
*

.options device debuglevel=2

* units for model parameters
* cMem = F/cm^2
* gMem = S/cm^2
* vRest = V
* eNa = V
* gNa = S/cm^2
* eK = V
* gK = S/cm^2
* r  = ohms cm
*
* NOTE: length scale is immaterial as long as it's always a consistent unit
* parameters from Dayan's book pg 173, 157, 155
* cMem  = 1.0 uF/cm^2   =>  1.0e-6 F/cm^2
* gMem  = 0.003 mS/mm^2 =>  0.000003 S/mm^2  => 0.0003 S/cm^2
* vRest = -17 mV        => -0.017 V
*
* cMem  = 10 nF/mm^2    =>  1.0e-8 F/mm^2    => 1.0e-6 F/cm^2 
* r     = 1 kOhm mm     =>  1000 Ohm mm      => 100 Ohm cm 
*
* gk    = 0.36 mS/mm^2  => 0.00036 S/mm^2    => 0.036 S/cm^2
* ek    = -77mV         => -0.077 V
* gna   = 1.2 mS/mm^2   => 0.0012 S/mm^2     => 0.12 S/cm^2
* ena   = 50 mV         => 0.050 V

.model udParams neuron level=6 ionchannelmodel=UD
+ cmem=1.0e-6   gmem=0.0003  vrest=-0.017
* Contribution to membrane current
+ MM_CURRENT={{gk * n**4 *(V-ek) + gna * m**3 * h * (V-ena)}}     
* Independent variables for ion channel equations
+ MM_INDVARS={{n}, {m}, {h}}
* Independent variables: F equations
*+ MM_INDFEQUS={ {an(V) * (1-n) + bn(V) * n}, {am(V) * (1-m) + bm(V) * m}, {ah(V) * (1-h) + bh(V) * h}}    
+ MM_INDFEQUS={ {an(V+0.017) * (1-n) + bn(V+0.017) * n}, {am(V+0.017) * (1-m) + bm(V+0.017) * m}, {ah(V+0.017) * (1-h) + bh(V+0.017) * h}}    
* Independent variables: Q equations
+ MM_INDQEQUS={{-n}, {-m}, {-h}}
* additional functions for membrane model
+ MM_FUNCTIONS={{an(V)},{1000*(0.01*(1000*V+55)/(1-exp(-0.1*(1000*V+55))))}, {bn(V)},{1000*(0.125*exp(-0.0125*(1000*V+65)))},
+               {am(V)},{1000*(0.1 *(1000*V+40)/(1-exp(-0.1*(1000*V+40))))}, {bm(V)},{1000*(4*exp(-0.0556*(1000*V+65)))},
+               {ah(V)},{1000*(0.07*exp(-0.05*(1000*V+65)))}, {bh(V)},{1000*(1/(1+exp(-0.1*(1000*V+35))))}}    
* additional parameters for membrane model
+ MM_PARAMETERS={{gk},{0.036}, {ek},{-0.077}, {gna},{0.12}, {ena},{0.050}}  




*
* Using the above neuron model
*

* This is a standard current pulse to start an activation
*          pulse( initial_value pulse_value delay_time rise_time fall_time pulse_width period)
Iin a 0 PULSE( 0 0.40e-7 1.0e-3 1.0e-6 1.0e-6 1.0e-5 1.0e10)
*Vin a 0 PULSE( 0 0.100 1.0e-3 1.0e-5 1.0e-5 1.0e-4 1.0e10)

* the parameters R (intra-cellular resistivity Ohm/cm), A= radius (cm), L = length (cm)
* can be specified in the .model statement or as part of the instance.  Instance level
* parameters override model level ones.  N = number of segments.

* intra cellular resistivity, rl,  is typically 1-3 kOhm mm.  Resistance along the long axis (longitudinal resistance Rl = rl L / (pi a^2)
* 1 kOhm mm = 1000 Ohm mm = 100 Ohm cm 

*yneuron neuron1  a b udParams R=1.0e2 A=1.0e-4 L=0.4 N=100 
yneuron neuron1  a b udParams R=1.0e2 A=1.0e-4 L=0.004 N=3

.tran 0 2.0e-2 
.print tran i(iin) V(a)
*n(y%neuron%neuron1_V10) n(y%neuron%neuron1_V20) n(y%neuron%neuron1_V30) 
*+ n(y%neuron%neuron1_V40) n(y%neuron%neuron1_V50) n(y%neuron%neuron1_V60) n(y%neuron%neuron1_V70)
*+ n(y%neuron%neuron1_V80) n(y%neuron%neuron1_V90) V(b)


.end


