* Small circuit demonstrating the fix for issue 575.
* Issue 575 was about Bsrc-based table models being 
* ineffient when the table is large and the table 
* entries are based on expressions.
*
* In older versions of Xyce this circuit takes many minutes to run.
* After the fix it takes seconds.  (about 25 seconds on my old 
* laptop as of this writing)

.param eric=0.9
.param vdd2={eric*2.0}
.param vdd=1.8

.param vss=0.1

.step eric list 0.5 0.9

.print tran v(in_S)

.tran 12000.100000ns 1550611.300000ns noop

RS in_S 0 1.0
BS in_S 0 V= {table(time,
+ 0.100000ns, VSS,
+ 960.800000ns, VSS,
+ 960.900000ns, VDD2,
+ 1441.200000ns, VDD2,
+ 1441.300000ns, VSS,
+ 1921.600000ns, VSS,
+ 1921.700000ns, VDD,
+ 2882.400000ns, VDD,
+ 2882.500000ns, VSS,
+ 3843.200000ns, VSS,
+ 3843.300000ns, VDD,
+ 4563.800000ns, VDD,
+ 4563.900000ns, VSS,
+ 4924.100000ns, VSS,
+ 4924.200000ns, VDD,
+ 6125.100000ns, VDD,
+ 6125.200000ns, VSS,
+ 6245.200000ns, VSS,
+ 6245.300000ns, VDD,
+ 7326.100000ns, VDD,
+ 7326.200000ns, VSS,
+ 7686.400000ns, VSS,
+ 7686.500000ns, VDD,
+ 7806.500000ns, VDD,
+ 7806.600000ns, VSS,
+ 7926.600000ns, VSS,
+ 7926.700000ns, VDD,
+ 9728.100000ns, VDD,
+ 9728.200000ns, VSS,
+ 10088.400000ns, VSS,
+ 10088.500000ns, VDD,
+ 10328.600000ns, VDD,
+ 10328.700000ns, VSS,
+ 10448.700000ns, VSS,
+ 10448.800000ns, VDD,
+ 10688.900000ns, VDD,
+ 10689.000000ns, VSS,
+ 10929.100000ns, VSS,
+ 10929.200000ns, VDD,
+ 11529.600000ns, VDD,
+ 11529.700000ns, VSS,
+ 11649.700000ns, VSS,
+ 11649.800000ns, VDD,
+ 12490.400000ns, VDD,
+ 12490.500000ns, VSS,
+ 12970.800000ns, VSS,
+ 12970.900000ns, VDD,
+ 13090.900000ns, VDD,
+ 13091.000000ns, VSS,
+ 13451.200000ns, VSS,
+ 13451.300000ns, VDD,
+ 13811.500000ns, VDD,
+ 13811.600000ns, VSS,
+ 14291.900000ns, VSS,
+ 14292.000000ns, VDD,
+ 14772.300000ns, VDD,
+ 14772.400000ns, VSS,
+ 15132.600000ns, VSS,
+ 15132.700000ns, VDD,
+ 15372.800000ns, VDD,
+ 15372.900000ns, VSS,
+ 15613.000000ns, VSS,
+ 15613.100000ns, VDD,
+ 16093.400000ns, VDD,
+ 16093.500000ns, VSS,
+ 16333.600000ns, VSS,
+ 16333.700000ns, VDD,
+ 18855.700000ns, VDD,
+ 18855.800000ns, VSS,
+ 19095.900000ns, VSS,
+ 19096.000000ns, VDD,
+ 19216.000000ns, VDD,
+ 19216.100000ns, VSS,
+ 19336.100000ns, VSS,
+ 19336.200000ns, VDD,
+ 20176.800000ns, VDD,
+ 20176.900000ns, VSS,
+ 20296.900000ns, VSS,
+ 20297.000000ns, VDD,
+ 20417.000000ns, VDD,
+ 20417.100000ns, VSS,
+ 21618.000000ns, VSS,
+ 21618.100000ns, VDD,
+ 21978.300000ns, VDD,
+ 21978.400000ns, VSS,
+ 22338.600000ns, VSS,
+ 22338.700000ns, VDD,
+ 23299.400000ns, VDD,
+ 23299.500000ns, VSS,
+ 23779.800000ns, VSS,
+ 23779.900000ns, VDD,
+ 24740.600000ns, VDD,
+ 24740.700000ns, VSS,
+ 25100.900000ns, VSS,
+ 25101.000000ns, VDD,
+ 25701.400000ns, VDD,
+ 25701.500000ns, VSS,
+ 26422.000000ns, VSS,
+ 26422.100000ns, VDD,
+ 26902.400000ns, VDD,
+ 26902.500000ns, VSS,
+ 27262.700000ns, VSS,
+ 27262.800000ns, VDD,
+ 27983.300000ns, VDD,
+ 27983.400000ns, VSS,
+ 28343.600000ns, VSS,
+ 28343.700000ns, VDD,
+ 28583.800000ns, VDD,
+ 28583.900000ns, VSS,
+ 29664.700000ns, VSS,
+ 29664.800000ns, VDD,
+ 30025.000000ns, VDD,
+ 30025.100000ns, VSS,
+ 31466.200000ns, VSS,
+ 31466.300000ns, VDD,
+ 32066.700000ns, VDD,
+ 32066.800000ns, VSS,
+ 32547.100000ns, VSS,
+ 32547.200000ns, VDD,
+ 33387.800000ns, VDD,
+ 33387.900000ns, VSS,
+ 33748.100000ns, VSS,
+ 33748.200000ns, VDD,
+ 35669.700000ns, VDD,
+ 35669.800000ns, VSS,
+ 36390.300000ns, VSS,
+ 36390.400000ns, VDD,
+ 37471.200000ns, VDD,
+ 37471.300000ns, VSS,
+ 38071.700000ns, VSS,
+ 38071.800000ns, VDD,
+ 38552.100000ns, VDD,
+ 38552.200000ns, VSS,
+ 38672.200000ns, VSS,
+ 38672.300000ns, VDD,
+ 38792.300000ns, VDD,
+ 38792.400000ns, VSS,
+ 38912.400000ns, VSS,
+ 38912.500000ns, VDD,
+ 39032.500000ns, VDD,
+ 39032.600000ns, VSS,
+ 41434.500000ns, VSS,
+ 41434.600000ns, VDD,
+ 42035.000000ns, VDD,
+ 42035.100000ns, VSS,
+ 42515.400000ns, VSS,
+ 42515.500000ns, VDD,
+ 44557.100000ns, VDD,
+ 44557.200000ns, VSS,
+ 45397.800000ns, VSS,
+ 45397.900000ns, VDD,
+ 45878.200000ns, VDD,
+ 45878.300000ns, VSS,
+ 46478.700000ns, VSS,
+ 46478.800000ns, VDD,
+ 47559.600000ns, VDD,
+ 47559.700000ns, VSS,
+ 47799.800000ns, VSS,
+ 47799.900000ns, VDD,
+ 50081.700000ns, VDD,
+ 50081.800000ns, VSS,
+ 50321.900000ns, VSS,
+ 50322.000000ns, VDD,
+ 50442.000000ns, VDD,
+ 50442.100000ns, VSS,
+ 50802.300000ns, VSS,
+ 50802.400000ns, VDD,
+ 50922.400000ns, VDD,
+ 50922.500000ns, VSS,
+ 51042.500000ns, VSS,
+ 51042.600000ns, VDD,
+ 52483.700000ns, VDD,
+ 52483.800000ns, VSS,
+ 52844.000000ns, VSS,
+ 52844.100000ns, VDD,
+ 53324.400000ns, VDD,
+ 53324.500000ns, VSS,
+ 53924.900000ns, VSS,
+ 53925.000000ns, VDD,
+ 55246.000000ns, VDD,
+ 55246.100000ns, VSS,
+ 55726.400000ns, VSS,
+ 55726.500000ns, VDD,
+ 56567.100000ns, VDD,
+ 56567.200000ns, VSS,
+ 56927.400000ns, VSS,
+ 56927.500000ns, VDD,
+ 57047.500000ns, VDD,
+ 57047.600000ns, VSS,
+ 57407.800000ns, VSS,
+ 57407.900000ns, VDD,
+ 58008.300000ns, VDD,
+ 58008.400000ns, VSS,
+ 58488.700000ns, VSS,
+ 58488.800000ns, VDD,
+ 58608.800000ns, VDD,
+ 58608.900000ns, VSS,
+ 58728.900000ns, VSS,
+ 58729.000000ns, VDD,
+ 60290.200000ns, VDD,
+ 60290.300000ns, VSS,
+ 60530.400000ns, VSS,
+ 60530.500000ns, VDD,
+ 60650.500000ns, VDD,
+ 60650.600000ns, VSS,
+ 61130.900000ns, VSS,
+ 61131.000000ns, VDD,
+ 61731.400000ns, VDD,
+ 61731.500000ns, VSS,
+ 62211.800000ns, VSS,
+ 62211.900000ns, VDD,
+ 63653.000000ns, VDD,
+ 63653.100000ns, VSS,
+ 63773.100000ns, VSS,
+ 63773.200000ns, VDD,
+ 63893.200000ns, VDD,
+ 63893.300000ns, VSS,
+ 65934.900000ns, VSS,
+ 65935.000000ns, VDD,
+ 67135.900000ns, VDD,
+ 67136.000000ns, VSS,
+ 67616.300000ns, VSS,
+ 67616.400000ns, VDD,
+ 68096.700000ns, VDD,
+ 68096.800000ns, VSS,
+ 68457.000000ns, VSS,
+ 68457.100000ns, VDD,
+ 68817.300000ns, VDD,
+ 68817.400000ns, VSS,
+ 70859.000000ns, VSS,
+ 70859.100000ns, VDD,
+ 70979.100000ns, VDD,
+ 70979.200000ns, VSS,
+ 71459.500000ns, VSS,
+ 71459.600000ns, VDD,
+ 72060.000000ns, VDD,
+ 72060.100000ns, VSS,
+ 72540.400000ns, VSS,
+ 72540.500000ns, VDD,
+ 73621.300000ns, VDD,
+ 73621.400000ns, VSS,
+ 73741.400000ns, VSS,
+ 73741.500000ns, VDD,
+ 74341.900000ns, VDD,
+ 74342.000000ns, VSS,
+ 76263.500000ns, VSS,
+ 76263.600000ns, VDD,
+ 76503.700000ns, VDD,
+ 76503.800000ns, VSS,
+ 76864.000000ns, VSS,
+ 76864.100000ns, VDD,
+ 76984.100000ns, VDD,
+ 76984.200000ns, VSS,
+ 77104.200000ns, VSS,
+ 77104.300000ns, VDD,
+ 77344.400000ns, VDD,
+ 77344.500000ns, VSS,
+ 77464.500000ns, VSS,
+ 77464.600000ns, VDD,
+ 77584.600000ns, VDD,
+ 77584.700000ns, VSS,
+ 79266.000000ns, VSS,
+ 79266.100000ns, VDD,
+ 81187.600000ns, VDD,
+ 81187.700000ns, VSS,
+ 81307.700000ns, VSS,
+ 81307.800000ns, VDD,
+ 81427.800000ns, VDD,
+ 81427.900000ns, VSS,
+ 83469.500000ns, VSS,
+ 83469.600000ns, VDD,
+ 83949.900000ns, VDD,
+ 83950.000000ns, VSS,
+ 85030.800000ns, VSS,
+ 85030.900000ns, VDD,
+ 86111.700000ns, VDD,
+ 86111.800000ns, VSS,
+ 86592.100000ns, VSS,
+ 86592.200000ns, VDD,
+ 86712.200000ns, VDD,
+ 86712.300000ns, VSS,
+ 86832.300000ns, VSS,
+ 86832.400000ns, VDD,
+ 87072.500000ns, VDD,
+ 87072.600000ns, VSS,
+ 88033.300000ns, VSS,
+ 88033.400000ns, VDD,
+ 88513.700000ns, VDD,
+ 88513.800000ns, VSS,
+ 88994.100000ns, VSS,
+ 88994.200000ns, VDD,
+ 90555.400000ns, VDD,
+ 90555.500000ns, VSS,
+ 90915.700000ns, VSS,
+ 90915.800000ns, VDD,
+ 91155.900000ns, VDD,
+ 91156.000000ns, VSS,
+ 91276.000000ns, VSS,
+ 91276.100000ns, VDD,
+ 92356.900000ns, VDD,
+ 92357.000000ns, VSS,
+ 92717.200000ns, VSS,
+ 92717.300000ns, VDD,
+ 93197.600000ns, VDD,
+ 93197.700000ns, VSS,
+ 95359.400000ns, VSS,
+ 95359.500000ns, VDD,
+ 95719.700000ns, VDD,
+ 95719.800000ns, VSS,
+ 96440.300000ns, VSS,
+ 96440.400000ns, VDD,
+ 98962.400000ns, VDD,
+ 98962.500000ns, VSS,
+ 99202.600000ns, VSS,
+ 99202.700000ns, VDD,
+ 99683.000000ns, VDD,
+ 99683.100000ns, VSS,
+ 100403.600000ns, VSS,
+ 100403.700000ns, VDD,
+ 100643.800000ns, VDD,
+ 100643.900000ns, VSS,
+ 101244.300000ns, VSS,
+ 101244.400000ns, VDD,
+ 102205.100000ns, VDD,
+ 102205.200000ns, VSS,
+ 102325.200000ns, VSS,
+ 102325.300000ns, VDD,
+ 102445.300000ns, VDD,
+ 102445.400000ns, VSS,
+ 102925.700000ns, VSS,
+ 102925.800000ns, VDD,
+ 103286.000000ns, VDD,
+ 103286.100000ns, VSS,
+ 104006.600000ns, VSS,
+ 104006.700000ns, VDD,
+ 104487.000000ns, VDD,
+ 104487.100000ns, VSS,
+ 104607.100000ns, VSS,
+ 104607.200000ns, VDD,
+ 105087.500000ns, VDD,
+ 105087.600000ns, VSS,
+ 105207.600000ns, VSS,
+ 105207.700000ns, VDD,
+ 105327.700000ns, VDD,
+ 105327.800000ns, VSS,
+ 106408.600000ns, VSS,
+ 106408.700000ns, VDD,
+ 106528.700000ns, VDD,
+ 106528.800000ns, VSS,
+ 107009.100000ns, VSS,
+ 107009.200000ns, VDD,
+ 107489.500000ns, VDD,
+ 107489.600000ns, VSS,
+ 108330.200000ns, VSS,
+ 108330.300000ns, VDD,
+ 108450.300000ns, VDD,
+ 108450.400000ns, VSS,
+ 108810.600000ns, VSS,
+ 108810.700000ns, VDD,
+ 109050.800000ns, VDD,
+ 109050.900000ns, VSS,
+ 109291.000000ns, VSS,
+ 109291.100000ns, VDD,
+ 111572.900000ns, VDD,
+ 111573.000000ns, VSS,
+ 112413.600000ns, VSS,
+ 112413.700000ns, VDD,
+ 112773.900000ns, VDD,
+ 112774.000000ns, VSS,
+ 113014.100000ns, VSS,
+ 113014.200000ns, VDD,
+ 113614.600000ns, VDD,
+ 113614.700000ns, VSS,
+ 114935.700000ns, VSS,
+ 114935.800000ns, VDD,
+ 115175.900000ns, VDD,
+ 115176.000000ns, VSS,
+ 116136.700000ns, VSS,
+ 116136.800000ns, VDD,
+ 116497.000000ns, VDD,
+ 116497.100000ns, VSS,
+ 116617.100000ns, VSS,
+ 116617.200000ns, VDD,
+ 116737.200000ns, VDD,
+ 116737.300000ns, VSS,
+ 116977.400000ns, VSS,
+ 116977.500000ns, VDD,
+ 118178.400000ns, VDD,
+ 118178.500000ns, VSS,
+ 118658.800000ns, VSS,
+ 118658.900000ns, VDD,
+ 118778.900000ns, VDD,
+ 118779.000000ns, VSS,
+ 118899.000000ns, VSS,
+ 118899.100000ns, VDD,
+ 119379.400000ns, VDD,
+ 119379.500000ns, VSS,
+ 120100.000000ns, VSS,
+ 120100.100000ns, VDD,
+ 120340.200000ns, VDD,
+ 120340.300000ns, VSS,
+ 120820.600000ns, VSS,
+ 120820.700000ns, VDD,
+ 121180.900000ns, VDD,
+ 121181.000000ns, VSS,
+ 121781.400000ns, VSS,
+ 121781.500000ns, VDD,
+ 121901.500000ns, VDD,
+ 121901.600000ns, VSS,
+ 122141.700000ns, VSS,
+ 122141.800000ns, VDD,
+ 122862.300000ns, VDD,
+ 122862.400000ns, VSS,
+ 123102.500000ns, VSS,
+ 123102.600000ns, VDD,
+ 123222.600000ns, VDD,
+ 123222.700000ns, VSS,
+ 124183.400000ns, VSS,
+ 124183.500000ns, VDD,
+ 124543.700000ns, VDD,
+ 124543.800000ns, VSS,
+ 124663.800000ns, VSS,
+ 124663.900000ns, VDD,
+ 125504.500000ns, VDD,
+ 125504.600000ns, VSS,
+ 125984.900000ns, VSS,
+ 125985.000000ns, VDD,
+ 127906.500000ns, VDD,
+ 127906.600000ns, VSS,
+ 128386.900000ns, VSS,
+ 128387.000000ns, VDD,
+ 128867.300000ns, VDD,
+ 128867.400000ns, VSS,
+ 128987.400000ns, VSS,
+ 128987.500000ns, VDD,
+ 129587.900000ns, VDD,
+ 129588.000000ns, VSS,
+ 130188.400000ns, VSS,
+ 130188.500000ns, VDD,
+ 131149.200000ns, VDD,
+ 131149.300000ns, VSS,
+ 131869.800000ns, VSS,
+ 131869.900000ns, VDD,
+ 132230.100000ns, VDD,
+ 132230.200000ns, VSS,
+ 133551.200000ns, VSS,
+ 133551.300000ns, VDD,
+ 134271.800000ns, VDD,
+ 134271.900000ns, VSS,
+ 135352.700000ns, VSS,
+ 135352.800000ns, VDD,
+ 135713.000000ns, VDD,
+ 135713.100000ns, VSS,
+ 138355.200000ns, VSS,
+ 138355.300000ns, VDD,
+ 138715.500000ns, VDD,
+ 138715.600000ns, VSS,
+ 139195.900000ns, VSS,
+ 139196.000000ns, VDD,
+ 140156.700000ns, VDD,
+ 140156.800000ns, VSS,
+ 140517.000000ns, VSS,
+ 140517.100000ns, VDD,
+ 140757.200000ns, VDD,
+ 140757.300000ns, VSS,
+ 141597.900000ns, VSS,
+ 141598.000000ns, VDD,
+ 141838.100000ns, VDD,
+ 141838.200000ns, VSS,
+ 142318.500000ns, VSS,
+ 142318.600000ns, VDD,
+ 143639.600000ns, VDD,
+ 143639.700000ns, VSS,
+ 144600.400000ns, VSS,
+ 144600.500000ns, VDD,
+ 145681.300000ns, VDD,
+ 145681.400000ns, VSS,
+ 146161.700000ns, VSS,
+ 146161.800000ns, VDD,
+ 146642.100000ns, VDD,
+ 146642.200000ns, VSS,
+ 148323.500000ns, VSS,
+ 148323.600000ns, VDD,
+ 148443.600000ns, VDD,
+ 148443.700000ns, VSS,
+ 150004.900000ns, VSS,
+ 150005.000000ns, VDD,
+ 150965.700000ns, VDD,
+ 150965.800000ns, VSS,
+ 152767.200000ns, VSS,
+ 152767.300000ns, VDD,
+ 153367.700000ns, VDD,
+ 153367.800000ns, VSS,
+ 153728.000000ns, VSS,
+ 153728.100000ns, VDD,
+ 154088.300000ns, VDD,
+ 154088.400000ns, VSS,
+ 154688.800000ns, VSS,
+ 154688.900000ns, VDD,
+ 155049.100000ns, VDD,
+ 155049.200000ns, VSS,
+ 155529.500000ns, VSS,
+ 155529.600000ns, VDD,
+ 155649.600000ns, VDD,
+ 155649.700000ns, VSS,
+ 157331.000000ns, VSS,
+ 157331.100000ns, VDD,
+ 159853.100000ns, VDD,
+ 159853.200000ns, VSS,
+ 160453.600000ns, VSS,
+ 160453.700000ns, VDD,
+ 160573.700000ns, VDD,
+ 160573.800000ns, VSS,
+ 160693.800000ns, VSS,
+ 160693.900000ns, VDD,
+ 161174.200000ns, VDD,
+ 161174.300000ns, VSS,
+ 161654.600000ns, VSS,
+ 161654.700000ns, VDD,
+ 162135.000000ns, VDD,
+ 162135.100000ns, VSS,
+ 162735.500000ns, VSS,
+ 162735.600000ns, VDD,
+ 162855.600000ns, VDD,
+ 162855.700000ns, VSS,
+ 163215.900000ns, VSS,
+ 163216.000000ns, VDD,
+ 163696.300000ns, VDD,
+ 163696.400000ns, VSS,
+ 164657.100000ns, VSS,
+ 164657.200000ns, VDD,
+ 165137.500000ns, VDD,
+ 165137.600000ns, VSS,
+ 165377.700000ns, VSS,
+ 165377.800000ns, VDD,
+ 165978.200000ns, VDD,
+ 165978.300000ns, VSS,
+ 166939.000000ns, VSS,
+ 166939.100000ns, VDD,
+ 167779.700000ns, VDD,
+ 167779.800000ns, VSS,
+ 169581.200000ns, VSS,
+ 169581.300000ns, VDD,
+ 169821.400000ns, VDD,
+ 169821.500000ns, VSS,
+ 170782.200000ns, VSS,
+ 170782.300000ns, VDD,
+ 171382.700000ns, VDD,
+ 171382.800000ns, VSS,
+ 171502.800000ns, VSS,
+ 171502.900000ns, VDD,
+ 172463.600000ns, VDD,
+ 172463.700000ns, VSS,
+ 172583.700000ns, VSS,
+ 172583.800000ns, VDD,
+ 172703.800000ns, VDD,
+ 172703.900000ns, VSS,
+ 173184.200000ns, VSS,
+ 173184.300000ns, VDD,
+ 174265.100000ns, VDD,
+ 174265.200000ns, VSS,
+ 174865.600000ns, VSS,
+ 174865.700000ns, VDD,
+ 176426.900000ns, VDD,
+ 176427.000000ns, VSS,
+ 177027.400000ns, VSS,
+ 177027.500000ns, VDD,
+ 177748.000000ns, VDD,
+ 177748.100000ns, VSS,
+ 178108.300000ns, VSS,
+ 178108.400000ns, VDD,
+ 178588.700000ns, VDD,
+ 178588.800000ns, VSS,
+ 178708.800000ns, VSS,
+ 178708.900000ns, VDD,
+ 179549.500000ns, VDD,
+ 179549.600000ns, VSS,
+ 180029.900000ns, VSS,
+ 180030.000000ns, VDD,
+ 181351.000000ns, VDD,
+ 181351.100000ns, VSS,
+ 182311.800000ns, VSS,
+ 182311.900000ns, VDD,
+ 182552.000000ns, VDD,
+ 182552.100000ns, VSS,
+ 183753.000000ns, VSS,
+ 183753.100000ns, VDD,
+ 183993.200000ns, VDD,
+ 183993.300000ns, VSS,
+ 184233.400000ns, VSS,
+ 184233.500000ns, VDD,
+ 184593.700000ns, VDD,
+ 184593.800000ns, VSS,
+ 185314.300000ns, VSS,
+ 185314.400000ns, VDD,
+ 185674.600000ns, VDD,
+ 185674.700000ns, VSS,
+ 186034.900000ns, VSS,
+ 186035.000000ns, VDD,
+ 186155.000000ns, VDD,
+ 186155.100000ns, VSS,
+ 186635.400000ns, VSS,
+ 186635.500000ns, VDD,
+ 186995.700000ns, VDD,
+ 186995.800000ns, VSS,
+ 187476.100000ns, VSS,
+ 187476.200000ns, VDD,
+ 189397.700000ns, VDD,
+ 189397.800000ns, VSS,
+ 190478.600000ns, VSS,
+ 190478.700000ns, VDD,
+ 190838.900000ns, VDD,
+ 190839.000000ns, VSS,
+ 190959.000000ns, VSS,
+ 190959.100000ns, VDD,
+ 191559.500000ns, VDD,
+ 191559.600000ns, VSS,
+ 191679.600000ns, VSS,
+ 191679.700000ns, VDD,
+ 192520.300000ns, VDD,
+ 192520.400000ns, VSS,
+ 192880.600000ns, VSS,
+ 192880.700000ns, VDD,
+ 193361.000000ns, VDD,
+ 193361.100000ns, VSS,
+ 193841.400000ns, VSS,
+ 193841.500000ns, VDD,
+ 196003.200000ns, VDD,
+ 196003.300000ns, VSS,
+ 196123.300000ns, VSS,
+ 196123.400000ns, VDD,
+ 197444.400000ns, VDD,
+ 197444.500000ns, VSS,
+ 198405.200000ns, VSS,
+ 198405.300000ns, VDD,
+ 198645.400000ns, VDD,
+ 198645.500000ns, VSS,
+ 199245.900000ns, VSS,
+ 199246.000000ns, VDD,
+ 199966.500000ns, VDD,
+ 199966.600000ns, VSS,
+ 200927.300000ns, VSS,
+ 200927.400000ns, VDD,
+ 201768.000000ns, VDD,
+ 201768.100000ns, VSS,
+ 202248.400000ns, VSS,
+ 202248.500000ns, VDD,
+ 203689.600000ns, VDD,
+ 203689.700000ns, VSS,
+ 204530.300000ns, VSS,
+ 204530.400000ns, VDD,
+ 204770.500000ns, VDD,
+ 204770.600000ns, VSS,
+ 207532.800000ns, VSS,
+ 207532.900000ns, VDD,
+ 207893.100000ns, VDD,
+ 207893.200000ns, VSS,
+ 208133.300000ns, VSS,
+ 208133.400000ns, VDD,
+ 208253.400000ns, VDD,
+ 208253.500000ns, VSS,
+ 208613.700000ns, VSS,
+ 208613.800000ns, VDD,
+ 209094.100000ns, VDD,
+ 209094.200000ns, VSS,
+ 209574.500000ns, VSS,
+ 209574.600000ns, VDD,
+ 210655.400000ns, VDD,
+ 210655.500000ns, VSS,
+ 211135.800000ns, VSS,
+ 211135.900000ns, VDD,
+ 211376.000000ns, VDD,
+ 211376.100000ns, VSS,
+ 211856.400000ns, VSS,
+ 211856.500000ns, VDD,
+ 215579.500000ns, VDD,
+ 215579.600000ns, VSS,
+ 215819.700000ns, VSS,
+ 215819.800000ns, VDD,
+ 216660.400000ns, VDD,
+ 216660.500000ns, VSS,
+ 216780.500000ns, VSS,
+ 216780.600000ns, VDD,
+ 217741.300000ns, VDD,
+ 217741.400000ns, VSS,
+ 217981.500000ns, VSS,
+ 217981.600000ns, VDD,
+ 219182.500000ns, VDD,
+ 219182.600000ns, VSS,
+ 219783.000000ns, VSS,
+ 219783.100000ns, VDD,
+ 220263.400000ns, VDD,
+ 220263.500000ns, VSS,
+ 220743.800000ns, VSS,
+ 220743.900000ns, VDD,
+ 221224.200000ns, VDD,
+ 221224.300000ns, VSS,
+ 221704.600000ns, VSS,
+ 221704.700000ns, VDD,
+ 222665.400000ns, VDD,
+ 222665.500000ns, VSS,
+ 223025.700000ns, VSS,
+ 223025.800000ns, VDD,
+ 223746.300000ns, VDD,
+ 223746.400000ns, VSS,
+ 224226.700000ns, VSS,
+ 224226.800000ns, VDD,
+ 224466.900000ns, VDD,
+ 224467.000000ns, VSS,
+ 224947.300000ns, VSS,
+ 224947.400000ns, VDD,
+ 225307.600000ns, VDD,
+ 225307.700000ns, VSS,
+ 225788.000000ns, VSS,
+ 225788.100000ns, VDD,
+ 226148.300000ns, VDD,
+ 226148.400000ns, VSS,
+ 226628.700000ns, VSS,
+ 226628.800000ns, VDD,
+ 227109.100000ns, VDD,
+ 227109.200000ns, VSS,
+ 228430.200000ns, VSS,
+ 228430.300000ns, VDD,
+ 229030.700000ns, VDD,
+ 229030.800000ns, VSS,
+ 229391.000000ns, VSS,
+ 229391.100000ns, VDD,
+ 229511.100000ns, VDD,
+ 229511.200000ns, VSS,
+ 230832.200000ns, VSS,
+ 230832.300000ns, VDD,
+ 231552.800000ns, VDD,
+ 231552.900000ns, VSS,
+ 232033.200000ns, VSS,
+ 232033.300000ns, VDD,
+ 232994.000000ns, VDD,
+ 232994.100000ns, VSS,
+ 233234.200000ns, VSS,
+ 233234.300000ns, VDD,
+ 233954.800000ns, VDD,
+ 233954.900000ns, VSS,
+ 234074.900000ns, VSS,
+ 234075.000000ns, VDD,
+ 234795.500000ns, VDD,
+ 234795.600000ns, VSS,
+ 235035.700000ns, VSS,
+ 235035.800000ns, VDD,
+ 235275.900000ns, VDD,
+ 235276.000000ns, VSS,
+ 235756.300000ns, VSS,
+ 235756.400000ns, VDD,
+ 235876.400000ns, VDD,
+ 235876.500000ns, VSS,
+ 237557.800000ns, VSS,
+ 237557.900000ns, VDD,
+ 239599.500000ns, VDD,
+ 239599.600000ns, VSS,
+ 239719.600000ns, VSS,
+ 239719.700000ns, VDD,
+ 239839.700000ns, VDD,
+ 239839.800000ns, VSS,
+ 241280.900000ns, VSS,
+ 241281.000000ns, VDD,
+ 242121.600000ns, VDD,
+ 242121.700000ns, VSS,
+ 242481.900000ns, VSS,
+ 242482.000000ns, VDD,
+ 243682.900000ns, VDD,
+ 243683.000000ns, VSS,
+ 244643.700000ns, VSS,
+ 244643.800000ns, VDD,
+ 246325.100000ns, VDD,
+ 246325.200000ns, VSS,
+ 247526.100000ns, VSS,
+ 247526.200000ns, VDD,
+ 249687.900000ns, VDD,
+ 249688.000000ns, VSS,
+ 250048.200000ns, VSS,
+ 250048.300000ns, VDD,
+ 250408.500000ns, VDD,
+ 250408.600000ns, VSS,
+ 250888.900000ns, VSS,
+ 250889.000000ns, VDD,
+ 251969.800000ns, VDD,
+ 251969.900000ns, VSS,
+ 253290.900000ns, VSS,
+ 253291.000000ns, VDD,
+ 253651.200000ns, VDD,
+ 253651.300000ns, VSS,
+ 253771.300000ns, VSS,
+ 253771.400000ns, VDD,
+ 253891.400000ns, VDD,
+ 253891.500000ns, VSS,
+ 254732.100000ns, VSS,
+ 254732.200000ns, VDD,
+ 255452.700000ns, VDD,
+ 255452.800000ns, VSS,
+ 255813.000000ns, VSS,
+ 255813.100000ns, VDD,
+ 256173.300000ns, VDD,
+ 256173.400000ns, VSS,
+ 256293.400000ns, VSS,
+ 256293.500000ns, VDD,
+ 256413.500000ns, VDD,
+ 256413.600000ns, VSS,
+ 257494.400000ns, VSS,
+ 257494.500000ns, VDD,
+ 258575.300000ns, VDD,
+ 258575.400000ns, VSS,
+ 259776.300000ns, VSS,
+ 259776.400000ns, VDD,
+ 260136.600000ns, VDD,
+ 260136.700000ns, VSS,
+ 260857.200000ns, VSS,
+ 260857.300000ns, VDD,
+ 261337.600000ns, VDD,
+ 261337.700000ns, VSS,
+ 262538.600000ns, VSS,
+ 262538.700000ns, VDD,
+ 263019.000000ns, VDD,
+ 263019.100000ns, VSS,
+ 263259.200000ns, VSS,
+ 263259.300000ns, VDD,
+ 264220.000000ns, VDD,
+ 264220.100000ns, VSS,
+ 265060.700000ns, VSS,
+ 265060.800000ns, VDD,
+ 265421.000000ns, VDD,
+ 265421.100000ns, VSS,
+ 266501.900000ns, VSS,
+ 266502.000000ns, VDD,
+ 267222.500000ns, VDD,
+ 267222.600000ns, VSS,
+ 267342.600000ns, VSS,
+ 267342.700000ns, VDD,
+ 267823.000000ns, VDD,
+ 267823.100000ns, VSS,
+ 267943.100000ns, VSS,
+ 267943.200000ns, VDD,
+ 268543.600000ns, VDD,
+ 268543.700000ns, VSS,
+ 270345.100000ns, VSS,
+ 270345.200000ns, VDD,
+ 270945.600000ns, VDD,
+ 270945.700000ns, VSS,
+ 272146.600000ns, VSS,
+ 272146.700000ns, VDD,
+ 272266.700000ns, VDD,
+ 272266.800000ns, VSS,
+ 272386.800000ns, VSS,
+ 272386.900000ns, VDD,
+ 273347.600000ns, VDD,
+ 273347.700000ns, VSS,
+ 273828.000000ns, VSS,
+ 273828.100000ns, VDD,
+ 274068.200000ns, VDD,
+ 274068.300000ns, VSS,
+ 274188.300000ns, VSS,
+ 274188.400000ns, VDD,
+ 275509.400000ns, VDD,
+ 275509.500000ns, VSS,
+ 275629.500000ns, VSS,
+ 275629.600000ns, VDD,
+ 276350.100000ns, VDD,
+ 276350.200000ns, VSS,
+ 277310.900000ns, VSS,
+ 277311.000000ns, VDD,
+ 277431.000000ns, VDD,
+ 277431.100000ns, VSS,
+ 277551.100000ns, VSS,
+ 277551.200000ns, VDD,
+ 277791.300000ns, VDD,
+ 277791.400000ns, VSS,
+ 278391.800000ns, VSS,
+ 278391.900000ns, VDD,
+ 279712.900000ns, VDD,
+ 279713.000000ns, VSS,
+ 280313.400000ns, VSS,
+ 280313.500000ns, VDD,
+ 280673.700000ns, VDD,
+ 280673.800000ns, VSS,
+ 281274.200000ns, VSS,
+ 281274.300000ns, VDD,
+ 282114.900000ns, VDD,
+ 282115.000000ns, VSS,
+ 282235.000000ns, VSS,
+ 282235.100000ns, VDD,
+ 283916.400000ns, VDD,
+ 283916.500000ns, VSS,
+ 284757.100000ns, VSS,
+ 284757.200000ns, VDD,
+ 284997.300000ns, VDD,
+ 284997.400000ns, VSS,
+ 285357.600000ns, VSS,
+ 285357.700000ns, VDD,
+ 286798.800000ns, VDD,
+ 286798.900000ns, VSS,
+ 287399.300000ns, VSS,
+ 287399.400000ns, VDD,
+ 288119.900000ns, VDD,
+ 288120.000000ns, VSS,
+ 288240.000000ns, VSS,
+ 288240.100000ns, VDD,
+ 288720.400000ns, VDD,
+ 288720.500000ns, VSS,
+ 289080.700000ns, VSS,
+ 289080.800000ns, VDD,
+ 290161.600000ns, VDD,
+ 290161.700000ns, VSS,
+ 290762.100000ns, VSS,
+ 290762.200000ns, VDD,
+ 291002.300000ns, VDD,
+ 291002.400000ns, VSS,
+ 291362.600000ns, VSS,
+ 291362.700000ns, VDD,
+ 291722.900000ns, VDD,
+ 291723.000000ns, VSS,
+ 292203.300000ns, VSS,
+ 292203.400000ns, VDD,
+ 292683.700000ns, VDD,
+ 292683.800000ns, VSS,
+ 293644.500000ns, VSS,
+ 293644.600000ns, VDD,
+ 294605.300000ns, VDD,
+ 294605.400000ns, VSS,
+ 294965.600000ns, VSS,
+ 294965.700000ns, VDD,
+ 296526.900000ns, VDD,
+ 296527.000000ns, VSS,
+ 297727.900000ns, VSS,
+ 297728.000000ns, VDD,
+ 298208.300000ns, VDD,
+ 298208.400000ns, VSS,
+ 298688.700000ns, VSS,
+ 298688.800000ns, VDD,
+ 299049.000000ns, VDD,
+ 299049.100000ns, VSS,
+ 301571.100000ns, VSS,
+ 301571.200000ns, VDD,
+ 302171.600000ns, VDD,
+ 302171.700000ns, VSS,
+ 303372.600000ns, VSS,
+ 303372.700000ns, VDD,
+ 304693.700000ns, VDD,
+ 304693.800000ns, VSS,
+ 305174.100000ns, VSS,
+ 305174.200000ns, VDD,
+ 305894.700000ns, VDD,
+ 305894.800000ns, VSS,
+ 306134.900000ns, VSS,
+ 306135.000000ns, VDD,
+ 306255.000000ns, VDD,
+ 306255.100000ns, VSS,
+ 306615.300000ns, VSS,
+ 306615.400000ns, VDD,
+ 306735.400000ns, VDD,
+ 306735.500000ns, VSS,
+ 309017.300000ns, VSS,
+ 309017.400000ns, VDD,
+ 310218.300000ns, VDD,
+ 310218.400000ns, VSS,
+ 311179.100000ns, VSS,
+ 311179.200000ns, VDD,
+ 311299.200000ns, VDD,
+ 311299.300000ns, VSS,
+ 311419.300000ns, VSS,
+ 311419.400000ns, VDD,
+ 313461.000000ns, VDD,
+ 313461.100000ns, VSS,
+ 314782.100000ns, VSS,
+ 314782.200000ns, VDD,
+ 315142.400000ns, VDD,
+ 315142.500000ns, VSS,
+ 315382.600000ns, VSS,
+ 315382.700000ns, VDD,
+ 315502.700000ns, VDD,
+ 315502.800000ns, VSS,
+ 315622.800000ns, VSS,
+ 315622.900000ns, VDD,
+ 316103.200000ns, VDD,
+ 316103.300000ns, VSS,
+ 316583.600000ns, VSS,
+ 316583.700000ns, VDD,
+ 317544.400000ns, VDD,
+ 317544.500000ns, VSS,
+ 317784.600000ns, VSS,
+ 317784.700000ns, VDD,
+ 318265.000000ns, VDD,
+ 318265.100000ns, VSS,
+ 319225.800000ns, VSS,
+ 319225.900000ns, VDD,
+ 319345.900000ns, VDD,
+ 319346.000000ns, VSS,
+ 319466.000000ns, VSS,
+ 319466.100000ns, VDD,
+ 319706.200000ns, VDD,
+ 319706.300000ns, VSS,
+ 320186.600000ns, VSS,
+ 320186.700000ns, VDD,
+ 320426.800000ns, VDD,
+ 320426.900000ns, VSS,
+ 320667.000000ns, VSS,
+ 320667.100000ns, VDD,
+ 321147.400000ns, VDD,
+ 321147.500000ns, VSS,
+ 321387.600000ns, VSS,
+ 321387.700000ns, VDD,
+ 321507.700000ns, VDD,
+ 321507.800000ns, VSS,
+ 321627.800000ns, VSS,
+ 321627.900000ns, VDD,
+ 322828.800000ns, VDD,
+ 322828.900000ns, VSS,
+ 323429.300000ns, VSS,
+ 323429.400000ns, VDD,
+ 323669.500000ns, VDD,
+ 323669.600000ns, VSS,
+ 323789.600000ns, VSS,
+ 323789.700000ns, VDD,
+ 324630.300000ns, VDD,
+ 324630.400000ns, VSS,
+ 327032.300000ns, VSS,
+ 327032.400000ns, VDD,
+ 327392.600000ns, VDD,
+ 327392.700000ns, VSS,
+ 327873.000000ns, VSS,
+ 327873.100000ns, VDD,
+ 329074.000000ns, VDD,
+ 329074.100000ns, VSS,
+ 331115.700000ns, VSS,
+ 331115.800000ns, VDD,
+ 331235.800000ns, VDD,
+ 331235.900000ns, VSS,
+ 331836.300000ns, VSS,
+ 331836.400000ns, VDD,
+ 334358.400000ns, VDD,
+ 334358.500000ns, VSS,
+ 334958.900000ns, VSS,
+ 334959.000000ns, VDD,
+ 335199.100000ns, VDD,
+ 335199.200000ns, VSS,
+ 335679.500000ns, VSS,
+ 335679.600000ns, VDD,
+ 336760.400000ns, VDD,
+ 336760.500000ns, VSS,
+ 337000.600000ns, VSS,
+ 337000.700000ns, VDD,
+ 337841.300000ns, VDD,
+ 337841.400000ns, VSS,
+ 338321.700000ns, VSS,
+ 338321.800000ns, VDD,
+ 339762.900000ns, VDD,
+ 339763.000000ns, VSS,
+ 340483.500000ns, VSS,
+ 340483.600000ns, VDD,
+ 340843.800000ns, VDD,
+ 340843.900000ns, VSS,
+ 341324.200000ns, VSS,
+ 341324.300000ns, VDD,
+ 343245.800000ns, VDD,
+ 343245.900000ns, VSS,
+ 344206.600000ns, VSS,
+ 344206.700000ns, VDD,
+ 344326.700000ns, VDD,
+ 344326.800000ns, VSS,
+ 344687.000000ns, VSS,
+ 344687.100000ns, VDD,
+ 345407.600000ns, VDD,
+ 345407.700000ns, VSS,
+ 346248.300000ns, VSS,
+ 346248.400000ns, VDD,
+ 346728.700000ns, VDD,
+ 346728.800000ns, VSS,
+ 348410.100000ns, VSS,
+ 348410.200000ns, VDD,
+ 348890.500000ns, VDD,
+ 348890.600000ns, VSS,
+ 349491.000000ns, VSS,
+ 349491.100000ns, VDD,
+ 349731.200000ns, VDD,
+ 349731.300000ns, VSS,
+ 350091.500000ns, VSS,
+ 350091.600000ns, VDD,
+ 350571.900000ns, VDD,
+ 350572.000000ns, VSS,
+ 350812.100000ns, VSS,
+ 350812.200000ns, VDD,
+ 351172.400000ns, VDD,
+ 351172.500000ns, VSS,
+ 351772.900000ns, VSS,
+ 351773.000000ns, VDD,
+ 351893.000000ns, VDD,
+ 351893.100000ns, VSS,
+ 352373.400000ns, VSS,
+ 352373.500000ns, VDD,
+ 352853.800000ns, VDD,
+ 352853.900000ns, VSS,
+ 356576.900000ns, VSS,
+ 356577.000000ns, VDD,
+ 358018.100000ns, VDD,
+ 358018.200000ns, VSS,
+ 358258.300000ns, VSS,
+ 358258.400000ns, VDD,
+ 358378.400000ns, VDD,
+ 358378.500000ns, VSS,
+ 358858.800000ns, VSS,
+ 358858.900000ns, VDD,
+ 359099.000000ns, VDD,
+ 359099.100000ns, VSS,
+ 360300.000000ns, VSS,
+ 360300.100000ns, VDD,
+ 361020.600000ns, VDD,
+ 361020.700000ns, VSS,
+ 361981.400000ns, VSS,
+ 361981.500000ns, VDD,
+ 363182.400000ns, VDD,
+ 363182.500000ns, VSS,
+ 363302.500000ns, VSS,
+ 363302.600000ns, VDD,
+ 363542.700000ns, VDD,
+ 363542.800000ns, VSS,
+ 364263.300000ns, VSS,
+ 364263.400000ns, VDD,
+ 364743.700000ns, VDD,
+ 364743.800000ns, VSS,
+ 366184.900000ns, VSS,
+ 366185.000000ns, VDD,
+ 366665.300000ns, VDD,
+ 366665.400000ns, VSS,
+ 367145.700000ns, VSS,
+ 367145.800000ns, VDD,
+ 368707.000000ns, VDD,
+ 368707.100000ns, VSS,
+ 369067.300000ns, VSS,
+ 369067.400000ns, VDD,
+ 370988.900000ns, VDD,
+ 370989.000000ns, VSS,
+ 372069.800000ns, VSS,
+ 372069.900000ns, VDD,
+ 374832.100000ns, VDD,
+ 374832.200000ns, VSS,
+ 376033.100000ns, VSS,
+ 376033.200000ns, VDD,
+ 376633.600000ns, VDD,
+ 376633.700000ns, VSS,
+ 376993.900000ns, VSS,
+ 376994.000000ns, VDD,
+ 377714.500000ns, VDD,
+ 377714.600000ns, VSS,
+ 378315.000000ns, VSS,
+ 378315.100000ns, VDD,
+ 378795.400000ns, VDD,
+ 378795.500000ns, VSS,
+ 379275.800000ns, VSS,
+ 379275.900000ns, VDD,
+ 379996.400000ns, VDD,
+ 379996.500000ns, VSS,
+ 382038.100000ns, VSS,
+ 382038.200000ns, VDD,
+ 383359.200000ns, VDD,
+ 383359.300000ns, VSS,
+ 384920.500000ns, VSS,
+ 384920.600000ns, VDD,
+ 385040.600000ns, VDD,
+ 385040.700000ns, VSS,
+ 386722.000000ns, VSS,
+ 386722.100000ns, VDD,
+ 388043.100000ns, VDD,
+ 388043.200000ns, VSS,
+ 388883.800000ns, VSS,
+ 388883.900000ns, VDD,
+ 389124.000000ns, VDD,
+ 389124.100000ns, VSS,
+ 389244.100000ns, VSS,
+ 389244.200000ns, VDD,
+ 389364.200000ns, VDD,
+ 389364.300000ns, VSS,
+ 389724.500000ns, VSS,
+ 389724.600000ns, VDD,
+ 390325.000000ns, VDD,
+ 390325.100000ns, VSS,
+ 390565.200000ns, VSS,
+ 390565.300000ns, VDD,
+ 392006.400000ns, VDD,
+ 392006.500000ns, VSS,
+ 392246.600000ns, VSS,
+ 392246.700000ns, VDD,
+ 392366.700000ns, VDD,
+ 392366.800000ns, VSS,
+ 392727.000000ns, VSS,
+ 392727.100000ns, VDD,
+ 392967.200000ns, VDD,
+ 392967.300000ns, VSS,
+ 393327.500000ns, VSS,
+ 393327.600000ns, VDD,
+ 393807.900000ns, VDD,
+ 393808.000000ns, VSS,
+ 394408.400000ns, VSS,
+ 394408.500000ns, VDD,
+ 395369.200000ns, VDD,
+ 395369.300000ns, VSS,
+ 396570.200000ns, VSS,
+ 396570.300000ns, VDD,
+ 396690.300000ns, VDD,
+ 396690.400000ns, VSS,
+ 396810.400000ns, VSS,
+ 396810.500000ns, VDD,
+ 397170.700000ns, VDD,
+ 397170.800000ns, VSS,
+ 397771.200000ns, VSS,
+ 397771.300000ns, VDD,
+ 398371.700000ns, VDD,
+ 398371.800000ns, VSS,
+ 400053.100000ns, VSS,
+ 400053.200000ns, VDD,
+ 401494.300000ns, VDD,
+ 401494.400000ns, VSS,
+ 402935.500000ns, VSS,
+ 402935.600000ns, VDD,
+ 403175.700000ns, VDD,
+ 403175.800000ns, VSS,
+ 404016.400000ns, VSS,
+ 404016.500000ns, VDD,
+ 405577.700000ns, VDD,
+ 405577.800000ns, VSS,
+ 406418.400000ns, VSS,
+ 406418.500000ns, VDD,
+ 406898.800000ns, VDD,
+ 406898.900000ns, VSS,
+ 407619.400000ns, VSS,
+ 407619.500000ns, VDD,
+ 407859.600000ns, VDD,
+ 407859.700000ns, VSS,
+ 409541.000000ns, VSS,
+ 409541.100000ns, VDD,
+ 410021.400000ns, VDD,
+ 410021.500000ns, VSS,
+ 410261.600000ns, VSS,
+ 410261.700000ns, VDD,
+ 410621.900000ns, VDD,
+ 410622.000000ns, VSS,
+ 410742.000000ns, VSS,
+ 410742.100000ns, VDD,
+ 410862.100000ns, VDD,
+ 410862.200000ns, VSS,
+ 411342.500000ns, VSS,
+ 411342.600000ns, VDD,
+ 412303.300000ns, VDD,
+ 412303.400000ns, VSS,
+ 413023.900000ns, VSS,
+ 413024.000000ns, VDD,
+ 414705.300000ns, VDD,
+ 414705.400000ns, VSS,
+ 415666.100000ns, VSS,
+ 415666.200000ns, VDD,
+ 416867.100000ns, VDD,
+ 416867.200000ns, VSS,
+ 417707.800000ns, VSS,
+ 417707.900000ns, VDD,
+ 418548.500000ns, VDD,
+ 418548.600000ns, VSS,
+ 419509.300000ns, VSS,
+ 419509.400000ns, VDD,
+ 419989.700000ns, VDD,
+ 419989.800000ns, VSS,
+ 420229.900000ns, VSS,
+ 420230.000000ns, VDD,
+ 420710.300000ns, VDD,
+ 420710.400000ns, VSS,
+ 421190.700000ns, VSS,
+ 421190.800000ns, VDD,
+ 421551.000000ns, VDD,
+ 421551.100000ns, VSS,
+ 422031.400000ns, VSS,
+ 422031.500000ns, VDD,
+ 422151.500000ns, VDD,
+ 422151.600000ns, VSS,
+ 422752.000000ns, VSS,
+ 422752.100000ns, VDD,
+ 423472.600000ns, VDD,
+ 423472.700000ns, VSS,
+ 423953.000000ns, VSS,
+ 423953.100000ns, VDD,
+ 424553.500000ns, VDD,
+ 424553.600000ns, VSS,
+ 425033.900000ns, VSS,
+ 425034.000000ns, VDD,
+ 426355.000000ns, VDD,
+ 426355.100000ns, VSS,
+ 427676.100000ns, VSS,
+ 427676.200000ns, VDD,
+ 429117.300000ns, VDD,
+ 429117.400000ns, VSS,
+ 431038.900000ns, VSS,
+ 431039.000000ns, VDD,
+ 431519.300000ns, VDD,
+ 431519.400000ns, VSS,
+ 431639.400000ns, VSS,
+ 431639.500000ns, VDD,
+ 431759.500000ns, VDD,
+ 431759.600000ns, VSS,
+ 434401.700000ns, VSS,
+ 434401.800000ns, VDD,
+ 434521.800000ns, VDD,
+ 434521.900000ns, VSS,
+ 435482.600000ns, VSS,
+ 435482.700000ns, VDD,
+ 436323.300000ns, VDD,
+ 436323.400000ns, VSS,
+ 436803.700000ns, VSS,
+ 436803.800000ns, VDD,
+ 436923.800000ns, VDD,
+ 436923.900000ns, VSS,
+ 437164.000000ns, VSS,
+ 437164.100000ns, VDD,
+ 437644.400000ns, VDD,
+ 437644.500000ns, VSS,
+ 438725.300000ns, VSS,
+ 438725.400000ns, VDD,
+ 438965.500000ns, VDD,
+ 438965.600000ns, VSS,
+ 439205.700000ns, VSS,
+ 439205.800000ns, VDD,
+ 439325.800000ns, VDD,
+ 439325.900000ns, VSS,
+ 441487.600000ns, VSS,
+ 441487.700000ns, VDD,
+ 442568.500000ns, VDD,
+ 442568.600000ns, VSS,
+ 442808.700000ns, VSS,
+ 442808.800000ns, VDD,
+ 444970.500000ns, VDD,
+ 444970.600000ns, VSS,
+ 445450.900000ns, VSS,
+ 445451.000000ns, VDD,
+ 446411.700000ns, VDD,
+ 446411.800000ns, VSS,
+ 446772.000000ns, VSS,
+ 446772.100000ns, VDD,
+ 447492.600000ns, VDD,
+ 447492.700000ns, VSS,
+ 448333.300000ns, VSS,
+ 448333.400000ns, VDD,
+ 448453.400000ns, VDD,
+ 448453.500000ns, VSS,
+ 448573.500000ns, VSS,
+ 448573.600000ns, VDD,
+ 449414.200000ns, VDD,
+ 449414.300000ns, VSS,
+ 451576.000000ns, VSS,
+ 451576.100000ns, VDD,
+ 452296.600000ns, VDD,
+ 452296.700000ns, VSS,
+ 453137.300000ns, VSS,
+ 453137.400000ns, VDD,
+ 453257.400000ns, VDD,
+ 453257.500000ns, VSS,
+ 453857.900000ns, VSS,
+ 453858.000000ns, VDD,
+ 453978.000000ns, VDD,
+ 453978.100000ns, VSS,
+ 454578.500000ns, VSS,
+ 454578.600000ns, VDD,
+ 454818.700000ns, VDD,
+ 454818.800000ns, VSS,
+ 456019.700000ns, VSS,
+ 456019.800000ns, VDD,
+ 456740.300000ns, VDD,
+ 456740.400000ns, VSS,
+ 457701.100000ns, VSS,
+ 457701.200000ns, VDD,
+ 458301.600000ns, VDD,
+ 458301.700000ns, VSS,
+ 458421.700000ns, VSS,
+ 458421.800000ns, VDD,
+ 458541.800000ns, VDD,
+ 458541.900000ns, VSS,
+ 458902.100000ns, VSS,
+ 458902.200000ns, VDD,
+ 459622.700000ns, VDD,
+ 459622.800000ns, VSS,
+ 459862.900000ns, VSS,
+ 459863.000000ns, VDD,
+ 459983.000000ns, VDD,
+ 459983.100000ns, VSS,
+ 460103.100000ns, VSS,
+ 460103.200000ns, VDD,
+ 460463.400000ns, VDD,
+ 460463.500000ns, VSS,
+ 462264.900000ns, VSS,
+ 462265.000000ns, VDD,
+ 462625.200000ns, VDD,
+ 462625.300000ns, VSS,
+ 463345.800000ns, VSS,
+ 463345.900000ns, VDD,
+ 463465.900000ns, VDD,
+ 463466.000000ns, VSS,
+ 464546.800000ns, VSS,
+ 464546.900000ns, VDD,
+ 464907.100000ns, VDD,
+ 464907.200000ns, VSS,
+ 465988.000000ns, VSS,
+ 465988.100000ns, VDD,
+ 468029.700000ns, VDD,
+ 468029.800000ns, VSS,
+ 470071.400000ns, VSS,
+ 470071.500000ns, VDD,
+ 470431.700000ns, VDD,
+ 470431.800000ns, VSS,
+ 471152.300000ns, VSS,
+ 471152.400000ns, VDD,
+ 471272.400000ns, VDD,
+ 471272.500000ns, VSS,
+ 471392.500000ns, VSS,
+ 471392.600000ns, VDD,
+ 471512.600000ns, VDD,
+ 471512.700000ns, VSS,
+ 472113.100000ns, VSS,
+ 472113.200000ns, VDD,
+ 472953.800000ns, VDD,
+ 472953.900000ns, VSS,
+ 473674.400000ns, VSS,
+ 473674.500000ns, VDD,
+ 475235.700000ns, VDD,
+ 475235.800000ns, VSS,
+ 476076.400000ns, VSS,
+ 476076.500000ns, VDD,
+ 476316.600000ns, VDD,
+ 476316.700000ns, VSS,
+ 476797.000000ns, VSS,
+ 476797.100000ns, VDD,
+ 477277.400000ns, VDD,
+ 477277.500000ns, VSS,
+ 477757.800000ns, VSS,
+ 477757.900000ns, VDD,
+ 478118.100000ns, VDD,
+ 478118.200000ns, VSS,
+ 478238.200000ns, VSS,
+ 478238.300000ns, VDD,
+ 478958.800000ns, VDD,
+ 478958.900000ns, VSS,
+ 480640.200000ns, VSS,
+ 480640.300000ns, VDD,
+ 481000.500000ns, VDD,
+ 481000.600000ns, VSS,
+ 481841.200000ns, VSS,
+ 481841.300000ns, VDD,
+ 482081.400000ns, VDD,
+ 482081.500000ns, VSS,
+ 483282.400000ns, VSS,
+ 483282.500000ns, VDD,
+ 483762.800000ns, VDD,
+ 483762.900000ns, VSS,
+ 484363.300000ns, VSS,
+ 484363.400000ns, VDD,
+ 485804.500000ns, VDD,
+ 485804.600000ns, VSS,
+ 486765.300000ns, VSS,
+ 486765.400000ns, VDD,
+ 489287.400000ns, VDD,
+ 489287.500000ns, VSS,
+ 490128.100000ns, VSS,
+ 490128.200000ns, VDD,
+ 490368.300000ns, VDD,
+ 490368.400000ns, VSS,
+ 490728.600000ns, VSS,
+ 490728.700000ns, VDD,
+ 491809.500000ns, VDD,
+ 491809.600000ns, VSS,
+ 493010.500000ns, VSS,
+ 493010.600000ns, VDD,
+ 494331.600000ns, VDD,
+ 494331.700000ns, VSS,
+ 494812.000000ns, VSS,
+ 494812.100000ns, VDD,
+ 495172.300000ns, VDD,
+ 495172.400000ns, VSS,
+ 495412.500000ns, VSS,
+ 495412.600000ns, VDD,
+ 496133.100000ns, VDD,
+ 496133.200000ns, VSS,
+ 497214.000000ns, VSS,
+ 497214.100000ns, VDD,
+ 498294.900000ns, VDD,
+ 498295.000000ns, VSS,
+ 499015.500000ns, VSS,
+ 499015.600000ns, VDD,
+ 500817.000000ns, VDD,
+ 500817.100000ns, VSS,
+ 501417.500000ns, VSS,
+ 501417.600000ns, VDD,
+ 502018.000000ns, VDD,
+ 502018.100000ns, VSS,
+ 502978.800000ns, VSS,
+ 502978.900000ns, VDD,
+ 503819.500000ns, VDD,
+ 503819.600000ns, VSS,
+ 505260.700000ns, VSS,
+ 505260.800000ns, VDD,
+ 505621.000000ns, VDD,
+ 505621.100000ns, VSS,
+ 505741.100000ns, VSS,
+ 505741.200000ns, VDD,
+ 506221.500000ns, VDD,
+ 506221.600000ns, VSS,
+ 507782.800000ns, VSS,
+ 507782.900000ns, VDD,
+ 508143.100000ns, VDD,
+ 508143.200000ns, VSS,
+ 509464.200000ns, VSS,
+ 509464.300000ns, VDD,
+ 510665.200000ns, VDD,
+ 510665.300000ns, VSS,
+ 510785.300000ns, VSS,
+ 510785.400000ns, VDD,
+ 511986.300000ns, VDD,
+ 511986.400000ns, VSS,
+ 512947.100000ns, VSS,
+ 512947.200000ns, VDD,
+ 513067.200000ns, VDD,
+ 513067.300000ns, VSS,
+ 514748.600000ns, VSS,
+ 514748.700000ns, VDD,
+ 514868.700000ns, VDD,
+ 514868.800000ns, VSS,
+ 515108.900000ns, VSS,
+ 515109.000000ns, VDD,
+ 516069.700000ns, VDD,
+ 516069.800000ns, VSS,
+ 516309.900000ns, VSS,
+ 516310.000000ns, VDD,
+ 517270.700000ns, VDD,
+ 517270.800000ns, VSS,
+ 518952.100000ns, VSS,
+ 518952.200000ns, VDD,
+ 519432.500000ns, VDD,
+ 519432.600000ns, VSS,
+ 519672.700000ns, VSS,
+ 519672.800000ns, VDD,
+ 520033.000000ns, VDD,
+ 520033.100000ns, VSS,
+ 520273.200000ns, VSS,
+ 520273.300000ns, VDD,
+ 521954.600000ns, VDD,
+ 521954.700000ns, VSS,
+ 522435.000000ns, VSS,
+ 522435.100000ns, VDD,
+ 522915.400000ns, VDD,
+ 522915.500000ns, VSS,
+ 523275.700000ns, VSS,
+ 523275.800000ns, VDD,
+ 523395.800000ns, VDD,
+ 523395.900000ns, VSS,
+ 523515.900000ns, VSS,
+ 523516.000000ns, VDD,
+ 523996.300000ns, VDD,
+ 523996.400000ns, VSS,
+ 524356.600000ns, VSS,
+ 524356.700000ns, VDD,
+ 525317.400000ns, VDD,
+ 525317.500000ns, VSS,
+ 525917.900000ns, VSS,
+ 525918.000000ns, VDD,
+ 526158.100000ns, VDD,
+ 526158.200000ns, VSS,
+ 526878.700000ns, VSS,
+ 526878.800000ns, VDD,
+ 526998.800000ns, VDD,
+ 526998.900000ns, VSS,
+ 527479.200000ns, VSS,
+ 527479.300000ns, VDD,
+ 528319.900000ns, VDD,
+ 528320.000000ns, VSS,
+ 528800.300000ns, VSS,
+ 528800.400000ns, VDD,
+ 529280.700000ns, VDD,
+ 529280.800000ns, VSS,
+ 531802.800000ns, VSS,
+ 531802.900000ns, VDD,
+ 533123.900000ns, VDD,
+ 533124.000000ns, VSS,
+ 533364.100000ns, VSS,
+ 533364.200000ns, VDD,
+ 533484.200000ns, VDD,
+ 533484.300000ns, VSS,
+ 534084.700000ns, VSS,
+ 534084.800000ns, VDD,
+ 535165.600000ns, VDD,
+ 535165.700000ns, VSS,
+ 535766.100000ns, VSS,
+ 535766.200000ns, VDD,
+ 536126.400000ns, VDD,
+ 536126.500000ns, VSS,
+ 536967.100000ns, VSS,
+ 536967.200000ns, VDD,
+ 537447.500000ns, VDD,
+ 537447.600000ns, VSS,
+ 537927.900000ns, VSS,
+ 537928.000000ns, VDD,
+ 538288.200000ns, VDD,
+ 538288.300000ns, VSS,
+ 539609.300000ns, VSS,
+ 539609.400000ns, VDD,
+ 541530.900000ns, VDD,
+ 541531.000000ns, VSS,
+ 541771.100000ns, VSS,
+ 541771.200000ns, VDD,
+ 542371.600000ns, VDD,
+ 542371.700000ns, VSS,
+ 542491.700000ns, VSS,
+ 542491.800000ns, VDD,
+ 543212.300000ns, VDD,
+ 543212.400000ns, VSS,
+ 544293.200000ns, VSS,
+ 544293.300000ns, VDD,
+ 544773.600000ns, VDD,
+ 544773.700000ns, VSS,
+ 545614.300000ns, VSS,
+ 545614.400000ns, VDD,
+ 546575.100000ns, VDD,
+ 546575.200000ns, VSS,
+ 547535.900000ns, VSS,
+ 547536.000000ns, VDD,
+ 548376.600000ns, VDD,
+ 548376.700000ns, VSS,
+ 550778.600000ns, VSS,
+ 550778.700000ns, VDD,
+ 551619.300000ns, VDD,
+ 551619.400000ns, VSS,
+ 552339.900000ns, VSS,
+ 552340.000000ns, VDD,
+ 553420.800000ns, VDD,
+ 553420.900000ns, VSS,
+ 553661.000000ns, VSS,
+ 553661.100000ns, VDD,
+ 554141.400000ns, VDD,
+ 554141.500000ns, VSS,
+ 554261.500000ns, VSS,
+ 554261.600000ns, VDD,
+ 556303.200000ns, VDD,
+ 556303.300000ns, VSS,
+ 557624.300000ns, VSS,
+ 557624.400000ns, VDD,
+ 558104.700000ns, VDD,
+ 558104.800000ns, VSS,
+ 558825.300000ns, VSS,
+ 558825.400000ns, VDD,
+ 558945.400000ns, VDD,
+ 558945.500000ns, VSS,
+ 559065.500000ns, VSS,
+ 559065.600000ns, VDD,
+ 560626.800000ns, VDD,
+ 560626.900000ns, VSS,
+ 560746.900000ns, VSS,
+ 560747.000000ns, VDD,
+ 560867.000000ns, VDD,
+ 560867.100000ns, VSS,
+ 561347.400000ns, VSS,
+ 561347.500000ns, VDD,
+ 562188.100000ns, VDD,
+ 562188.200000ns, VSS,
+ 564470.000000ns, VSS,
+ 564470.100000ns, VDD,
+ 564590.100000ns, VDD,
+ 564590.200000ns, VSS,
+ 565310.700000ns, VSS,
+ 565310.800000ns, VDD,
+ 566031.300000ns, VDD,
+ 566031.400000ns, VSS,
+ 566511.700000ns, VSS,
+ 566511.800000ns, VDD,
+ 567952.900000ns, VDD,
+ 567953.000000ns, VSS,
+ 568073.000000ns, VSS,
+ 568073.100000ns, VDD,
+ 568193.100000ns, VDD,
+ 568193.200000ns, VSS,
+ 568433.300000ns, VSS,
+ 568433.400000ns, VDD,
+ 570354.900000ns, VDD,
+ 570355.000000ns, VSS,
+ 570595.100000ns, VSS,
+ 570595.200000ns, VDD,
+ 571195.600000ns, VDD,
+ 571195.700000ns, VSS,
+ 572156.400000ns, VSS,
+ 572156.500000ns, VDD,
+ 572276.500000ns, VDD,
+ 572276.600000ns, VSS,
+ 572396.600000ns, VSS,
+ 572396.700000ns, VDD,
+ 572877.000000ns, VDD,
+ 572877.100000ns, VSS,
+ 573357.400000ns, VSS,
+ 573357.500000ns, VDD,
+ 573837.800000ns, VDD,
+ 573837.900000ns, VSS,
+ 574078.000000ns, VSS,
+ 574078.100000ns, VDD,
+ 574438.300000ns, VDD,
+ 574438.400000ns, VSS,
+ 574558.400000ns, VSS,
+ 574558.500000ns, VDD,
+ 576239.800000ns, VDD,
+ 576239.900000ns, VSS,
+ 577200.600000ns, VSS,
+ 577200.700000ns, VDD,
+ 577681.000000ns, VDD,
+ 577681.100000ns, VSS,
+ 578281.500000ns, VSS,
+ 578281.600000ns, VDD,
+ 579362.400000ns, VDD,
+ 579362.500000ns, VSS,
+ 580803.600000ns, VSS,
+ 580803.700000ns, VDD,
+ 581884.500000ns, VDD,
+ 581884.600000ns, VSS,
+ 582364.900000ns, VSS,
+ 582365.000000ns, VDD,
+ 582845.300000ns, VDD,
+ 582845.400000ns, VSS,
+ 583085.500000ns, VSS,
+ 583085.600000ns, VDD,
+ 584286.500000ns, VDD,
+ 584286.600000ns, VSS,
+ 584766.900000ns, VSS,
+ 584767.000000ns, VDD,
+ 585127.200000ns, VDD,
+ 585127.300000ns, VSS,
+ 585487.500000ns, VSS,
+ 585487.600000ns, VDD,
+ 586208.100000ns, VDD,
+ 586208.200000ns, VSS,
+ 587649.300000ns, VSS,
+ 587649.400000ns, VDD,
+ 587769.400000ns, VDD,
+ 587769.500000ns, VSS,
+ 589450.800000ns, VSS,
+ 589450.900000ns, VDD,
+ 589570.900000ns, VDD,
+ 589571.000000ns, VSS,
+ 589931.200000ns, VSS,
+ 589931.300000ns, VDD,
+ 592453.300000ns, VDD,
+ 592453.400000ns, VSS,
+ 593053.800000ns, VSS,
+ 593053.900000ns, VDD,
+ 593534.200000ns, VDD,
+ 593534.300000ns, VSS,
+ 593894.500000ns, VSS,
+ 593894.600000ns, VDD,
+ 594615.100000ns, VDD,
+ 594615.200000ns, VSS,
+ 594855.300000ns, VSS,
+ 594855.400000ns, VDD,
+ 595696.000000ns, VDD,
+ 595696.100000ns, VSS,
+ 595816.100000ns, VSS,
+ 595816.200000ns, VDD,
+ 595936.200000ns, VDD,
+ 595936.300000ns, VSS,
+ 596776.900000ns, VSS,
+ 596777.000000ns, VDD,
+ 597257.300000ns, VDD,
+ 597257.400000ns, VSS,
+ 598098.000000ns, VSS,
+ 598098.100000ns, VDD,
+ 598338.200000ns, VDD,
+ 598338.300000ns, VSS,
+ 598578.400000ns, VSS,
+ 598578.500000ns, VDD,
+ 598938.700000ns, VDD,
+ 598938.800000ns, VSS,
+ 600019.600000ns, VSS,
+ 600019.700000ns, VDD,
+ 600139.700000ns, VDD,
+ 600139.800000ns, VSS,
+ 600259.800000ns, VSS,
+ 600259.900000ns, VDD,
+ 600379.900000ns, VDD,
+ 600380.000000ns, VSS,
+ 602421.600000ns, VSS,
+ 602421.700000ns, VDD,
+ 603022.100000ns, VDD,
+ 603022.200000ns, VSS,
+ 603142.200000ns, VSS,
+ 603142.300000ns, VDD,
+ 603862.800000ns, VDD,
+ 603862.900000ns, VSS,
+ 604583.400000ns, VSS,
+ 604583.500000ns, VDD,
+ 605304.000000ns, VDD,
+ 605304.100000ns, VSS,
+ 605544.200000ns, VSS,
+ 605544.300000ns, VDD,
+ 605664.300000ns, VDD,
+ 605664.400000ns, VSS,
+ 605784.400000ns, VSS,
+ 605784.500000ns, VDD,
+ 606144.700000ns, VDD,
+ 606144.800000ns, VSS,
+ 606625.100000ns, VSS,
+ 606625.200000ns, VDD,
+ 607585.900000ns, VDD,
+ 607586.000000ns, VSS,
+ 608066.300000ns, VSS,
+ 608066.400000ns, VDD,
+ 608186.400000ns, VDD,
+ 608186.500000ns, VSS,
+ 609267.300000ns, VSS,
+ 609267.400000ns, VDD,
+ 610348.200000ns, VDD,
+ 610348.300000ns, VSS,
+ 610948.700000ns, VSS,
+ 610948.800000ns, VDD,
+ 613110.500000ns, VDD,
+ 613110.600000ns, VSS,
+ 613230.600000ns, VSS,
+ 613230.700000ns, VDD,
+ 613350.700000ns, VDD,
+ 613350.800000ns, VSS,
+ 614671.800000ns, VSS,
+ 614671.900000ns, VDD,
+ 614912.000000ns, VDD,
+ 614912.100000ns, VSS,
+ 616473.300000ns, VSS,
+ 616473.400000ns, VDD,
+ 617554.200000ns, VDD,
+ 617554.300000ns, VSS,
+ 618394.900000ns, VSS,
+ 618395.000000ns, VDD,
+ 619475.800000ns, VDD,
+ 619475.900000ns, VSS,
+ 620556.700000ns, VSS,
+ 620556.800000ns, VDD,
+ 621277.300000ns, VDD,
+ 621277.400000ns, VSS,
+ 621637.600000ns, VSS,
+ 621637.700000ns, VDD,
+ 622118.000000ns, VDD,
+ 622118.100000ns, VSS,
+ 622958.700000ns, VSS,
+ 622958.800000ns, VDD,
+ 623679.300000ns, VDD,
+ 623679.400000ns, VSS,
+ 624039.600000ns, VSS,
+ 624039.700000ns, VDD,
+ 625120.500000ns, VDD,
+ 625120.600000ns, VSS,
+ 627882.800000ns, VSS,
+ 627882.900000ns, VDD,
+ 629684.300000ns, VDD,
+ 629684.400000ns, VSS,
+ 630284.800000ns, VSS,
+ 630284.900000ns, VDD,
+ 630404.900000ns, VDD,
+ 630405.000000ns, VSS,
+ 630525.000000ns, VSS,
+ 630525.100000ns, VDD,
+ 630885.300000ns, VDD,
+ 630885.400000ns, VSS,
+ 631125.500000ns, VSS,
+ 631125.600000ns, VDD,
+ 633167.200000ns, VDD,
+ 633167.300000ns, VSS,
+ 634368.200000ns, VSS,
+ 634368.300000ns, VDD,
+ 634608.400000ns, VDD,
+ 634608.500000ns, VSS,
+ 634728.500000ns, VSS,
+ 634728.600000ns, VDD,
+ 636169.700000ns, VDD,
+ 636169.800000ns, VSS,
+ 636890.300000ns, VSS,
+ 636890.400000ns, VDD,
+ 637250.600000ns, VDD,
+ 637250.700000ns, VSS,
+ 637490.800000ns, VSS,
+ 637490.900000ns, VDD,
+ 638211.400000ns, VDD,
+ 638211.500000ns, VSS,
+ 638451.600000ns, VSS,
+ 638451.700000ns, VDD,
+ 638691.800000ns, VDD,
+ 638691.900000ns, VSS,
+ 638811.900000ns, VSS,
+ 638812.000000ns, VDD,
+ 641934.500000ns, VDD,
+ 641934.600000ns, VSS,
+ 642414.900000ns, VSS,
+ 642415.000000ns, VDD,
+ 642655.100000ns, VDD,
+ 642655.200000ns, VSS,
+ 642895.300000ns, VSS,
+ 642895.400000ns, VDD,
+ 643375.700000ns, VDD,
+ 643375.800000ns, VSS,
+ 643976.200000ns, VSS,
+ 643976.300000ns, VDD,
+ 644456.600000ns, VDD,
+ 644456.700000ns, VSS,
+ 644816.900000ns, VSS,
+ 644817.000000ns, VDD,
+ 645297.300000ns, VDD,
+ 645297.400000ns, VSS,
+ 645897.800000ns, VSS,
+ 645897.900000ns, VDD,
+ 646258.100000ns, VDD,
+ 646258.200000ns, VSS,
+ 646618.400000ns, VSS,
+ 646618.500000ns, VDD,
+ 646978.700000ns, VDD,
+ 646978.800000ns, VSS,
+ 647098.800000ns, VSS,
+ 647098.900000ns, VDD,
+ 648419.900000ns, VDD,
+ 648420.000000ns, VSS,
+ 649260.600000ns, VSS,
+ 649260.700000ns, VDD,
+ 649741.000000ns, VDD,
+ 649741.100000ns, VSS,
+ 650701.800000ns, VSS,
+ 650701.900000ns, VDD,
+ 652623.400000ns, VDD,
+ 652623.500000ns, VSS,
+ 653103.800000ns, VSS,
+ 653103.900000ns, VDD,
+ 653584.200000ns, VDD,
+ 653584.300000ns, VSS,
+ 653704.300000ns, VSS,
+ 653704.400000ns, VDD,
+ 653824.400000ns, VDD,
+ 653824.500000ns, VSS,
+ 653944.500000ns, VSS,
+ 653944.600000ns, VDD,
+ 654304.800000ns, VDD,
+ 654304.900000ns, VSS,
+ 655025.400000ns, VSS,
+ 655025.500000ns, VDD,
+ 655265.600000ns, VDD,
+ 655265.700000ns, VSS,
+ 655746.000000ns, VSS,
+ 655746.100000ns, VDD,
+ 656106.300000ns, VDD,
+ 656106.400000ns, VSS,
+ 656586.700000ns, VSS,
+ 656586.800000ns, VDD,
+ 657547.500000ns, VDD,
+ 657547.600000ns, VSS,
+ 657787.700000ns, VSS,
+ 657787.800000ns, VDD,
+ 659108.800000ns, VDD,
+ 659108.900000ns, VSS,
+ 659228.900000ns, VSS,
+ 659229.000000ns, VDD,
+ 659349.000000ns, VDD,
+ 659349.100000ns, VSS,
+ 661150.500000ns, VSS,
+ 661150.600000ns, VDD,
+ 662831.900000ns, VDD,
+ 662832.000000ns, VSS,
+ 665233.900000ns, VSS,
+ 665234.000000ns, VDD,
+ 665834.400000ns, VDD,
+ 665834.500000ns, VSS,
+ 666314.800000ns, VSS,
+ 666314.900000ns, VDD,
+ 667395.700000ns, VDD,
+ 667395.800000ns, VSS,
+ 667876.100000ns, VSS,
+ 667876.200000ns, VDD,
+ 668716.800000ns, VDD,
+ 668716.900000ns, VSS,
+ 669317.300000ns, VSS,
+ 669317.400000ns, VDD,
+ 669677.600000ns, VDD,
+ 669677.700000ns, VSS,
+ 671599.200000ns, VSS,
+ 671599.300000ns, VDD,
+ 671839.400000ns, VDD,
+ 671839.500000ns, VSS,
+ 672079.600000ns, VSS,
+ 672079.700000ns, VDD,
+ 672800.200000ns, VDD,
+ 672800.300000ns, VSS,
+ 673040.400000ns, VSS,
+ 673040.500000ns, VDD,
+ 673160.500000ns, VDD,
+ 673160.600000ns, VSS,
+ 674241.400000ns, VSS,
+ 674241.500000ns, VDD,
+ 675322.300000ns, VDD,
+ 675322.400000ns, VSS,
+ 675922.800000ns, VSS,
+ 675922.900000ns, VDD,
+ 676283.100000ns, VDD,
+ 676283.200000ns, VSS,
+ 676643.400000ns, VSS,
+ 676643.500000ns, VDD,
+ 677604.200000ns, VDD,
+ 677604.300000ns, VSS,
+ 678925.300000ns, VSS,
+ 678925.400000ns, VDD,
+ 679886.100000ns, VDD,
+ 679886.200000ns, VSS,
+ 680486.600000ns, VSS,
+ 680486.700000ns, VDD,
+ 681207.200000ns, VDD,
+ 681207.300000ns, VSS,
+ 682288.100000ns, VSS,
+ 682288.200000ns, VDD,
+ 682528.300000ns, VDD,
+ 682528.400000ns, VSS,
+ 683128.800000ns, VSS,
+ 683128.900000ns, VDD,
+ 683609.200000ns, VDD,
+ 683609.300000ns, VSS,
+ 684570.000000ns, VSS,
+ 684570.100000ns, VDD,
+ 684690.100000ns, VDD,
+ 684690.200000ns, VSS,
+ 685290.600000ns, VSS,
+ 685290.700000ns, VDD,
+ 685410.700000ns, VDD,
+ 685410.800000ns, VSS,
+ 685530.800000ns, VSS,
+ 685530.900000ns, VDD,
+ 687932.800000ns, VDD,
+ 687932.900000ns, VSS,
+ 690214.700000ns, VSS,
+ 690214.800000ns, VDD,
+ 690935.300000ns, VDD,
+ 690935.400000ns, VSS,
+ 692016.200000ns, VSS,
+ 692016.300000ns, VDD,
+ 692136.300000ns, VDD,
+ 692136.400000ns, VSS,
+ 692496.600000ns, VSS,
+ 692496.700000ns, VDD,
+ 692616.700000ns, VDD,
+ 692616.800000ns, VSS,
+ 693457.400000ns, VSS,
+ 693457.500000ns, VDD,
+ 693937.800000ns, VDD,
+ 693937.900000ns, VSS,
+ 694418.200000ns, VSS,
+ 694418.300000ns, VDD,
+ 695499.100000ns, VDD,
+ 695499.200000ns, VSS,
+ 696700.100000ns, VSS,
+ 696700.200000ns, VDD,
+ 696940.300000ns, VDD,
+ 696940.400000ns, VSS,
+ 697540.800000ns, VSS,
+ 697540.900000ns, VDD,
+ 697901.100000ns, VDD,
+ 697901.200000ns, VSS,
+ 698261.400000ns, VSS,
+ 698261.500000ns, VDD,
+ 698982.000000ns, VDD,
+ 698982.100000ns, VSS,
+ 699822.700000ns, VSS,
+ 699822.800000ns, VDD,
+ 700303.100000ns, VDD,
+ 700303.200000ns, VSS,
+ 700783.500000ns, VSS,
+ 700783.600000ns, VDD,
+ 701143.800000ns, VDD,
+ 701143.900000ns, VSS,
+ 702464.900000ns, VSS,
+ 702465.000000ns, VDD,
+ 703065.400000ns, VDD,
+ 703065.500000ns, VSS,
+ 703305.600000ns, VSS,
+ 703305.700000ns, VDD,
+ 704386.500000ns, VDD,
+ 704386.600000ns, VSS,
+ 704506.600000ns, VSS,
+ 704506.700000ns, VDD,
+ 704626.700000ns, VDD,
+ 704626.800000ns, VSS,
+ 705107.100000ns, VSS,
+ 705107.200000ns, VDD,
+ 705467.400000ns, VDD,
+ 705467.500000ns, VSS,
+ 705827.700000ns, VSS,
+ 705827.800000ns, VDD,
+ 705947.800000ns, VDD,
+ 705947.900000ns, VSS,
+ 706308.100000ns, VSS,
+ 706308.200000ns, VDD,
+ 708349.800000ns, VDD,
+ 708349.900000ns, VSS,
+ 709070.400000ns, VSS,
+ 709070.500000ns, VDD,
+ 710031.200000ns, VDD,
+ 710031.300000ns, VSS,
+ 710871.900000ns, VSS,
+ 710872.000000ns, VDD,
+ 710992.000000ns, VDD,
+ 710992.100000ns, VSS,
+ 711112.100000ns, VSS,
+ 711112.200000ns, VDD,
+ 711352.300000ns, VDD,
+ 711352.400000ns, VSS,
+ 711472.400000ns, VSS,
+ 711472.500000ns, VDD,
+ 711592.500000ns, VDD,
+ 711592.600000ns, VSS,
+ 712673.400000ns, VSS,
+ 712673.500000ns, VDD,
+ 713153.800000ns, VDD,
+ 713153.900000ns, VSS,
+ 714114.600000ns, VSS,
+ 714114.700000ns, VDD,
+ 715195.500000ns, VDD,
+ 715195.600000ns, VSS,
+ 715435.700000ns, VSS,
+ 715435.800000ns, VDD,
+ 715675.900000ns, VDD,
+ 715676.000000ns, VSS,
+ 715796.000000ns, VSS,
+ 715796.100000ns, VDD,
+ 715916.100000ns, VDD,
+ 715916.200000ns, VSS,
+ 716636.700000ns, VSS,
+ 716636.800000ns, VDD,
+ 717717.600000ns, VDD,
+ 717717.700000ns, VSS,
+ 718198.000000ns, VSS,
+ 718198.100000ns, VDD,
+ 718558.300000ns, VDD,
+ 718558.400000ns, VSS,
+ 720960.300000ns, VSS,
+ 720960.400000ns, VDD,
+ 721320.600000ns, VDD,
+ 721320.700000ns, VSS,
+ 722041.200000ns, VSS,
+ 722041.300000ns, VDD,
+ 722521.600000ns, VDD,
+ 722521.700000ns, VSS,
+ 723362.300000ns, VSS,
+ 723362.400000ns, VDD,
+ 723842.700000ns, VDD,
+ 723842.800000ns, VSS,
+ 723962.800000ns, VSS,
+ 723962.900000ns, VDD,
+ 724082.900000ns, VDD,
+ 724083.000000ns, VSS,
+ 724323.100000ns, VSS,
+ 724323.200000ns, VDD,
+ 724443.200000ns, VDD,
+ 724443.300000ns, VSS,
+ 725163.800000ns, VSS,
+ 725163.900000ns, VDD,
+ 725644.200000ns, VDD,
+ 725644.300000ns, VSS,
+ 726364.800000ns, VSS,
+ 726364.900000ns, VDD,
+ 726725.100000ns, VDD,
+ 726725.200000ns, VSS,
+ 727325.600000ns, VSS,
+ 727325.700000ns, VDD,
+ 729847.700000ns, VDD,
+ 729847.800000ns, VSS,
+ 730568.300000ns, VSS,
+ 730568.400000ns, VDD,
+ 731288.900000ns, VDD,
+ 731289.000000ns, VSS,
+ 731649.200000ns, VSS,
+ 731649.300000ns, VDD,
+ 731769.300000ns, VDD,
+ 731769.400000ns, VSS,
+ 732249.700000ns, VSS,
+ 732249.800000ns, VDD,
+ 733330.600000ns, VDD,
+ 733330.700000ns, VSS,
+ 734171.300000ns, VSS,
+ 734171.400000ns, VDD,
+ 734291.400000ns, VDD,
+ 734291.500000ns, VSS,
+ 735132.100000ns, VSS,
+ 735132.200000ns, VDD,
+ 735252.200000ns, VDD,
+ 735252.300000ns, VSS,
+ 735372.300000ns, VSS,
+ 735372.400000ns, VDD,
+ 735492.400000ns, VDD,
+ 735492.500000ns, VSS,
+ 736453.200000ns, VSS,
+ 736453.300000ns, VDD,
+ 736573.300000ns, VDD,
+ 736573.400000ns, VSS,
+ 737774.300000ns, VSS,
+ 737774.400000ns, VDD,
+ 738134.600000ns, VDD,
+ 738134.700000ns, VSS,
+ 738615.000000ns, VSS,
+ 738615.100000ns, VDD,
+ 739215.500000ns, VDD,
+ 739215.600000ns, VSS,
+ 740176.300000ns, VSS,
+ 740176.400000ns, VDD,
+ 741857.700000ns, VDD,
+ 741857.800000ns, VSS,
+ 742338.100000ns, VSS,
+ 742338.200000ns, VDD,
+ 743298.900000ns, VDD,
+ 743299.000000ns, VSS,
+ 743659.200000ns, VSS,
+ 743659.300000ns, VDD,
+ 744620.000000ns, VDD,
+ 744620.100000ns, VSS,
+ 745340.600000ns, VSS,
+ 745340.700000ns, VDD,
+ 745821.000000ns, VDD,
+ 745821.100000ns, VSS,
+ 746181.300000ns, VSS,
+ 746181.400000ns, VDD,
+ 746301.400000ns, VDD,
+ 746301.500000ns, VSS,
+ 746541.600000ns, VSS,
+ 746541.700000ns, VDD,
+ 747022.000000ns, VDD,
+ 747022.100000ns, VSS,
+ 747142.100000ns, VSS,
+ 747142.200000ns, VDD,
+ 747262.200000ns, VDD,
+ 747262.300000ns, VSS,
+ 747502.400000ns, VSS,
+ 747502.500000ns, VDD,
+ 747622.500000ns, VDD,
+ 747622.600000ns, VSS,
+ 748583.300000ns, VSS,
+ 748583.400000ns, VDD,
+ 748823.500000ns, VDD,
+ 748823.600000ns, VSS,
+ 748943.600000ns, VSS,
+ 748943.700000ns, VDD,
+ 749183.800000ns, VDD,
+ 749183.900000ns, VSS,
+ 749303.900000ns, VSS,
+ 749304.000000ns, VDD,
+ 750745.100000ns, VDD,
+ 750745.200000ns, VSS,
+ 751585.800000ns, VSS,
+ 751585.900000ns, VDD,
+ 751946.100000ns, VDD,
+ 751946.200000ns, VSS,
+ 752906.900000ns, VSS,
+ 752907.000000ns, VDD,
+ 753627.500000ns, VDD,
+ 753627.600000ns, VSS,
+ 753747.600000ns, VSS,
+ 753747.700000ns, VDD,
+ 754228.000000ns, VDD,
+ 754228.100000ns, VSS,
+ 754348.100000ns, VSS,
+ 754348.200000ns, VDD,
+ 754708.400000ns, VDD,
+ 754708.500000ns, VSS,
+ 754828.500000ns, VSS,
+ 754828.600000ns, VDD,
+ 754948.600000ns, VDD,
+ 754948.700000ns, VSS,
+ 755068.700000ns, VSS,
+ 755068.800000ns, VDD,
+ 755429.000000ns, VDD,
+ 755429.100000ns, VSS,
+ 756029.500000ns, VSS,
+ 756029.600000ns, VDD,
+ 756630.000000ns, VDD,
+ 756630.100000ns, VSS,
+ 756750.100000ns, VSS,
+ 756750.200000ns, VDD,
+ 757590.800000ns, VDD,
+ 757590.900000ns, VSS,
+ 758191.300000ns, VSS,
+ 758191.400000ns, VDD,
+ 759152.100000ns, VDD,
+ 759152.200000ns, VSS,
+ 759992.800000ns, VSS,
+ 759992.900000ns, VDD,
+ 760473.200000ns, VDD,
+ 760473.300000ns, VSS,
+ 760953.600000ns, VSS,
+ 760953.700000ns, VDD,
+ 761434.000000ns, VDD,
+ 761434.100000ns, VSS,
+ 763956.100000ns, VSS,
+ 763956.200000ns, VDD,
+ 764076.200000ns, VDD,
+ 764076.300000ns, VSS,
+ 764316.400000ns, VSS,
+ 764316.500000ns, VDD,
+ 764436.500000ns, VDD,
+ 764436.600000ns, VSS,
+ 764916.900000ns, VSS,
+ 764917.000000ns, VDD,
+ 765277.200000ns, VDD,
+ 765277.300000ns, VSS,
+ 765637.500000ns, VSS,
+ 765637.600000ns, VDD,
+ 765877.700000ns, VDD,
+ 765877.800000ns, VSS,
+ 766718.400000ns, VSS,
+ 766718.500000ns, VDD,
+ 766958.600000ns, VDD,
+ 766958.700000ns, VSS,
+ 767198.800000ns, VSS,
+ 767198.900000ns, VDD,
+ 767439.000000ns, VDD,
+ 767439.100000ns, VSS,
+ 767559.100000ns, VSS,
+ 767559.200000ns, VDD,
+ 768279.700000ns, VDD,
+ 768279.800000ns, VSS,
+ 768760.100000ns, VSS,
+ 768760.200000ns, VDD,
+ 769120.400000ns, VDD,
+ 769120.500000ns, VSS,
+ 769600.800000ns, VSS,
+ 769600.900000ns, VDD,
+ 771282.200000ns, VDD,
+ 771282.300000ns, VSS,
+ 771882.700000ns, VSS,
+ 771882.800000ns, VDD,
+ 772483.200000ns, VDD,
+ 772483.300000ns, VSS,
+ 772723.400000ns, VSS,
+ 772723.500000ns, VDD,
+ 773203.800000ns, VDD,
+ 773203.900000ns, VSS,
+ 773684.200000ns, VSS,
+ 773684.300000ns, VDD,
+ 774524.900000ns, VDD,
+ 774525.000000ns, VSS,
+ 775605.800000ns, VSS,
+ 775605.900000ns, VDD,
+ 775846.000000ns, VDD,
+ 775846.100000ns, VSS,
+ 775966.100000ns, VSS,
+ 775966.200000ns, VDD,
+ 776686.700000ns, VDD,
+ 776686.800000ns, VSS,
+ 777887.700000ns, VSS,
+ 777887.800000ns, VDD,
+ 778248.000000ns, VDD,
+ 778248.100000ns, VSS,
+ 778848.500000ns, VSS,
+ 778848.600000ns, VDD,
+ 782571.600000ns, VDD,
+ 782571.700000ns, VSS,
+ 783292.200000ns, VSS,
+ 783292.300000ns, VDD,
+ 785093.700000ns, VDD,
+ 785093.800000ns, VSS,
+ 786895.200000ns, VSS,
+ 786895.300000ns, VDD,
+ 788696.700000ns, VDD,
+ 788696.800000ns, VSS,
+ 788816.800000ns, VSS,
+ 788816.900000ns, VDD,
+ 788936.900000ns, VDD,
+ 788937.000000ns, VSS,
+ 789177.100000ns, VSS,
+ 789177.200000ns, VDD,
+ 789297.200000ns, VDD,
+ 789297.300000ns, VSS,
+ 791579.100000ns, VSS,
+ 791579.200000ns, VDD,
+ 791819.300000ns, VDD,
+ 791819.400000ns, VSS,
+ 792900.200000ns, VSS,
+ 792900.300000ns, VDD,
+ 794341.400000ns, VDD,
+ 794341.500000ns, VSS,
+ 794701.700000ns, VSS,
+ 794701.800000ns, VDD,
+ 795182.100000ns, VDD,
+ 795182.200000ns, VSS,
+ 795302.200000ns, VSS,
+ 795302.300000ns, VDD,
+ 795422.300000ns, VDD,
+ 795422.400000ns, VSS,
+ 796142.900000ns, VSS,
+ 796143.000000ns, VDD,
+ 796863.500000ns, VDD,
+ 796863.600000ns, VSS,
+ 797584.100000ns, VSS,
+ 797584.200000ns, VDD,
+ 798064.500000ns, VDD,
+ 798064.600000ns, VSS,
+ 798184.600000ns, VSS,
+ 798184.700000ns, VDD,
+ 800826.800000ns, VDD,
+ 800826.900000ns, VSS,
+ 801787.600000ns, VSS,
+ 801787.700000ns, VDD,
+ 802268.000000ns, VDD,
+ 802268.100000ns, VSS,
+ 802508.200000ns, VSS,
+ 802508.300000ns, VDD,
+ 803348.900000ns, VDD,
+ 803349.000000ns, VSS,
+ 803829.300000ns, VSS,
+ 803829.400000ns, VDD,
+ 804429.800000ns, VDD,
+ 804429.900000ns, VSS,
+ 804790.100000ns, VSS,
+ 804790.200000ns, VDD,
+ 805390.600000ns, VDD,
+ 805390.700000ns, VSS,
+ 806231.300000ns, VSS,
+ 806231.400000ns, VDD,
+ 807432.300000ns, VDD,
+ 807432.400000ns, VSS,
+ 808753.400000ns, VSS,
+ 808753.500000ns, VDD,
+ 809353.900000ns, VDD,
+ 809354.000000ns, VSS,
+ 810194.600000ns, VSS,
+ 810194.700000ns, VDD,
+ 810314.700000ns, VDD,
+ 810314.800000ns, VSS,
+ 811635.800000ns, VSS,
+ 811635.900000ns, VDD,
+ 812116.200000ns, VDD,
+ 812116.300000ns, VSS,
+ 812956.900000ns, VSS,
+ 812957.000000ns, VDD,
+ 813077.000000ns, VDD,
+ 813077.100000ns, VSS,
+ 813437.300000ns, VSS,
+ 813437.400000ns, VDD,
+ 813677.500000ns, VDD,
+ 813677.600000ns, VSS,
+ 813917.700000ns, VSS,
+ 813917.800000ns, VDD,
+ 814878.500000ns, VDD,
+ 814878.600000ns, VSS,
+ 815479.000000ns, VSS,
+ 815479.100000ns, VDD,
+ 816199.600000ns, VDD,
+ 816199.700000ns, VSS,
+ 816800.100000ns, VSS,
+ 816800.200000ns, VDD,
+ 819562.400000ns, VDD,
+ 819562.500000ns, VSS,
+ 819802.600000ns, VSS,
+ 819802.700000ns, VDD,
+ 820042.800000ns, VDD,
+ 820042.900000ns, VSS,
+ 821003.600000ns, VSS,
+ 821003.700000ns, VDD,
+ 821964.400000ns, VDD,
+ 821964.500000ns, VSS,
+ 822084.500000ns, VSS,
+ 822084.600000ns, VDD,
+ 822685.000000ns, VDD,
+ 822685.100000ns, VSS,
+ 823165.400000ns, VSS,
+ 823165.500000ns, VDD,
+ 823886.000000ns, VDD,
+ 823886.100000ns, VSS,
+ 824006.100000ns, VSS,
+ 824006.200000ns, VDD,
+ 824126.200000ns, VDD,
+ 824126.300000ns, VSS,
+ 824486.500000ns, VSS,
+ 824486.600000ns, VDD,
+ 824726.700000ns, VDD,
+ 824726.800000ns, VSS,
+ 824846.800000ns, VSS,
+ 824846.900000ns, VDD,
+ 824966.900000ns, VDD,
+ 824967.000000ns, VSS,
+ 826528.200000ns, VSS,
+ 826528.300000ns, VDD,
+ 827008.600000ns, VDD,
+ 827008.700000ns, VSS,
+ 827128.700000ns, VSS,
+ 827128.800000ns, VDD,
+ 827248.800000ns, VDD,
+ 827248.900000ns, VSS,
+ 827969.400000ns, VSS,
+ 827969.500000ns, VDD,
+ 828329.700000ns, VDD,
+ 828329.800000ns, VSS,
+ 828690.000000ns, VSS,
+ 828690.100000ns, VDD,
+ 828930.200000ns, VDD,
+ 828930.300000ns, VSS,
+ 829050.300000ns, VSS,
+ 829050.400000ns, VDD,
+ 829170.400000ns, VDD,
+ 829170.500000ns, VSS,
+ 829530.700000ns, VSS,
+ 829530.800000ns, VDD,
+ 829650.800000ns, VDD,
+ 829650.900000ns, VSS,
+ 829770.900000ns, VSS,
+ 829771.000000ns, VDD,
+ 830731.700000ns, VDD,
+ 830731.800000ns, VSS,
+ 833013.600000ns, VSS,
+ 833013.700000ns, VDD,
+ 833734.200000ns, VDD,
+ 833734.300000ns, VSS,
+ 834935.200000ns, VSS,
+ 834935.300000ns, VDD,
+ 835415.600000ns, VDD,
+ 835415.700000ns, VSS,
+ 836496.500000ns, VSS,
+ 836496.600000ns, VDD,
+ 837097.000000ns, VDD,
+ 837097.100000ns, VSS,
+ 838298.000000ns, VSS,
+ 838298.100000ns, VDD,
+ 838778.400000ns, VDD,
+ 838778.500000ns, VSS,
+ 839018.600000ns, VSS,
+ 839018.700000ns, VDD,
+ 839739.200000ns, VDD,
+ 839739.300000ns, VSS,
+ 839979.400000ns, VSS,
+ 839979.500000ns, VDD,
+ 840700.000000ns, VDD,
+ 840700.100000ns, VSS,
+ 841540.700000ns, VSS,
+ 841540.800000ns, VDD,
+ 842021.100000ns, VDD,
+ 842021.200000ns, VSS,
+ 842261.300000ns, VSS,
+ 842261.400000ns, VDD,
+ 842861.800000ns, VDD,
+ 842861.900000ns, VSS,
+ 844182.900000ns, VSS,
+ 844183.000000ns, VDD,
+ 844663.300000ns, VDD,
+ 844663.400000ns, VSS,
+ 845383.900000ns, VSS,
+ 845384.000000ns, VDD,
+ 845984.400000ns, VDD,
+ 845984.500000ns, VSS,
+ 846464.800000ns, VSS,
+ 846464.900000ns, VDD,
+ 847785.900000ns, VDD,
+ 847786.000000ns, VSS,
+ 848626.600000ns, VSS,
+ 848626.700000ns, VDD,
+ 849107.000000ns, VDD,
+ 849107.100000ns, VSS,
+ 849587.400000ns, VSS,
+ 849587.500000ns, VDD,
+ 850668.300000ns, VDD,
+ 850668.400000ns, VSS,
+ 851869.300000ns, VSS,
+ 851869.400000ns, VDD,
+ 852830.100000ns, VDD,
+ 852830.200000ns, VSS,
+ 853070.300000ns, VSS,
+ 853070.400000ns, VDD,
+ 853911.000000ns, VDD,
+ 853911.100000ns, VSS,
+ 854511.500000ns, VSS,
+ 854511.600000ns, VDD,
+ 855592.400000ns, VDD,
+ 855592.500000ns, VSS,
+ 855832.600000ns, VSS,
+ 855832.700000ns, VDD,
+ 855952.700000ns, VDD,
+ 855952.800000ns, VSS,
+ 856553.200000ns, VSS,
+ 856553.300000ns, VDD,
+ 857153.700000ns, VDD,
+ 857153.800000ns, VSS,
+ 857634.100000ns, VSS,
+ 857634.200000ns, VDD,
+ 858234.600000ns, VDD,
+ 858234.700000ns, VSS,
+ 859195.400000ns, VSS,
+ 859195.500000ns, VDD,
+ 860996.900000ns, VDD,
+ 860997.000000ns, VSS,
+ 862077.800000ns, VSS,
+ 862077.900000ns, VDD,
+ 862318.000000ns, VDD,
+ 862318.100000ns, VSS,
+ 863038.600000ns, VSS,
+ 863038.700000ns, VDD,
+ 863519.000000ns, VDD,
+ 863519.100000ns, VSS,
+ 864239.600000ns, VSS,
+ 864239.700000ns, VDD,
+ 864960.200000ns, VDD,
+ 864960.300000ns, VSS,
+ 865680.800000ns, VSS,
+ 865680.900000ns, VDD,
+ 868082.800000ns, VDD,
+ 868082.900000ns, VSS,
+ 870244.600000ns, VSS,
+ 870244.700000ns, VDD,
+ 871685.800000ns, VDD,
+ 871685.900000ns, VSS,
+ 872766.700000ns, VSS,
+ 872766.800000ns, VDD,
+ 873247.100000ns, VDD,
+ 873247.200000ns, VSS,
+ 873487.300000ns, VSS,
+ 873487.400000ns, VDD,
+ 874688.300000ns, VDD,
+ 874688.400000ns, VSS,
+ 876489.800000ns, VSS,
+ 876489.900000ns, VDD,
+ 877090.300000ns, VDD,
+ 877090.400000ns, VSS,
+ 877810.900000ns, VSS,
+ 877811.000000ns, VDD,
+ 878171.200000ns, VDD,
+ 878171.300000ns, VSS,
+ 878411.400000ns, VSS,
+ 878411.500000ns, VDD,
+ 878531.500000ns, VDD,
+ 878531.600000ns, VSS,
+ 878771.700000ns, VSS,
+ 878771.800000ns, VDD,
+ 878891.800000ns, VDD,
+ 878891.900000ns, VSS,
+ 879372.200000ns, VSS,
+ 879372.300000ns, VDD,
+ 880092.800000ns, VDD,
+ 880092.900000ns, VSS,
+ 880212.900000ns, VSS,
+ 880213.000000ns, VDD,
+ 880333.000000ns, VDD,
+ 880333.100000ns, VSS,
+ 880693.300000ns, VSS,
+ 880693.400000ns, VDD,
+ 881173.700000ns, VDD,
+ 881173.800000ns, VSS,
+ 881534.000000ns, VSS,
+ 881534.100000ns, VDD,
+ 881894.300000ns, VDD,
+ 881894.400000ns, VSS,
+ 883215.400000ns, VSS,
+ 883215.500000ns, VDD,
+ 883815.900000ns, VDD,
+ 883816.000000ns, VSS,
+ 884776.700000ns, VSS,
+ 884776.800000ns, VDD,
+ 885377.200000ns, VDD,
+ 885377.300000ns, VSS,
+ 885857.600000ns, VSS,
+ 885857.700000ns, VDD,
+ 886578.200000ns, VDD,
+ 886578.300000ns, VSS,
+ 887659.100000ns, VSS,
+ 887659.200000ns, VDD,
+ 888259.600000ns, VDD,
+ 888259.700000ns, VSS,
+ 888619.900000ns, VSS,
+ 888620.000000ns, VDD,
+ 888980.200000ns, VDD,
+ 888980.300000ns, VSS,
+ 889580.700000ns, VSS,
+ 889580.800000ns, VDD,
+ 891382.200000ns, VDD,
+ 891382.300000ns, VSS,
+ 891502.300000ns, VSS,
+ 891502.400000ns, VDD,
+ 891622.400000ns, VDD,
+ 891622.500000ns, VSS,
+ 892222.900000ns, VSS,
+ 892223.000000ns, VDD,
+ 892823.400000ns, VDD,
+ 892823.500000ns, VSS,
+ 893183.700000ns, VSS,
+ 893183.800000ns, VDD,
+ 893664.100000ns, VDD,
+ 893664.200000ns, VSS,
+ 893904.300000ns, VSS,
+ 893904.400000ns, VDD,
+ 894384.700000ns, VDD,
+ 894384.800000ns, VSS,
+ 895946.000000ns, VSS,
+ 895946.100000ns, VDD,
+ 896066.100000ns, VDD,
+ 896066.200000ns, VSS,
+ 896426.400000ns, VSS,
+ 896426.500000ns, VDD,
+ 897387.200000ns, VDD,
+ 897387.300000ns, VSS,
+ 899068.600000ns, VSS,
+ 899068.700000ns, VDD,
+ 899549.000000ns, VDD,
+ 899549.100000ns, VSS,
+ 899669.100000ns, VSS,
+ 899669.200000ns, VDD,
+ 900269.600000ns, VDD,
+ 900269.700000ns, VSS,
+ 900509.800000ns, VSS,
+ 900509.900000ns, VDD,
+ 900629.900000ns, VDD,
+ 900630.000000ns, VSS,
+ 901230.400000ns, VSS,
+ 901230.500000ns, VDD,
+ 901951.000000ns, VDD,
+ 901951.100000ns, VSS,
+ 903031.900000ns, VSS,
+ 903032.000000ns, VDD,
+ 903272.100000ns, VDD,
+ 903272.200000ns, VSS,
+ 905554.000000ns, VSS,
+ 905554.100000ns, VDD,
+ 905674.100000ns, VDD,
+ 905674.200000ns, VSS,
+ 905794.200000ns, VSS,
+ 905794.300000ns, VDD,
+ 907595.700000ns, VDD,
+ 907595.800000ns, VSS,
+ 908076.100000ns, VSS,
+ 908076.200000ns, VDD,
+ 908796.700000ns, VDD,
+ 908796.800000ns, VSS,
+ 910478.100000ns, VSS,
+ 910478.200000ns, VDD,
+ 910838.400000ns, VDD,
+ 910838.500000ns, VSS,
+ 911679.100000ns, VSS,
+ 911679.200000ns, VDD,
+ 912880.100000ns, VDD,
+ 912880.200000ns, VSS,
+ 913360.500000ns, VSS,
+ 913360.600000ns, VDD,
+ 914321.300000ns, VDD,
+ 914321.400000ns, VSS,
+ 915162.000000ns, VSS,
+ 915162.100000ns, VDD,
+ 915402.200000ns, VDD,
+ 915402.300000ns, VSS,
+ 915642.400000ns, VSS,
+ 915642.500000ns, VDD,
+ 916843.400000ns, VDD,
+ 916843.500000ns, VSS,
+ 917083.600000ns, VSS,
+ 917083.700000ns, VDD,
+ 917443.900000ns, VDD,
+ 917444.000000ns, VSS,
+ 918044.400000ns, VSS,
+ 918044.500000ns, VDD,
+ 919125.300000ns, VDD,
+ 919125.400000ns, VSS,
+ 919365.500000ns, VSS,
+ 919365.600000ns, VDD,
+ 919485.600000ns, VDD,
+ 919485.700000ns, VSS,
+ 920566.500000ns, VSS,
+ 920566.600000ns, VDD,
+ 920806.700000ns, VDD,
+ 920806.800000ns, VSS,
+ 922007.700000ns, VSS,
+ 922007.800000ns, VDD,
+ 922488.100000ns, VDD,
+ 922488.200000ns, VSS,
+ 923809.200000ns, VSS,
+ 923809.300000ns, VDD,
+ 924169.500000ns, VDD,
+ 924169.600000ns, VSS,
+ 924529.800000ns, VSS,
+ 924529.900000ns, VDD,
+ 924649.900000ns, VDD,
+ 924650.000000ns, VSS,
+ 925971.000000ns, VSS,
+ 925971.100000ns, VDD,
+ 926691.600000ns, VDD,
+ 926691.700000ns, VSS,
+ 928132.800000ns, VSS,
+ 928132.900000ns, VDD,
+ 929453.900000ns, VDD,
+ 929454.000000ns, VSS,
+ 929934.300000ns, VSS,
+ 929934.400000ns, VDD,
+ 930775.000000ns, VDD,
+ 930775.100000ns, VSS,
+ 931495.600000ns, VSS,
+ 931495.700000ns, VDD,
+ 932336.300000ns, VDD,
+ 932336.400000ns, VSS,
+ 933777.500000ns, VSS,
+ 933777.600000ns, VDD,
+ 934378.000000ns, VDD,
+ 934378.100000ns, VSS,
+ 934498.100000ns, VSS,
+ 934498.200000ns, VDD,
+ 934858.400000ns, VDD,
+ 934858.500000ns, VSS,
+ 935098.600000ns, VSS,
+ 935098.700000ns, VDD,
+ 935338.800000ns, VDD,
+ 935338.900000ns, VSS,
+ 935579.000000ns, VSS,
+ 935579.100000ns, VDD,
+ 935819.200000ns, VDD,
+ 935819.300000ns, VSS,
+ 936539.800000ns, VSS,
+ 936539.900000ns, VDD,
+ 937020.200000ns, VDD,
+ 937020.300000ns, VSS,
+ 937380.500000ns, VSS,
+ 937380.600000ns, VDD,
+ 937860.900000ns, VDD,
+ 937861.000000ns, VSS,
+ 938341.300000ns, VSS,
+ 938341.400000ns, VDD,
+ 939422.200000ns, VDD,
+ 939422.300000ns, VSS,
+ 940022.700000ns, VSS,
+ 940022.800000ns, VDD,
+ 940383.000000ns, VDD,
+ 940383.100000ns, VSS,
+ 943745.800000ns, VSS,
+ 943745.900000ns, VDD,
+ 944586.500000ns, VDD,
+ 944586.600000ns, VSS,
+ 945187.000000ns, VSS,
+ 945187.100000ns, VDD,
+ 945667.400000ns, VDD,
+ 945667.500000ns, VSS,
+ 948669.900000ns, VSS,
+ 948670.000000ns, VDD,
+ 949870.900000ns, VDD,
+ 949871.000000ns, VSS,
+ 950951.800000ns, VSS,
+ 950951.900000ns, VDD,
+ 951312.100000ns, VDD,
+ 951312.200000ns, VSS,
+ 951432.200000ns, VSS,
+ 951432.300000ns, VDD,
+ 951672.400000ns, VDD,
+ 951672.500000ns, VSS,
+ 952032.700000ns, VSS,
+ 952032.800000ns, VDD,
+ 952753.300000ns, VDD,
+ 952753.400000ns, VSS,
+ 953233.700000ns, VSS,
+ 953233.800000ns, VDD,
+ 953954.300000ns, VDD,
+ 953954.400000ns, VSS,
+ 954194.500000ns, VSS,
+ 954194.600000ns, VDD,
+ 954314.600000ns, VDD,
+ 954314.700000ns, VSS,
+ 954915.100000ns, VSS,
+ 954915.200000ns, VDD,
+ 955515.600000ns, VDD,
+ 955515.700000ns, VSS,
+ 957076.900000ns, VSS,
+ 957077.000000ns, VDD,
+ 957917.600000ns, VDD,
+ 957917.700000ns, VSS,
+ 958398.000000ns, VSS,
+ 958398.100000ns, VDD,
+ 958998.500000ns, VDD,
+ 958998.600000ns, VSS,
+ 959599.000000ns, VSS,
+ 959599.100000ns, VDD,
+ 960920.100000ns, VDD,
+ 960920.200000ns, VSS,
+ 961280.400000ns, VSS,
+ 961280.500000ns, VDD,
+ 961760.800000ns, VDD,
+ 961760.900000ns, VSS,
+ 962241.200000ns, VSS,
+ 962241.300000ns, VDD,
+ 962721.600000ns, VDD,
+ 962721.700000ns, VSS,
+ 963081.900000ns, VSS,
+ 963082.000000ns, VDD,
+ 963202.000000ns, VDD,
+ 963202.100000ns, VSS,
+ 963802.500000ns, VSS,
+ 963802.600000ns, VDD,
+ 964403.000000ns, VDD,
+ 964403.100000ns, VSS,
+ 965724.100000ns, VSS,
+ 965724.200000ns, VDD,
+ 966204.500000ns, VDD,
+ 966204.600000ns, VSS,
+ 967045.200000ns, VSS,
+ 967045.300000ns, VDD,
+ 967885.900000ns, VDD,
+ 967886.000000ns, VSS,
+ 968606.500000ns, VSS,
+ 968606.600000ns, VDD,
+ 969207.000000ns, VDD,
+ 969207.100000ns, VSS,
+ 969687.400000ns, VSS,
+ 969687.500000ns, VDD,
+ 970648.200000ns, VDD,
+ 970648.300000ns, VSS,
+ 971128.600000ns, VSS,
+ 971128.700000ns, VDD,
+ 971729.100000ns, VDD,
+ 971729.200000ns, VSS,
+ 972089.400000ns, VSS,
+ 972089.500000ns, VDD,
+ 972329.600000ns, VDD,
+ 972329.700000ns, VSS,
+ 972810.000000ns, VSS,
+ 972810.100000ns, VDD,
+ 973170.300000ns, VDD,
+ 973170.400000ns, VSS,
+ 973650.700000ns, VSS,
+ 973650.800000ns, VDD,
+ 974131.100000ns, VDD,
+ 974131.200000ns, VSS,
+ 974611.500000ns, VSS,
+ 974611.600000ns, VDD,
+ 974851.700000ns, VDD,
+ 974851.800000ns, VSS,
+ 974971.800000ns, VSS,
+ 974971.900000ns, VDD,
+ 975572.300000ns, VDD,
+ 975572.400000ns, VSS,
+ 975932.600000ns, VSS,
+ 975932.700000ns, VDD,
+ 976052.700000ns, VDD,
+ 976052.800000ns, VSS,
+ 976773.300000ns, VSS,
+ 976773.400000ns, VDD,
+ 977614.000000ns, VDD,
+ 977614.100000ns, VSS,
+ 977734.100000ns, VSS,
+ 977734.200000ns, VDD,
+ 978214.500000ns, VDD,
+ 978214.600000ns, VSS,
+ 978574.800000ns, VSS,
+ 978574.900000ns, VDD,
+ 979415.500000ns, VDD,
+ 979415.600000ns, VSS,
+ 979775.800000ns, VSS,
+ 979775.900000ns, VDD,
+ 980736.600000ns, VDD,
+ 980736.700000ns, VSS,
+ 981817.500000ns, VSS,
+ 981817.600000ns, VDD,
+ 982057.700000ns, VDD,
+ 982057.800000ns, VSS,
+ 982297.900000ns, VSS,
+ 982298.000000ns, VDD,
+ 984219.500000ns, VDD,
+ 984219.600000ns, VSS,
+ 984699.900000ns, VSS,
+ 984700.000000ns, VDD,
+ 987702.400000ns, VDD,
+ 987702.500000ns, VSS,
+ 987942.600000ns, VSS,
+ 987942.700000ns, VDD,
+ 988182.800000ns, VDD,
+ 988182.900000ns, VSS,
+ 988543.100000ns, VSS,
+ 988543.200000ns, VDD,
+ 990224.500000ns, VDD,
+ 990224.600000ns, VSS,
+ 990344.600000ns, VSS,
+ 990344.700000ns, VDD,
+ 990584.800000ns, VDD,
+ 990584.900000ns, VSS,
+ 990704.900000ns, VSS,
+ 990705.000000ns, VDD,
+ 991185.300000ns, VDD,
+ 991185.400000ns, VSS,
+ 991665.700000ns, VSS,
+ 991665.800000ns, VDD,
+ 992266.200000ns, VDD,
+ 992266.300000ns, VSS,
+ 992386.300000ns, VSS,
+ 992386.400000ns, VDD,
+ 993707.400000ns, VDD,
+ 993707.500000ns, VSS,
+ 993947.600000ns, VSS,
+ 993947.700000ns, VDD,
+ 994428.000000ns, VDD,
+ 994428.100000ns, VSS,
+ 995148.600000ns, VSS,
+ 995148.700000ns, VDD,
+ 997070.200000ns, VDD,
+ 997070.300000ns, VSS,
+ 997670.700000ns, VSS,
+ 997670.800000ns, VDD,
+ 998151.100000ns, VDD,
+ 998151.200000ns, VSS,
+ 998991.800000ns, VSS,
+ 998991.900000ns, VDD,
+ 999111.900000ns, VDD,
+ 999112.000000ns, VSS,
+ 999232.000000ns, VSS,
+ 999232.100000ns, VDD,
+ 1000072.700000ns, VDD,
+ 1000072.800000ns, VSS,
+ 1000192.800000ns, VSS,
+ 1000192.900000ns, VDD,
+ 1001754.100000ns, VDD,
+ 1001754.200000ns, VSS,
+ 1002354.600000ns, VSS,
+ 1002354.700000ns, VDD,
+ 1002594.800000ns, VDD,
+ 1002594.900000ns, VSS,
+ 1002955.100000ns, VSS,
+ 1002955.200000ns, VDD,
+ 1003195.300000ns, VDD,
+ 1003195.400000ns, VSS,
+ 1003435.500000ns, VSS,
+ 1003435.600000ns, VDD,
+ 1005237.000000ns, VDD,
+ 1005237.100000ns, VSS,
+ 1006077.700000ns, VSS,
+ 1006077.800000ns, VDD,
+ 1007398.800000ns, VDD,
+ 1007398.900000ns, VSS,
+ 1008359.600000ns, VSS,
+ 1008359.700000ns, VDD,
+ 1009080.200000ns, VDD,
+ 1009080.300000ns, VSS,
+ 1009920.900000ns, VSS,
+ 1009921.000000ns, VDD,
+ 1010281.200000ns, VDD,
+ 1010281.300000ns, VSS,
+ 1010641.500000ns, VSS,
+ 1010641.600000ns, VDD,
+ 1011121.900000ns, VDD,
+ 1011122.000000ns, VSS,
+ 1011362.100000ns, VSS,
+ 1011362.200000ns, VDD,
+ 1011482.200000ns, VDD,
+ 1011482.300000ns, VSS,
+ 1012803.300000ns, VSS,
+ 1012803.400000ns, VDD,
+ 1013283.700000ns, VDD,
+ 1013283.800000ns, VSS,
+ 1014364.600000ns, VSS,
+ 1014364.700000ns, VDD,
+ 1014724.900000ns, VDD,
+ 1014725.000000ns, VSS,
+ 1015685.700000ns, VSS,
+ 1015685.800000ns, VDD,
+ 1016166.100000ns, VDD,
+ 1016166.200000ns, VSS,
+ 1017126.900000ns, VSS,
+ 1017127.000000ns, VDD,
+ 1019408.800000ns, VDD,
+ 1019408.900000ns, VSS,
+ 1020970.100000ns, VSS,
+ 1020970.200000ns, VDD,
+ 1021210.300000ns, VDD,
+ 1021210.400000ns, VSS,
+ 1021690.700000ns, VSS,
+ 1021690.800000ns, VDD,
+ 1023732.400000ns, VDD,
+ 1023732.500000ns, VSS,
+ 1024453.000000ns, VSS,
+ 1024453.100000ns, VDD,
+ 1025293.700000ns, VDD,
+ 1025293.800000ns, VSS,
+ 1026014.300000ns, VSS,
+ 1026014.400000ns, VDD,
+ 1027095.200000ns, VDD,
+ 1027095.300000ns, VSS,
+ 1027575.600000ns, VSS,
+ 1027575.700000ns, VDD,
+ 1027935.900000ns, VDD,
+ 1027936.000000ns, VSS,
+ 1030578.100000ns, VSS,
+ 1030578.200000ns, VDD,
+ 1030698.200000ns, VDD,
+ 1030698.300000ns, VSS,
+ 1030938.400000ns, VSS,
+ 1030938.500000ns, VDD,
+ 1032139.400000ns, VDD,
+ 1032139.500000ns, VSS,
+ 1032499.700000ns, VSS,
+ 1032499.800000ns, VDD,
+ 1032739.900000ns, VDD,
+ 1032740.000000ns, VSS,
+ 1033580.600000ns, VSS,
+ 1033580.700000ns, VDD,
+ 1034181.100000ns, VDD,
+ 1034181.200000ns, VSS,
+ 1034301.200000ns, VSS,
+ 1034301.300000ns, VDD,
+ 1035141.900000ns, VDD,
+ 1035142.000000ns, VSS,
+ 1036102.700000ns, VSS,
+ 1036102.800000ns, VDD,
+ 1036342.900000ns, VDD,
+ 1036343.000000ns, VSS,
+ 1036463.000000ns, VSS,
+ 1036463.100000ns, VDD,
+ 1037183.600000ns, VDD,
+ 1037183.700000ns, VSS,
+ 1037664.000000ns, VSS,
+ 1037664.100000ns, VDD,
+ 1039225.300000ns, VDD,
+ 1039225.400000ns, VSS,
+ 1039945.900000ns, VSS,
+ 1039946.000000ns, VDD,
+ 1040186.100000ns, VDD,
+ 1040186.200000ns, VSS,
+ 1040306.200000ns, VSS,
+ 1040306.300000ns, VDD,
+ 1040426.300000ns, VDD,
+ 1040426.400000ns, VSS,
+ 1041987.600000ns, VSS,
+ 1041987.700000ns, VDD,
+ 1042107.700000ns, VDD,
+ 1042107.800000ns, VSS,
+ 1042828.300000ns, VSS,
+ 1042828.400000ns, VDD,
+ 1043068.500000ns, VDD,
+ 1043068.600000ns, VSS,
+ 1043428.800000ns, VSS,
+ 1043428.900000ns, VDD,
+ 1044870.000000ns, VDD,
+ 1044870.100000ns, VSS,
+ 1046551.400000ns, VSS,
+ 1046551.500000ns, VDD,
+ 1047031.800000ns, VDD,
+ 1047031.900000ns, VSS,
+ 1047392.100000ns, VSS,
+ 1047392.200000ns, VDD,
+ 1047872.500000ns, VDD,
+ 1047872.600000ns, VSS,
+ 1048473.000000ns, VSS,
+ 1048473.100000ns, VDD,
+ 1049433.800000ns, VDD,
+ 1049433.900000ns, VSS,
+ 1050394.600000ns, VSS,
+ 1050394.700000ns, VDD,
+ 1052436.300000ns, VDD,
+ 1052436.400000ns, VSS,
+ 1052916.700000ns, VSS,
+ 1052916.800000ns, VDD,
+ 1053277.000000ns, VDD,
+ 1053277.100000ns, VSS,
+ 1053877.500000ns, VSS,
+ 1053877.600000ns, VDD,
+ 1054357.900000ns, VDD,
+ 1054358.000000ns, VSS,
+ 1055318.700000ns, VSS,
+ 1055318.800000ns, VDD,
+ 1055679.000000ns, VDD,
+ 1055679.100000ns, VSS,
+ 1056159.400000ns, VSS,
+ 1056159.500000ns, VDD,
+ 1056279.500000ns, VDD,
+ 1056279.600000ns, VSS,
+ 1056399.600000ns, VSS,
+ 1056399.700000ns, VDD,
+ 1056880.000000ns, VDD,
+ 1056880.100000ns, VSS,
+ 1058801.600000ns, VSS,
+ 1058801.700000ns, VDD,
+ 1059282.000000ns, VDD,
+ 1059282.100000ns, VSS,
+ 1059762.400000ns, VSS,
+ 1059762.500000ns, VDD,
+ 1060242.800000ns, VDD,
+ 1060242.900000ns, VSS,
+ 1060843.300000ns, VSS,
+ 1060843.400000ns, VDD,
+ 1060963.400000ns, VDD,
+ 1060963.500000ns, VSS,
+ 1061203.600000ns, VSS,
+ 1061203.700000ns, VDD,
+ 1061323.700000ns, VDD,
+ 1061323.800000ns, VSS,
+ 1063125.200000ns, VSS,
+ 1063125.300000ns, VDD,
+ 1064686.500000ns, VDD,
+ 1064686.600000ns, VSS,
+ 1065287.000000ns, VSS,
+ 1065287.100000ns, VDD,
+ 1065767.400000ns, VDD,
+ 1065767.500000ns, VSS,
+ 1065887.500000ns, VSS,
+ 1065887.600000ns, VDD,
+ 1067328.700000ns, VDD,
+ 1067328.800000ns, VSS,
+ 1068649.800000ns, VSS,
+ 1068649.900000ns, VDD,
+ 1069730.700000ns, VDD,
+ 1069730.800000ns, VSS,
+ 1070931.700000ns, VSS,
+ 1070931.800000ns, VDD,
+ 1071051.800000ns, VDD,
+ 1071051.900000ns, VSS,
+ 1072132.700000ns, VSS,
+ 1072132.800000ns, VDD,
+ 1072613.100000ns, VDD,
+ 1072613.200000ns, VSS,
+ 1074054.300000ns, VSS,
+ 1074054.400000ns, VDD,
+ 1074174.400000ns, VDD,
+ 1074174.500000ns, VSS,
+ 1074294.500000ns, VSS,
+ 1074294.600000ns, VDD,
+ 1074774.900000ns, VDD,
+ 1074775.000000ns, VSS,
+ 1075135.200000ns, VSS,
+ 1075135.300000ns, VDD,
+ 1076336.200000ns, VDD,
+ 1076336.300000ns, VSS,
+ 1077297.000000ns, VSS,
+ 1077297.100000ns, VDD,
+ 1077417.100000ns, VDD,
+ 1077417.200000ns, VSS,
+ 1077777.400000ns, VSS,
+ 1077777.500000ns, VDD,
+ 1078738.200000ns, VDD,
+ 1078738.300000ns, VSS,
+ 1079338.700000ns, VSS,
+ 1079338.800000ns, VDD,
+ 1079578.900000ns, VDD,
+ 1079579.000000ns, VSS,
+ 1079819.100000ns, VSS,
+ 1079819.200000ns, VDD,
+ 1080419.600000ns, VDD,
+ 1080419.700000ns, VSS,
+ 1080659.800000ns, VSS,
+ 1080659.900000ns, VDD,
+ 1081140.200000ns, VDD,
+ 1081140.300000ns, VSS,
+ 1081620.600000ns, VSS,
+ 1081620.700000ns, VDD,
+ 1081860.800000ns, VDD,
+ 1081860.900000ns, VSS,
+ 1081980.900000ns, VSS,
+ 1081981.000000ns, VDD,
+ 1082221.100000ns, VDD,
+ 1082221.200000ns, VSS,
+ 1082581.400000ns, VSS,
+ 1082581.500000ns, VDD,
+ 1083302.000000ns, VDD,
+ 1083302.100000ns, VSS,
+ 1083542.200000ns, VSS,
+ 1083542.300000ns, VDD,
+ 1083662.300000ns, VDD,
+ 1083662.400000ns, VSS,
+ 1084262.800000ns, VSS,
+ 1084262.900000ns, VDD,
+ 1085704.000000ns, VDD,
+ 1085704.100000ns, VSS,
+ 1086424.600000ns, VSS,
+ 1086424.700000ns, VDD,
+ 1087145.200000ns, VDD,
+ 1087145.300000ns, VSS,
+ 1087385.400000ns, VSS,
+ 1087385.500000ns, VDD,
+ 1087865.800000ns, VDD,
+ 1087865.900000ns, VSS,
+ 1088706.500000ns, VSS,
+ 1088706.600000ns, VDD,
+ 1089787.400000ns, VDD,
+ 1089787.500000ns, VSS,
+ 1090027.600000ns, VSS,
+ 1090027.700000ns, VDD,
+ 1090267.800000ns, VDD,
+ 1090267.900000ns, VSS,
+ 1090387.900000ns, VSS,
+ 1090388.000000ns, VDD,
+ 1090508.000000ns, VDD,
+ 1090508.100000ns, VSS,
+ 1090988.400000ns, VSS,
+ 1090988.500000ns, VDD,
+ 1091108.500000ns, VDD,
+ 1091108.600000ns, VSS,
+ 1092429.600000ns, VSS,
+ 1092429.700000ns, VDD,
+ 1094591.400000ns, VDD,
+ 1094591.500000ns, VSS,
+ 1096272.800000ns, VSS,
+ 1096272.900000ns, VDD,
+ 1096392.900000ns, VDD,
+ 1096393.000000ns, VSS,
+ 1096633.100000ns, VSS,
+ 1096633.200000ns, VDD,
+ 1097233.600000ns, VDD,
+ 1097233.700000ns, VSS,
+ 1097353.700000ns, VSS,
+ 1097353.800000ns, VDD,
+ 1097834.100000ns, VDD,
+ 1097834.200000ns, VSS,
+ 1098194.400000ns, VSS,
+ 1098194.500000ns, VDD,
+ 1098314.500000ns, VDD,
+ 1098314.600000ns, VSS,
+ 1098674.800000ns, VSS,
+ 1098674.900000ns, VDD,
+ 1099635.600000ns, VDD,
+ 1099635.700000ns, VSS,
+ 1099875.800000ns, VSS,
+ 1099875.900000ns, VDD,
+ 1099995.900000ns, VDD,
+ 1099996.000000ns, VSS,
+ 1100836.600000ns, VSS,
+ 1100836.700000ns, VDD,
+ 1101196.900000ns, VDD,
+ 1101197.000000ns, VSS,
+ 1102157.700000ns, VSS,
+ 1102157.800000ns, VDD,
+ 1102518.000000ns, VDD,
+ 1102518.100000ns, VSS,
+ 1103598.900000ns, VSS,
+ 1103599.000000ns, VDD,
+ 1103839.100000ns, VDD,
+ 1103839.200000ns, VSS,
+ 1103959.200000ns, VSS,
+ 1103959.300000ns, VDD,
+ 1104079.300000ns, VDD,
+ 1104079.400000ns, VSS,
+ 1104799.900000ns, VSS,
+ 1104800.000000ns, VDD,
+ 1105040.100000ns, VDD,
+ 1105040.200000ns, VSS,
+ 1106241.100000ns, VSS,
+ 1106241.200000ns, VDD,
+ 1107322.000000ns, VDD,
+ 1107322.100000ns, VSS,
+ 1107922.500000ns, VSS,
+ 1107922.600000ns, VDD,
+ 1108282.800000ns, VDD,
+ 1108282.900000ns, VSS,
+ 1109003.400000ns, VSS,
+ 1109003.500000ns, VDD,
+ 1110684.800000ns, VDD,
+ 1110684.900000ns, VSS,
+ 1111765.700000ns, VSS,
+ 1111765.800000ns, VDD,
+ 1112126.000000ns, VDD,
+ 1112126.100000ns, VSS,
+ 1113567.200000ns, VSS,
+ 1113567.300000ns, VDD,
+ 1114167.700000ns, VDD,
+ 1114167.800000ns, VSS,
+ 1114648.100000ns, VSS,
+ 1114648.200000ns, VDD,
+ 1115128.500000ns, VDD,
+ 1115128.600000ns, VSS,
+ 1115969.200000ns, VSS,
+ 1115969.300000ns, VDD,
+ 1116689.800000ns, VDD,
+ 1116689.900000ns, VSS,
+ 1116930.000000ns, VSS,
+ 1116930.100000ns, VDD,
+ 1117050.100000ns, VDD,
+ 1117050.200000ns, VSS,
+ 1117170.200000ns, VSS,
+ 1117170.300000ns, VDD,
+ 1118010.900000ns, VDD,
+ 1118011.000000ns, VSS,
+ 1118371.200000ns, VSS,
+ 1118371.300000ns, VDD,
+ 1119572.200000ns, VDD,
+ 1119572.300000ns, VSS,
+ 1120052.600000ns, VSS,
+ 1120052.700000ns, VDD,
+ 1120653.100000ns, VDD,
+ 1120653.200000ns, VSS,
+ 1120893.300000ns, VSS,
+ 1120893.400000ns, VDD,
+ 1121013.400000ns, VDD,
+ 1121013.500000ns, VSS,
+ 1122094.300000ns, VSS,
+ 1122094.400000ns, VDD,
+ 1123655.600000ns, VDD,
+ 1123655.700000ns, VSS,
+ 1123895.800000ns, VSS,
+ 1123895.900000ns, VDD,
+ 1124616.400000ns, VDD,
+ 1124616.500000ns, VSS,
+ 1125337.000000ns, VSS,
+ 1125337.100000ns, VDD,
+ 1127018.400000ns, VDD,
+ 1127018.500000ns, VSS,
+ 1127859.100000ns, VSS,
+ 1127859.200000ns, VDD,
+ 1128579.700000ns, VDD,
+ 1128579.800000ns, VSS,
+ 1130141.000000ns, VSS,
+ 1130141.100000ns, VDD,
+ 1130381.200000ns, VDD,
+ 1130381.300000ns, VSS,
+ 1130501.300000ns, VSS,
+ 1130501.400000ns, VDD,
+ 1130621.400000ns, VDD,
+ 1130621.500000ns, VSS,
+ 1131942.500000ns, VSS,
+ 1131942.600000ns, VDD,
+ 1132903.300000ns, VDD,
+ 1132903.400000ns, VSS,
+ 1133984.200000ns, VSS,
+ 1133984.300000ns, VDD,
+ 1134704.800000ns, VDD,
+ 1134704.900000ns, VSS,
+ 1136025.900000ns, VSS,
+ 1136026.000000ns, VDD,
+ 1136866.600000ns, VDD,
+ 1136866.700000ns, VSS,
+ 1137106.800000ns, VSS,
+ 1137106.900000ns, VDD,
+ 1137226.900000ns, VDD,
+ 1137227.000000ns, VSS,
+ 1137587.200000ns, VSS,
+ 1137587.300000ns, VDD,
+ 1137707.300000ns, VDD,
+ 1137707.400000ns, VSS,
+ 1139508.800000ns, VSS,
+ 1139508.900000ns, VDD,
+ 1140109.300000ns, VDD,
+ 1140109.400000ns, VSS,
+ 1140229.400000ns, VSS,
+ 1140229.500000ns, VDD,
+ 1141310.300000ns, VDD,
+ 1141310.400000ns, VSS,
+ 1142391.200000ns, VSS,
+ 1142391.300000ns, VDD,
+ 1142751.500000ns, VDD,
+ 1142751.600000ns, VSS,
+ 1142871.600000ns, VSS,
+ 1142871.700000ns, VDD,
+ 1143712.300000ns, VDD,
+ 1143712.400000ns, VSS,
+ 1143832.400000ns, VSS,
+ 1143832.500000ns, VDD,
+ 1144432.900000ns, VDD,
+ 1144433.000000ns, VSS,
+ 1145393.700000ns, VSS,
+ 1145393.800000ns, VDD,
+ 1146354.500000ns, VDD,
+ 1146354.600000ns, VSS,
+ 1146474.600000ns, VSS,
+ 1146474.700000ns, VDD,
+ 1146594.700000ns, VDD,
+ 1146594.800000ns, VSS,
+ 1147075.100000ns, VSS,
+ 1147075.200000ns, VDD,
+ 1148035.900000ns, VDD,
+ 1148036.000000ns, VSS,
+ 1148156.000000ns, VSS,
+ 1148156.100000ns, VDD,
+ 1149116.800000ns, VDD,
+ 1149116.900000ns, VSS,
+ 1149236.900000ns, VSS,
+ 1149237.000000ns, VDD,
+ 1150077.600000ns, VDD,
+ 1150077.700000ns, VSS,
+ 1150197.700000ns, VSS,
+ 1150197.800000ns, VDD,
+ 1150317.800000ns, VDD,
+ 1150317.900000ns, VSS,
+ 1150798.200000ns, VSS,
+ 1150798.300000ns, VDD,
+ 1151158.500000ns, VDD,
+ 1151158.600000ns, VSS,
+ 1151759.000000ns, VSS,
+ 1151759.100000ns, VDD,
+ 1152239.400000ns, VDD,
+ 1152239.500000ns, VSS,
+ 1152839.900000ns, VSS,
+ 1152840.000000ns, VDD,
+ 1153440.400000ns, VDD,
+ 1153440.500000ns, VSS,
+ 1154521.300000ns, VSS,
+ 1154521.400000ns, VDD,
+ 1154761.500000ns, VDD,
+ 1154761.600000ns, VSS,
+ 1155001.700000ns, VSS,
+ 1155001.800000ns, VDD,
+ 1155121.800000ns, VDD,
+ 1155121.900000ns, VSS,
+ 1156082.600000ns, VSS,
+ 1156082.700000ns, VDD,
+ 1156563.000000ns, VDD,
+ 1156563.100000ns, VSS,
+ 1156803.200000ns, VSS,
+ 1156803.300000ns, VDD,
+ 1156923.300000ns, VDD,
+ 1156923.400000ns, VSS,
+ 1157043.400000ns, VSS,
+ 1157043.500000ns, VDD,
+ 1157283.600000ns, VDD,
+ 1157283.700000ns, VSS,
+ 1157764.000000ns, VSS,
+ 1157764.100000ns, VDD,
+ 1158124.300000ns, VDD,
+ 1158124.400000ns, VSS,
+ 1159445.400000ns, VSS,
+ 1159445.500000ns, VDD,
+ 1159565.500000ns, VDD,
+ 1159565.600000ns, VSS,
+ 1159685.600000ns, VSS,
+ 1159685.700000ns, VDD,
+ 1160526.300000ns, VDD,
+ 1160526.400000ns, VSS,
+ 1162327.800000ns, VSS,
+ 1162327.900000ns, VDD,
+ 1162808.200000ns, VDD,
+ 1162808.300000ns, VSS,
+ 1163769.000000ns, VSS,
+ 1163769.100000ns, VDD,
+ 1165450.400000ns, VDD,
+ 1165450.500000ns, VSS,
+ 1166050.900000ns, VSS,
+ 1166051.000000ns, VDD,
+ 1166171.000000ns, VDD,
+ 1166171.100000ns, VSS,
+ 1166291.100000ns, VSS,
+ 1166291.200000ns, VDD,
+ 1166531.300000ns, VDD,
+ 1166531.400000ns, VSS,
+ 1166651.400000ns, VSS,
+ 1166651.500000ns, VDD,
+ 1167011.700000ns, VDD,
+ 1167011.800000ns, VSS,
+ 1167131.800000ns, VSS,
+ 1167131.900000ns, VDD,
+ 1167852.400000ns, VDD,
+ 1167852.500000ns, VSS,
+ 1168332.800000ns, VSS,
+ 1168332.900000ns, VDD,
+ 1170374.500000ns, VDD,
+ 1170374.600000ns, VSS,
+ 1170975.000000ns, VSS,
+ 1170975.100000ns, VDD,
+ 1173016.700000ns, VDD,
+ 1173016.800000ns, VSS,
+ 1174578.000000ns, VSS,
+ 1174578.100000ns, VDD,
+ 1174698.100000ns, VDD,
+ 1174698.200000ns, VSS,
+ 1174818.200000ns, VSS,
+ 1174818.300000ns, VDD,
+ 1175298.600000ns, VDD,
+ 1175298.700000ns, VSS,
+ 1175658.900000ns, VSS,
+ 1175659.000000ns, VDD,
+ 1177100.100000ns, VDD,
+ 1177100.200000ns, VSS,
+ 1177220.200000ns, VSS,
+ 1177220.300000ns, VDD,
+ 1177340.300000ns, VDD,
+ 1177340.400000ns, VSS,
+ 1178421.200000ns, VSS,
+ 1178421.300000ns, VDD,
+ 1179982.500000ns, VDD,
+ 1179982.600000ns, VSS,
+ 1180462.900000ns, VSS,
+ 1180463.000000ns, VDD,
+ 1180823.200000ns, VDD,
+ 1180823.300000ns, VSS,
+ 1181303.600000ns, VSS,
+ 1181303.700000ns, VDD,
+ 1181904.100000ns, VDD,
+ 1181904.200000ns, VSS,
+ 1182384.500000ns, VSS,
+ 1182384.600000ns, VDD,
+ 1183585.500000ns, VDD,
+ 1183585.600000ns, VSS,
+ 1183945.800000ns, VSS,
+ 1183945.900000ns, VDD,
+ 1184426.200000ns, VDD,
+ 1184426.300000ns, VSS,
+ 1184666.400000ns, VSS,
+ 1184666.500000ns, VDD,
+ 1185747.300000ns, VDD,
+ 1185747.400000ns, VSS,
+ 1188389.500000ns, VSS,
+ 1188389.600000ns, VDD,
+ 1189470.400000ns, VDD,
+ 1189470.500000ns, VSS,
+ 1191512.100000ns, VSS,
+ 1191512.200000ns, VDD,
+ 1192112.600000ns, VDD,
+ 1192112.700000ns, VSS,
+ 1192352.800000ns, VSS,
+ 1192352.900000ns, VDD,
+ 1192593.000000ns, VDD,
+ 1192593.100000ns, VSS,
+ 1192713.100000ns, VSS,
+ 1192713.200000ns, VDD,
+ 1193914.100000ns, VDD,
+ 1193914.200000ns, VSS,
+ 1194154.300000ns, VSS,
+ 1194154.400000ns, VDD,
+ 1194514.600000ns, VDD,
+ 1194514.700000ns, VSS,
+ 1194995.000000ns, VSS,
+ 1194995.100000ns, VDD,
+ 1195115.100000ns, VDD,
+ 1195115.200000ns, VSS,
+ 1197877.400000ns, VSS,
+ 1197877.500000ns, VDD,
+ 1199438.700000ns, VDD,
+ 1199438.800000ns, VSS,
+ 1200159.300000ns, VSS,
+ 1200159.400000ns, VDD,
+ 1200639.700000ns, VDD,
+ 1200639.800000ns, VSS,
+ 1200879.900000ns, VSS,
+ 1200880.000000ns, VDD,
+ 1202201.000000ns, VDD,
+ 1202201.100000ns, VSS,
+ 1202561.300000ns, VSS,
+ 1202561.400000ns, VDD,
+ 1203041.700000ns, VDD,
+ 1203041.800000ns, VSS,
+ 1203882.400000ns, VSS,
+ 1203882.500000ns, VDD,
+ 1205083.400000ns, VDD,
+ 1205083.500000ns, VSS,
+ 1205563.800000ns, VSS,
+ 1205563.900000ns, VDD,
+ 1206164.300000ns, VDD,
+ 1206164.400000ns, VSS,
+ 1206524.600000ns, VSS,
+ 1206524.700000ns, VDD,
+ 1206644.700000ns, VDD,
+ 1206644.800000ns, VSS,
+ 1206884.900000ns, VSS,
+ 1206885.000000ns, VDD,
+ 1207005.000000ns, VDD,
+ 1207005.100000ns, VSS,
+ 1207125.100000ns, VSS,
+ 1207125.200000ns, VDD,
+ 1207245.200000ns, VDD,
+ 1207245.300000ns, VSS,
+ 1207365.300000ns, VSS,
+ 1207365.400000ns, VDD,
+ 1207845.700000ns, VDD,
+ 1207845.800000ns, VSS,
+ 1207965.800000ns, VSS,
+ 1207965.900000ns, VDD,
+ 1208326.100000ns, VDD,
+ 1208326.200000ns, VSS,
+ 1208566.300000ns, VSS,
+ 1208566.400000ns, VDD,
+ 1209166.800000ns, VDD,
+ 1209166.900000ns, VSS,
+ 1209527.100000ns, VSS,
+ 1209527.200000ns, VDD,
+ 1209767.300000ns, VDD,
+ 1209767.400000ns, VSS,
+ 1210007.500000ns, VSS,
+ 1210007.600000ns, VDD,
+ 1210968.300000ns, VDD,
+ 1210968.400000ns, VSS,
+ 1212409.500000ns, VSS,
+ 1212409.600000ns, VDD,
+ 1212889.900000ns, VDD,
+ 1212890.000000ns, VSS,
+ 1213250.200000ns, VSS,
+ 1213250.300000ns, VDD,
+ 1213370.300000ns, VDD,
+ 1213370.400000ns, VSS,
+ 1213610.500000ns, VSS,
+ 1213610.600000ns, VDD,
+ 1213850.700000ns, VDD,
+ 1213850.800000ns, VSS,
+ 1214811.500000ns, VSS,
+ 1214811.600000ns, VDD,
+ 1215051.700000ns, VDD,
+ 1215051.800000ns, VSS,
+ 1215532.100000ns, VSS,
+ 1215532.200000ns, VDD,
+ 1216132.600000ns, VDD,
+ 1216132.700000ns, VSS,
+ 1216492.900000ns, VSS,
+ 1216493.000000ns, VDD,
+ 1216733.100000ns, VDD,
+ 1216733.200000ns, VSS,
+ 1218774.800000ns, VSS,
+ 1218774.900000ns, VDD,
+ 1220336.100000ns, VDD,
+ 1220336.200000ns, VSS,
+ 1220816.500000ns, VSS,
+ 1220816.600000ns, VDD,
+ 1221657.200000ns, VDD,
+ 1221657.300000ns, VSS,
+ 1222257.700000ns, VSS,
+ 1222257.800000ns, VDD,
+ 1224539.600000ns, VDD,
+ 1224539.700000ns, VSS,
+ 1225260.200000ns, VSS,
+ 1225260.300000ns, VDD,
+ 1225860.700000ns, VDD,
+ 1225860.800000ns, VSS,
+ 1226341.100000ns, VSS,
+ 1226341.200000ns, VDD,
+ 1226581.300000ns, VDD,
+ 1226581.400000ns, VSS,
+ 1227782.300000ns, VSS,
+ 1227782.400000ns, VDD,
+ 1228743.100000ns, VDD,
+ 1228743.200000ns, VSS,
+ 1229223.500000ns, VSS,
+ 1229223.600000ns, VDD,
+ 1229944.100000ns, VDD,
+ 1229944.200000ns, VSS,
+ 1230784.800000ns, VSS,
+ 1230784.900000ns, VDD,
+ 1232826.500000ns, VDD,
+ 1232826.600000ns, VSS,
+ 1233306.900000ns, VSS,
+ 1233307.000000ns, VDD,
+ 1234267.700000ns, VDD,
+ 1234267.800000ns, VSS,
+ 1234387.800000ns, VSS,
+ 1234387.900000ns, VDD,
+ 1236549.600000ns, VDD,
+ 1236549.700000ns, VSS,
+ 1237750.600000ns, VSS,
+ 1237750.700000ns, VDD,
+ 1238231.000000ns, VDD,
+ 1238231.100000ns, VSS,
+ 1238711.400000ns, VSS,
+ 1238711.500000ns, VDD,
+ 1240272.700000ns, VDD,
+ 1240272.800000ns, VSS,
+ 1240753.100000ns, VSS,
+ 1240753.200000ns, VDD,
+ 1241113.400000ns, VDD,
+ 1241113.500000ns, VSS,
+ 1242794.800000ns, VSS,
+ 1242794.900000ns, VDD,
+ 1244596.300000ns, VDD,
+ 1244596.400000ns, VSS,
+ 1244716.400000ns, VSS,
+ 1244716.500000ns, VDD,
+ 1245076.700000ns, VDD,
+ 1245076.800000ns, VSS,
+ 1245557.100000ns, VSS,
+ 1245557.200000ns, VDD,
+ 1246758.100000ns, VDD,
+ 1246758.200000ns, VSS,
+ 1247238.500000ns, VSS,
+ 1247238.600000ns, VDD,
+ 1249160.100000ns, VDD,
+ 1249160.200000ns, VSS,
+ 1249880.700000ns, VSS,
+ 1249880.800000ns, VDD,
+ 1250961.600000ns, VDD,
+ 1250961.700000ns, VSS,
+ 1251201.800000ns, VSS,
+ 1251201.900000ns, VDD,
+ 1251682.200000ns, VDD,
+ 1251682.300000ns, VSS,
+ 1253723.900000ns, VSS,
+ 1253724.000000ns, VDD,
+ 1254204.300000ns, VDD,
+ 1254204.400000ns, VSS,
+ 1254444.500000ns, VSS,
+ 1254444.600000ns, VDD,
+ 1254924.900000ns, VDD,
+ 1254925.000000ns, VSS,
+ 1255285.200000ns, VSS,
+ 1255285.300000ns, VDD,
+ 1255405.300000ns, VDD,
+ 1255405.400000ns, VSS,
+ 1256366.100000ns, VSS,
+ 1256366.200000ns, VDD,
+ 1257807.300000ns, VDD,
+ 1257807.400000ns, VSS,
+ 1259008.300000ns, VSS,
+ 1259008.400000ns, VDD,
+ 1259248.500000ns, VDD,
+ 1259248.600000ns, VSS,
+ 1260209.300000ns, VSS,
+ 1260209.400000ns, VDD,
+ 1260569.600000ns, VDD,
+ 1260569.700000ns, VSS,
+ 1262491.200000ns, VSS,
+ 1262491.300000ns, VDD,
+ 1262611.300000ns, VDD,
+ 1262611.400000ns, VSS,
+ 1263211.800000ns, VSS,
+ 1263211.900000ns, VDD,
+ 1264292.700000ns, VDD,
+ 1264292.800000ns, VSS,
+ 1264532.900000ns, VSS,
+ 1264533.000000ns, VDD,
+ 1264653.000000ns, VDD,
+ 1264653.100000ns, VSS,
+ 1265133.400000ns, VSS,
+ 1265133.500000ns, VDD,
+ 1265373.600000ns, VDD,
+ 1265373.700000ns, VSS,
+ 1266934.900000ns, VSS,
+ 1266935.000000ns, VDD,
+ 1267775.600000ns, VDD,
+ 1267775.700000ns, VSS,
+ 1268256.000000ns, VSS,
+ 1268256.100000ns, VDD,
+ 1268736.400000ns, VDD,
+ 1268736.500000ns, VSS,
+ 1269697.200000ns, VSS,
+ 1269697.300000ns, VDD,
+ 1270297.700000ns, VDD,
+ 1270297.800000ns, VSS,
+ 1272219.300000ns, VSS,
+ 1272219.400000ns, VDD,
+ 1272579.600000ns, VDD,
+ 1272579.700000ns, VSS,
+ 1273180.100000ns, VSS,
+ 1273180.200000ns, VDD,
+ 1273540.400000ns, VDD,
+ 1273540.500000ns, VSS,
+ 1273780.600000ns, VSS,
+ 1273780.700000ns, VDD,
+ 1275582.100000ns, VDD,
+ 1275582.200000ns, VSS,
+ 1275702.200000ns, VSS,
+ 1275702.300000ns, VDD,
+ 1275822.300000ns, VDD,
+ 1275822.400000ns, VSS,
+ 1276783.100000ns, VSS,
+ 1276783.200000ns, VDD,
+ 1276903.200000ns, VDD,
+ 1276903.300000ns, VSS,
+ 1277023.300000ns, VSS,
+ 1277023.400000ns, VDD,
+ 1277984.100000ns, VDD,
+ 1277984.200000ns, VSS,
+ 1278104.200000ns, VSS,
+ 1278104.300000ns, VDD,
+ 1278224.300000ns, VDD,
+ 1278224.400000ns, VSS,
+ 1278344.400000ns, VSS,
+ 1278344.500000ns, VDD,
+ 1278584.600000ns, VDD,
+ 1278584.700000ns, VSS,
+ 1278944.900000ns, VSS,
+ 1278945.000000ns, VDD,
+ 1279065.000000ns, VDD,
+ 1279065.100000ns, VSS,
+ 1280746.400000ns, VSS,
+ 1280746.500000ns, VDD,
+ 1280866.500000ns, VDD,
+ 1280866.600000ns, VSS,
+ 1282427.800000ns, VSS,
+ 1282427.900000ns, VDD,
+ 1283028.300000ns, VDD,
+ 1283028.400000ns, VSS,
+ 1283388.600000ns, VSS,
+ 1283388.700000ns, VDD,
+ 1283989.100000ns, VDD,
+ 1283989.200000ns, VSS,
+ 1284589.600000ns, VSS,
+ 1284589.700000ns, VDD,
+ 1284949.900000ns, VDD,
+ 1284950.000000ns, VSS,
+ 1285190.100000ns, VSS,
+ 1285190.200000ns, VDD,
+ 1285310.200000ns, VDD,
+ 1285310.300000ns, VSS,
+ 1285430.300000ns, VSS,
+ 1285430.400000ns, VDD,
+ 1286271.000000ns, VDD,
+ 1286271.100000ns, VSS,
+ 1286631.300000ns, VSS,
+ 1286631.400000ns, VDD,
+ 1287111.700000ns, VDD,
+ 1287111.800000ns, VSS,
+ 1288192.600000ns, VSS,
+ 1288192.700000ns, VDD,
+ 1288552.900000ns, VDD,
+ 1288553.000000ns, VSS,
+ 1289994.100000ns, VSS,
+ 1289994.200000ns, VDD,
+ 1290234.300000ns, VDD,
+ 1290234.400000ns, VSS,
+ 1290834.800000ns, VSS,
+ 1290834.900000ns, VDD,
+ 1291795.600000ns, VDD,
+ 1291795.700000ns, VSS,
+ 1292516.200000ns, VSS,
+ 1292516.300000ns, VDD,
+ 1292876.500000ns, VDD,
+ 1292876.600000ns, VSS,
+ 1293356.900000ns, VSS,
+ 1293357.000000ns, VDD,
+ 1293597.100000ns, VDD,
+ 1293597.200000ns, VSS,
+ 1294437.800000ns, VSS,
+ 1294437.900000ns, VDD,
+ 1295758.900000ns, VDD,
+ 1295759.000000ns, VSS,
+ 1296359.400000ns, VSS,
+ 1296359.500000ns, VDD,
+ 1297560.400000ns, VDD,
+ 1297560.500000ns, VSS,
+ 1297680.500000ns, VSS,
+ 1297680.600000ns, VDD,
+ 1297800.600000ns, VDD,
+ 1297800.700000ns, VSS,
+ 1298281.000000ns, VSS,
+ 1298281.100000ns, VDD,
+ 1300322.700000ns, VDD,
+ 1300322.800000ns, VSS,
+ 1300442.800000ns, VSS,
+ 1300442.900000ns, VDD,
+ 1300562.900000ns, VDD,
+ 1300563.000000ns, VSS,
+ 1301523.700000ns, VSS,
+ 1301523.800000ns, VDD,
+ 1302844.800000ns, VDD,
+ 1302844.900000ns, VSS,
+ 1304286.000000ns, VSS,
+ 1304286.100000ns, VDD,
+ 1304406.100000ns, VDD,
+ 1304406.200000ns, VSS,
+ 1304886.500000ns, VSS,
+ 1304886.600000ns, VDD,
+ 1305366.900000ns, VDD,
+ 1305367.000000ns, VSS,
+ 1305607.100000ns, VSS,
+ 1305607.200000ns, VDD,
+ 1305727.200000ns, VDD,
+ 1305727.300000ns, VSS,
+ 1306087.500000ns, VSS,
+ 1306087.600000ns, VDD,
+ 1307648.800000ns, VDD,
+ 1307648.900000ns, VSS,
+ 1308609.600000ns, VSS,
+ 1308609.700000ns, VDD,
+ 1308969.900000ns, VDD,
+ 1308970.000000ns, VSS,
+ 1309570.400000ns, VSS,
+ 1309570.500000ns, VDD,
+ 1309810.600000ns, VDD,
+ 1309810.700000ns, VSS,
+ 1309930.700000ns, VSS,
+ 1309930.800000ns, VDD,
+ 1310891.500000ns, VDD,
+ 1310891.600000ns, VSS,
+ 1311732.200000ns, VSS,
+ 1311732.300000ns, VDD,
+ 1312092.500000ns, VDD,
+ 1312092.600000ns, VSS,
+ 1312572.900000ns, VSS,
+ 1312573.000000ns, VDD,
+ 1312933.200000ns, VDD,
+ 1312933.300000ns, VSS,
+ 1313773.900000ns, VSS,
+ 1313774.000000ns, VDD,
+ 1314614.600000ns, VDD,
+ 1314614.700000ns, VSS,
+ 1314974.900000ns, VSS,
+ 1314975.000000ns, VDD,
+ 1315215.100000ns, VDD,
+ 1315215.200000ns, VSS,
+ 1315335.200000ns, VSS,
+ 1315335.300000ns, VDD,
+ 1315935.700000ns, VDD,
+ 1315935.800000ns, VSS,
+ 1317256.800000ns, VSS,
+ 1317256.900000ns, VDD,
+ 1317376.900000ns, VDD,
+ 1317377.000000ns, VSS,
+ 1317497.000000ns, VSS,
+ 1317497.100000ns, VDD,
+ 1317857.300000ns, VDD,
+ 1317857.400000ns, VSS,
+ 1319058.300000ns, VSS,
+ 1319058.400000ns, VDD,
+ 1320019.100000ns, VDD,
+ 1320019.200000ns, VSS,
+ 1321220.100000ns, VSS,
+ 1321220.200000ns, VDD,
+ 1321460.300000ns, VDD,
+ 1321460.400000ns, VSS,
+ 1322901.500000ns, VSS,
+ 1322901.600000ns, VDD,
+ 1323502.000000ns, VDD,
+ 1323502.100000ns, VSS,
+ 1323982.400000ns, VSS,
+ 1323982.500000ns, VDD,
+ 1324462.800000ns, VDD,
+ 1324462.900000ns, VSS,
+ 1324823.100000ns, VSS,
+ 1324823.200000ns, VDD,
+ 1325303.500000ns, VDD,
+ 1325303.600000ns, VSS,
+ 1325543.700000ns, VSS,
+ 1325543.800000ns, VDD,
+ 1325904.000000ns, VDD,
+ 1325904.100000ns, VSS,
+ 1326144.200000ns, VSS,
+ 1326144.300000ns, VDD,
+ 1326264.300000ns, VDD,
+ 1326264.400000ns, VSS,
+ 1326984.900000ns, VSS,
+ 1326985.000000ns, VDD,
+ 1327465.300000ns, VDD,
+ 1327465.400000ns, VSS,
+ 1328546.200000ns, VSS,
+ 1328546.300000ns, VDD,
+ 1328786.400000ns, VDD,
+ 1328786.500000ns, VSS,
+ 1329507.000000ns, VSS,
+ 1329507.100000ns, VDD,
+ 1330467.800000ns, VDD,
+ 1330467.900000ns, VSS,
+ 1330587.900000ns, VSS,
+ 1330588.000000ns, VDD,
+ 1331428.600000ns, VDD,
+ 1331428.700000ns, VSS,
+ 1332629.600000ns, VSS,
+ 1332629.700000ns, VDD,
+ 1332869.800000ns, VDD,
+ 1332869.900000ns, VSS,
+ 1332989.900000ns, VSS,
+ 1332990.000000ns, VDD,
+ 1333110.000000ns, VDD,
+ 1333110.100000ns, VSS,
+ 1333350.200000ns, VSS,
+ 1333350.300000ns, VDD,
+ 1333950.700000ns, VDD,
+ 1333950.800000ns, VSS,
+ 1334190.900000ns, VSS,
+ 1334191.000000ns, VDD,
+ 1335031.600000ns, VDD,
+ 1335031.700000ns, VSS,
+ 1335271.800000ns, VSS,
+ 1335271.900000ns, VDD,
+ 1335752.200000ns, VDD,
+ 1335752.300000ns, VSS,
+ 1336232.600000ns, VSS,
+ 1336232.700000ns, VDD,
+ 1336953.200000ns, VDD,
+ 1336953.300000ns, VSS,
+ 1337313.500000ns, VSS,
+ 1337313.600000ns, VDD,
+ 1337553.700000ns, VDD,
+ 1337553.800000ns, VSS,
+ 1338514.500000ns, VSS,
+ 1338514.600000ns, VDD,
+ 1339115.000000ns, VDD,
+ 1339115.100000ns, VSS,
+ 1339595.400000ns, VSS,
+ 1339595.500000ns, VDD,
+ 1340075.800000ns, VDD,
+ 1340075.900000ns, VSS,
+ 1340796.400000ns, VSS,
+ 1340796.500000ns, VDD,
+ 1341997.400000ns, VDD,
+ 1341997.500000ns, VSS,
+ 1342477.800000ns, VSS,
+ 1342477.900000ns, VDD,
+ 1342597.900000ns, VDD,
+ 1342598.000000ns, VSS,
+ 1343318.500000ns, VSS,
+ 1343318.600000ns, VDD,
+ 1343558.700000ns, VDD,
+ 1343558.800000ns, VSS,
+ 1343798.900000ns, VSS,
+ 1343799.000000ns, VDD,
+ 1344039.100000ns, VDD,
+ 1344039.200000ns, VSS,
+ 1344879.800000ns, VSS,
+ 1344879.900000ns, VDD,
+ 1345600.400000ns, VDD,
+ 1345600.500000ns, VSS,
+ 1345720.500000ns, VSS,
+ 1345720.600000ns, VDD,
+ 1346321.000000ns, VDD,
+ 1346321.100000ns, VSS,
+ 1347041.600000ns, VSS,
+ 1347041.700000ns, VDD,
+ 1347401.900000ns, VDD,
+ 1347402.000000ns, VSS,
+ 1347762.200000ns, VSS,
+ 1347762.300000ns, VDD,
+ 1349323.500000ns, VDD,
+ 1349323.600000ns, VSS,
+ 1349683.800000ns, VSS,
+ 1349683.900000ns, VDD,
+ 1350284.300000ns, VDD,
+ 1350284.400000ns, VSS,
+ 1350884.800000ns, VSS,
+ 1350884.900000ns, VDD,
+ 1351004.900000ns, VDD,
+ 1351005.000000ns, VSS,
+ 1352446.100000ns, VSS,
+ 1352446.200000ns, VDD,
+ 1352566.200000ns, VDD,
+ 1352566.300000ns, VSS,
+ 1352686.300000ns, VSS,
+ 1352686.400000ns, VDD,
+ 1353166.700000ns, VDD,
+ 1353166.800000ns, VSS,
+ 1353286.800000ns, VSS,
+ 1353286.900000ns, VDD,
+ 1353406.900000ns, VDD,
+ 1353407.000000ns, VSS,
+ 1355929.000000ns, VSS,
+ 1355929.100000ns, VDD,
+ 1357370.200000ns, VDD,
+ 1357370.300000ns, VSS,
+ 1358451.100000ns, VSS,
+ 1358451.200000ns, VDD,
+ 1360252.600000ns, VDD,
+ 1360252.700000ns, VSS,
+ 1360492.800000ns, VSS,
+ 1360492.900000ns, VDD,
+ 1360612.900000ns, VDD,
+ 1360613.000000ns, VSS,
+ 1361093.300000ns, VSS,
+ 1361093.400000ns, VDD,
+ 1361453.600000ns, VDD,
+ 1361453.700000ns, VSS,
+ 1361573.700000ns, VSS,
+ 1361573.800000ns, VDD,
+ 1361934.000000ns, VDD,
+ 1361934.100000ns, VSS,
+ 1362174.200000ns, VSS,
+ 1362174.300000ns, VDD,
+ 1362534.500000ns, VDD,
+ 1362534.600000ns, VSS,
+ 1363255.100000ns, VSS,
+ 1363255.200000ns, VDD,
+ 1364696.300000ns, VDD,
+ 1364696.400000ns, VSS,
+ 1365537.000000ns, VSS,
+ 1365537.100000ns, VDD,
+ 1366017.400000ns, VDD,
+ 1366017.500000ns, VSS,
+ 1366257.600000ns, VSS,
+ 1366257.700000ns, VDD,
+ 1366978.200000ns, VDD,
+ 1366978.300000ns, VSS,
+ 1367698.800000ns, VSS,
+ 1367698.900000ns, VDD,
+ 1368419.400000ns, VDD,
+ 1368419.500000ns, VSS,
+ 1368899.800000ns, VSS,
+ 1368899.900000ns, VDD,
+ 1369019.900000ns, VDD,
+ 1369020.000000ns, VSS,
+ 1369140.000000ns, VSS,
+ 1369140.100000ns, VDD,
+ 1369620.400000ns, VDD,
+ 1369620.500000ns, VSS,
+ 1370581.200000ns, VSS,
+ 1370581.300000ns, VDD,
+ 1370821.400000ns, VDD,
+ 1370821.500000ns, VSS,
+ 1371301.800000ns, VSS,
+ 1371301.900000ns, VDD,
+ 1371542.000000ns, VDD,
+ 1371542.100000ns, VSS,
+ 1371662.100000ns, VSS,
+ 1371662.200000ns, VDD,
+ 1371902.300000ns, VDD,
+ 1371902.400000ns, VSS,
+ 1372983.200000ns, VSS,
+ 1372983.300000ns, VDD,
+ 1373463.600000ns, VDD,
+ 1373463.700000ns, VSS,
+ 1373703.800000ns, VSS,
+ 1373703.900000ns, VDD,
+ 1373823.900000ns, VDD,
+ 1373824.000000ns, VSS,
+ 1374064.100000ns, VSS,
+ 1374064.200000ns, VDD,
+ 1374304.300000ns, VDD,
+ 1374304.400000ns, VSS,
+ 1374904.800000ns, VSS,
+ 1374904.900000ns, VDD,
+ 1375985.700000ns, VDD,
+ 1375985.800000ns, VSS,
+ 1377667.100000ns, VSS,
+ 1377667.200000ns, VDD,
+ 1379708.800000ns, VDD,
+ 1379708.900000ns, VSS,
+ 1381270.100000ns, VSS,
+ 1381270.200000ns, VDD,
+ 1381750.500000ns, VDD,
+ 1381750.600000ns, VSS,
+ 1381870.600000ns, VSS,
+ 1381870.700000ns, VDD,
+ 1382110.800000ns, VDD,
+ 1382110.900000ns, VSS,
+ 1382230.900000ns, VSS,
+ 1382231.000000ns, VDD,
+ 1382831.400000ns, VDD,
+ 1382831.500000ns, VSS,
+ 1383191.700000ns, VSS,
+ 1383191.800000ns, VDD,
+ 1383311.800000ns, VDD,
+ 1383311.900000ns, VSS,
+ 1383431.900000ns, VSS,
+ 1383432.000000ns, VDD,
+ 1383552.000000ns, VDD,
+ 1383552.100000ns, VSS,
+ 1383672.100000ns, VSS,
+ 1383672.200000ns, VDD,
+ 1384152.500000ns, VDD,
+ 1384152.600000ns, VSS,
+ 1384753.000000ns, VSS,
+ 1384753.100000ns, VDD,
+ 1385233.400000ns, VDD,
+ 1385233.500000ns, VSS,
+ 1385473.600000ns, VSS,
+ 1385473.700000ns, VDD,
+ 1385593.700000ns, VDD,
+ 1385593.800000ns, VSS,
+ 1387034.900000ns, VSS,
+ 1387035.000000ns, VDD,
+ 1387875.600000ns, VDD,
+ 1387875.700000ns, VSS,
+ 1388235.900000ns, VSS,
+ 1388236.000000ns, VDD,
+ 1388956.500000ns, VDD,
+ 1388956.600000ns, VSS,
+ 1389076.600000ns, VSS,
+ 1389076.700000ns, VDD,
+ 1389196.700000ns, VDD,
+ 1389196.800000ns, VSS,
+ 1389557.000000ns, VSS,
+ 1389557.100000ns, VDD,
+ 1389677.100000ns, VDD,
+ 1389677.200000ns, VSS,
+ 1391238.400000ns, VSS,
+ 1391238.500000ns, VDD,
+ 1391838.900000ns, VDD,
+ 1391839.000000ns, VSS,
+ 1391959.000000ns, VSS,
+ 1391959.100000ns, VDD,
+ 1392319.300000ns, VDD,
+ 1392319.400000ns, VSS,
+ 1392919.800000ns, VSS,
+ 1392919.900000ns, VDD,
+ 1393880.600000ns, VDD,
+ 1393880.700000ns, VSS,
+ 1394120.800000ns, VSS,
+ 1394120.900000ns, VDD,
+ 1397003.200000ns, VDD,
+ 1397003.300000ns, VSS,
+ 1397843.900000ns, VSS,
+ 1397844.000000ns, VDD,
+ 1398324.300000ns, VDD,
+ 1398324.400000ns, VSS,
+ 1398564.500000ns, VSS,
+ 1398564.600000ns, VDD,
+ 1398684.600000ns, VDD,
+ 1398684.700000ns, VSS,
+ 1403248.400000ns, VSS,
+ 1403248.500000ns, VDD,
+ 1404329.300000ns, VDD,
+ 1404329.400000ns, VSS,
+ 1404449.400000ns, VSS,
+ 1404449.500000ns, VDD,
+ 1404569.500000ns, VDD,
+ 1404569.600000ns, VSS,
+ 1405049.900000ns, VSS,
+ 1405050.000000ns, VDD,
+ 1405650.400000ns, VDD,
+ 1405650.500000ns, VSS,
+ 1406130.800000ns, VSS,
+ 1406130.900000ns, VDD,
+ 1406731.300000ns, VDD,
+ 1406731.400000ns, VSS,
+ 1408412.700000ns, VSS,
+ 1408412.800000ns, VDD,
+ 1410214.200000ns, VDD,
+ 1410214.300000ns, VSS,
+ 1410814.700000ns, VSS,
+ 1410814.800000ns, VDD,
+ 1411295.100000ns, VDD,
+ 1411295.200000ns, VSS,
+ 1411775.500000ns, VSS,
+ 1411775.600000ns, VDD,
+ 1412255.900000ns, VDD,
+ 1412256.000000ns, VSS,
+ 1412856.400000ns, VSS,
+ 1412856.500000ns, VDD,
+ 1414057.400000ns, VDD,
+ 1414057.500000ns, VSS,
+ 1414537.800000ns, VSS,
+ 1414537.900000ns, VDD,
+ 1414778.000000ns, VDD,
+ 1414778.100000ns, VSS,
+ 1415498.600000ns, VSS,
+ 1415498.700000ns, VDD,
+ 1416219.200000ns, VDD,
+ 1416219.300000ns, VSS,
+ 1417420.200000ns, VSS,
+ 1417420.300000ns, VDD,
+ 1417660.400000ns, VDD,
+ 1417660.500000ns, VSS,
+ 1418140.800000ns, VSS,
+ 1418140.900000ns, VDD,
+ 1419582.000000ns, VDD,
+ 1419582.100000ns, VSS,
+ 1419822.200000ns, VSS,
+ 1419822.300000ns, VDD,
+ 1419942.300000ns, VDD,
+ 1419942.400000ns, VSS,
+ 1420062.400000ns, VSS,
+ 1420062.500000ns, VDD,
+ 1420542.800000ns, VDD,
+ 1420542.900000ns, VSS,
+ 1421984.000000ns, VSS,
+ 1421984.100000ns, VDD,
+ 1423064.900000ns, VDD,
+ 1423065.000000ns, VSS,
+ 1425947.300000ns, VSS,
+ 1425947.400000ns, VDD,
+ 1427268.400000ns, VDD,
+ 1427268.500000ns, VSS,
+ 1428229.200000ns, VSS,
+ 1428229.300000ns, VDD,
+ 1429190.000000ns, VDD,
+ 1429190.100000ns, VSS,
+ 1430631.200000ns, VSS,
+ 1430631.300000ns, VDD,
+ 1431712.100000ns, VDD,
+ 1431712.200000ns, VSS,
+ 1431832.200000ns, VSS,
+ 1431832.300000ns, VDD,
+ 1432793.000000ns, VDD,
+ 1432793.100000ns, VSS,
+ 1433873.900000ns, VSS,
+ 1433874.000000ns, VDD,
+ 1435675.400000ns, VDD,
+ 1435675.500000ns, VSS,
+ 1436275.900000ns, VSS,
+ 1436276.000000ns, VDD,
+ 1436636.200000ns, VDD,
+ 1436636.300000ns, VSS,
+ 1438317.600000ns, VSS,
+ 1438317.700000ns, VDD,
+ 1439518.600000ns, VDD,
+ 1439518.700000ns, VSS,
+ 1440359.300000ns, VSS,
+ 1440359.400000ns, VDD,
+ 1442280.900000ns, VDD,
+ 1442281.000000ns, VSS,
+ 1443121.600000ns, VSS,
+ 1443121.700000ns, VDD,
+ 1443361.800000ns, VDD,
+ 1443361.900000ns, VSS,
+ 1444322.600000ns, VSS,
+ 1444322.700000ns, VDD,
+ 1444923.100000ns, VDD,
+ 1444923.200000ns, VSS,
+ 1445643.700000ns, VSS,
+ 1445643.800000ns, VDD,
+ 1445763.800000ns, VDD,
+ 1445763.900000ns, VSS,
+ 1446364.300000ns, VSS,
+ 1446364.400000ns, VDD,
+ 1446844.700000ns, VDD,
+ 1446844.800000ns, VSS,
+ 1447084.900000ns, VSS,
+ 1447085.000000ns, VDD,
+ 1448165.800000ns, VDD,
+ 1448165.900000ns, VSS,
+ 1448886.400000ns, VSS,
+ 1448886.500000ns, VDD,
+ 1449727.100000ns, VDD,
+ 1449727.200000ns, VSS,
+ 1449847.200000ns, VSS,
+ 1449847.300000ns, VDD,
+ 1450808.000000ns, VDD,
+ 1450808.100000ns, VSS,
+ 1450928.100000ns, VSS,
+ 1450928.200000ns, VDD,
+ 1451048.200000ns, VDD,
+ 1451048.300000ns, VSS,
+ 1451528.600000ns, VSS,
+ 1451528.700000ns, VDD,
+ 1452129.100000ns, VDD,
+ 1452129.200000ns, VSS,
+ 1452849.700000ns, VSS,
+ 1452849.800000ns, VDD,
+ 1453690.400000ns, VDD,
+ 1453690.500000ns, VSS,
+ 1454411.000000ns, VSS,
+ 1454411.100000ns, VDD,
+ 1455612.000000ns, VDD,
+ 1455612.100000ns, VSS,
+ 1457293.400000ns, VSS,
+ 1457293.500000ns, VDD,
+ 1459215.000000ns, VDD,
+ 1459215.100000ns, VSS,
+ 1459695.400000ns, VSS,
+ 1459695.500000ns, VDD,
+ 1460416.000000ns, VDD,
+ 1460416.100000ns, VSS,
+ 1460536.100000ns, VSS,
+ 1460536.200000ns, VDD,
+ 1462217.500000ns, VDD,
+ 1462217.600000ns, VSS,
+ 1462818.000000ns, VSS,
+ 1462818.100000ns, VDD,
+ 1463658.700000ns, VDD,
+ 1463658.800000ns, VSS,
+ 1465700.400000ns, VSS,
+ 1465700.500000ns, VDD,
+ 1466661.200000ns, VDD,
+ 1466661.300000ns, VSS,
+ 1467141.600000ns, VSS,
+ 1467141.700000ns, VDD,
+ 1468342.600000ns, VDD,
+ 1468342.700000ns, VSS,
+ 1468702.900000ns, VSS,
+ 1468703.000000ns, VDD,
+ 1468943.100000ns, VDD,
+ 1468943.200000ns, VSS,
+ 1469303.400000ns, VSS,
+ 1469303.500000ns, VDD,
+ 1469903.900000ns, VDD,
+ 1469904.000000ns, VSS,
+ 1471225.000000ns, VSS,
+ 1471225.100000ns, VDD,
+ 1471825.500000ns, VDD,
+ 1471825.600000ns, VSS,
+ 1472426.000000ns, VSS,
+ 1472426.100000ns, VDD,
+ 1472546.100000ns, VDD,
+ 1472546.200000ns, VSS,
+ 1472666.200000ns, VSS,
+ 1472666.300000ns, VDD,
+ 1473747.100000ns, VDD,
+ 1473747.200000ns, VSS,
+ 1474227.500000ns, VSS,
+ 1474227.600000ns, VDD,
+ 1474467.700000ns, VDD,
+ 1474467.800000ns, VSS,
+ 1474707.900000ns, VSS,
+ 1474708.000000ns, VDD,
+ 1475188.300000ns, VDD,
+ 1475188.400000ns, VSS,
+ 1475308.400000ns, VSS,
+ 1475308.500000ns, VDD,
+ 1476629.500000ns, VDD,
+ 1476629.600000ns, VSS,
+ 1477950.600000ns, VSS,
+ 1477950.700000ns, VDD,
+ 1478310.900000ns, VDD,
+ 1478311.000000ns, VSS,
+ 1478791.300000ns, VSS,
+ 1478791.400000ns, VDD,
+ 1479872.200000ns, VDD,
+ 1479872.300000ns, VSS,
+ 1481433.500000ns, VSS,
+ 1481433.600000ns, VDD,
+ 1481673.700000ns, VDD,
+ 1481673.800000ns, VSS,
+ 1481793.800000ns, VSS,
+ 1481793.900000ns, VDD,
+ 1481913.900000ns, VDD,
+ 1481914.000000ns, VSS,
+ 1484436.000000ns, VSS,
+ 1484436.100000ns, VDD,
+ 1486597.800000ns, VDD,
+ 1486597.900000ns, VSS,
+ 1486958.100000ns, VSS,
+ 1486958.200000ns, VDD,
+ 1487678.700000ns, VDD,
+ 1487678.800000ns, VSS,
+ 1488519.400000ns, VSS,
+ 1488519.500000ns, VDD,
+ 1488999.800000ns, VDD,
+ 1488999.900000ns, VSS,
+ 1489840.500000ns, VSS,
+ 1489840.600000ns, VDD,
+ 1491521.900000ns, VDD,
+ 1491522.000000ns, VSS,
+ 1491642.000000ns, VSS,
+ 1491642.100000ns, VDD,
+ 1492602.800000ns, VDD,
+ 1492602.900000ns, VSS,
+ 1492722.900000ns, VSS,
+ 1492723.000000ns, VDD,
+ 1492843.000000ns, VDD,
+ 1492843.100000ns, VSS,
+ 1494644.500000ns, VSS,
+ 1494644.600000ns, VDD,
+ 1494764.600000ns, VDD,
+ 1494764.700000ns, VSS,
+ 1495124.900000ns, VSS,
+ 1495125.000000ns, VDD,
+ 1495365.100000ns, VDD,
+ 1495365.200000ns, VSS,
+ 1495725.400000ns, VSS,
+ 1495725.500000ns, VDD,
+ 1495845.500000ns, VDD,
+ 1495845.600000ns, VSS,
+ 1496085.700000ns, VSS,
+ 1496085.800000ns, VDD,
+ 1496205.800000ns, VDD,
+ 1496205.900000ns, VSS,
+ 1496926.400000ns, VSS,
+ 1496926.500000ns, VDD,
+ 1497526.900000ns, VDD,
+ 1497527.000000ns, VSS,
+ 1497767.100000ns, VSS,
+ 1497767.200000ns, VDD,
+ 1498007.300000ns, VDD,
+ 1498007.400000ns, VSS,
+ 1498487.700000ns, VSS,
+ 1498487.800000ns, VDD,
+ 1498968.100000ns, VDD,
+ 1498968.200000ns, VSS,
+ 1499688.700000ns, VSS,
+ 1499688.800000ns, VDD,
+ 1499928.900000ns, VDD,
+ 1499929.000000ns, VSS,
+ 1501250.000000ns, VSS,
+ 1501250.100000ns, VDD,
+ 1502330.900000ns, VDD,
+ 1502331.000000ns, VSS,
+ 1502811.300000ns, VSS,
+ 1502811.400000ns, VDD,
+ 1503291.700000ns, VDD,
+ 1503291.800000ns, VSS,
+ 1504252.500000ns, VSS,
+ 1504252.600000ns, VDD,
+ 1504612.800000ns, VDD,
+ 1504612.900000ns, VSS,
+ 1504853.000000ns, VSS,
+ 1504853.100000ns, VDD,
+ 1505453.500000ns, VDD,
+ 1505453.600000ns, VSS,
+ 1505573.600000ns, VSS,
+ 1505573.700000ns, VDD,
+ 1505693.700000ns, VDD,
+ 1505693.800000ns, VSS,
+ 1506054.000000ns, VSS,
+ 1506054.100000ns, VDD,
+ 1507975.600000ns, VDD,
+ 1507975.700000ns, VSS,
+ 1509416.800000ns, VSS,
+ 1509416.900000ns, VDD,
+ 1509657.000000ns, VDD,
+ 1509657.100000ns, VSS,
+ 1510137.400000ns, VSS,
+ 1510137.500000ns, VDD,
+ 1512059.000000ns, VDD,
+ 1512059.100000ns, VSS,
+ 1512419.300000ns, VSS,
+ 1512419.400000ns, VDD,
+ 1513620.300000ns, VDD,
+ 1513620.400000ns, VSS,
+ 1514461.000000ns, VSS,
+ 1514461.100000ns, VDD,
+ 1515662.000000ns, VDD,
+ 1515662.100000ns, VSS,
+ 1516262.500000ns, VSS,
+ 1516262.600000ns, VDD,
+ 1516382.600000ns, VDD,
+ 1516382.700000ns, VSS,
+ 1516502.700000ns, VSS,
+ 1516502.800000ns, VDD,
+ 1516622.800000ns, VDD,
+ 1516622.900000ns, VSS,
+ 1516742.900000ns, VSS,
+ 1516743.000000ns, VDD,
+ 1517943.900000ns, VDD,
+ 1517944.000000ns, VSS,
+ 1518424.300000ns, VSS,
+ 1518424.400000ns, VDD,
+ 1519144.900000ns, VDD,
+ 1519145.000000ns, VSS,
+ 1519625.300000ns, VSS,
+ 1519625.400000ns, VDD,
+ 1519745.400000ns, VDD,
+ 1519745.500000ns, VSS,
+ 1520105.700000ns, VSS,
+ 1520105.800000ns, VDD,
+ 1520826.300000ns, VDD,
+ 1520826.400000ns, VSS,
+ 1522147.400000ns, VSS,
+ 1522147.500000ns, VDD,
+ 1523348.400000ns, VDD,
+ 1523348.500000ns, VSS,
+ 1523708.700000ns, VSS,
+ 1523708.800000ns, VDD,
+ 1525029.800000ns, VDD,
+ 1525029.900000ns, VSS,
+ 1526591.100000ns, VSS,
+ 1526591.200000ns, VDD,
+ 1526711.200000ns, VDD,
+ 1526711.300000ns, VSS,
+ 1526831.300000ns, VSS,
+ 1526831.400000ns, VDD,
+ 1527071.500000ns, VDD,
+ 1527071.600000ns, VSS,
+ 1527191.600000ns, VSS,
+ 1527191.700000ns, VDD,
+ 1528272.500000ns, VDD,
+ 1528272.600000ns, VSS,
+ 1528752.900000ns, VSS,
+ 1528753.000000ns, VDD,
+ 1528873.000000ns, VDD,
+ 1528873.100000ns, VSS,
+ 1529113.200000ns, VSS,
+ 1529113.300000ns, VDD,
+ 1529233.300000ns, VDD,
+ 1529233.400000ns, VSS,
+ 1529353.400000ns, VSS,
+ 1529353.500000ns, VDD,
+ 1529473.500000ns, VDD,
+ 1529473.600000ns, VSS,
+ 1529593.600000ns, VSS,
+ 1529593.700000ns, VDD,
+ 1529953.900000ns, VDD,
+ 1529954.000000ns, VSS,
+ 1530194.100000ns, VSS,
+ 1530194.200000ns, VDD,
+ 1530314.200000ns, VDD,
+ 1530314.300000ns, VSS,
+ 1530554.400000ns, VSS,
+ 1530554.500000ns, VDD,
+ 1531395.100000ns, VDD,
+ 1531395.200000ns, VSS,
+ 1531635.300000ns, VSS,
+ 1531635.400000ns, VDD,
+ 1531755.400000ns, VDD,
+ 1531755.500000ns, VSS,
+ 1532235.800000ns, VSS,
+ 1532235.900000ns, VDD,
+ 1532716.200000ns, VDD,
+ 1532716.300000ns, VSS,
+ 1533196.600000ns, VSS,
+ 1533196.700000ns, VDD,
+ 1533677.000000ns, VDD,
+ 1533677.100000ns, VSS,
+ 1534397.600000ns, VSS,
+ 1534397.700000ns, VDD,
+ 1535238.300000ns, VDD,
+ 1535238.400000ns, VSS,
+ 1535478.500000ns, VSS,
+ 1535478.600000ns, VDD,
+ 1535718.700000ns, VDD,
+ 1535718.800000ns, VSS,
+ 1536559.400000ns, VSS,
+ 1536559.500000ns, VDD,
+ 1537640.300000ns, VDD,
+ 1537640.400000ns, VSS,
+ 1538000.600000ns, VSS,
+ 1538000.700000ns, VDD,
+ 1539561.900000ns, VDD,
+ 1539562.000000ns, VSS,
+ 1539682.000000ns, VSS,
+ 1539682.100000ns, VDD,
+ 1540642.800000ns, VDD,
+ 1540642.900000ns, VSS,
+ 1541603.600000ns, VSS,
+ 1541603.700000ns, VDD,
+ 1541723.700000ns, VDD,
+ 1541723.800000ns, VSS,
+ 1542324.200000ns, VSS,
+ 1542324.300000ns, VDD,
+ 1543285.000000ns, VDD,
+ 1543285.100000ns, VSS,
+ 1544365.900000ns, VSS,
+ 1544366.000000ns, VDD,
+ 1544486.000000ns, VDD,
+ 1544486.100000ns, VSS,
+ 1545807.100000ns, VSS,
+ 1545807.200000ns, VDD,
+ 1547128.200000ns, VDD,
+ 1547128.300000ns, VSS,
+ 1548689.500000ns, VSS,
+ 1548689.600000ns, VDD,
+ 1549530.200000ns, VDD,
+ 1549530.300000ns, VSS
+)}


rCP in_CP 0 1.0
BCP in_CP 0 V={table(time,
+ 0.100000ns, VDD,
+ 120.100000ns, VDD,
+ 120.200000ns, VSS,
+ 240.200000ns, VSS,
+ 240.300000ns, VDD,
+ 600.500000ns, VDD,
+ 600.600000ns, VSS,
+ 1441.200000ns, VSS,
+ 1441.300000ns, VDD,
+ 1921.600000ns, VDD,
+ 1921.700000ns, VSS,
+ 2041.700000ns, VSS,
+ 2041.800000ns, VDD,
+ 2402.000000ns, VDD,
+ 2402.100000ns, VSS,
+ 2882.400000ns, VSS,
+ 2882.500000ns, VDD,
+ 3122.600000ns, VDD,
+ 3122.700000ns, VSS,
+ 3362.800000ns, VSS,
+ 3362.900000ns, VDD,
+ 3963.300000ns, VDD,
+ 3963.400000ns, VSS,
+ 4683.900000ns, VSS,
+ 4684.000000ns, VDD,
+ 4924.100000ns, VDD,
+ 4924.200000ns, VSS,
+ 5524.600000ns, VSS,
+ 5524.700000ns, VDD,
+ 6125.100000ns, VDD,
+ 6125.200000ns, VSS,
+ 6485.400000ns, VSS,
+ 6485.500000ns, VDD,
+ 6965.800000ns, VDD,
+ 6965.900000ns, VSS,
+ 8407.000000ns, VSS,
+ 8407.100000ns, VDD,
+ 8767.300000ns, VDD,
+ 8767.400000ns, VSS,
+ 8887.400000ns, VSS,
+ 8887.500000ns, VDD,
+ 10208.500000ns, VDD,
+ 10208.600000ns, VSS,
+ 10448.700000ns, VSS,
+ 10448.800000ns, VDD,
+ 11049.200000ns, VDD,
+ 11049.300000ns, VSS,
+ 11409.500000ns, VSS,
+ 11409.600000ns, VDD,
+ 12130.100000ns, VDD,
+ 12130.200000ns, VSS,
+ 12490.400000ns, VSS,
+ 12490.500000ns, VDD,
+ 12730.600000ns, VDD,
+ 12730.700000ns, VSS,
+ 12850.700000ns, VSS,
+ 12850.800000ns, VDD,
+ 13931.600000ns, VDD,
+ 13931.700000ns, VSS,
+ 14412.000000ns, VSS,
+ 14412.100000ns, VDD,
+ 14652.200000ns, VDD,
+ 14652.300000ns, VSS,
+ 15012.500000ns, VSS,
+ 15012.600000ns, VDD,
+ 15132.600000ns, VDD,
+ 15132.700000ns, VSS,
+ 15252.700000ns, VSS,
+ 15252.800000ns, VDD,
+ 15613.000000ns, VDD,
+ 15613.100000ns, VSS,
+ 15733.100000ns, VSS,
+ 15733.200000ns, VDD,
+ 16093.400000ns, VDD,
+ 16093.500000ns, VSS,
+ 16693.900000ns, VSS,
+ 16694.000000ns, VDD,
+ 16934.100000ns, VDD,
+ 16934.200000ns, VSS,
+ 17294.400000ns, VSS,
+ 17294.500000ns, VDD,
+ 17414.500000ns, VDD,
+ 17414.600000ns, VSS,
+ 17534.600000ns, VSS,
+ 17534.700000ns, VDD,
+ 18015.000000ns, VDD,
+ 18015.100000ns, VSS,
+ 18135.100000ns, VSS,
+ 18135.200000ns, VDD,
+ 18375.300000ns, VDD,
+ 18375.400000ns, VSS,
+ 18735.600000ns, VSS,
+ 18735.700000ns, VDD,
+ 18855.700000ns, VDD,
+ 18855.800000ns, VSS,
+ 19456.200000ns, VSS,
+ 19456.300000ns, VDD,
+ 19816.500000ns, VDD,
+ 19816.600000ns, VSS,
+ 20176.800000ns, VSS,
+ 20176.900000ns, VDD,
+ 20417.000000ns, VDD,
+ 20417.100000ns, VSS,
+ 20777.300000ns, VSS,
+ 20777.400000ns, VDD,
+ 21618.000000ns, VDD,
+ 21618.100000ns, VSS,
+ 21738.100000ns, VSS,
+ 21738.200000ns, VDD,
+ 22098.400000ns, VDD,
+ 22098.500000ns, VSS,
+ 22458.700000ns, VSS,
+ 22458.800000ns, VDD,
+ 22698.900000ns, VDD,
+ 22699.000000ns, VSS,
+ 23899.900000ns, VSS,
+ 23900.000000ns, VDD,
+ 24380.300000ns, VDD,
+ 24380.400000ns, VSS,
+ 24500.400000ns, VSS,
+ 24500.500000ns, VDD,
+ 24860.700000ns, VDD,
+ 24860.800000ns, VSS,
+ 25100.900000ns, VSS,
+ 25101.000000ns, VDD,
+ 25221.000000ns, VDD,
+ 25221.100000ns, VSS,
+ 25581.300000ns, VSS,
+ 25581.400000ns, VDD,
+ 25821.500000ns, VDD,
+ 25821.600000ns, VSS,
+ 26902.400000ns, VSS,
+ 26902.500000ns, VDD,
+ 27022.500000ns, VDD,
+ 27022.600000ns, VSS,
+ 27382.800000ns, VSS,
+ 27382.900000ns, VDD,
+ 28103.400000ns, VDD,
+ 28103.500000ns, VSS,
+ 28343.600000ns, VSS,
+ 28343.700000ns, VDD,
+ 28463.700000ns, VDD,
+ 28463.800000ns, VSS,
+ 28703.900000ns, VSS,
+ 28704.000000ns, VDD,
+ 28944.100000ns, VDD,
+ 28944.200000ns, VSS,
+ 29304.400000ns, VSS,
+ 29304.500000ns, VDD,
+ 29544.600000ns, VDD,
+ 29544.700000ns, VSS,
+ 29784.800000ns, VSS,
+ 29784.900000ns, VDD,
+ 30025.000000ns, VDD,
+ 30025.100000ns, VSS,
+ 30985.800000ns, VSS,
+ 30985.900000ns, VDD,
+ 31826.500000ns, VDD,
+ 31826.600000ns, VSS,
+ 32066.700000ns, VSS,
+ 32066.800000ns, VDD,
+ 32547.100000ns, VDD,
+ 32547.200000ns, VSS,
+ 33868.200000ns, VSS,
+ 33868.300000ns, VDD,
+ 34108.400000ns, VDD,
+ 34108.500000ns, VSS,
+ 34348.600000ns, VSS,
+ 34348.700000ns, VDD,
+ 34829.000000ns, VDD,
+ 34829.100000ns, VSS,
+ 34949.100000ns, VSS,
+ 34949.200000ns, VDD,
+ 36390.300000ns, VDD,
+ 36390.400000ns, VSS,
+ 36510.400000ns, VSS,
+ 36510.500000ns, VDD,
+ 36750.600000ns, VDD,
+ 36750.700000ns, VSS,
+ 37231.000000ns, VSS,
+ 37231.100000ns, VDD,
+ 37471.200000ns, VDD,
+ 37471.300000ns, VSS,
+ 37591.300000ns, VSS,
+ 37591.400000ns, VDD,
+ 37831.500000ns, VDD,
+ 37831.600000ns, VSS,
+ 38191.800000ns, VSS,
+ 38191.900000ns, VDD,
+ 39032.500000ns, VDD,
+ 39032.600000ns, VSS,
+ 39152.600000ns, VSS,
+ 39152.700000ns, VDD,
+ 40113.400000ns, VDD,
+ 40113.500000ns, VSS,
+ 40233.500000ns, VSS,
+ 40233.600000ns, VDD,
+ 40593.800000ns, VDD,
+ 40593.900000ns, VSS,
+ 40713.900000ns, VSS,
+ 40714.000000ns, VDD,
+ 42035.000000ns, VDD,
+ 42035.100000ns, VSS,
+ 42515.400000ns, VSS,
+ 42515.500000ns, VDD,
+ 42635.500000ns, VDD,
+ 42635.600000ns, VSS,
+ 43836.500000ns, VSS,
+ 43836.600000ns, VDD,
+ 44076.700000ns, VDD,
+ 44076.800000ns, VSS,
+ 44437.000000ns, VSS,
+ 44437.100000ns, VDD,
+ 44557.100000ns, VDD,
+ 44557.200000ns, VSS,
+ 45517.900000ns, VSS,
+ 45518.000000ns, VDD,
+ 45878.200000ns, VDD,
+ 45878.300000ns, VSS,
+ 45998.300000ns, VSS,
+ 45998.400000ns, VDD,
+ 46478.700000ns, VDD,
+ 46478.800000ns, VSS,
+ 46718.900000ns, VSS,
+ 46719.000000ns, VDD,
+ 46839.000000ns, VDD,
+ 46839.100000ns, VSS,
+ 47199.300000ns, VSS,
+ 47199.400000ns, VDD,
+ 47319.400000ns, VDD,
+ 47319.500000ns, VSS,
+ 47799.800000ns, VSS,
+ 47799.900000ns, VDD,
+ 48400.300000ns, VDD,
+ 48400.400000ns, VSS,
+ 48520.400000ns, VSS,
+ 48520.500000ns, VDD,
+ 48640.500000ns, VDD,
+ 48640.600000ns, VSS,
+ 48760.600000ns, VSS,
+ 48760.700000ns, VDD,
+ 49000.800000ns, VDD,
+ 49000.900000ns, VSS,
+ 49361.100000ns, VSS,
+ 49361.200000ns, VDD,
+ 49481.200000ns, VDD,
+ 49481.300000ns, VSS,
+ 49961.600000ns, VSS,
+ 49961.700000ns, VDD,
+ 50081.700000ns, VDD,
+ 50081.800000ns, VSS,
+ 50201.800000ns, VSS,
+ 50201.900000ns, VDD,
+ 50442.000000ns, VDD,
+ 50442.100000ns, VSS,
+ 51162.600000ns, VSS,
+ 51162.700000ns, VDD,
+ 52363.600000ns, VDD,
+ 52363.700000ns, VSS,
+ 52964.100000ns, VSS,
+ 52964.200000ns, VDD,
+ 53324.400000ns, VDD,
+ 53324.500000ns, VSS,
+ 53804.800000ns, VSS,
+ 53804.900000ns, VDD,
+ 53924.900000ns, VDD,
+ 53925.000000ns, VSS,
+ 54045.000000ns, VSS,
+ 54045.100000ns, VDD,
+ 54405.300000ns, VDD,
+ 54405.400000ns, VSS,
+ 54885.700000ns, VSS,
+ 54885.800000ns, VDD,
+ 55125.900000ns, VDD,
+ 55126.000000ns, VSS,
+ 55486.200000ns, VSS,
+ 55486.300000ns, VDD,
+ 55606.300000ns, VDD,
+ 55606.400000ns, VSS,
+ 55726.400000ns, VSS,
+ 55726.500000ns, VDD,
+ 56086.700000ns, VDD,
+ 56086.800000ns, VSS,
+ 56206.800000ns, VSS,
+ 56206.900000ns, VDD,
+ 56567.100000ns, VDD,
+ 56567.200000ns, VSS,
+ 57047.500000ns, VSS,
+ 57047.600000ns, VDD,
+ 57527.900000ns, VDD,
+ 57528.000000ns, VSS,
+ 58128.400000ns, VSS,
+ 58128.500000ns, VDD,
+ 58849.000000ns, VDD,
+ 58849.100000ns, VSS,
+ 59209.300000ns, VSS,
+ 59209.400000ns, VDD,
+ 59689.700000ns, VDD,
+ 59689.800000ns, VSS,
+ 60290.200000ns, VSS,
+ 60290.300000ns, VDD,
+ 60410.300000ns, VDD,
+ 60410.400000ns, VSS,
+ 61010.800000ns, VSS,
+ 61010.900000ns, VDD,
+ 61130.900000ns, VDD,
+ 61131.000000ns, VSS,
+ 61251.000000ns, VSS,
+ 61251.100000ns, VDD,
+ 62331.900000ns, VDD,
+ 62332.000000ns, VSS,
+ 62692.200000ns, VSS,
+ 62692.300000ns, VDD,
+ 63292.700000ns, VDD,
+ 63292.800000ns, VSS,
+ 64253.500000ns, VSS,
+ 64253.600000ns, VDD,
+ 64373.600000ns, VDD,
+ 64373.700000ns, VSS,
+ 64974.100000ns, VSS,
+ 64974.200000ns, VDD,
+ 65694.700000ns, VDD,
+ 65694.800000ns, VSS,
+ 66055.000000ns, VSS,
+ 66055.100000ns, VDD,
+ 66535.400000ns, VDD,
+ 66535.500000ns, VSS,
+ 66655.500000ns, VSS,
+ 66655.600000ns, VDD,
+ 66775.600000ns, VDD,
+ 66775.700000ns, VSS,
+ 67256.000000ns, VSS,
+ 67256.100000ns, VDD,
+ 67496.200000ns, VDD,
+ 67496.300000ns, VSS,
+ 67856.500000ns, VSS,
+ 67856.600000ns, VDD,
+ 67976.600000ns, VDD,
+ 67976.700000ns, VSS,
+ 68096.700000ns, VSS,
+ 68096.800000ns, VDD,
+ 68457.000000ns, VDD,
+ 68457.100000ns, VSS,
+ 68577.100000ns, VSS,
+ 68577.200000ns, VDD,
+ 69177.600000ns, VDD,
+ 69177.700000ns, VSS,
+ 69297.700000ns, VSS,
+ 69297.800000ns, VDD,
+ 70018.300000ns, VDD,
+ 70018.400000ns, VSS,
+ 71099.200000ns, VSS,
+ 71099.300000ns, VDD,
+ 71579.600000ns, VDD,
+ 71579.700000ns, VSS,
+ 72540.400000ns, VSS,
+ 72540.500000ns, VDD,
+ 73261.000000ns, VDD,
+ 73261.100000ns, VSS,
+ 73861.500000ns, VSS,
+ 73861.600000ns, VDD,
+ 74341.900000ns, VDD,
+ 74342.000000ns, VSS,
+ 75663.000000ns, VSS,
+ 75663.100000ns, VDD,
+ 75783.100000ns, VDD,
+ 75783.200000ns, VSS,
+ 76263.500000ns, VSS,
+ 76263.600000ns, VDD,
+ 76503.700000ns, VDD,
+ 76503.800000ns, VSS,
+ 77104.200000ns, VSS,
+ 77104.300000ns, VDD,
+ 77224.300000ns, VDD,
+ 77224.400000ns, VSS,
+ 77704.700000ns, VSS,
+ 77704.800000ns, VDD,
+ 78305.200000ns, VDD,
+ 78305.300000ns, VSS,
+ 78425.300000ns, VSS,
+ 78425.400000ns, VDD,
+ 78665.500000ns, VDD,
+ 78665.600000ns, VSS,
+ 78905.700000ns, VSS,
+ 78905.800000ns, VDD,
+ 79145.900000ns, VDD,
+ 79146.000000ns, VSS,
+ 79266.000000ns, VSS,
+ 79266.100000ns, VDD,
+ 79626.300000ns, VDD,
+ 79626.400000ns, VSS,
+ 79866.500000ns, VSS,
+ 79866.600000ns, VDD,
+ 80106.700000ns, VDD,
+ 80106.800000ns, VSS,
+ 80226.800000ns, VSS,
+ 80226.900000ns, VDD,
+ 80707.200000ns, VDD,
+ 80707.300000ns, VSS,
+ 81067.500000ns, VSS,
+ 81067.600000ns, VDD,
+ 81547.900000ns, VDD,
+ 81548.000000ns, VSS,
+ 82028.300000ns, VSS,
+ 82028.400000ns, VDD,
+ 82388.600000ns, VDD,
+ 82388.700000ns, VSS,
+ 82748.900000ns, VSS,
+ 82749.000000ns, VDD,
+ 82989.100000ns, VDD,
+ 82989.200000ns, VSS,
+ 83109.200000ns, VSS,
+ 83109.300000ns, VDD,
+ 84430.300000ns, VDD,
+ 84430.400000ns, VSS,
+ 85030.800000ns, VSS,
+ 85030.900000ns, VDD,
+ 85150.900000ns, VDD,
+ 85151.000000ns, VSS,
+ 85631.300000ns, VSS,
+ 85631.400000ns, VDD,
+ 86231.800000ns, VDD,
+ 86231.900000ns, VSS,
+ 86952.400000ns, VSS,
+ 86952.500000ns, VDD,
+ 87552.900000ns, VDD,
+ 87553.000000ns, VSS,
+ 88153.400000ns, VSS,
+ 88153.500000ns, VDD,
+ 88513.700000ns, VDD,
+ 88513.800000ns, VSS,
+ 89474.500000ns, VSS,
+ 89474.600000ns, VDD,
+ 89594.600000ns, VDD,
+ 89594.700000ns, VSS,
+ 90075.000000ns, VSS,
+ 90075.100000ns, VDD,
+ 90195.100000ns, VDD,
+ 90195.200000ns, VSS,
+ 90315.200000ns, VSS,
+ 90315.300000ns, VDD,
+ 90555.400000ns, VDD,
+ 90555.500000ns, VSS,
+ 90675.500000ns, VSS,
+ 90675.600000ns, VDD,
+ 91035.800000ns, VDD,
+ 91035.900000ns, VSS,
+ 91876.500000ns, VSS,
+ 91876.600000ns, VDD,
+ 92477.000000ns, VDD,
+ 92477.100000ns, VSS,
+ 92597.100000ns, VSS,
+ 92597.200000ns, VDD,
+ 92717.200000ns, VDD,
+ 92717.300000ns, VSS,
+ 93077.500000ns, VSS,
+ 93077.600000ns, VDD,
+ 93317.700000ns, VDD,
+ 93317.800000ns, VSS,
+ 93437.800000ns, VSS,
+ 93437.900000ns, VDD,
+ 93678.000000ns, VDD,
+ 93678.100000ns, VSS,
+ 94038.300000ns, VSS,
+ 94038.400000ns, VDD,
+ 94879.000000ns, VDD,
+ 94879.100000ns, VSS,
+ 94999.100000ns, VSS,
+ 94999.200000ns, VDD,
+ 95239.300000ns, VDD,
+ 95239.400000ns, VSS,
+ 95599.600000ns, VSS,
+ 95599.700000ns, VDD,
+ 95719.700000ns, VDD,
+ 95719.800000ns, VSS,
+ 95839.800000ns, VSS,
+ 95839.900000ns, VDD,
+ 96440.300000ns, VDD,
+ 96440.400000ns, VSS,
+ 96560.400000ns, VSS,
+ 96560.500000ns, VDD,
+ 97040.800000ns, VDD,
+ 97040.900000ns, VSS,
+ 97401.100000ns, VSS,
+ 97401.200000ns, VDD,
+ 97641.300000ns, VDD,
+ 97641.400000ns, VSS,
+ 97881.500000ns, VSS,
+ 97881.600000ns, VDD,
+ 98241.800000ns, VDD,
+ 98241.900000ns, VSS,
+ 98482.000000ns, VSS,
+ 98482.100000ns, VDD,
+ 98722.200000ns, VDD,
+ 98722.300000ns, VSS,
+ 99562.900000ns, VSS,
+ 99563.000000ns, VDD,
+ 100163.400000ns, VDD,
+ 100163.500000ns, VSS,
+ 100283.500000ns, VSS,
+ 100283.600000ns, VDD,
+ 101124.200000ns, VDD,
+ 101124.300000ns, VSS,
+ 101244.300000ns, VSS,
+ 101244.400000ns, VDD,
+ 103286.000000ns, VDD,
+ 103286.100000ns, VSS,
+ 103406.100000ns, VSS,
+ 103406.200000ns, VDD,
+ 103766.400000ns, VDD,
+ 103766.500000ns, VSS,
+ 104366.900000ns, VSS,
+ 104367.000000ns, VDD,
+ 104727.200000ns, VDD,
+ 104727.300000ns, VSS,
+ 105327.700000ns, VSS,
+ 105327.800000ns, VDD,
+ 105928.200000ns, VDD,
+ 105928.300000ns, VSS,
+ 106648.800000ns, VSS,
+ 106648.900000ns, VDD,
+ 107009.100000ns, VDD,
+ 107009.200000ns, VSS,
+ 107489.500000ns, VSS,
+ 107489.600000ns, VDD,
+ 108450.300000ns, VDD,
+ 108450.400000ns, VSS,
+ 109050.800000ns, VSS,
+ 109050.900000ns, VDD,
+ 109170.900000ns, VDD,
+ 109171.000000ns, VSS,
+ 109531.200000ns, VSS,
+ 109531.300000ns, VDD,
+ 110131.700000ns, VDD,
+ 110131.800000ns, VSS,
+ 110852.300000ns, VSS,
+ 110852.400000ns, VDD,
+ 111212.600000ns, VDD,
+ 111212.700000ns, VSS,
+ 111693.000000ns, VSS,
+ 111693.100000ns, VDD,
+ 112413.600000ns, VDD,
+ 112413.700000ns, VSS,
+ 112533.700000ns, VSS,
+ 112533.800000ns, VDD,
+ 112773.900000ns, VDD,
+ 112774.000000ns, VSS,
+ 113614.600000ns, VSS,
+ 113614.700000ns, VDD,
+ 113734.700000ns, VDD,
+ 113734.800000ns, VSS,
+ 113974.900000ns, VSS,
+ 113975.000000ns, VDD,
+ 114095.000000ns, VDD,
+ 114095.100000ns, VSS,
+ 115175.900000ns, VSS,
+ 115176.000000ns, VDD,
+ 115416.100000ns, VDD,
+ 115416.200000ns, VSS,
+ 115536.200000ns, VSS,
+ 115536.300000ns, VDD,
+ 115656.300000ns, VDD,
+ 115656.400000ns, VSS,
+ 115896.500000ns, VSS,
+ 115896.600000ns, VDD,
+ 116737.200000ns, VDD,
+ 116737.300000ns, VSS,
+ 116977.400000ns, VSS,
+ 116977.500000ns, VDD,
+ 117097.500000ns, VDD,
+ 117097.600000ns, VSS,
+ 117457.800000ns, VSS,
+ 117457.900000ns, VDD,
+ 117938.200000ns, VDD,
+ 117938.300000ns, VSS,
+ 118298.500000ns, VSS,
+ 118298.600000ns, VDD,
+ 118899.000000ns, VDD,
+ 118899.100000ns, VSS,
+ 119379.400000ns, VSS,
+ 119379.500000ns, VDD,
+ 119499.500000ns, VDD,
+ 119499.600000ns, VSS,
+ 120100.000000ns, VSS,
+ 120100.100000ns, VDD,
+ 120460.300000ns, VDD,
+ 120460.400000ns, VSS,
+ 120820.600000ns, VSS,
+ 120820.700000ns, VDD,
+ 121421.100000ns, VDD,
+ 121421.200000ns, VSS,
+ 122261.800000ns, VSS,
+ 122261.900000ns, VDD,
+ 123342.700000ns, VDD,
+ 123342.800000ns, VSS,
+ 123462.800000ns, VSS,
+ 123462.900000ns, VDD,
+ 123823.100000ns, VDD,
+ 123823.200000ns, VSS,
+ 124063.300000ns, VSS,
+ 124063.400000ns, VDD,
+ 124183.400000ns, VDD,
+ 124183.500000ns, VSS,
+ 124423.600000ns, VSS,
+ 124423.700000ns, VDD,
+ 125024.100000ns, VDD,
+ 125024.200000ns, VSS,
+ 125504.500000ns, VSS,
+ 125504.600000ns, VDD,
+ 125624.600000ns, VDD,
+ 125624.700000ns, VSS,
+ 126705.500000ns, VSS,
+ 126705.600000ns, VDD,
+ 126825.600000ns, VDD,
+ 126825.700000ns, VSS,
+ 126945.700000ns, VSS,
+ 126945.800000ns, VDD,
+ 127185.900000ns, VDD,
+ 127186.000000ns, VSS,
+ 127306.000000ns, VSS,
+ 127306.100000ns, VDD,
+ 127666.300000ns, VDD,
+ 127666.400000ns, VSS,
+ 128026.600000ns, VSS,
+ 128026.700000ns, VDD,
+ 128266.800000ns, VDD,
+ 128266.900000ns, VSS,
+ 128386.900000ns, VSS,
+ 128387.000000ns, VDD,
+ 129587.900000ns, VDD,
+ 129588.000000ns, VSS,
+ 129708.000000ns, VSS,
+ 129708.100000ns, VDD,
+ 130188.400000ns, VDD,
+ 130188.500000ns, VSS,
+ 131149.200000ns, VSS,
+ 131149.300000ns, VDD,
+ 131269.300000ns, VDD,
+ 131269.400000ns, VSS,
+ 131749.700000ns, VSS,
+ 131749.800000ns, VDD,
+ 132230.100000ns, VDD,
+ 132230.200000ns, VSS,
+ 132350.200000ns, VSS,
+ 132350.300000ns, VDD,
+ 132710.500000ns, VDD,
+ 132710.600000ns, VSS,
+ 133070.800000ns, VSS,
+ 133070.900000ns, VDD,
+ 133671.300000ns, VDD,
+ 133671.400000ns, VSS,
+ 134271.800000ns, VSS,
+ 134271.900000ns, VDD,
+ 134391.900000ns, VDD,
+ 134392.000000ns, VSS,
+ 134752.200000ns, VSS,
+ 134752.300000ns, VDD,
+ 134992.400000ns, VDD,
+ 134992.500000ns, VSS,
+ 135112.500000ns, VSS,
+ 135112.600000ns, VDD,
+ 135352.700000ns, VDD,
+ 135352.800000ns, VSS,
+ 135833.100000ns, VSS,
+ 135833.200000ns, VDD,
+ 137274.300000ns, VDD,
+ 137274.400000ns, VSS,
+ 137394.400000ns, VSS,
+ 137394.500000ns, VDD,
+ 137634.600000ns, VDD,
+ 137634.700000ns, VSS,
+ 137754.700000ns, VSS,
+ 137754.800000ns, VDD,
+ 138235.100000ns, VDD,
+ 138235.200000ns, VSS,
+ 138355.200000ns, VSS,
+ 138355.300000ns, VDD,
+ 138475.300000ns, VDD,
+ 138475.400000ns, VSS,
+ 138715.500000ns, VSS,
+ 138715.600000ns, VDD,
+ 138835.600000ns, VDD,
+ 138835.700000ns, VSS,
+ 139075.800000ns, VSS,
+ 139075.900000ns, VDD,
+ 139195.900000ns, VDD,
+ 139196.000000ns, VSS,
+ 139316.000000ns, VSS,
+ 139316.100000ns, VDD,
+ 139556.200000ns, VDD,
+ 139556.300000ns, VSS,
+ 139916.500000ns, VSS,
+ 139916.600000ns, VDD,
+ 140517.000000ns, VDD,
+ 140517.100000ns, VSS,
+ 141597.900000ns, VSS,
+ 141598.000000ns, VDD,
+ 142438.600000ns, VDD,
+ 142438.700000ns, VSS,
+ 142919.000000ns, VSS,
+ 142919.100000ns, VDD,
+ 143159.200000ns, VDD,
+ 143159.300000ns, VSS,
+ 143399.400000ns, VSS,
+ 143399.500000ns, VDD,
+ 143639.600000ns, VDD,
+ 143639.700000ns, VSS,
+ 144960.700000ns, VSS,
+ 144960.800000ns, VDD,
+ 145441.100000ns, VDD,
+ 145441.200000ns, VSS,
+ 145561.200000ns, VSS,
+ 145561.300000ns, VDD,
+ 145801.400000ns, VDD,
+ 145801.500000ns, VSS,
+ 146281.800000ns, VSS,
+ 146281.900000ns, VDD,
+ 146522.000000ns, VDD,
+ 146522.100000ns, VSS,
+ 147362.700000ns, VSS,
+ 147362.800000ns, VDD,
+ 147723.000000ns, VDD,
+ 147723.100000ns, VSS,
+ 147963.200000ns, VSS,
+ 147963.300000ns, VDD,
+ 148443.600000ns, VDD,
+ 148443.700000ns, VSS,
+ 148563.700000ns, VSS,
+ 148563.800000ns, VDD,
+ 148803.900000ns, VDD,
+ 148804.000000ns, VSS,
+ 149164.200000ns, VSS,
+ 149164.300000ns, VDD,
+ 149524.500000ns, VDD,
+ 149524.600000ns, VSS,
+ 150004.900000ns, VSS,
+ 150005.000000ns, VDD,
+ 150485.300000ns, VDD,
+ 150485.400000ns, VSS,
+ 150605.400000ns, VSS,
+ 150605.500000ns, VDD,
+ 150965.700000ns, VDD,
+ 150965.800000ns, VSS,
+ 151566.200000ns, VSS,
+ 151566.300000ns, VDD,
+ 151806.400000ns, VDD,
+ 151806.500000ns, VSS,
+ 152166.700000ns, VSS,
+ 152166.800000ns, VDD,
+ 152647.100000ns, VDD,
+ 152647.200000ns, VSS,
+ 152767.200000ns, VSS,
+ 152767.300000ns, VDD,
+ 153247.600000ns, VDD,
+ 153247.700000ns, VSS,
+ 153487.800000ns, VSS,
+ 153487.900000ns, VDD,
+ 153728.000000ns, VDD,
+ 153728.100000ns, VSS,
+ 153968.200000ns, VSS,
+ 153968.300000ns, VDD,
+ 154088.300000ns, VDD,
+ 154088.400000ns, VSS,
+ 154688.800000ns, VSS,
+ 154688.900000ns, VDD,
+ 154808.900000ns, VDD,
+ 154809.000000ns, VSS,
+ 155169.200000ns, VSS,
+ 155169.300000ns, VDD,
+ 155769.700000ns, VDD,
+ 155769.800000ns, VSS,
+ 155889.800000ns, VSS,
+ 155889.900000ns, VDD,
+ 156250.100000ns, VDD,
+ 156250.200000ns, VSS,
+ 156370.200000ns, VSS,
+ 156370.300000ns, VDD,
+ 156610.400000ns, VDD,
+ 156610.500000ns, VSS,
+ 156970.700000ns, VSS,
+ 156970.800000ns, VDD,
+ 157090.800000ns, VDD,
+ 157090.900000ns, VSS,
+ 157571.200000ns, VSS,
+ 157571.300000ns, VDD,
+ 158171.700000ns, VDD,
+ 158171.800000ns, VSS,
+ 158291.800000ns, VSS,
+ 158291.900000ns, VDD,
+ 158411.900000ns, VDD,
+ 158412.000000ns, VSS,
+ 158532.000000ns, VSS,
+ 158532.100000ns, VDD,
+ 158652.100000ns, VDD,
+ 158652.200000ns, VSS,
+ 159132.500000ns, VSS,
+ 159132.600000ns, VDD,
+ 159612.900000ns, VDD,
+ 159613.000000ns, VSS,
+ 159733.000000ns, VSS,
+ 159733.100000ns, VDD,
+ 160093.300000ns, VDD,
+ 160093.400000ns, VSS,
+ 160813.900000ns, VSS,
+ 160814.000000ns, VDD,
+ 161054.100000ns, VDD,
+ 161054.200000ns, VSS,
+ 161894.800000ns, VSS,
+ 161894.900000ns, VDD,
+ 162255.100000ns, VDD,
+ 162255.200000ns, VSS,
+ 162615.400000ns, VSS,
+ 162615.500000ns, VDD,
+ 163456.100000ns, VDD,
+ 163456.200000ns, VSS,
+ 163816.400000ns, VSS,
+ 163816.500000ns, VDD,
+ 164056.600000ns, VDD,
+ 164056.700000ns, VSS,
+ 164296.800000ns, VSS,
+ 164296.900000ns, VDD,
+ 164897.300000ns, VDD,
+ 164897.400000ns, VSS,
+ 165497.800000ns, VSS,
+ 165497.900000ns, VDD,
+ 166098.300000ns, VDD,
+ 166098.400000ns, VSS,
+ 167059.100000ns, VSS,
+ 167059.200000ns, VDD,
+ 167419.400000ns, VDD,
+ 167419.500000ns, VSS,
+ 167539.500000ns, VSS,
+ 167539.600000ns, VDD,
+ 167779.700000ns, VDD,
+ 167779.800000ns, VSS,
+ 168260.100000ns, VSS,
+ 168260.200000ns, VDD,
+ 168500.300000ns, VDD,
+ 168500.400000ns, VSS,
+ 168620.400000ns, VSS,
+ 168620.500000ns, VDD,
+ 168860.600000ns, VDD,
+ 168860.700000ns, VSS,
+ 168980.700000ns, VSS,
+ 168980.800000ns, VDD,
+ 170061.600000ns, VDD,
+ 170061.700000ns, VSS,
+ 170542.000000ns, VSS,
+ 170542.100000ns, VDD,
+ 171022.400000ns, VDD,
+ 171022.500000ns, VSS,
+ 171622.900000ns, VSS,
+ 171623.000000ns, VDD,
+ 171983.200000ns, VDD,
+ 171983.300000ns, VSS,
+ 172103.300000ns, VSS,
+ 172103.400000ns, VDD,
+ 172703.800000ns, VDD,
+ 172703.900000ns, VSS,
+ 172823.900000ns, VSS,
+ 172824.000000ns, VDD,
+ 173184.200000ns, VDD,
+ 173184.300000ns, VSS,
+ 173304.300000ns, VSS,
+ 173304.400000ns, VDD,
+ 173544.500000ns, VDD,
+ 173544.600000ns, VSS,
+ 173904.800000ns, VSS,
+ 173904.900000ns, VDD,
+ 174385.200000ns, VDD,
+ 174385.300000ns, VSS,
+ 174745.500000ns, VSS,
+ 174745.600000ns, VDD,
+ 174865.600000ns, VDD,
+ 174865.700000ns, VSS,
+ 175225.900000ns, VSS,
+ 175226.000000ns, VDD,
+ 175826.400000ns, VDD,
+ 175826.500000ns, VSS,
+ 176426.900000ns, VSS,
+ 176427.000000ns, VDD,
+ 176547.000000ns, VDD,
+ 176547.100000ns, VSS,
+ 177387.700000ns, VSS,
+ 177387.800000ns, VDD,
+ 177507.800000ns, VDD,
+ 177507.900000ns, VSS,
+ 177868.100000ns, VSS,
+ 177868.200000ns, VDD,
+ 177988.200000ns, VDD,
+ 177988.300000ns, VSS,
+ 178108.300000ns, VSS,
+ 178108.400000ns, VDD,
+ 178228.400000ns, VDD,
+ 178228.500000ns, VSS,
+ 178708.800000ns, VSS,
+ 178708.900000ns, VDD,
+ 179429.400000ns, VDD,
+ 179429.500000ns, VSS,
+ 180150.000000ns, VSS,
+ 180150.100000ns, VDD,
+ 180630.400000ns, VDD,
+ 180630.500000ns, VSS,
+ 181110.800000ns, VSS,
+ 181110.900000ns, VDD,
+ 182311.800000ns, VDD,
+ 182311.900000ns, VSS,
+ 182431.900000ns, VSS,
+ 182432.000000ns, VDD,
+ 182672.100000ns, VDD,
+ 182672.200000ns, VSS,
+ 182792.200000ns, VSS,
+ 182792.300000ns, VDD,
+ 183152.500000ns, VDD,
+ 183152.600000ns, VSS,
+ 183512.800000ns, VSS,
+ 183512.900000ns, VDD,
+ 183632.900000ns, VDD,
+ 183633.000000ns, VSS,
+ 183753.000000ns, VSS,
+ 183753.100000ns, VDD,
+ 184353.500000ns, VDD,
+ 184353.600000ns, VSS,
+ 184473.600000ns, VSS,
+ 184473.700000ns, VDD,
+ 184713.800000ns, VDD,
+ 184713.900000ns, VSS,
+ 185074.100000ns, VSS,
+ 185074.200000ns, VDD,
+ 185434.400000ns, VDD,
+ 185434.500000ns, VSS,
+ 185674.600000ns, VSS,
+ 185674.700000ns, VDD,
+ 186155.000000ns, VDD,
+ 186155.100000ns, VSS,
+ 186275.100000ns, VSS,
+ 186275.200000ns, VDD,
+ 186635.400000ns, VDD,
+ 186635.500000ns, VSS,
+ 186755.500000ns, VSS,
+ 186755.600000ns, VDD,
+ 186995.700000ns, VDD,
+ 186995.800000ns, VSS,
+ 187235.900000ns, VSS,
+ 187236.000000ns, VDD,
+ 187476.100000ns, VDD,
+ 187476.200000ns, VSS,
+ 187596.200000ns, VSS,
+ 187596.300000ns, VDD,
+ 187956.500000ns, VDD,
+ 187956.600000ns, VSS,
+ 188677.100000ns, VSS,
+ 188677.200000ns, VDD,
+ 188917.300000ns, VDD,
+ 188917.400000ns, VSS,
+ 189277.600000ns, VSS,
+ 189277.700000ns, VDD,
+ 189998.200000ns, VDD,
+ 189998.300000ns, VSS,
+ 190118.300000ns, VSS,
+ 190118.400000ns, VDD,
+ 190238.400000ns, VDD,
+ 190238.500000ns, VSS,
+ 190358.500000ns, VSS,
+ 190358.600000ns, VDD,
+ 190598.700000ns, VDD,
+ 190598.800000ns, VSS,
+ 190718.800000ns, VSS,
+ 190718.900000ns, VDD,
+ 191799.700000ns, VDD,
+ 191799.800000ns, VSS,
+ 191919.800000ns, VSS,
+ 191919.900000ns, VDD,
+ 192520.300000ns, VDD,
+ 192520.400000ns, VSS,
+ 192640.400000ns, VSS,
+ 192640.500000ns, VDD,
+ 192880.600000ns, VDD,
+ 192880.700000ns, VSS,
+ 193361.000000ns, VSS,
+ 193361.100000ns, VDD,
+ 193841.400000ns, VDD,
+ 193841.500000ns, VSS,
+ 194321.800000ns, VSS,
+ 194321.900000ns, VDD,
+ 194802.200000ns, VDD,
+ 194802.300000ns, VSS,
+ 195282.600000ns, VSS,
+ 195282.700000ns, VDD,
+ 196243.400000ns, VDD,
+ 196243.500000ns, VSS,
+ 196723.800000ns, VSS,
+ 196723.900000ns, VDD,
+ 196843.900000ns, VDD,
+ 196844.000000ns, VSS,
+ 196964.000000ns, VSS,
+ 196964.100000ns, VDD,
+ 198165.000000ns, VDD,
+ 198165.100000ns, VSS,
+ 198285.100000ns, VSS,
+ 198285.200000ns, VDD,
+ 199606.200000ns, VDD,
+ 199606.300000ns, VSS,
+ 200326.800000ns, VSS,
+ 200326.900000ns, VDD,
+ 200927.300000ns, VDD,
+ 200927.400000ns, VSS,
+ 201047.400000ns, VSS,
+ 201047.500000ns, VDD,
+ 201287.600000ns, VDD,
+ 201287.700000ns, VSS,
+ 201647.900000ns, VSS,
+ 201648.000000ns, VDD,
+ 201768.000000ns, VDD,
+ 201768.100000ns, VSS,
+ 201888.100000ns, VSS,
+ 201888.200000ns, VDD,
+ 202488.600000ns, VDD,
+ 202488.700000ns, VSS,
+ 202848.900000ns, VSS,
+ 202849.000000ns, VDD,
+ 203809.700000ns, VDD,
+ 203809.800000ns, VSS,
+ 204170.000000ns, VSS,
+ 204170.100000ns, VDD,
+ 204650.400000ns, VDD,
+ 204650.500000ns, VSS,
+ 205010.700000ns, VSS,
+ 205010.800000ns, VDD,
+ 205250.900000ns, VDD,
+ 205251.000000ns, VSS,
+ 205491.100000ns, VSS,
+ 205491.200000ns, VDD,
+ 205731.300000ns, VDD,
+ 205731.400000ns, VSS,
+ 207172.500000ns, VSS,
+ 207172.600000ns, VDD,
+ 207292.600000ns, VDD,
+ 207292.700000ns, VSS,
+ 207412.700000ns, VSS,
+ 207412.800000ns, VDD,
+ 207652.900000ns, VDD,
+ 207653.000000ns, VSS,
+ 207773.000000ns, VSS,
+ 207773.100000ns, VDD,
+ 208253.400000ns, VDD,
+ 208253.500000ns, VSS,
+ 208373.500000ns, VSS,
+ 208373.600000ns, VDD,
+ 208733.800000ns, VDD,
+ 208733.900000ns, VSS,
+ 209214.200000ns, VSS,
+ 209214.300000ns, VDD,
+ 209574.500000ns, VDD,
+ 209574.600000ns, VSS,
+ 209694.600000ns, VSS,
+ 209694.700000ns, VDD,
+ 210535.300000ns, VDD,
+ 210535.400000ns, VSS,
+ 210655.400000ns, VSS,
+ 210655.500000ns, VDD,
+ 211135.800000ns, VDD,
+ 211135.900000ns, VSS,
+ 211255.900000ns, VSS,
+ 211256.000000ns, VDD,
+ 211736.300000ns, VDD,
+ 211736.400000ns, VSS,
+ 211856.400000ns, VSS,
+ 211856.500000ns, VDD,
+ 211976.500000ns, VDD,
+ 211976.600000ns, VSS,
+ 212336.800000ns, VSS,
+ 212336.900000ns, VDD,
+ 212577.000000ns, VDD,
+ 212577.100000ns, VSS,
+ 212697.100000ns, VSS,
+ 212697.200000ns, VDD,
+ 212937.300000ns, VDD,
+ 212937.400000ns, VSS,
+ 213057.400000ns, VSS,
+ 213057.500000ns, VDD,
+ 213657.900000ns, VDD,
+ 213658.000000ns, VSS,
+ 213778.000000ns, VSS,
+ 213778.100000ns, VDD,
+ 214378.500000ns, VDD,
+ 214378.600000ns, VSS,
+ 214498.600000ns, VSS,
+ 214498.700000ns, VDD,
+ 215099.100000ns, VDD,
+ 215099.200000ns, VSS,
+ 215459.400000ns, VSS,
+ 215459.500000ns, VDD,
+ 215579.500000ns, VDD,
+ 215579.600000ns, VSS,
+ 215699.600000ns, VSS,
+ 215699.700000ns, VDD,
+ 216059.900000ns, VDD,
+ 216060.000000ns, VSS,
+ 216180.000000ns, VSS,
+ 216180.100000ns, VDD,
+ 216900.600000ns, VDD,
+ 216900.700000ns, VSS,
+ 217741.300000ns, VSS,
+ 217741.400000ns, VDD,
+ 218221.700000ns, VDD,
+ 218221.800000ns, VSS,
+ 218822.200000ns, VSS,
+ 218822.300000ns, VDD,
+ 219182.500000ns, VDD,
+ 219182.600000ns, VSS,
+ 219302.600000ns, VSS,
+ 219302.700000ns, VDD,
+ 219783.000000ns, VDD,
+ 219783.100000ns, VSS,
+ 221104.100000ns, VSS,
+ 221104.200000ns, VDD,
+ 221224.200000ns, VDD,
+ 221224.300000ns, VSS,
+ 221824.700000ns, VSS,
+ 221824.800000ns, VDD,
+ 222064.900000ns, VDD,
+ 222065.000000ns, VSS,
+ 222665.400000ns, VSS,
+ 222665.500000ns, VDD,
+ 222785.500000ns, VDD,
+ 222785.600000ns, VSS,
+ 223746.300000ns, VSS,
+ 223746.400000ns, VDD,
+ 224226.700000ns, VDD,
+ 224226.800000ns, VSS,
+ 224466.900000ns, VSS,
+ 224467.000000ns, VDD,
+ 224947.300000ns, VDD,
+ 224947.400000ns, VSS,
+ 225067.400000ns, VSS,
+ 225067.500000ns, VDD,
+ 225427.700000ns, VDD,
+ 225427.800000ns, VSS,
+ 225788.000000ns, VSS,
+ 225788.100000ns, VDD,
+ 226388.500000ns, VDD,
+ 226388.600000ns, VSS,
+ 226748.800000ns, VSS,
+ 226748.900000ns, VDD,
+ 226989.000000ns, VDD,
+ 226989.100000ns, VSS,
+ 227109.100000ns, VSS,
+ 227109.200000ns, VDD,
+ 227229.200000ns, VDD,
+ 227229.300000ns, VSS,
+ 227589.500000ns, VSS,
+ 227589.600000ns, VDD,
+ 227949.800000ns, VDD,
+ 227949.900000ns, VSS,
+ 228069.900000ns, VSS,
+ 228070.000000ns, VDD,
+ 228310.100000ns, VDD,
+ 228310.200000ns, VSS,
+ 228670.400000ns, VSS,
+ 228670.500000ns, VDD,
+ 228910.600000ns, VDD,
+ 228910.700000ns, VSS,
+ 229270.900000ns, VSS,
+ 229271.000000ns, VDD,
+ 229631.200000ns, VDD,
+ 229631.300000ns, VSS,
+ 229751.300000ns, VSS,
+ 229751.400000ns, VDD,
+ 231552.800000ns, VDD,
+ 231552.900000ns, VSS,
+ 231672.900000ns, VSS,
+ 231673.000000ns, VDD,
+ 232033.200000ns, VDD,
+ 232033.300000ns, VSS,
+ 232393.500000ns, VSS,
+ 232393.600000ns, VDD,
+ 233234.200000ns, VDD,
+ 233234.300000ns, VSS,
+ 233354.300000ns, VSS,
+ 233354.400000ns, VDD,
+ 234074.900000ns, VDD,
+ 234075.000000ns, VSS,
+ 234795.500000ns, VSS,
+ 234795.600000ns, VDD,
+ 235035.700000ns, VDD,
+ 235035.800000ns, VSS,
+ 235275.900000ns, VSS,
+ 235276.000000ns, VDD,
+ 235396.000000ns, VDD,
+ 235396.100000ns, VSS,
+ 235996.500000ns, VSS,
+ 235996.600000ns, VDD,
+ 236236.700000ns, VDD,
+ 236236.800000ns, VSS,
+ 236356.800000ns, VSS,
+ 236356.900000ns, VDD,
+ 237317.600000ns, VDD,
+ 237317.700000ns, VSS,
+ 238038.200000ns, VSS,
+ 238038.300000ns, VDD,
+ 238158.300000ns, VDD,
+ 238158.400000ns, VSS,
+ 238398.500000ns, VSS,
+ 238398.600000ns, VDD,
+ 238638.700000ns, VDD,
+ 238638.800000ns, VSS,
+ 238878.900000ns, VSS,
+ 238879.000000ns, VDD,
+ 239839.700000ns, VDD,
+ 239839.800000ns, VSS,
+ 239959.800000ns, VSS,
+ 239959.900000ns, VDD,
+ 240200.000000ns, VDD,
+ 240200.100000ns, VSS,
+ 240440.200000ns, VSS,
+ 240440.300000ns, VDD,
+ 240680.400000ns, VDD,
+ 240680.500000ns, VSS,
+ 241040.700000ns, VSS,
+ 241040.800000ns, VDD,
+ 241401.000000ns, VDD,
+ 241401.100000ns, VSS,
+ 241641.200000ns, VSS,
+ 241641.300000ns, VDD,
+ 241761.300000ns, VDD,
+ 241761.400000ns, VSS,
+ 241881.400000ns, VSS,
+ 241881.500000ns, VDD,
+ 242121.600000ns, VDD,
+ 242121.700000ns, VSS,
+ 242481.900000ns, VSS,
+ 242482.000000ns, VDD,
+ 243082.400000ns, VDD,
+ 243082.500000ns, VSS,
+ 243202.500000ns, VSS,
+ 243202.600000ns, VDD,
+ 243442.700000ns, VDD,
+ 243442.800000ns, VSS,
+ 243803.000000ns, VSS,
+ 243803.100000ns, VDD,
+ 244403.500000ns, VDD,
+ 244403.600000ns, VSS,
+ 244763.800000ns, VSS,
+ 244763.900000ns, VDD,
+ 245244.200000ns, VDD,
+ 245244.300000ns, VSS,
+ 245724.600000ns, VSS,
+ 245724.700000ns, VDD,
+ 246084.900000ns, VDD,
+ 246085.000000ns, VSS,
+ 246325.100000ns, VSS,
+ 246325.200000ns, VDD,
+ 246445.200000ns, VDD,
+ 246445.300000ns, VSS,
+ 247045.700000ns, VSS,
+ 247045.800000ns, VDD,
+ 247526.100000ns, VDD,
+ 247526.200000ns, VSS,
+ 247886.400000ns, VSS,
+ 247886.500000ns, VDD,
+ 248126.600000ns, VDD,
+ 248126.700000ns, VSS,
+ 248246.700000ns, VSS,
+ 248246.800000ns, VDD,
+ 248486.900000ns, VDD,
+ 248487.000000ns, VSS,
+ 248607.000000ns, VSS,
+ 248607.100000ns, VDD,
+ 248847.200000ns, VDD,
+ 248847.300000ns, VSS,
+ 249207.500000ns, VSS,
+ 249207.600000ns, VDD,
+ 249447.700000ns, VDD,
+ 249447.800000ns, VSS,
+ 249808.000000ns, VSS,
+ 249808.100000ns, VDD,
+ 250048.200000ns, VDD,
+ 250048.300000ns, VSS,
+ 250408.500000ns, VSS,
+ 250408.600000ns, VDD,
+ 250528.600000ns, VDD,
+ 250528.700000ns, VSS,
+ 251129.100000ns, VSS,
+ 251129.200000ns, VDD,
+ 251369.300000ns, VDD,
+ 251369.400000ns, VSS,
+ 251729.600000ns, VSS,
+ 251729.700000ns, VDD,
+ 251849.700000ns, VDD,
+ 251849.800000ns, VSS,
+ 252089.900000ns, VSS,
+ 252090.000000ns, VDD,
+ 252330.100000ns, VDD,
+ 252330.200000ns, VSS,
+ 252690.400000ns, VSS,
+ 252690.500000ns, VDD,
+ 252810.500000ns, VDD,
+ 252810.600000ns, VSS,
+ 252930.600000ns, VSS,
+ 252930.700000ns, VDD,
+ 253531.100000ns, VDD,
+ 253531.200000ns, VSS,
+ 254131.600000ns, VSS,
+ 254131.700000ns, VDD,
+ 254251.700000ns, VDD,
+ 254251.800000ns, VSS,
+ 254852.200000ns, VSS,
+ 254852.300000ns, VDD,
+ 255092.400000ns, VDD,
+ 255092.500000ns, VSS,
+ 255452.700000ns, VSS,
+ 255452.800000ns, VDD,
+ 255572.800000ns, VDD,
+ 255572.900000ns, VSS,
+ 256533.600000ns, VSS,
+ 256533.700000ns, VDD,
+ 256893.900000ns, VDD,
+ 256894.000000ns, VSS,
+ 257254.200000ns, VSS,
+ 257254.300000ns, VDD,
+ 258815.500000ns, VDD,
+ 258815.600000ns, VSS,
+ 258935.600000ns, VSS,
+ 258935.700000ns, VDD,
+ 259175.800000ns, VDD,
+ 259175.900000ns, VSS,
+ 259536.100000ns, VSS,
+ 259536.200000ns, VDD,
+ 259656.200000ns, VDD,
+ 259656.300000ns, VSS,
+ 259776.300000ns, VSS,
+ 259776.400000ns, VDD,
+ 260136.600000ns, VDD,
+ 260136.700000ns, VSS,
+ 260256.700000ns, VSS,
+ 260256.800000ns, VDD,
+ 260857.200000ns, VDD,
+ 260857.300000ns, VSS,
+ 260977.300000ns, VSS,
+ 260977.400000ns, VDD,
+ 261217.500000ns, VDD,
+ 261217.600000ns, VSS,
+ 261457.700000ns, VSS,
+ 261457.800000ns, VDD,
+ 261697.900000ns, VDD,
+ 261698.000000ns, VSS,
+ 261938.100000ns, VSS,
+ 261938.200000ns, VDD,
+ 263019.000000ns, VDD,
+ 263019.100000ns, VSS,
+ 263499.400000ns, VSS,
+ 263499.500000ns, VDD,
+ 263979.800000ns, VDD,
+ 263979.900000ns, VSS,
+ 264220.000000ns, VSS,
+ 264220.100000ns, VDD,
+ 264820.500000ns, VDD,
+ 264820.600000ns, VSS,
+ 265300.900000ns, VSS,
+ 265301.000000ns, VDD,
+ 266021.500000ns, VDD,
+ 266021.600000ns, VSS,
+ 266501.900000ns, VSS,
+ 266502.000000ns, VDD,
+ 266982.300000ns, VDD,
+ 266982.400000ns, VSS,
+ 267702.900000ns, VSS,
+ 267703.000000ns, VDD,
+ 269384.300000ns, VDD,
+ 269384.400000ns, VSS,
+ 269744.600000ns, VSS,
+ 269744.700000ns, VDD,
+ 270465.200000ns, VDD,
+ 270465.300000ns, VSS,
+ 270945.600000ns, VSS,
+ 270945.700000ns, VDD,
+ 271065.700000ns, VDD,
+ 271065.800000ns, VSS,
+ 271786.300000ns, VSS,
+ 271786.400000ns, VDD,
+ 272386.800000ns, VDD,
+ 272386.900000ns, VSS,
+ 272506.900000ns, VSS,
+ 272507.000000ns, VDD,
+ 272987.300000ns, VDD,
+ 272987.400000ns, VSS,
+ 273227.500000ns, VSS,
+ 273227.600000ns, VDD,
+ 273347.600000ns, VDD,
+ 273347.700000ns, VSS,
+ 273587.800000ns, VSS,
+ 273587.900000ns, VDD,
+ 273828.000000ns, VDD,
+ 273828.100000ns, VSS,
+ 273948.100000ns, VSS,
+ 273948.200000ns, VDD,
+ 274788.800000ns, VDD,
+ 274788.900000ns, VSS,
+ 274908.900000ns, VSS,
+ 274909.000000ns, VDD,
+ 275149.100000ns, VDD,
+ 275149.200000ns, VSS,
+ 275389.300000ns, VSS,
+ 275389.400000ns, VDD,
+ 275629.500000ns, VDD,
+ 275629.600000ns, VSS,
+ 275749.600000ns, VSS,
+ 275749.700000ns, VDD,
+ 276230.000000ns, VDD,
+ 276230.100000ns, VSS,
+ 276350.100000ns, VSS,
+ 276350.200000ns, VDD,
+ 276470.200000ns, VDD,
+ 276470.300000ns, VSS,
+ 276950.600000ns, VSS,
+ 276950.700000ns, VDD,
+ 277190.800000ns, VDD,
+ 277190.900000ns, VSS,
+ 277671.200000ns, VSS,
+ 277671.300000ns, VDD,
+ 277911.400000ns, VDD,
+ 277911.500000ns, VSS,
+ 278271.700000ns, VSS,
+ 278271.800000ns, VDD,
+ 278391.800000ns, VDD,
+ 278391.900000ns, VSS,
+ 278511.900000ns, VSS,
+ 278512.000000ns, VDD,
+ 279112.400000ns, VDD,
+ 279112.500000ns, VSS,
+ 279232.500000ns, VSS,
+ 279232.600000ns, VDD,
+ 279712.900000ns, VDD,
+ 279713.000000ns, VSS,
+ 279833.000000ns, VSS,
+ 279833.100000ns, VDD,
+ 280073.200000ns, VDD,
+ 280073.300000ns, VSS,
+ 280313.400000ns, VSS,
+ 280313.500000ns, VDD,
+ 280673.700000ns, VDD,
+ 280673.800000ns, VSS,
+ 280793.800000ns, VSS,
+ 280793.900000ns, VDD,
+ 281034.000000ns, VDD,
+ 281034.100000ns, VSS,
+ 281754.600000ns, VSS,
+ 281754.700000ns, VDD,
+ 282355.100000ns, VDD,
+ 282355.200000ns, VSS,
+ 283556.100000ns, VSS,
+ 283556.200000ns, VDD,
+ 283796.300000ns, VDD,
+ 283796.400000ns, VSS,
+ 284516.900000ns, VSS,
+ 284517.000000ns, VDD,
+ 286438.500000ns, VDD,
+ 286438.600000ns, VSS,
+ 287039.000000ns, VSS,
+ 287039.100000ns, VDD,
+ 287999.800000ns, VDD,
+ 287999.900000ns, VSS,
+ 288360.100000ns, VSS,
+ 288360.200000ns, VDD,
+ 288840.500000ns, VDD,
+ 288840.600000ns, VSS,
+ 289441.000000ns, VSS,
+ 289441.100000ns, VDD,
+ 289561.100000ns, VDD,
+ 289561.200000ns, VSS,
+ 289681.200000ns, VSS,
+ 289681.300000ns, VDD,
+ 289921.400000ns, VDD,
+ 289921.500000ns, VSS,
+ 290041.500000ns, VSS,
+ 290041.600000ns, VDD,
+ 290161.600000ns, VDD,
+ 290161.700000ns, VSS,
+ 290281.700000ns, VSS,
+ 290281.800000ns, VDD,
+ 291002.300000ns, VDD,
+ 291002.400000ns, VSS,
+ 291482.700000ns, VSS,
+ 291482.800000ns, VDD,
+ 291722.900000ns, VDD,
+ 291723.000000ns, VSS,
+ 292803.800000ns, VSS,
+ 292803.900000ns, VDD,
+ 293044.000000ns, VDD,
+ 293044.100000ns, VSS,
+ 293284.200000ns, VSS,
+ 293284.300000ns, VDD,
+ 293524.400000ns, VDD,
+ 293524.500000ns, VSS,
+ 293644.500000ns, VSS,
+ 293644.600000ns, VDD,
+ 293764.600000ns, VDD,
+ 293764.700000ns, VSS,
+ 294605.300000ns, VSS,
+ 294605.400000ns, VDD,
+ 295205.800000ns, VDD,
+ 295205.900000ns, VSS,
+ 296166.600000ns, VSS,
+ 296166.700000ns, VDD,
+ 296526.900000ns, VDD,
+ 296527.000000ns, VSS,
+ 297848.000000ns, VSS,
+ 297848.100000ns, VDD,
+ 298568.600000ns, VDD,
+ 298568.700000ns, VSS,
+ 298808.800000ns, VSS,
+ 298808.900000ns, VDD,
+ 298928.900000ns, VDD,
+ 298929.000000ns, VSS,
+ 299289.200000ns, VSS,
+ 299289.300000ns, VDD,
+ 300009.800000ns, VDD,
+ 300009.900000ns, VSS,
+ 300490.200000ns, VSS,
+ 300490.300000ns, VDD,
+ 301090.700000ns, VDD,
+ 301090.800000ns, VSS,
+ 301811.300000ns, VSS,
+ 301811.400000ns, VDD,
+ 302171.600000ns, VDD,
+ 302171.700000ns, VSS,
+ 302772.100000ns, VSS,
+ 302772.200000ns, VDD,
+ 303612.800000ns, VDD,
+ 303612.900000ns, VSS,
+ 303732.900000ns, VSS,
+ 303733.000000ns, VDD,
+ 304213.300000ns, VDD,
+ 304213.400000ns, VSS,
+ 304693.700000ns, VSS,
+ 304693.800000ns, VDD,
+ 305174.100000ns, VDD,
+ 305174.200000ns, VSS,
+ 305534.400000ns, VSS,
+ 305534.500000ns, VDD,
+ 306735.400000ns, VDD,
+ 306735.500000ns, VSS,
+ 307095.700000ns, VSS,
+ 307095.800000ns, VDD,
+ 307215.800000ns, VDD,
+ 307215.900000ns, VSS,
+ 307335.900000ns, VSS,
+ 307336.000000ns, VDD,
+ 307576.100000ns, VDD,
+ 307576.200000ns, VSS,
+ 307816.300000ns, VSS,
+ 307816.400000ns, VDD,
+ 308176.600000ns, VDD,
+ 308176.700000ns, VSS,
+ 309017.300000ns, VSS,
+ 309017.400000ns, VDD,
+ 309137.400000ns, VDD,
+ 309137.500000ns, VSS,
+ 310098.200000ns, VSS,
+ 310098.300000ns, VDD,
+ 310218.300000ns, VDD,
+ 310218.400000ns, VSS,
+ 310698.700000ns, VSS,
+ 310698.800000ns, VDD,
+ 310818.800000ns, VDD,
+ 310818.900000ns, VSS,
+ 312019.800000ns, VSS,
+ 312019.900000ns, VDD,
+ 312260.000000ns, VDD,
+ 312260.100000ns, VSS,
+ 312380.100000ns, VSS,
+ 312380.200000ns, VDD,
+ 313220.800000ns, VDD,
+ 313220.900000ns, VSS,
+ 313701.200000ns, VSS,
+ 313701.300000ns, VDD,
+ 313941.400000ns, VDD,
+ 313941.500000ns, VSS,
+ 314782.100000ns, VSS,
+ 314782.200000ns, VDD,
+ 315142.400000ns, VDD,
+ 315142.500000ns, VSS,
+ 316223.300000ns, VSS,
+ 316223.400000ns, VDD,
+ 316823.800000ns, VDD,
+ 316823.900000ns, VSS,
+ 316943.900000ns, VSS,
+ 316944.000000ns, VDD,
+ 317184.100000ns, VDD,
+ 317184.200000ns, VSS,
+ 317424.300000ns, VSS,
+ 317424.400000ns, VDD,
+ 317664.500000ns, VDD,
+ 317664.600000ns, VSS,
+ 318385.100000ns, VSS,
+ 318385.200000ns, VDD,
+ 318745.400000ns, VDD,
+ 318745.500000ns, VSS,
+ 318865.500000ns, VSS,
+ 318865.600000ns, VDD,
+ 319466.000000ns, VDD,
+ 319466.100000ns, VSS,
+ 320787.100000ns, VSS,
+ 320787.200000ns, VDD,
+ 321027.300000ns, VDD,
+ 321027.400000ns, VSS,
+ 321147.400000ns, VSS,
+ 321147.500000ns, VDD,
+ 321868.000000ns, VDD,
+ 321868.100000ns, VSS,
+ 322108.200000ns, VSS,
+ 322108.300000ns, VDD,
+ 322588.600000ns, VDD,
+ 322588.700000ns, VSS,
+ 322708.700000ns, VSS,
+ 322708.800000ns, VDD,
+ 322828.800000ns, VDD,
+ 322828.900000ns, VSS,
+ 322948.900000ns, VSS,
+ 322949.000000ns, VDD,
+ 323189.100000ns, VDD,
+ 323189.200000ns, VSS,
+ 323549.400000ns, VSS,
+ 323549.500000ns, VDD,
+ 324029.800000ns, VDD,
+ 324029.900000ns, VSS,
+ 324510.200000ns, VSS,
+ 324510.300000ns, VDD,
+ 324870.500000ns, VDD,
+ 324870.600000ns, VSS,
+ 325110.700000ns, VSS,
+ 325110.800000ns, VDD,
+ 325350.900000ns, VDD,
+ 325351.000000ns, VSS,
+ 325711.200000ns, VSS,
+ 325711.300000ns, VDD,
+ 326071.500000ns, VDD,
+ 326071.600000ns, VSS,
+ 326191.600000ns, VSS,
+ 326191.700000ns, VDD,
+ 327632.800000ns, VDD,
+ 327632.900000ns, VSS,
+ 327993.100000ns, VSS,
+ 327993.200000ns, VDD,
+ 328833.800000ns, VDD,
+ 328833.900000ns, VSS,
+ 329194.100000ns, VSS,
+ 329194.200000ns, VDD,
+ 329794.600000ns, VDD,
+ 329794.700000ns, VSS,
+ 329914.700000ns, VSS,
+ 329914.800000ns, VDD,
+ 330154.900000ns, VDD,
+ 330155.000000ns, VSS,
+ 330275.000000ns, VSS,
+ 330275.100000ns, VDD,
+ 330515.200000ns, VDD,
+ 330515.300000ns, VSS,
+ 330755.400000ns, VSS,
+ 330755.500000ns, VDD,
+ 330995.600000ns, VDD,
+ 330995.700000ns, VSS,
+ 331235.800000ns, VSS,
+ 331235.900000ns, VDD,
+ 331355.900000ns, VDD,
+ 331356.000000ns, VSS,
+ 331836.300000ns, VSS,
+ 331836.400000ns, VDD,
+ 332316.700000ns, VDD,
+ 332316.800000ns, VSS,
+ 332436.800000ns, VSS,
+ 332436.900000ns, VDD,
+ 332677.000000ns, VDD,
+ 332677.100000ns, VSS,
+ 332797.100000ns, VSS,
+ 332797.200000ns, VDD,
+ 332917.200000ns, VDD,
+ 332917.300000ns, VSS,
+ 333037.300000ns, VSS,
+ 333037.400000ns, VDD,
+ 333517.700000ns, VDD,
+ 333517.800000ns, VSS,
+ 333637.800000ns, VSS,
+ 333637.900000ns, VDD,
+ 333878.000000ns, VDD,
+ 333878.100000ns, VSS,
+ 334238.300000ns, VSS,
+ 334238.400000ns, VDD,
+ 334718.700000ns, VDD,
+ 334718.800000ns, VSS,
+ 335439.300000ns, VSS,
+ 335439.400000ns, VDD,
+ 335679.500000ns, VDD,
+ 335679.600000ns, VSS,
+ 336400.100000ns, VSS,
+ 336400.200000ns, VDD,
+ 337240.800000ns, VDD,
+ 337240.900000ns, VSS,
+ 337481.000000ns, VSS,
+ 337481.100000ns, VDD,
+ 337961.400000ns, VDD,
+ 337961.500000ns, VSS,
+ 338682.000000ns, VSS,
+ 338682.100000ns, VDD,
+ 339762.900000ns, VDD,
+ 339763.000000ns, VSS,
+ 339883.000000ns, VSS,
+ 339883.100000ns, VDD,
+ 340483.500000ns, VDD,
+ 340483.600000ns, VSS,
+ 340603.600000ns, VSS,
+ 340603.700000ns, VDD,
+ 340843.800000ns, VDD,
+ 340843.900000ns, VSS,
+ 341204.100000ns, VSS,
+ 341204.200000ns, VDD,
+ 341804.600000ns, VDD,
+ 341804.700000ns, VSS,
+ 341924.700000ns, VSS,
+ 341924.800000ns, VDD,
+ 342405.100000ns, VDD,
+ 342405.200000ns, VSS,
+ 342765.400000ns, VSS,
+ 342765.500000ns, VDD,
+ 343365.900000ns, VDD,
+ 343366.000000ns, VSS,
+ 343966.400000ns, VSS,
+ 343966.500000ns, VDD,
+ 344446.800000ns, VDD,
+ 344446.900000ns, VSS,
+ 344687.000000ns, VSS,
+ 344687.100000ns, VDD,
+ 344927.200000ns, VDD,
+ 344927.300000ns, VSS,
+ 345407.600000ns, VSS,
+ 345407.700000ns, VDD,
+ 345527.700000ns, VDD,
+ 345527.800000ns, VSS,
+ 345888.000000ns, VSS,
+ 345888.100000ns, VDD,
+ 346128.200000ns, VDD,
+ 346128.300000ns, VSS,
+ 346488.500000ns, VSS,
+ 346488.600000ns, VDD,
+ 346848.800000ns, VDD,
+ 346848.900000ns, VSS,
+ 347329.200000ns, VSS,
+ 347329.300000ns, VDD,
+ 348169.900000ns, VDD,
+ 348170.000000ns, VSS,
+ 348410.100000ns, VSS,
+ 348410.200000ns, VDD,
+ 348650.300000ns, VDD,
+ 348650.400000ns, VSS,
+ 348770.400000ns, VSS,
+ 348770.500000ns, VDD,
+ 349851.300000ns, VDD,
+ 349851.400000ns, VSS,
+ 351052.300000ns, VSS,
+ 351052.400000ns, VDD,
+ 351172.400000ns, VDD,
+ 351172.500000ns, VSS,
+ 351412.600000ns, VSS,
+ 351412.700000ns, VDD,
+ 351652.800000ns, VDD,
+ 351652.900000ns, VSS,
+ 352013.100000ns, VSS,
+ 352013.200000ns, VDD,
+ 352373.400000ns, VDD,
+ 352373.500000ns, VSS,
+ 352493.500000ns, VSS,
+ 352493.600000ns, VDD,
+ 352973.900000ns, VDD,
+ 352974.000000ns, VSS,
+ 353454.300000ns, VSS,
+ 353454.400000ns, VDD,
+ 353694.500000ns, VDD,
+ 353694.600000ns, VSS,
+ 353814.600000ns, VSS,
+ 353814.700000ns, VDD,
+ 355135.700000ns, VDD,
+ 355135.800000ns, VSS,
+ 355375.900000ns, VSS,
+ 355376.000000ns, VDD,
+ 356216.600000ns, VDD,
+ 356216.700000ns, VSS,
+ 356456.800000ns, VSS,
+ 356456.900000ns, VDD,
+ 357057.300000ns, VDD,
+ 357057.400000ns, VSS,
+ 357177.400000ns, VSS,
+ 357177.500000ns, VDD,
+ 357417.600000ns, VDD,
+ 357417.700000ns, VSS,
+ 357657.800000ns, VSS,
+ 357657.900000ns, VDD,
+ 357898.000000ns, VDD,
+ 357898.100000ns, VSS,
+ 358138.200000ns, VSS,
+ 358138.300000ns, VDD,
+ 358378.400000ns, VDD,
+ 358378.500000ns, VSS,
+ 358858.800000ns, VSS,
+ 358858.900000ns, VDD,
+ 359219.100000ns, VDD,
+ 359219.200000ns, VSS,
+ 359339.200000ns, VSS,
+ 359339.300000ns, VDD,
+ 360420.100000ns, VDD,
+ 360420.200000ns, VSS,
+ 361380.900000ns, VSS,
+ 361381.000000ns, VDD,
+ 361981.400000ns, VDD,
+ 361981.500000ns, VSS,
+ 362101.500000ns, VSS,
+ 362101.600000ns, VDD,
+ 362822.100000ns, VDD,
+ 362822.200000ns, VSS,
+ 364143.200000ns, VSS,
+ 364143.300000ns, VDD,
+ 364743.700000ns, VDD,
+ 364743.800000ns, VSS,
+ 364863.800000ns, VSS,
+ 364863.900000ns, VDD,
+ 365104.000000ns, VDD,
+ 365104.100000ns, VSS,
+ 365464.300000ns, VSS,
+ 365464.400000ns, VDD,
+ 365584.400000ns, VDD,
+ 365584.500000ns, VSS,
+ 365704.500000ns, VSS,
+ 365704.600000ns, VDD,
+ 366184.900000ns, VDD,
+ 366185.000000ns, VSS,
+ 366665.300000ns, VSS,
+ 366665.400000ns, VDD,
+ 367025.600000ns, VDD,
+ 367025.700000ns, VSS,
+ 367145.700000ns, VSS,
+ 367145.800000ns, VDD,
+ 367265.800000ns, VDD,
+ 367265.900000ns, VSS,
+ 367866.300000ns, VSS,
+ 367866.400000ns, VDD,
+ 369187.400000ns, VDD,
+ 369187.500000ns, VSS,
+ 369547.700000ns, VSS,
+ 369547.800000ns, VDD,
+ 369667.800000ns, VDD,
+ 369667.900000ns, VSS,
+ 369908.000000ns, VSS,
+ 369908.100000ns, VDD,
+ 370628.600000ns, VDD,
+ 370628.700000ns, VSS,
+ 370748.700000ns, VSS,
+ 370748.800000ns, VDD,
+ 371469.300000ns, VDD,
+ 371469.400000ns, VSS,
+ 371589.400000ns, VSS,
+ 371589.500000ns, VDD,
+ 371709.500000ns, VDD,
+ 371709.600000ns, VSS,
+ 372189.900000ns, VSS,
+ 372190.000000ns, VDD,
+ 372310.000000ns, VDD,
+ 372310.100000ns, VSS,
+ 372910.500000ns, VSS,
+ 372910.600000ns, VDD,
+ 373390.900000ns, VDD,
+ 373391.000000ns, VSS,
+ 373871.300000ns, VSS,
+ 373871.400000ns, VDD,
+ 374351.700000ns, VDD,
+ 374351.800000ns, VSS,
+ 374471.800000ns, VSS,
+ 374471.900000ns, VDD,
+ 374712.000000ns, VDD,
+ 374712.100000ns, VSS,
+ 375072.300000ns, VSS,
+ 375072.400000ns, VDD,
+ 375192.400000ns, VDD,
+ 375192.500000ns, VSS,
+ 375312.500000ns, VSS,
+ 375312.600000ns, VDD,
+ 376033.100000ns, VDD,
+ 376033.200000ns, VSS,
+ 376153.200000ns, VSS,
+ 376153.300000ns, VDD,
+ 376393.400000ns, VDD,
+ 376393.500000ns, VSS,
+ 376753.700000ns, VSS,
+ 376753.800000ns, VDD,
+ 376873.800000ns, VDD,
+ 376873.900000ns, VSS,
+ 376993.900000ns, VSS,
+ 376994.000000ns, VDD,
+ 377234.100000ns, VDD,
+ 377234.200000ns, VSS,
+ 377354.200000ns, VSS,
+ 377354.300000ns, VDD,
+ 378315.000000ns, VDD,
+ 378315.100000ns, VSS,
+ 378795.400000ns, VSS,
+ 378795.500000ns, VDD,
+ 379395.900000ns, VDD,
+ 379396.000000ns, VSS,
+ 380116.500000ns, VSS,
+ 380116.600000ns, VDD,
+ 380717.000000ns, VDD,
+ 380717.100000ns, VSS,
+ 381317.500000ns, VSS,
+ 381317.600000ns, VDD,
+ 381557.700000ns, VDD,
+ 381557.800000ns, VSS,
+ 381918.000000ns, VSS,
+ 381918.100000ns, VDD,
+ 382038.100000ns, VDD,
+ 382038.200000ns, VSS,
+ 382158.200000ns, VSS,
+ 382158.300000ns, VDD,
+ 382398.400000ns, VDD,
+ 382398.500000ns, VSS,
+ 382518.500000ns, VSS,
+ 382518.600000ns, VDD,
+ 382758.700000ns, VDD,
+ 382758.800000ns, VSS,
+ 382998.900000ns, VSS,
+ 382999.000000ns, VDD,
+ 383239.100000ns, VDD,
+ 383239.200000ns, VSS,
+ 383479.300000ns, VSS,
+ 383479.400000ns, VDD,
+ 383719.500000ns, VDD,
+ 383719.600000ns, VSS,
+ 384079.800000ns, VSS,
+ 384079.900000ns, VDD,
+ 384199.900000ns, VDD,
+ 384200.000000ns, VSS,
+ 384320.000000ns, VSS,
+ 384320.100000ns, VDD,
+ 384440.100000ns, VDD,
+ 384440.200000ns, VSS,
+ 384800.400000ns, VSS,
+ 384800.500000ns, VDD,
+ 385040.600000ns, VDD,
+ 385040.700000ns, VSS,
+ 385400.900000ns, VSS,
+ 385401.000000ns, VDD,
+ 385521.000000ns, VDD,
+ 385521.100000ns, VSS,
+ 386361.700000ns, VSS,
+ 386361.800000ns, VDD,
+ 386601.900000ns, VDD,
+ 386602.000000ns, VSS,
+ 386962.200000ns, VSS,
+ 386962.300000ns, VDD,
+ 387082.300000ns, VDD,
+ 387082.400000ns, VSS,
+ 387202.400000ns, VSS,
+ 387202.500000ns, VDD,
+ 387562.700000ns, VDD,
+ 387562.800000ns, VSS,
+ 387682.800000ns, VSS,
+ 387682.900000ns, VDD,
+ 388043.100000ns, VDD,
+ 388043.200000ns, VSS,
+ 388163.200000ns, VSS,
+ 388163.300000ns, VDD,
+ 388883.800000ns, VDD,
+ 388883.900000ns, VSS,
+ 389003.900000ns, VSS,
+ 389004.000000ns, VDD,
+ 389364.200000ns, VDD,
+ 389364.300000ns, VSS,
+ 389724.500000ns, VSS,
+ 389724.600000ns, VDD,
+ 391285.800000ns, VDD,
+ 391285.900000ns, VSS,
+ 391886.300000ns, VSS,
+ 391886.400000ns, VDD,
+ 392246.600000ns, VDD,
+ 392246.700000ns, VSS,
+ 392486.800000ns, VSS,
+ 392486.900000ns, VDD,
+ 393807.900000ns, VDD,
+ 393808.000000ns, VSS,
+ 394408.400000ns, VSS,
+ 394408.500000ns, VDD,
+ 394888.800000ns, VDD,
+ 394888.900000ns, VSS,
+ 395008.900000ns, VSS,
+ 395009.000000ns, VDD,
+ 395249.100000ns, VDD,
+ 395249.200000ns, VSS,
+ 395609.400000ns, VSS,
+ 395609.500000ns, VDD,
+ 395729.500000ns, VDD,
+ 395729.600000ns, VSS,
+ 395849.600000ns, VSS,
+ 395849.700000ns, VDD,
+ 396089.800000ns, VDD,
+ 396089.900000ns, VSS,
+ 396450.100000ns, VSS,
+ 396450.200000ns, VDD,
+ 396810.400000ns, VDD,
+ 396810.500000ns, VSS,
+ 397410.900000ns, VSS,
+ 397411.000000ns, VDD,
+ 397891.300000ns, VDD,
+ 397891.400000ns, VSS,
+ 398972.200000ns, VSS,
+ 398972.300000ns, VDD,
+ 399212.400000ns, VDD,
+ 399212.500000ns, VSS,
+ 399452.600000ns, VSS,
+ 399452.700000ns, VDD,
+ 399812.900000ns, VDD,
+ 399813.000000ns, VSS,
+ 400533.500000ns, VSS,
+ 400533.600000ns, VDD,
+ 403415.900000ns, VDD,
+ 403416.000000ns, VSS,
+ 403536.000000ns, VSS,
+ 403536.100000ns, VDD,
+ 404857.100000ns, VDD,
+ 404857.200000ns, VSS,
+ 404977.200000ns, VSS,
+ 404977.300000ns, VDD,
+ 405217.400000ns, VDD,
+ 405217.500000ns, VSS,
+ 405457.600000ns, VSS,
+ 405457.700000ns, VDD,
+ 406298.300000ns, VDD,
+ 406298.400000ns, VSS,
+ 406418.400000ns, VSS,
+ 406418.500000ns, VDD,
+ 406538.500000ns, VDD,
+ 406538.600000ns, VSS,
+ 406898.800000ns, VSS,
+ 406898.900000ns, VDD,
+ 407379.200000ns, VDD,
+ 407379.300000ns, VSS,
+ 407499.300000ns, VSS,
+ 407499.400000ns, VDD,
+ 408219.900000ns, VDD,
+ 408220.000000ns, VSS,
+ 408580.200000ns, VSS,
+ 408580.300000ns, VDD,
+ 409300.800000ns, VDD,
+ 409300.900000ns, VSS,
+ 410021.400000ns, VSS,
+ 410021.500000ns, VDD,
+ 410381.700000ns, VDD,
+ 410381.800000ns, VSS,
+ 411342.500000ns, VSS,
+ 411342.600000ns, VDD,
+ 411462.600000ns, VDD,
+ 411462.700000ns, VSS,
+ 411702.800000ns, VSS,
+ 411702.900000ns, VDD,
+ 411822.900000ns, VDD,
+ 411823.000000ns, VSS,
+ 412663.600000ns, VSS,
+ 412663.700000ns, VDD,
+ 412903.800000ns, VDD,
+ 412903.900000ns, VSS,
+ 413144.000000ns, VSS,
+ 413144.100000ns, VDD,
+ 414345.000000ns, VDD,
+ 414345.100000ns, VSS,
+ 415185.700000ns, VSS,
+ 415185.800000ns, VDD,
+ 415666.100000ns, VDD,
+ 415666.200000ns, VSS,
+ 416026.400000ns, VSS,
+ 416026.500000ns, VDD,
+ 416266.600000ns, VDD,
+ 416266.700000ns, VSS,
+ 416506.800000ns, VSS,
+ 416506.900000ns, VDD,
+ 416747.000000ns, VDD,
+ 416747.100000ns, VSS,
+ 417347.500000ns, VSS,
+ 417347.600000ns, VDD,
+ 417707.800000ns, VDD,
+ 417707.900000ns, VSS,
+ 419149.000000ns, VSS,
+ 419149.100000ns, VDD,
+ 419749.500000ns, VDD,
+ 419749.600000ns, VSS,
+ 420229.900000ns, VSS,
+ 420230.000000ns, VDD,
+ 420830.400000ns, VDD,
+ 420830.500000ns, VSS,
+ 421671.100000ns, VSS,
+ 421671.200000ns, VDD,
+ 422271.600000ns, VDD,
+ 422271.700000ns, VSS,
+ 423112.300000ns, VSS,
+ 423112.400000ns, VDD,
+ 423352.500000ns, VDD,
+ 423352.600000ns, VSS,
+ 423592.700000ns, VSS,
+ 423592.800000ns, VDD,
+ 423953.000000ns, VDD,
+ 423953.100000ns, VSS,
+ 424073.100000ns, VSS,
+ 424073.200000ns, VDD,
+ 424433.400000ns, VDD,
+ 424433.500000ns, VSS,
+ 424553.500000ns, VSS,
+ 424553.600000ns, VDD,
+ 425033.900000ns, VDD,
+ 425034.000000ns, VSS,
+ 425154.000000ns, VSS,
+ 425154.100000ns, VDD,
+ 425754.500000ns, VDD,
+ 425754.600000ns, VSS,
+ 425874.600000ns, VSS,
+ 425874.700000ns, VDD,
+ 426114.800000ns, VDD,
+ 426114.900000ns, VSS,
+ 426475.100000ns, VSS,
+ 426475.200000ns, VDD,
+ 426835.400000ns, VDD,
+ 426835.500000ns, VSS,
+ 427075.600000ns, VSS,
+ 427075.700000ns, VDD,
+ 427195.700000ns, VDD,
+ 427195.800000ns, VSS,
+ 427916.300000ns, VSS,
+ 427916.400000ns, VDD,
+ 428396.700000ns, VDD,
+ 428396.800000ns, VSS,
+ 428757.000000ns, VSS,
+ 428757.100000ns, VDD,
+ 429117.300000ns, VDD,
+ 429117.400000ns, VSS,
+ 429837.900000ns, VSS,
+ 429838.000000ns, VDD,
+ 430438.400000ns, VDD,
+ 430438.500000ns, VSS,
+ 430558.500000ns, VSS,
+ 430558.600000ns, VDD,
+ 431159.000000ns, VDD,
+ 431159.100000ns, VSS,
+ 431759.500000ns, VSS,
+ 431759.600000ns, VDD,
+ 432360.000000ns, VDD,
+ 432360.100000ns, VSS,
+ 432840.400000ns, VSS,
+ 432840.500000ns, VDD,
+ 433320.800000ns, VDD,
+ 433320.900000ns, VSS,
+ 433440.900000ns, VSS,
+ 433441.000000ns, VDD,
+ 433681.100000ns, VDD,
+ 433681.200000ns, VSS,
+ 433801.200000ns, VSS,
+ 433801.300000ns, VDD,
+ 434641.900000ns, VDD,
+ 434642.000000ns, VSS,
+ 434762.000000ns, VSS,
+ 434762.100000ns, VDD,
+ 435122.300000ns, VDD,
+ 435122.400000ns, VSS,
+ 435722.800000ns, VSS,
+ 435722.900000ns, VDD,
+ 436323.300000ns, VDD,
+ 436323.400000ns, VSS,
+ 437284.100000ns, VSS,
+ 437284.200000ns, VDD,
+ 437404.200000ns, VDD,
+ 437404.300000ns, VSS,
+ 437644.400000ns, VSS,
+ 437644.500000ns, VDD,
+ 438365.000000ns, VDD,
+ 438365.100000ns, VSS,
+ 438725.300000ns, VSS,
+ 438725.400000ns, VDD,
+ 439686.100000ns, VDD,
+ 439686.200000ns, VSS,
+ 439926.300000ns, VSS,
+ 439926.400000ns, VDD,
+ 441007.200000ns, VDD,
+ 441007.300000ns, VSS,
+ 441247.400000ns, VSS,
+ 441247.500000ns, VDD,
+ 441487.600000ns, VDD,
+ 441487.700000ns, VSS,
+ 441847.900000ns, VSS,
+ 441848.000000ns, VDD,
+ 442328.300000ns, VDD,
+ 442328.400000ns, VSS,
+ 442568.500000ns, VSS,
+ 442568.600000ns, VDD,
+ 442808.700000ns, VDD,
+ 442808.800000ns, VSS,
+ 443289.100000ns, VSS,
+ 443289.200000ns, VDD,
+ 444009.700000ns, VDD,
+ 444009.800000ns, VSS,
+ 444249.900000ns, VSS,
+ 444250.000000ns, VDD,
+ 444490.100000ns, VDD,
+ 444490.200000ns, VSS,
+ 444850.400000ns, VSS,
+ 444850.500000ns, VDD,
+ 446411.700000ns, VDD,
+ 446411.800000ns, VSS,
+ 446651.900000ns, VSS,
+ 446652.000000ns, VDD,
+ 446892.100000ns, VDD,
+ 446892.200000ns, VSS,
+ 448333.300000ns, VSS,
+ 448333.400000ns, VDD,
+ 448573.500000ns, VDD,
+ 448573.600000ns, VSS,
+ 448813.700000ns, VSS,
+ 448813.800000ns, VDD,
+ 448933.800000ns, VDD,
+ 448933.900000ns, VSS,
+ 449053.900000ns, VSS,
+ 449054.000000ns, VDD,
+ 449414.200000ns, VDD,
+ 449414.300000ns, VSS,
+ 449774.500000ns, VSS,
+ 449774.600000ns, VDD,
+ 450014.700000ns, VDD,
+ 450014.800000ns, VSS,
+ 450375.000000ns, VSS,
+ 450375.100000ns, VDD,
+ 450615.200000ns, VDD,
+ 450615.300000ns, VSS,
+ 451215.700000ns, VSS,
+ 451215.800000ns, VDD,
+ 451576.000000ns, VDD,
+ 451576.100000ns, VSS,
+ 451936.300000ns, VSS,
+ 451936.400000ns, VDD,
+ 452056.400000ns, VDD,
+ 452056.500000ns, VSS,
+ 452897.100000ns, VSS,
+ 452897.200000ns, VDD,
+ 453017.200000ns, VDD,
+ 453017.300000ns, VSS,
+ 453137.300000ns, VSS,
+ 453137.400000ns, VDD,
+ 453978.000000ns, VDD,
+ 453978.100000ns, VSS,
+ 455058.900000ns, VSS,
+ 455059.000000ns, VDD,
+ 455779.500000ns, VDD,
+ 455779.600000ns, VSS,
+ 456019.700000ns, VSS,
+ 456019.800000ns, VDD,
+ 456380.000000ns, VDD,
+ 456380.100000ns, VSS,
+ 457340.800000ns, VSS,
+ 457340.900000ns, VDD,
+ 457581.000000ns, VDD,
+ 457581.100000ns, VSS,
+ 458061.400000ns, VSS,
+ 458061.500000ns, VDD,
+ 458541.800000ns, VDD,
+ 458541.900000ns, VSS,
+ 458661.900000ns, VSS,
+ 458662.000000ns, VDD,
+ 458902.100000ns, VDD,
+ 458902.200000ns, VSS,
+ 459262.400000ns, VSS,
+ 459262.500000ns, VDD,
+ 459742.800000ns, VDD,
+ 459742.900000ns, VSS,
+ 460103.100000ns, VSS,
+ 460103.200000ns, VDD,
+ 460223.200000ns, VDD,
+ 460223.300000ns, VSS,
+ 460463.400000ns, VSS,
+ 460463.500000ns, VDD,
+ 460583.500000ns, VDD,
+ 460583.600000ns, VSS,
+ 461184.000000ns, VSS,
+ 461184.100000ns, VDD,
+ 461664.400000ns, VDD,
+ 461664.500000ns, VSS,
+ 461784.500000ns, VSS,
+ 461784.600000ns, VDD,
+ 462625.200000ns, VDD,
+ 462625.300000ns, VSS,
+ 462745.300000ns, VSS,
+ 462745.400000ns, VDD,
+ 463105.600000ns, VDD,
+ 463105.700000ns, VSS,
+ 463225.700000ns, VSS,
+ 463225.800000ns, VDD,
+ 464426.700000ns, VDD,
+ 464426.800000ns, VSS,
+ 464546.800000ns, VSS,
+ 464546.900000ns, VDD,
+ 464907.100000ns, VDD,
+ 464907.200000ns, VSS,
+ 465267.400000ns, VSS,
+ 465267.500000ns, VDD,
+ 465507.600000ns, VDD,
+ 465507.700000ns, VSS,
+ 466588.500000ns, VSS,
+ 466588.600000ns, VDD,
+ 466948.800000ns, VDD,
+ 466948.900000ns, VSS,
+ 468630.200000ns, VSS,
+ 468630.300000ns, VDD,
+ 468870.400000ns, VDD,
+ 468870.500000ns, VSS,
+ 469110.600000ns, VSS,
+ 469110.700000ns, VDD,
+ 469230.700000ns, VDD,
+ 469230.800000ns, VSS,
+ 469711.100000ns, VSS,
+ 469711.200000ns, VDD,
+ 469951.300000ns, VDD,
+ 469951.400000ns, VSS,
+ 470311.600000ns, VSS,
+ 470311.700000ns, VDD,
+ 470431.700000ns, VDD,
+ 470431.800000ns, VSS,
+ 470551.800000ns, VSS,
+ 470551.900000ns, VDD,
+ 470912.100000ns, VDD,
+ 470912.200000ns, VSS,
+ 471392.500000ns, VSS,
+ 471392.600000ns, VDD,
+ 472113.100000ns, VDD,
+ 472113.200000ns, VSS,
+ 473194.000000ns, VSS,
+ 473194.100000ns, VDD,
+ 473314.100000ns, VDD,
+ 473314.200000ns, VSS,
+ 473794.500000ns, VSS,
+ 473794.600000ns, VDD,
+ 474154.800000ns, VDD,
+ 474154.900000ns, VSS,
+ 474515.100000ns, VSS,
+ 474515.200000ns, VDD,
+ 474635.200000ns, VDD,
+ 474635.300000ns, VSS,
+ 474755.300000ns, VSS,
+ 474755.400000ns, VDD,
+ 474995.500000ns, VDD,
+ 474995.600000ns, VSS,
+ 475355.800000ns, VSS,
+ 475355.900000ns, VDD,
+ 476316.600000ns, VDD,
+ 476316.700000ns, VSS,
+ 476797.000000ns, VSS,
+ 476797.100000ns, VDD,
+ 476917.100000ns, VDD,
+ 476917.200000ns, VSS,
+ 477397.500000ns, VSS,
+ 477397.600000ns, VDD,
+ 477757.800000ns, VDD,
+ 477757.900000ns, VSS,
+ 478718.600000ns, VSS,
+ 478718.700000ns, VDD,
+ 479439.200000ns, VDD,
+ 479439.300000ns, VSS,
+ 480520.100000ns, VSS,
+ 480520.200000ns, VDD,
+ 481000.500000ns, VDD,
+ 481000.600000ns, VSS,
+ 481120.600000ns, VSS,
+ 481120.700000ns, VDD,
+ 481360.800000ns, VDD,
+ 481360.900000ns, VSS,
+ 481721.100000ns, VSS,
+ 481721.200000ns, VDD,
+ 482081.400000ns, VDD,
+ 482081.500000ns, VSS,
+ 482201.500000ns, VSS,
+ 482201.600000ns, VDD,
+ 482561.800000ns, VDD,
+ 482561.900000ns, VSS,
+ 482681.900000ns, VSS,
+ 482682.000000ns, VDD,
+ 483402.500000ns, VDD,
+ 483402.600000ns, VSS,
+ 483762.800000ns, VSS,
+ 483762.900000ns, VDD,
+ 483882.900000ns, VDD,
+ 483883.000000ns, VSS,
+ 484243.200000ns, VSS,
+ 484243.300000ns, VDD,
+ 484363.300000ns, VDD,
+ 484363.400000ns, VSS,
+ 484963.800000ns, VSS,
+ 484963.900000ns, VDD,
+ 485083.900000ns, VDD,
+ 485084.000000ns, VSS,
+ 485444.200000ns, VSS,
+ 485444.300000ns, VDD,
+ 485564.300000ns, VDD,
+ 485564.400000ns, VSS,
+ 485804.500000ns, VSS,
+ 485804.600000ns, VDD,
+ 485924.600000ns, VDD,
+ 485924.700000ns, VSS,
+ 486164.800000ns, VSS,
+ 486164.900000ns, VDD,
+ 486525.100000ns, VDD,
+ 486525.200000ns, VSS,
+ 486885.400000ns, VSS,
+ 486885.500000ns, VDD,
+ 487606.000000ns, VDD,
+ 487606.100000ns, VSS,
+ 487726.100000ns, VSS,
+ 487726.200000ns, VDD,
+ 488566.800000ns, VDD,
+ 488566.900000ns, VSS,
+ 488807.000000ns, VSS,
+ 488807.100000ns, VDD,
+ 489047.200000ns, VDD,
+ 489047.300000ns, VSS,
+ 489167.300000ns, VSS,
+ 489167.400000ns, VDD,
+ 489527.600000ns, VDD,
+ 489527.700000ns, VSS,
+ 489647.700000ns, VSS,
+ 489647.800000ns, VDD,
+ 489887.900000ns, VDD,
+ 489888.000000ns, VSS,
+ 490128.100000ns, VSS,
+ 490128.200000ns, VDD,
+ 490728.600000ns, VDD,
+ 490728.700000ns, VSS,
+ 490848.700000ns, VSS,
+ 490848.800000ns, VDD,
+ 491088.900000ns, VDD,
+ 491089.000000ns, VSS,
+ 491329.100000ns, VSS,
+ 491329.200000ns, VDD,
+ 492289.900000ns, VDD,
+ 492290.000000ns, VSS,
+ 492890.400000ns, VSS,
+ 492890.500000ns, VDD,
+ 493010.500000ns, VDD,
+ 493010.600000ns, VSS,
+ 493130.600000ns, VSS,
+ 493130.700000ns, VDD,
+ 493611.000000ns, VDD,
+ 493611.100000ns, VSS,
+ 493731.100000ns, VSS,
+ 493731.200000ns, VDD,
+ 493971.300000ns, VDD,
+ 493971.400000ns, VSS,
+ 494571.800000ns, VSS,
+ 494571.900000ns, VDD,
+ 494812.000000ns, VDD,
+ 494812.100000ns, VSS,
+ 495052.200000ns, VSS,
+ 495052.300000ns, VDD,
+ 495292.400000ns, VDD,
+ 495292.500000ns, VSS,
+ 495652.700000ns, VSS,
+ 495652.800000ns, VDD,
+ 495892.900000ns, VDD,
+ 495893.000000ns, VSS,
+ 496253.200000ns, VSS,
+ 496253.300000ns, VDD,
+ 496733.600000ns, VDD,
+ 496733.700000ns, VSS,
+ 497334.100000ns, VSS,
+ 497334.200000ns, VDD,
+ 497574.300000ns, VDD,
+ 497574.400000ns, VSS,
+ 497694.400000ns, VSS,
+ 497694.500000ns, VDD,
+ 498294.900000ns, VDD,
+ 498295.000000ns, VSS,
+ 498655.200000ns, VSS,
+ 498655.300000ns, VDD,
+ 498775.300000ns, VDD,
+ 498775.400000ns, VSS,
+ 499015.500000ns, VSS,
+ 499015.600000ns, VDD,
+ 500096.400000ns, VDD,
+ 500096.500000ns, VSS,
+ 500216.500000ns, VSS,
+ 500216.600000ns, VDD,
+ 500696.900000ns, VDD,
+ 500697.000000ns, VSS,
+ 500817.000000ns, VSS,
+ 500817.100000ns, VDD,
+ 500937.100000ns, VDD,
+ 500937.200000ns, VSS,
+ 501297.400000ns, VSS,
+ 501297.500000ns, VDD,
+ 502018.000000ns, VDD,
+ 502018.100000ns, VSS,
+ 502138.100000ns, VSS,
+ 502138.200000ns, VDD,
+ 502498.400000ns, VDD,
+ 502498.500000ns, VSS,
+ 502618.500000ns, VSS,
+ 502618.600000ns, VDD,
+ 502858.700000ns, VDD,
+ 502858.800000ns, VSS,
+ 502978.800000ns, VSS,
+ 502978.900000ns, VDD,
+ 503098.900000ns, VDD,
+ 503099.000000ns, VSS,
+ 503699.400000ns, VSS,
+ 503699.500000ns, VDD,
+ 503819.500000ns, VDD,
+ 503819.600000ns, VSS,
+ 504660.200000ns, VSS,
+ 504660.300000ns, VDD,
+ 504780.300000ns, VDD,
+ 504780.400000ns, VSS,
+ 505861.200000ns, VSS,
+ 505861.300000ns, VDD,
+ 505981.300000ns, VDD,
+ 505981.400000ns, VSS,
+ 506221.500000ns, VSS,
+ 506221.600000ns, VDD,
+ 506341.600000ns, VDD,
+ 506341.700000ns, VSS,
+ 506581.800000ns, VSS,
+ 506581.900000ns, VDD,
+ 507062.200000ns, VDD,
+ 507062.300000ns, VSS,
+ 507182.300000ns, VSS,
+ 507182.400000ns, VDD,
+ 507542.600000ns, VDD,
+ 507542.700000ns, VSS,
+ 507782.800000ns, VSS,
+ 507782.900000ns, VDD,
+ 508263.200000ns, VDD,
+ 508263.300000ns, VSS,
+ 508623.500000ns, VSS,
+ 508623.600000ns, VDD,
+ 508743.600000ns, VDD,
+ 508743.700000ns, VSS,
+ 509704.400000ns, VSS,
+ 509704.500000ns, VDD,
+ 510184.800000ns, VDD,
+ 510184.900000ns, VSS,
+ 510304.900000ns, VSS,
+ 510305.000000ns, VDD,
+ 510905.400000ns, VDD,
+ 510905.500000ns, VSS,
+ 511385.800000ns, VSS,
+ 511385.900000ns, VDD,
+ 511866.200000ns, VDD,
+ 511866.300000ns, VSS,
+ 512346.600000ns, VSS,
+ 512346.700000ns, VDD,
+ 512586.800000ns, VDD,
+ 512586.900000ns, VSS,
+ 512706.900000ns, VSS,
+ 512707.000000ns, VDD,
+ 513667.700000ns, VDD,
+ 513667.800000ns, VSS,
+ 514028.000000ns, VSS,
+ 514028.100000ns, VDD,
+ 514628.500000ns, VDD,
+ 514628.600000ns, VSS,
+ 514988.800000ns, VSS,
+ 514988.900000ns, VDD,
+ 515349.100000ns, VDD,
+ 515349.200000ns, VSS,
+ 516430.000000ns, VSS,
+ 516430.100000ns, VDD,
+ 516670.200000ns, VDD,
+ 516670.300000ns, VSS,
+ 517030.500000ns, VSS,
+ 517030.600000ns, VDD,
+ 517150.600000ns, VDD,
+ 517150.700000ns, VSS,
+ 517270.700000ns, VSS,
+ 517270.800000ns, VDD,
+ 517510.900000ns, VDD,
+ 517511.000000ns, VSS,
+ 517751.100000ns, VSS,
+ 517751.200000ns, VDD,
+ 519432.500000ns, VDD,
+ 519432.600000ns, VSS,
+ 519552.600000ns, VSS,
+ 519552.700000ns, VDD,
+ 520033.000000ns, VDD,
+ 520033.100000ns, VSS,
+ 520393.300000ns, VSS,
+ 520393.400000ns, VDD,
+ 520753.600000ns, VDD,
+ 520753.700000ns, VSS,
+ 521354.100000ns, VSS,
+ 521354.200000ns, VDD,
+ 521954.600000ns, VDD,
+ 521954.700000ns, VSS,
+ 522194.800000ns, VSS,
+ 522194.900000ns, VDD,
+ 522435.000000ns, VDD,
+ 522435.100000ns, VSS,
+ 522555.100000ns, VSS,
+ 522555.200000ns, VDD,
+ 523515.900000ns, VDD,
+ 523516.000000ns, VSS,
+ 523996.300000ns, VSS,
+ 523996.400000ns, VDD,
+ 524356.600000ns, VDD,
+ 524356.700000ns, VSS,
+ 524476.700000ns, VSS,
+ 524476.800000ns, VDD,
+ 524716.900000ns, VDD,
+ 524717.000000ns, VSS,
+ 526158.100000ns, VSS,
+ 526158.200000ns, VDD,
+ 527599.300000ns, VDD,
+ 527599.400000ns, VSS,
+ 527959.600000ns, VSS,
+ 527959.700000ns, VDD,
+ 528560.100000ns, VDD,
+ 528560.200000ns, VSS,
+ 528800.300000ns, VSS,
+ 528800.400000ns, VDD,
+ 528920.400000ns, VDD,
+ 528920.500000ns, VSS,
+ 529520.900000ns, VSS,
+ 529521.000000ns, VDD,
+ 530121.400000ns, VDD,
+ 530121.500000ns, VSS,
+ 530241.500000ns, VSS,
+ 530241.600000ns, VDD,
+ 531082.200000ns, VDD,
+ 531082.300000ns, VSS,
+ 531202.300000ns, VSS,
+ 531202.400000ns, VDD,
+ 531802.800000ns, VDD,
+ 531802.900000ns, VSS,
+ 532163.100000ns, VSS,
+ 532163.200000ns, VDD,
+ 532643.500000ns, VDD,
+ 532643.600000ns, VSS,
+ 532763.600000ns, VSS,
+ 532763.700000ns, VDD,
+ 533123.900000ns, VDD,
+ 533124.000000ns, VSS,
+ 533364.100000ns, VSS,
+ 533364.200000ns, VDD,
+ 533604.300000ns, VDD,
+ 533604.400000ns, VSS,
+ 533724.400000ns, VSS,
+ 533724.500000ns, VDD,
+ 534204.800000ns, VDD,
+ 534204.900000ns, VSS,
+ 535045.500000ns, VSS,
+ 535045.600000ns, VDD,
+ 535285.700000ns, VDD,
+ 535285.800000ns, VSS,
+ 535405.800000ns, VSS,
+ 535405.900000ns, VDD,
+ 535646.000000ns, VDD,
+ 535646.100000ns, VSS,
+ 536006.300000ns, VSS,
+ 536006.400000ns, VDD,
+ 536246.500000ns, VDD,
+ 536246.600000ns, VSS,
+ 536606.800000ns, VSS,
+ 536606.900000ns, VDD,
+ 537087.200000ns, VDD,
+ 537087.300000ns, VSS,
+ 537447.500000ns, VSS,
+ 537447.600000ns, VDD,
+ 537567.600000ns, VDD,
+ 537567.700000ns, VSS,
+ 537807.800000ns, VSS,
+ 537807.900000ns, VDD,
+ 537927.900000ns, VDD,
+ 537928.000000ns, VSS,
+ 538408.300000ns, VSS,
+ 538408.400000ns, VDD,
+ 538648.500000ns, VDD,
+ 538648.600000ns, VSS,
+ 538768.600000ns, VSS,
+ 538768.700000ns, VDD,
+ 539008.800000ns, VDD,
+ 539008.900000ns, VSS,
+ 539369.100000ns, VSS,
+ 539369.200000ns, VDD,
+ 539489.200000ns, VDD,
+ 539489.300000ns, VSS,
+ 539609.300000ns, VSS,
+ 539609.400000ns, VDD,
+ 539729.400000ns, VDD,
+ 539729.500000ns, VSS,
+ 540089.700000ns, VSS,
+ 540089.800000ns, VDD,
+ 540329.900000ns, VDD,
+ 540330.000000ns, VSS,
+ 540570.100000ns, VSS,
+ 540570.200000ns, VDD,
+ 540690.200000ns, VDD,
+ 540690.300000ns, VSS,
+ 541651.000000ns, VSS,
+ 541651.100000ns, VDD,
+ 541891.200000ns, VDD,
+ 541891.300000ns, VSS,
+ 542011.300000ns, VSS,
+ 542011.400000ns, VDD,
+ 542611.800000ns, VDD,
+ 542611.900000ns, VSS,
+ 543812.800000ns, VSS,
+ 543812.900000ns, VDD,
+ 544293.200000ns, VDD,
+ 544293.300000ns, VSS,
+ 544413.300000ns, VSS,
+ 544413.400000ns, VDD,
+ 544653.500000ns, VDD,
+ 544653.600000ns, VSS,
+ 545013.800000ns, VSS,
+ 545013.900000ns, VDD,
+ 545254.000000ns, VDD,
+ 545254.100000ns, VSS,
+ 545854.500000ns, VSS,
+ 545854.600000ns, VDD,
+ 546214.800000ns, VDD,
+ 546214.900000ns, VSS,
+ 546334.900000ns, VSS,
+ 546335.000000ns, VDD,
+ 546575.100000ns, VDD,
+ 546575.200000ns, VSS,
+ 546695.200000ns, VSS,
+ 546695.300000ns, VDD,
+ 546935.400000ns, VDD,
+ 546935.500000ns, VSS,
+ 547656.000000ns, VSS,
+ 547656.100000ns, VDD,
+ 547896.200000ns, VDD,
+ 547896.300000ns, VSS,
+ 548256.500000ns, VSS,
+ 548256.600000ns, VDD,
+ 548496.700000ns, VDD,
+ 548496.800000ns, VSS,
+ 549337.400000ns, VSS,
+ 549337.500000ns, VDD,
+ 549457.500000ns, VDD,
+ 549457.600000ns, VSS,
+ 549937.900000ns, VSS,
+ 549938.000000ns, VDD,
+ 550898.700000ns, VDD,
+ 550898.800000ns, VSS,
+ 551259.000000ns, VSS,
+ 551259.100000ns, VDD,
+ 553420.800000ns, VDD,
+ 553420.900000ns, VSS,
+ 554021.300000ns, VSS,
+ 554021.400000ns, VDD,
+ 554381.600000ns, VDD,
+ 554381.700000ns, VSS,
+ 554741.900000ns, VSS,
+ 554742.000000ns, VDD,
+ 555582.600000ns, VDD,
+ 555582.700000ns, VSS,
+ 555702.700000ns, VSS,
+ 555702.800000ns, VDD,
+ 555822.800000ns, VDD,
+ 555822.900000ns, VSS,
+ 555942.900000ns, VSS,
+ 555943.000000ns, VDD,
+ 556183.100000ns, VDD,
+ 556183.200000ns, VSS,
+ 556543.400000ns, VSS,
+ 556543.500000ns, VDD,
+ 557264.000000ns, VDD,
+ 557264.100000ns, VSS,
+ 557624.300000ns, VSS,
+ 557624.400000ns, VDD,
+ 557744.400000ns, VDD,
+ 557744.500000ns, VSS,
+ 557984.600000ns, VSS,
+ 557984.700000ns, VDD,
+ 558825.300000ns, VDD,
+ 558825.400000ns, VSS,
+ 559065.500000ns, VSS,
+ 559065.600000ns, VDD,
+ 559185.600000ns, VDD,
+ 559185.700000ns, VSS,
+ 560266.500000ns, VSS,
+ 560266.600000ns, VDD,
+ 560867.000000ns, VDD,
+ 560867.100000ns, VSS,
+ 561227.300000ns, VSS,
+ 561227.400000ns, VDD,
+ 561467.500000ns, VDD,
+ 561467.600000ns, VSS,
+ 561587.600000ns, VSS,
+ 561587.700000ns, VDD,
+ 561827.800000ns, VDD,
+ 561827.900000ns, VSS,
+ 562068.000000ns, VSS,
+ 562068.100000ns, VDD,
+ 562188.100000ns, VDD,
+ 562188.200000ns, VSS,
+ 563028.800000ns, VSS,
+ 563028.900000ns, VDD,
+ 563989.600000ns, VDD,
+ 563989.700000ns, VSS,
+ 564109.700000ns, VSS,
+ 564109.800000ns, VDD,
+ 565430.800000ns, VDD,
+ 565430.900000ns, VSS,
+ 565791.100000ns, VSS,
+ 565791.200000ns, VDD,
+ 566031.300000ns, VDD,
+ 566031.400000ns, VSS,
+ 566151.400000ns, VSS,
+ 566151.500000ns, VDD,
+ 566511.700000ns, VDD,
+ 566511.800000ns, VSS,
+ 566631.800000ns, VSS,
+ 566631.900000ns, VDD,
+ 566872.000000ns, VDD,
+ 566872.100000ns, VSS,
+ 566992.100000ns, VSS,
+ 566992.200000ns, VDD,
+ 567232.300000ns, VDD,
+ 567232.400000ns, VSS,
+ 567472.500000ns, VSS,
+ 567472.600000ns, VDD,
+ 567592.600000ns, VDD,
+ 567592.700000ns, VSS,
+ 568433.300000ns, VSS,
+ 568433.400000ns, VDD,
+ 568913.700000ns, VDD,
+ 568913.800000ns, VSS,
+ 569033.800000ns, VSS,
+ 569033.900000ns, VDD,
+ 569394.100000ns, VDD,
+ 569394.200000ns, VSS,
+ 570114.700000ns, VSS,
+ 570114.800000ns, VDD,
+ 570835.300000ns, VDD,
+ 570835.400000ns, VSS,
+ 570955.400000ns, VSS,
+ 570955.500000ns, VDD,
+ 571796.100000ns, VDD,
+ 571796.200000ns, VSS,
+ 572997.100000ns, VSS,
+ 572997.200000ns, VDD,
+ 573357.400000ns, VDD,
+ 573357.500000ns, VSS,
+ 573477.500000ns, VSS,
+ 573477.600000ns, VDD,
+ 573837.800000ns, VDD,
+ 573837.900000ns, VSS,
+ 575279.000000ns, VSS,
+ 575279.100000ns, VDD,
+ 576359.900000ns, VDD,
+ 576360.000000ns, VSS,
+ 576720.200000ns, VSS,
+ 576720.300000ns, VDD,
+ 577200.600000ns, VDD,
+ 577200.700000ns, VSS,
+ 577801.100000ns, VSS,
+ 577801.200000ns, VDD,
+ 578401.600000ns, VDD,
+ 578401.700000ns, VSS,
+ 578882.000000ns, VSS,
+ 578882.100000ns, VDD,
+ 579362.400000ns, VDD,
+ 579362.500000ns, VSS,
+ 580083.000000ns, VSS,
+ 580083.100000ns, VDD,
+ 580323.200000ns, VDD,
+ 580323.300000ns, VSS,
+ 580683.500000ns, VSS,
+ 580683.600000ns, VDD,
+ 581284.000000ns, VDD,
+ 581284.100000ns, VSS,
+ 581404.100000ns, VSS,
+ 581404.200000ns, VDD,
+ 582364.900000ns, VDD,
+ 582365.000000ns, VSS,
+ 582485.000000ns, VSS,
+ 582485.100000ns, VDD,
+ 582845.300000ns, VDD,
+ 582845.400000ns, VSS,
+ 583085.500000ns, VSS,
+ 583085.600000ns, VDD,
+ 583205.600000ns, VDD,
+ 583205.700000ns, VSS,
+ 583565.900000ns, VSS,
+ 583566.000000ns, VDD,
+ 583926.200000ns, VDD,
+ 583926.300000ns, VSS,
+ 584406.600000ns, VSS,
+ 584406.700000ns, VDD,
+ 584646.800000ns, VDD,
+ 584646.900000ns, VSS,
+ 585007.100000ns, VSS,
+ 585007.200000ns, VDD,
+ 585247.300000ns, VDD,
+ 585247.400000ns, VSS,
+ 585487.500000ns, VSS,
+ 585487.600000ns, VDD,
+ 585967.900000ns, VDD,
+ 585968.000000ns, VSS,
+ 586208.100000ns, VSS,
+ 586208.200000ns, VDD,
+ 586688.500000ns, VDD,
+ 586688.600000ns, VSS,
+ 586808.600000ns, VSS,
+ 586808.700000ns, VDD,
+ 586928.700000ns, VDD,
+ 586928.800000ns, VSS,
+ 587289.000000ns, VSS,
+ 587289.100000ns, VDD,
+ 587529.200000ns, VDD,
+ 587529.300000ns, VSS,
+ 587889.500000ns, VSS,
+ 587889.600000ns, VDD,
+ 588249.800000ns, VDD,
+ 588249.900000ns, VSS,
+ 588610.100000ns, VSS,
+ 588610.200000ns, VDD,
+ 589691.000000ns, VDD,
+ 589691.100000ns, VSS,
+ 589931.200000ns, VSS,
+ 589931.300000ns, VDD,
+ 590291.500000ns, VDD,
+ 590291.600000ns, VSS,
+ 590651.800000ns, VSS,
+ 590651.900000ns, VDD,
+ 590892.000000ns, VDD,
+ 590892.100000ns, VSS,
+ 591252.300000ns, VSS,
+ 591252.400000ns, VDD,
+ 591612.600000ns, VDD,
+ 591612.700000ns, VSS,
+ 591732.700000ns, VSS,
+ 591732.800000ns, VDD,
+ 592093.000000ns, VDD,
+ 592093.100000ns, VSS,
+ 592213.100000ns, VSS,
+ 592213.200000ns, VDD,
+ 592453.300000ns, VDD,
+ 592453.400000ns, VSS,
+ 593053.800000ns, VSS,
+ 593053.900000ns, VDD,
+ 593534.200000ns, VDD,
+ 593534.300000ns, VSS,
+ 593654.300000ns, VSS,
+ 593654.400000ns, VDD,
+ 593894.500000ns, VDD,
+ 593894.600000ns, VSS,
+ 594134.700000ns, VSS,
+ 594134.800000ns, VDD,
+ 594855.300000ns, VDD,
+ 594855.400000ns, VSS,
+ 595335.700000ns, VSS,
+ 595335.800000ns, VDD,
+ 595455.800000ns, VDD,
+ 595455.900000ns, VSS,
+ 596536.700000ns, VSS,
+ 596536.800000ns, VDD,
+ 596776.900000ns, VDD,
+ 596777.000000ns, VSS,
+ 597737.700000ns, VSS,
+ 597737.800000ns, VDD,
+ 598098.000000ns, VDD,
+ 598098.100000ns, VSS,
+ 599419.100000ns, VSS,
+ 599419.200000ns, VDD,
+ 599779.400000ns, VDD,
+ 599779.500000ns, VSS,
+ 599899.500000ns, VSS,
+ 599899.600000ns, VDD,
+ 600259.800000ns, VDD,
+ 600259.900000ns, VSS,
+ 600500.000000ns, VSS,
+ 600500.100000ns, VDD,
+ 600620.100000ns, VDD,
+ 600620.200000ns, VSS,
+ 601100.500000ns, VSS,
+ 601100.600000ns, VDD,
+ 601701.000000ns, VDD,
+ 601701.100000ns, VSS,
+ 601941.200000ns, VSS,
+ 601941.300000ns, VDD,
+ 602061.300000ns, VDD,
+ 602061.400000ns, VSS,
+ 602181.400000ns, VSS,
+ 602181.500000ns, VDD,
+ 602902.000000ns, VDD,
+ 602902.100000ns, VSS,
+ 603622.600000ns, VSS,
+ 603622.700000ns, VDD,
+ 604103.000000ns, VDD,
+ 604103.100000ns, VSS,
+ 604583.400000ns, VSS,
+ 604583.500000ns, VDD,
+ 604703.500000ns, VDD,
+ 604703.600000ns, VSS,
+ 605183.900000ns, VSS,
+ 605184.000000ns, VDD,
+ 605424.100000ns, VDD,
+ 605424.200000ns, VSS,
+ 606024.600000ns, VSS,
+ 606024.700000ns, VDD,
+ 606144.700000ns, VDD,
+ 606144.800000ns, VSS,
+ 607345.700000ns, VSS,
+ 607345.800000ns, VDD,
+ 607585.900000ns, VDD,
+ 607586.000000ns, VSS,
+ 608306.500000ns, VSS,
+ 608306.600000ns, VDD,
+ 608426.600000ns, VDD,
+ 608426.700000ns, VSS,
+ 609027.100000ns, VSS,
+ 609027.200000ns, VDD,
+ 609267.300000ns, VDD,
+ 609267.400000ns, VSS,
+ 609627.600000ns, VSS,
+ 609627.700000ns, VDD,
+ 609867.800000ns, VDD,
+ 609867.900000ns, VSS,
+ 610228.100000ns, VSS,
+ 610228.200000ns, VDD,
+ 610348.200000ns, VDD,
+ 610348.300000ns, VSS,
+ 610468.300000ns, VSS,
+ 610468.400000ns, VDD,
+ 610948.700000ns, VDD,
+ 610948.800000ns, VSS,
+ 611068.800000ns, VSS,
+ 611068.900000ns, VDD,
+ 611549.200000ns, VDD,
+ 611549.300000ns, VSS,
+ 612029.600000ns, VSS,
+ 612029.700000ns, VDD,
+ 612149.700000ns, VDD,
+ 612149.800000ns, VSS,
+ 612630.100000ns, VSS,
+ 612630.200000ns, VDD,
+ 614071.300000ns, VDD,
+ 614071.400000ns, VSS,
+ 614551.700000ns, VSS,
+ 614551.800000ns, VDD,
+ 614671.800000ns, VDD,
+ 614671.900000ns, VSS,
+ 614791.900000ns, VSS,
+ 614792.000000ns, VDD,
+ 615032.100000ns, VDD,
+ 615032.200000ns, VSS,
+ 615392.400000ns, VSS,
+ 615392.500000ns, VDD,
+ 615752.700000ns, VDD,
+ 615752.800000ns, VSS,
+ 615992.900000ns, VSS,
+ 615993.000000ns, VDD,
+ 616113.000000ns, VDD,
+ 616113.100000ns, VSS,
+ 616593.400000ns, VSS,
+ 616593.500000ns, VDD,
+ 616833.600000ns, VDD,
+ 616833.700000ns, VSS,
+ 617073.800000ns, VSS,
+ 617073.900000ns, VDD,
+ 617434.100000ns, VDD,
+ 617434.200000ns, VSS,
+ 617674.300000ns, VSS,
+ 617674.400000ns, VDD,
+ 618154.700000ns, VDD,
+ 618154.800000ns, VSS,
+ 618394.900000ns, VSS,
+ 618395.000000ns, VDD,
+ 618995.400000ns, VDD,
+ 618995.500000ns, VSS,
+ 619475.800000ns, VSS,
+ 619475.900000ns, VDD,
+ 619595.900000ns, VDD,
+ 619596.000000ns, VSS,
+ 619956.200000ns, VSS,
+ 619956.300000ns, VDD,
+ 620196.400000ns, VDD,
+ 620196.500000ns, VSS,
+ 620436.600000ns, VSS,
+ 620436.700000ns, VDD,
+ 620676.800000ns, VDD,
+ 620676.900000ns, VSS,
+ 621637.600000ns, VSS,
+ 621637.700000ns, VDD,
+ 621877.800000ns, VDD,
+ 621877.900000ns, VSS,
+ 622118.000000ns, VSS,
+ 622118.100000ns, VDD,
+ 622958.700000ns, VDD,
+ 622958.800000ns, VSS,
+ 623198.900000ns, VSS,
+ 623199.000000ns, VDD,
+ 623319.000000ns, VDD,
+ 623319.100000ns, VSS,
+ 623439.100000ns, VSS,
+ 623439.200000ns, VDD,
+ 623679.300000ns, VDD,
+ 623679.400000ns, VSS,
+ 624880.300000ns, VSS,
+ 624880.400000ns, VDD,
+ 625120.500000ns, VDD,
+ 625120.600000ns, VSS,
+ 625240.600000ns, VSS,
+ 625240.700000ns, VDD,
+ 625600.900000ns, VDD,
+ 625601.000000ns, VSS,
+ 625721.000000ns, VSS,
+ 625721.100000ns, VDD,
+ 626201.400000ns, VDD,
+ 626201.500000ns, VSS,
+ 626321.500000ns, VSS,
+ 626321.600000ns, VDD,
+ 626922.000000ns, VDD,
+ 626922.100000ns, VSS,
+ 627042.100000ns, VSS,
+ 627042.200000ns, VDD,
+ 627882.800000ns, VDD,
+ 627882.900000ns, VSS,
+ 629083.800000ns, VSS,
+ 629083.900000ns, VDD,
+ 629324.000000ns, VDD,
+ 629324.100000ns, VSS,
+ 629684.300000ns, VSS,
+ 629684.400000ns, VDD,
+ 629804.400000ns, VDD,
+ 629804.500000ns, VSS,
+ 630044.600000ns, VSS,
+ 630044.700000ns, VDD,
+ 630164.700000ns, VDD,
+ 630164.800000ns, VSS,
+ 630525.000000ns, VSS,
+ 630525.100000ns, VDD,
+ 631125.500000ns, VDD,
+ 631125.600000ns, VSS,
+ 631245.600000ns, VSS,
+ 631245.700000ns, VDD,
+ 631485.800000ns, VDD,
+ 631485.900000ns, VSS,
+ 632326.500000ns, VSS,
+ 632326.600000ns, VDD,
+ 633287.300000ns, VDD,
+ 633287.400000ns, VSS,
+ 633647.600000ns, VSS,
+ 633647.700000ns, VDD,
+ 633887.800000ns, VDD,
+ 633887.900000ns, VSS,
+ 635088.800000ns, VSS,
+ 635088.900000ns, VDD,
+ 635449.100000ns, VDD,
+ 635449.200000ns, VSS,
+ 635569.200000ns, VSS,
+ 635569.300000ns, VDD,
+ 636169.700000ns, VDD,
+ 636169.800000ns, VSS,
+ 636289.800000ns, VSS,
+ 636289.900000ns, VDD,
+ 636530.000000ns, VDD,
+ 636530.100000ns, VSS,
+ 636770.200000ns, VSS,
+ 636770.300000ns, VDD,
+ 637010.400000ns, VDD,
+ 637010.500000ns, VSS,
+ 637130.500000ns, VSS,
+ 637130.600000ns, VDD,
+ 638932.000000ns, VDD,
+ 638932.100000ns, VSS,
+ 639532.500000ns, VSS,
+ 639532.600000ns, VDD,
+ 639772.700000ns, VDD,
+ 639772.800000ns, VSS,
+ 640133.000000ns, VSS,
+ 640133.100000ns, VDD,
+ 640493.300000ns, VDD,
+ 640493.400000ns, VSS,
+ 640973.700000ns, VSS,
+ 640973.800000ns, VDD,
+ 641454.100000ns, VDD,
+ 641454.200000ns, VSS,
+ 641934.500000ns, VSS,
+ 641934.600000ns, VDD,
+ 642054.600000ns, VDD,
+ 642054.700000ns, VSS,
+ 642414.900000ns, VSS,
+ 642415.000000ns, VDD,
+ 642895.300000ns, VDD,
+ 642895.400000ns, VSS,
+ 643015.400000ns, VSS,
+ 643015.500000ns, VDD,
+ 643615.900000ns, VDD,
+ 643616.000000ns, VSS,
+ 644096.300000ns, VSS,
+ 644096.400000ns, VDD,
+ 644456.600000ns, VDD,
+ 644456.700000ns, VSS,
+ 644576.700000ns, VSS,
+ 644576.800000ns, VDD,
+ 644816.900000ns, VDD,
+ 644817.000000ns, VSS,
+ 644937.000000ns, VSS,
+ 644937.100000ns, VDD,
+ 645537.500000ns, VDD,
+ 645537.600000ns, VSS,
+ 646017.900000ns, VSS,
+ 646018.000000ns, VDD,
+ 646258.100000ns, VDD,
+ 646258.200000ns, VSS,
+ 646498.300000ns, VSS,
+ 646498.400000ns, VDD,
+ 646618.400000ns, VDD,
+ 646618.500000ns, VSS,
+ 646738.500000ns, VSS,
+ 646738.600000ns, VDD,
+ 647339.000000ns, VDD,
+ 647339.100000ns, VSS,
+ 647699.300000ns, VSS,
+ 647699.400000ns, VDD,
+ 648179.700000ns, VDD,
+ 648179.800000ns, VSS,
+ 648419.900000ns, VSS,
+ 648420.000000ns, VDD,
+ 648540.000000ns, VDD,
+ 648540.100000ns, VSS,
+ 649020.400000ns, VSS,
+ 649020.500000ns, VDD,
+ 649861.100000ns, VDD,
+ 649861.200000ns, VSS,
+ 650221.400000ns, VSS,
+ 650221.500000ns, VDD,
+ 650461.600000ns, VDD,
+ 650461.700000ns, VSS,
+ 650581.700000ns, VSS,
+ 650581.800000ns, VDD,
+ 650701.800000ns, VDD,
+ 650701.900000ns, VSS,
+ 651302.300000ns, VSS,
+ 651302.400000ns, VDD,
+ 651542.500000ns, VDD,
+ 651542.600000ns, VSS,
+ 651902.800000ns, VSS,
+ 651902.900000ns, VDD,
+ 652143.000000ns, VDD,
+ 652143.100000ns, VSS,
+ 652503.300000ns, VSS,
+ 652503.400000ns, VDD,
+ 652623.400000ns, VDD,
+ 652623.500000ns, VSS,
+ 652743.500000ns, VSS,
+ 652743.600000ns, VDD,
+ 652983.700000ns, VDD,
+ 652983.800000ns, VSS,
+ 653223.900000ns, VSS,
+ 653224.000000ns, VDD,
+ 654064.600000ns, VDD,
+ 654064.700000ns, VSS,
+ 654424.900000ns, VSS,
+ 654425.000000ns, VDD,
+ 654665.100000ns, VDD,
+ 654665.200000ns, VSS,
+ 655025.400000ns, VSS,
+ 655025.500000ns, VDD,
+ 655145.500000ns, VDD,
+ 655145.600000ns, VSS,
+ 655385.700000ns, VSS,
+ 655385.800000ns, VDD,
+ 656106.300000ns, VDD,
+ 656106.400000ns, VSS,
+ 656586.700000ns, VSS,
+ 656586.800000ns, VDD,
+ 656706.800000ns, VDD,
+ 656706.900000ns, VSS,
+ 657067.100000ns, VSS,
+ 657067.200000ns, VDD,
+ 657307.300000ns, VDD,
+ 657307.400000ns, VSS,
+ 657427.400000ns, VSS,
+ 657427.500000ns, VDD,
+ 657547.500000ns, VDD,
+ 657547.600000ns, VSS,
+ 657667.600000ns, VSS,
+ 657667.700000ns, VDD,
+ 657787.700000ns, VDD,
+ 657787.800000ns, VSS,
+ 657907.800000ns, VSS,
+ 657907.900000ns, VDD,
+ 658148.000000ns, VDD,
+ 658148.100000ns, VSS,
+ 658508.300000ns, VSS,
+ 658508.400000ns, VDD,
+ 658628.400000ns, VDD,
+ 658628.500000ns, VSS,
+ 658748.500000ns, VSS,
+ 658748.600000ns, VDD,
+ 659349.000000ns, VDD,
+ 659349.100000ns, VSS,
+ 659469.100000ns, VSS,
+ 659469.200000ns, VDD,
+ 660189.700000ns, VDD,
+ 660189.800000ns, VSS,
+ 660309.800000ns, VSS,
+ 660309.900000ns, VDD,
+ 660670.100000ns, VDD,
+ 660670.200000ns, VSS,
+ 660790.200000ns, VSS,
+ 660790.300000ns, VDD,
+ 661030.400000ns, VDD,
+ 661030.500000ns, VSS,
+ 662351.500000ns, VSS,
+ 662351.600000ns, VDD,
+ 662591.700000ns, VDD,
+ 662591.800000ns, VSS,
+ 662831.900000ns, VSS,
+ 662832.000000ns, VDD,
+ 663072.100000ns, VDD,
+ 663072.200000ns, VSS,
+ 663192.200000ns, VSS,
+ 663192.300000ns, VDD,
+ 663432.400000ns, VDD,
+ 663432.500000ns, VSS,
+ 664153.000000ns, VSS,
+ 664153.100000ns, VDD,
+ 664513.300000ns, VDD,
+ 664513.400000ns, VSS,
+ 664873.600000ns, VSS,
+ 664873.700000ns, VDD,
+ 665233.900000ns, VDD,
+ 665234.000000ns, VSS,
+ 666194.700000ns, VSS,
+ 666194.800000ns, VDD,
+ 666314.800000ns, VDD,
+ 666314.900000ns, VSS,
+ 666555.000000ns, VSS,
+ 666555.100000ns, VDD,
+ 666795.200000ns, VDD,
+ 666795.300000ns, VSS,
+ 666915.300000ns, VSS,
+ 666915.400000ns, VDD,
+ 667035.400000ns, VDD,
+ 667035.500000ns, VSS,
+ 667515.800000ns, VSS,
+ 667515.900000ns, VDD,
+ 667756.000000ns, VDD,
+ 667756.100000ns, VSS,
+ 667876.100000ns, VSS,
+ 667876.200000ns, VDD,
+ 668236.400000ns, VDD,
+ 668236.500000ns, VSS,
+ 668356.500000ns, VSS,
+ 668356.600000ns, VDD,
+ 668716.800000ns, VDD,
+ 668716.900000ns, VSS,
+ 669437.400000ns, VSS,
+ 669437.500000ns, VDD,
+ 670278.100000ns, VDD,
+ 670278.200000ns, VSS,
+ 670998.700000ns, VSS,
+ 670998.800000ns, VDD,
+ 671599.200000ns, VDD,
+ 671599.300000ns, VSS,
+ 671719.300000ns, VSS,
+ 671719.400000ns, VDD,
+ 672079.600000ns, VDD,
+ 672079.700000ns, VSS,
+ 672199.700000ns, VSS,
+ 672199.800000ns, VDD,
+ 672319.800000ns, VDD,
+ 672319.900000ns, VSS,
+ 672800.200000ns, VSS,
+ 672800.300000ns, VDD,
+ 672920.300000ns, VDD,
+ 672920.400000ns, VSS,
+ 673280.600000ns, VSS,
+ 673280.700000ns, VDD,
+ 673881.100000ns, VDD,
+ 673881.200000ns, VSS,
+ 674361.500000ns, VSS,
+ 674361.600000ns, VDD,
+ 675442.400000ns, VDD,
+ 675442.500000ns, VSS,
+ 675682.600000ns, VSS,
+ 675682.700000ns, VDD,
+ 676042.900000ns, VDD,
+ 676043.000000ns, VSS,
+ 676283.100000ns, VSS,
+ 676283.200000ns, VDD,
+ 676763.500000ns, VDD,
+ 676763.600000ns, VSS,
+ 677364.000000ns, VSS,
+ 677364.100000ns, VDD,
+ 677604.200000ns, VDD,
+ 677604.300000ns, VSS,
+ 677724.300000ns, VSS,
+ 677724.400000ns, VDD,
+ 677964.500000ns, VDD,
+ 677964.600000ns, VSS,
+ 678324.800000ns, VSS,
+ 678324.900000ns, VDD,
+ 678444.900000ns, VDD,
+ 678445.000000ns, VSS,
+ 678565.000000ns, VSS,
+ 678565.100000ns, VDD,
+ 678805.200000ns, VDD,
+ 678805.300000ns, VSS,
+ 679165.500000ns, VSS,
+ 679165.600000ns, VDD,
+ 679285.600000ns, VDD,
+ 679285.700000ns, VSS,
+ 679645.900000ns, VSS,
+ 679646.000000ns, VDD,
+ 680006.200000ns, VDD,
+ 680006.300000ns, VSS,
+ 680486.600000ns, VSS,
+ 680486.700000ns, VDD,
+ 681327.300000ns, VDD,
+ 681327.400000ns, VSS,
+ 681447.400000ns, VSS,
+ 681447.500000ns, VDD,
+ 681807.700000ns, VDD,
+ 681807.800000ns, VSS,
+ 682408.200000ns, VSS,
+ 682408.300000ns, VDD,
+ 682648.400000ns, VDD,
+ 682648.500000ns, VSS,
+ 683008.700000ns, VSS,
+ 683008.800000ns, VDD,
+ 683128.800000ns, VDD,
+ 683128.900000ns, VSS,
+ 683248.900000ns, VSS,
+ 683249.000000ns, VDD,
+ 683609.200000ns, VDD,
+ 683609.300000ns, VSS,
+ 683729.300000ns, VSS,
+ 683729.400000ns, VDD,
+ 684089.600000ns, VDD,
+ 684089.700000ns, VSS,
+ 684209.700000ns, VSS,
+ 684209.800000ns, VDD,
+ 684449.900000ns, VDD,
+ 684450.000000ns, VSS,
+ 684690.100000ns, VSS,
+ 684690.200000ns, VDD,
+ 684810.200000ns, VDD,
+ 684810.300000ns, VSS,
+ 685170.500000ns, VSS,
+ 685170.600000ns, VDD,
+ 686011.200000ns, VDD,
+ 686011.300000ns, VSS,
+ 686131.300000ns, VSS,
+ 686131.400000ns, VDD,
+ 687332.300000ns, VDD,
+ 687332.400000ns, VSS,
+ 687452.400000ns, VSS,
+ 687452.500000ns, VDD,
+ 687932.800000ns, VDD,
+ 687932.900000ns, VSS,
+ 688052.900000ns, VSS,
+ 688053.000000ns, VDD,
+ 688413.200000ns, VDD,
+ 688413.300000ns, VSS,
+ 689013.700000ns, VSS,
+ 689013.800000ns, VDD,
+ 689494.100000ns, VDD,
+ 689494.200000ns, VSS,
+ 689854.400000ns, VSS,
+ 689854.500000ns, VDD,
+ 690214.700000ns, VDD,
+ 690214.800000ns, VSS,
+ 690695.100000ns, VSS,
+ 690695.200000ns, VDD,
+ 691055.400000ns, VDD,
+ 691055.500000ns, VSS,
+ 691415.700000ns, VSS,
+ 691415.800000ns, VDD,
+ 691535.800000ns, VDD,
+ 691535.900000ns, VSS,
+ 691776.000000ns, VSS,
+ 691776.100000ns, VDD,
+ 691896.100000ns, VDD,
+ 691896.200000ns, VSS,
+ 692256.400000ns, VSS,
+ 692256.500000ns, VDD,
+ 692376.500000ns, VDD,
+ 692376.600000ns, VSS,
+ 692856.900000ns, VSS,
+ 692857.000000ns, VDD,
+ 693937.800000ns, VDD,
+ 693937.900000ns, VSS,
+ 694057.900000ns, VSS,
+ 694058.000000ns, VDD,
+ 694418.200000ns, VDD,
+ 694418.300000ns, VSS,
+ 694778.500000ns, VSS,
+ 694778.600000ns, VDD,
+ 694898.600000ns, VDD,
+ 694898.700000ns, VSS,
+ 695619.200000ns, VSS,
+ 695619.300000ns, VDD,
+ 696099.600000ns, VDD,
+ 696099.700000ns, VSS,
+ 696580.000000ns, VSS,
+ 696580.100000ns, VDD,
+ 697060.400000ns, VDD,
+ 697060.500000ns, VSS,
+ 697540.800000ns, VSS,
+ 697540.900000ns, VDD,
+ 697660.900000ns, VDD,
+ 697661.000000ns, VSS,
+ 697901.100000ns, VSS,
+ 697901.200000ns, VDD,
+ 698141.300000ns, VDD,
+ 698141.400000ns, VSS,
+ 698261.400000ns, VSS,
+ 698261.500000ns, VDD,
+ 698621.700000ns, VDD,
+ 698621.800000ns, VSS,
+ 698982.000000ns, VSS,
+ 698982.100000ns, VDD,
+ 699342.300000ns, VDD,
+ 699342.400000ns, VSS,
+ 699702.600000ns, VSS,
+ 699702.700000ns, VDD,
+ 699822.700000ns, VDD,
+ 699822.800000ns, VSS,
+ 699942.800000ns, VSS,
+ 699942.900000ns, VDD,
+ 700183.000000ns, VDD,
+ 700183.100000ns, VSS,
+ 700543.300000ns, VSS,
+ 700543.400000ns, VDD,
+ 700663.400000ns, VDD,
+ 700663.500000ns, VSS,
+ 700783.500000ns, VSS,
+ 700783.600000ns, VDD,
+ 701143.800000ns, VDD,
+ 701143.900000ns, VSS,
+ 701864.400000ns, VSS,
+ 701864.500000ns, VDD,
+ 702464.900000ns, VDD,
+ 702465.000000ns, VSS,
+ 702585.000000ns, VSS,
+ 702585.100000ns, VDD,
+ 703425.700000ns, VDD,
+ 703425.800000ns, VSS,
+ 703906.100000ns, VSS,
+ 703906.200000ns, VDD,
+ 704266.400000ns, VDD,
+ 704266.500000ns, VSS,
+ 704626.700000ns, VSS,
+ 704626.800000ns, VDD,
+ 706308.100000ns, VDD,
+ 706308.200000ns, VSS,
+ 706548.300000ns, VSS,
+ 706548.400000ns, VDD,
+ 707268.900000ns, VDD,
+ 707269.000000ns, VSS,
+ 707629.200000ns, VSS,
+ 707629.300000ns, VDD,
+ 707869.400000ns, VDD,
+ 707869.500000ns, VSS,
+ 708229.700000ns, VSS,
+ 708229.800000ns, VDD,
+ 708830.200000ns, VDD,
+ 708830.300000ns, VSS,
+ 709190.500000ns, VSS,
+ 709190.600000ns, VDD,
+ 709430.700000ns, VDD,
+ 709430.800000ns, VSS,
+ 709791.000000ns, VSS,
+ 709791.100000ns, VDD,
+ 709911.100000ns, VDD,
+ 709911.200000ns, VSS,
+ 710151.300000ns, VSS,
+ 710151.400000ns, VDD,
+ 711592.500000ns, VDD,
+ 711592.600000ns, VSS,
+ 712433.200000ns, VSS,
+ 712433.300000ns, VDD,
+ 713153.800000ns, VDD,
+ 713153.900000ns, VSS,
+ 713273.900000ns, VSS,
+ 713274.000000ns, VDD,
+ 713754.300000ns, VDD,
+ 713754.400000ns, VSS,
+ 714234.700000ns, VSS,
+ 714234.800000ns, VDD,
+ 715195.500000ns, VDD,
+ 715195.600000ns, VSS,
+ 715555.800000ns, VSS,
+ 715555.900000ns, VDD,
+ 716036.200000ns, VDD,
+ 716036.300000ns, VSS,
+ 716276.400000ns, VSS,
+ 716276.500000ns, VDD,
+ 716636.700000ns, VDD,
+ 716636.800000ns, VSS,
+ 716756.800000ns, VSS,
+ 716756.900000ns, VDD,
+ 717117.100000ns, VDD,
+ 717117.200000ns, VSS,
+ 717837.700000ns, VSS,
+ 717837.800000ns, VDD,
+ 718198.000000ns, VDD,
+ 718198.100000ns, VSS,
+ 718558.300000ns, VSS,
+ 718558.400000ns, VDD,
+ 718678.400000ns, VDD,
+ 718678.500000ns, VSS,
+ 719158.800000ns, VSS,
+ 719158.900000ns, VDD,
+ 719999.500000ns, VDD,
+ 719999.600000ns, VSS,
+ 720720.100000ns, VSS,
+ 720720.200000ns, VDD,
+ 720960.300000ns, VDD,
+ 720960.400000ns, VSS,
+ 721200.500000ns, VSS,
+ 721200.600000ns, VDD,
+ 721440.700000ns, VDD,
+ 721440.800000ns, VSS,
+ 721560.800000ns, VSS,
+ 721560.900000ns, VDD,
+ 721801.000000ns, VDD,
+ 721801.100000ns, VSS,
+ 722041.200000ns, VSS,
+ 722041.300000ns, VDD,
+ 722521.600000ns, VDD,
+ 722521.700000ns, VSS,
+ 722641.700000ns, VSS,
+ 722641.800000ns, VDD,
+ 722881.900000ns, VDD,
+ 722882.000000ns, VSS,
+ 723362.300000ns, VSS,
+ 723362.400000ns, VDD,
+ 723482.400000ns, VDD,
+ 723482.500000ns, VSS,
+ 724203.000000ns, VSS,
+ 724203.100000ns, VDD,
+ 724443.200000ns, VDD,
+ 724443.300000ns, VSS,
+ 724563.300000ns, VSS,
+ 724563.400000ns, VDD,
+ 724803.500000ns, VDD,
+ 724803.600000ns, VSS,
+ 725283.900000ns, VSS,
+ 725284.000000ns, VDD,
+ 725524.100000ns, VDD,
+ 725524.200000ns, VSS,
+ 725884.400000ns, VSS,
+ 725884.500000ns, VDD,
+ 726124.600000ns, VDD,
+ 726124.700000ns, VSS,
+ 727205.500000ns, VSS,
+ 727205.600000ns, VDD,
+ 727325.600000ns, VDD,
+ 727325.700000ns, VSS,
+ 727806.000000ns, VSS,
+ 727806.100000ns, VDD,
+ 727926.100000ns, VDD,
+ 727926.200000ns, VSS,
+ 728286.400000ns, VSS,
+ 728286.500000ns, VDD,
+ 728526.600000ns, VDD,
+ 728526.700000ns, VSS,
+ 728886.900000ns, VSS,
+ 728887.000000ns, VDD,
+ 729007.000000ns, VDD,
+ 729007.100000ns, VSS,
+ 729127.100000ns, VSS,
+ 729127.200000ns, VDD,
+ 729367.300000ns, VDD,
+ 729367.400000ns, VSS,
+ 729607.500000ns, VSS,
+ 729607.600000ns, VDD,
+ 729727.600000ns, VDD,
+ 729727.700000ns, VSS,
+ 729967.800000ns, VSS,
+ 729967.900000ns, VDD,
+ 731409.000000ns, VDD,
+ 731409.100000ns, VSS,
+ 731529.100000ns, VSS,
+ 731529.200000ns, VDD,
+ 732489.900000ns, VDD,
+ 732490.000000ns, VSS,
+ 732970.300000ns, VSS,
+ 732970.400000ns, VDD,
+ 733090.400000ns, VDD,
+ 733090.500000ns, VSS,
+ 733811.000000ns, VSS,
+ 733811.100000ns, VDD,
+ 734411.500000ns, VDD,
+ 734411.600000ns, VSS,
+ 736092.900000ns, VSS,
+ 736093.000000ns, VDD,
+ 736333.100000ns, VDD,
+ 736333.200000ns, VSS,
+ 736693.400000ns, VSS,
+ 736693.500000ns, VDD,
+ 736933.600000ns, VDD,
+ 736933.700000ns, VSS,
+ 737293.900000ns, VSS,
+ 737294.000000ns, VDD,
+ 737414.000000ns, VDD,
+ 737414.100000ns, VSS,
+ 737654.200000ns, VSS,
+ 737654.300000ns, VDD,
+ 738615.000000ns, VDD,
+ 738615.100000ns, VSS,
+ 738855.200000ns, VSS,
+ 738855.300000ns, VDD,
+ 738975.300000ns, VDD,
+ 738975.400000ns, VSS,
+ 739335.600000ns, VSS,
+ 739335.700000ns, VDD,
+ 739575.800000ns, VDD,
+ 739575.900000ns, VSS,
+ 739695.900000ns, VSS,
+ 739696.000000ns, VDD,
+ 739936.100000ns, VDD,
+ 739936.200000ns, VSS,
+ 740776.800000ns, VSS,
+ 740776.900000ns, VDD,
+ 740896.900000ns, VDD,
+ 740897.000000ns, VSS,
+ 741257.200000ns, VSS,
+ 741257.300000ns, VDD,
+ 741617.500000ns, VDD,
+ 741617.600000ns, VSS,
+ 741977.800000ns, VSS,
+ 741977.900000ns, VDD,
+ 742458.200000ns, VDD,
+ 742458.300000ns, VSS,
+ 742578.300000ns, VSS,
+ 742578.400000ns, VDD,
+ 743298.900000ns, VDD,
+ 743299.000000ns, VSS,
+ 743419.000000ns, VSS,
+ 743419.100000ns, VDD,
+ 744019.500000ns, VDD,
+ 744019.600000ns, VSS,
+ 744620.000000ns, VSS,
+ 744620.100000ns, VDD,
+ 744740.100000ns, VDD,
+ 744740.200000ns, VSS,
+ 745460.700000ns, VSS,
+ 745460.800000ns, VDD,
+ 745700.900000ns, VDD,
+ 745701.000000ns, VSS,
+ 746061.200000ns, VSS,
+ 746061.300000ns, VDD,
+ 746541.600000ns, VDD,
+ 746541.700000ns, VSS,
+ 746781.800000ns, VSS,
+ 746781.900000ns, VDD,
+ 747382.300000ns, VDD,
+ 747382.400000ns, VSS,
+ 747742.600000ns, VSS,
+ 747742.700000ns, VDD,
+ 747982.800000ns, VDD,
+ 747982.900000ns, VSS,
+ 748343.100000ns, VSS,
+ 748343.200000ns, VDD,
+ 748463.200000ns, VDD,
+ 748463.300000ns, VSS,
+ 748583.300000ns, VSS,
+ 748583.400000ns, VDD,
+ 748703.400000ns, VDD,
+ 748703.500000ns, VSS,
+ 748943.600000ns, VSS,
+ 748943.700000ns, VDD,
+ 749784.300000ns, VDD,
+ 749784.400000ns, VSS,
+ 750264.700000ns, VSS,
+ 750264.800000ns, VDD,
+ 750384.800000ns, VDD,
+ 750384.900000ns, VSS,
+ 750625.000000ns, VSS,
+ 750625.100000ns, VDD,
+ 750865.200000ns, VDD,
+ 750865.300000ns, VSS,
+ 750985.300000ns, VSS,
+ 750985.400000ns, VDD,
+ 751225.500000ns, VDD,
+ 751225.600000ns, VSS,
+ 751585.800000ns, VSS,
+ 751585.900000ns, VDD,
+ 752546.600000ns, VDD,
+ 752546.700000ns, VSS,
+ 752906.900000ns, VSS,
+ 752907.000000ns, VDD,
+ 753387.300000ns, VDD,
+ 753387.400000ns, VSS,
+ 754468.200000ns, VSS,
+ 754468.300000ns, VDD,
+ 754588.300000ns, VDD,
+ 754588.400000ns, VSS,
+ 754828.500000ns, VSS,
+ 754828.600000ns, VDD,
+ 755188.800000ns, VDD,
+ 755188.900000ns, VSS,
+ 755549.100000ns, VSS,
+ 755549.200000ns, VDD,
+ 756029.500000ns, VDD,
+ 756029.600000ns, VSS,
+ 756149.600000ns, VSS,
+ 756149.700000ns, VDD,
+ 756389.800000ns, VDD,
+ 756389.900000ns, VSS,
+ 756509.900000ns, VSS,
+ 756510.000000ns, VDD,
+ 756750.100000ns, VDD,
+ 756750.200000ns, VSS,
+ 757710.900000ns, VSS,
+ 757711.000000ns, VDD,
+ 758191.300000ns, VDD,
+ 758191.400000ns, VSS,
+ 758791.800000ns, VSS,
+ 758791.900000ns, VDD,
+ 759032.000000ns, VDD,
+ 759032.100000ns, VSS,
+ 759632.500000ns, VSS,
+ 759632.600000ns, VDD,
+ 759992.800000ns, VDD,
+ 759992.900000ns, VSS,
+ 760112.900000ns, VSS,
+ 760113.000000ns, VDD,
+ 760473.200000ns, VDD,
+ 760473.300000ns, VSS,
+ 760593.300000ns, VSS,
+ 760593.400000ns, VDD,
+ 760833.500000ns, VDD,
+ 760833.600000ns, VSS,
+ 760953.600000ns, VSS,
+ 760953.700000ns, VDD,
+ 761434.000000ns, VDD,
+ 761434.100000ns, VSS,
+ 761554.100000ns, VSS,
+ 761554.200000ns, VDD,
+ 761794.300000ns, VDD,
+ 761794.400000ns, VSS,
+ 762514.900000ns, VSS,
+ 762515.000000ns, VDD,
+ 762755.100000ns, VDD,
+ 762755.200000ns, VSS,
+ 763115.400000ns, VSS,
+ 763115.500000ns, VDD,
+ 763355.600000ns, VDD,
+ 763355.700000ns, VSS,
+ 763956.100000ns, VSS,
+ 763956.200000ns, VDD,
+ 764556.600000ns, VDD,
+ 764556.700000ns, VSS,
+ 765397.300000ns, VSS,
+ 765397.400000ns, VDD,
+ 765877.700000ns, VDD,
+ 765877.800000ns, VSS,
+ 765997.800000ns, VSS,
+ 765997.900000ns, VDD,
+ 766238.000000ns, VDD,
+ 766238.100000ns, VSS,
+ 766598.300000ns, VSS,
+ 766598.400000ns, VDD,
+ 766718.400000ns, VDD,
+ 766718.500000ns, VSS,
+ 768039.500000ns, VSS,
+ 768039.600000ns, VDD,
+ 769000.300000ns, VDD,
+ 769000.400000ns, VSS,
+ 769240.500000ns, VSS,
+ 769240.600000ns, VDD,
+ 769600.800000ns, VDD,
+ 769600.900000ns, VSS,
+ 769720.900000ns, VSS,
+ 769721.000000ns, VDD,
+ 770201.300000ns, VDD,
+ 770201.400000ns, VSS,
+ 770801.800000ns, VSS,
+ 770801.900000ns, VDD,
+ 771282.200000ns, VDD,
+ 771282.300000ns, VSS,
+ 772243.000000ns, VSS,
+ 772243.100000ns, VDD,
+ 772483.200000ns, VDD,
+ 772483.300000ns, VSS,
+ 772603.300000ns, VSS,
+ 772603.400000ns, VDD,
+ 772723.400000ns, VDD,
+ 772723.500000ns, VSS,
+ 772963.600000ns, VSS,
+ 772963.700000ns, VDD,
+ 773203.800000ns, VDD,
+ 773203.900000ns, VSS,
+ 773564.100000ns, VSS,
+ 773564.200000ns, VDD,
+ 774284.700000ns, VDD,
+ 774284.800000ns, VSS,
+ 774645.000000ns, VSS,
+ 774645.100000ns, VDD,
+ 774885.200000ns, VDD,
+ 774885.300000ns, VSS,
+ 775245.500000ns, VSS,
+ 775245.600000ns, VDD,
+ 775725.900000ns, VDD,
+ 775726.000000ns, VSS,
+ 776206.300000ns, VSS,
+ 776206.400000ns, VDD,
+ 776686.700000ns, VDD,
+ 776686.800000ns, VSS,
+ 776806.800000ns, VSS,
+ 776806.900000ns, VDD,
+ 777047.000000ns, VDD,
+ 777047.100000ns, VSS,
+ 777647.500000ns, VSS,
+ 777647.600000ns, VDD,
+ 777887.700000ns, VDD,
+ 777887.800000ns, VSS,
+ 778007.800000ns, VSS,
+ 778007.900000ns, VDD,
+ 778248.000000ns, VDD,
+ 778248.100000ns, VSS,
+ 778368.100000ns, VSS,
+ 778368.200000ns, VDD,
+ 778728.400000ns, VDD,
+ 778728.500000ns, VSS,
+ 778968.600000ns, VSS,
+ 778968.700000ns, VDD,
+ 779088.700000ns, VDD,
+ 779088.800000ns, VSS,
+ 779569.100000ns, VSS,
+ 779569.200000ns, VDD,
+ 779809.300000ns, VDD,
+ 779809.400000ns, VSS,
+ 780049.500000ns, VSS,
+ 780049.600000ns, VDD,
+ 780169.600000ns, VDD,
+ 780169.700000ns, VSS,
+ 780289.700000ns, VSS,
+ 780289.800000ns, VDD,
+ 780529.900000ns, VDD,
+ 780530.000000ns, VSS,
+ 781250.500000ns, VSS,
+ 781250.600000ns, VDD,
+ 781610.800000ns, VDD,
+ 781610.900000ns, VSS,
+ 782091.200000ns, VSS,
+ 782091.300000ns, VDD,
+ 782811.800000ns, VDD,
+ 782811.900000ns, VSS,
+ 782931.900000ns, VSS,
+ 782932.000000ns, VDD,
+ 783652.500000ns, VDD,
+ 783652.600000ns, VSS,
+ 783772.600000ns, VSS,
+ 783772.700000ns, VDD,
+ 784132.900000ns, VDD,
+ 784133.000000ns, VSS,
+ 784253.000000ns, VSS,
+ 784253.100000ns, VDD,
+ 784493.200000ns, VDD,
+ 784493.300000ns, VSS,
+ 784733.400000ns, VSS,
+ 784733.500000ns, VDD,
+ 784973.600000ns, VDD,
+ 784973.700000ns, VSS,
+ 785574.100000ns, VSS,
+ 785574.200000ns, VDD,
+ 785814.300000ns, VDD,
+ 785814.400000ns, VSS,
+ 786174.600000ns, VSS,
+ 786174.700000ns, VDD,
+ 787255.500000ns, VDD,
+ 787255.600000ns, VSS,
+ 787375.600000ns, VSS,
+ 787375.700000ns, VDD,
+ 787615.800000ns, VDD,
+ 787615.900000ns, VSS,
+ 787856.000000ns, VSS,
+ 787856.100000ns, VDD,
+ 788096.200000ns, VDD,
+ 788096.300000ns, VSS,
+ 788216.300000ns, VSS,
+ 788216.400000ns, VDD,
+ 788336.400000ns, VDD,
+ 788336.500000ns, VSS,
+ 788696.700000ns, VSS,
+ 788696.800000ns, VDD,
+ 790017.800000ns, VDD,
+ 790017.900000ns, VSS,
+ 790618.300000ns, VSS,
+ 790618.400000ns, VDD,
+ 790738.400000ns, VDD,
+ 790738.500000ns, VSS,
+ 791459.000000ns, VSS,
+ 791459.100000ns, VDD,
+ 791819.300000ns, VDD,
+ 791819.400000ns, VSS,
+ 792539.900000ns, VSS,
+ 792540.000000ns, VDD,
+ 793620.800000ns, VDD,
+ 793620.900000ns, VSS,
+ 793740.900000ns, VSS,
+ 793741.000000ns, VDD,
+ 793861.000000ns, VDD,
+ 793861.100000ns, VSS,
+ 793981.100000ns, VSS,
+ 793981.200000ns, VDD,
+ 794221.300000ns, VDD,
+ 794221.400000ns, VSS,
+ 794581.600000ns, VSS,
+ 794581.700000ns, VDD,
+ 794821.800000ns, VDD,
+ 794821.900000ns, VSS,
+ 795182.100000ns, VSS,
+ 795182.200000ns, VDD,
+ 795422.300000ns, VDD,
+ 795422.400000ns, VSS,
+ 795542.400000ns, VSS,
+ 795542.500000ns, VDD,
+ 795902.700000ns, VDD,
+ 795902.800000ns, VSS,
+ 796022.800000ns, VSS,
+ 796022.900000ns, VDD,
+ 796142.900000ns, VDD,
+ 796143.000000ns, VSS,
+ 796263.000000ns, VSS,
+ 796263.100000ns, VDD,
+ 796623.300000ns, VDD,
+ 796623.400000ns, VSS,
+ 796983.600000ns, VSS,
+ 796983.700000ns, VDD,
+ 797223.800000ns, VDD,
+ 797223.900000ns, VSS,
+ 797464.000000ns, VSS,
+ 797464.100000ns, VDD,
+ 797584.100000ns, VDD,
+ 797584.200000ns, VSS,
+ 798064.500000ns, VSS,
+ 798064.600000ns, VDD,
+ 798665.000000ns, VDD,
+ 798665.100000ns, VSS,
+ 798905.200000ns, VSS,
+ 798905.300000ns, VDD,
+ 799385.600000ns, VDD,
+ 799385.700000ns, VSS,
+ 799625.800000ns, VSS,
+ 799625.900000ns, VDD,
+ 800226.300000ns, VDD,
+ 800226.400000ns, VSS,
+ 800346.400000ns, VSS,
+ 800346.500000ns, VDD,
+ 800586.600000ns, VDD,
+ 800586.700000ns, VSS,
+ 800826.800000ns, VSS,
+ 800826.900000ns, VDD,
+ 801307.200000ns, VDD,
+ 801307.300000ns, VSS,
+ 801427.300000ns, VSS,
+ 801427.400000ns, VDD,
+ 801787.600000ns, VDD,
+ 801787.700000ns, VSS,
+ 801907.700000ns, VSS,
+ 801907.800000ns, VDD,
+ 802508.200000ns, VDD,
+ 802508.300000ns, VSS,
+ 802628.300000ns, VSS,
+ 802628.400000ns, VDD,
+ 802868.500000ns, VDD,
+ 802868.600000ns, VSS,
+ 803228.800000ns, VSS,
+ 803228.900000ns, VDD,
+ 804429.800000ns, VDD,
+ 804429.900000ns, VSS,
+ 804549.900000ns, VSS,
+ 804550.000000ns, VDD,
+ 805630.800000ns, VDD,
+ 805630.900000ns, VSS,
+ 805871.000000ns, VSS,
+ 805871.100000ns, VDD,
+ 806951.900000ns, VDD,
+ 806952.000000ns, VSS,
+ 807072.000000ns, VSS,
+ 807072.100000ns, VDD,
+ 807432.300000ns, VDD,
+ 807432.400000ns, VSS,
+ 808032.800000ns, VSS,
+ 808032.900000ns, VDD,
+ 808993.600000ns, VDD,
+ 808993.700000ns, VSS,
+ 809233.800000ns, VSS,
+ 809233.900000ns, VDD,
+ 809714.200000ns, VDD,
+ 809714.300000ns, VSS,
+ 809834.300000ns, VSS,
+ 809834.400000ns, VDD,
+ 810314.700000ns, VDD,
+ 810314.800000ns, VSS,
+ 811035.300000ns, VSS,
+ 811035.400000ns, VDD,
+ 811635.800000ns, VDD,
+ 811635.900000ns, VSS,
+ 812116.200000ns, VSS,
+ 812116.300000ns, VDD,
+ 813197.100000ns, VDD,
+ 813197.200000ns, VSS,
+ 814518.200000ns, VSS,
+ 814518.300000ns, VDD,
+ 814638.300000ns, VDD,
+ 814638.400000ns, VSS,
+ 814878.500000ns, VSS,
+ 814878.600000ns, VDD,
+ 815479.000000ns, VDD,
+ 815479.100000ns, VSS,
+ 815599.100000ns, VSS,
+ 815599.200000ns, VDD,
+ 816199.600000ns, VDD,
+ 816199.700000ns, VSS,
+ 816319.700000ns, VSS,
+ 816319.800000ns, VDD,
+ 816800.100000ns, VDD,
+ 816800.200000ns, VSS,
+ 817160.400000ns, VSS,
+ 817160.500000ns, VDD,
+ 817280.500000ns, VDD,
+ 817280.600000ns, VSS,
+ 817640.800000ns, VSS,
+ 817640.900000ns, VDD,
+ 817881.000000ns, VDD,
+ 817881.100000ns, VSS,
+ 818721.700000ns, VSS,
+ 818721.800000ns, VDD,
+ 818841.800000ns, VDD,
+ 818841.900000ns, VSS,
+ 819202.100000ns, VSS,
+ 819202.200000ns, VDD,
+ 819562.400000ns, VDD,
+ 819562.500000ns, VSS,
+ 819682.500000ns, VSS,
+ 819682.600000ns, VDD,
+ 820042.800000ns, VDD,
+ 820042.900000ns, VSS,
+ 820283.000000ns, VSS,
+ 820283.100000ns, VDD,
+ 820523.200000ns, VDD,
+ 820523.300000ns, VSS,
+ 820643.300000ns, VSS,
+ 820643.400000ns, VDD,
+ 821844.300000ns, VDD,
+ 821844.400000ns, VSS,
+ 822204.600000ns, VSS,
+ 822204.700000ns, VDD,
+ 823285.500000ns, VDD,
+ 823285.600000ns, VSS,
+ 823886.000000ns, VSS,
+ 823886.100000ns, VDD,
+ 825447.300000ns, VDD,
+ 825447.400000ns, VSS,
+ 825927.700000ns, VSS,
+ 825927.800000ns, VDD,
+ 826528.200000ns, VDD,
+ 826528.300000ns, VSS,
+ 826888.500000ns, VSS,
+ 826888.600000ns, VDD,
+ 827248.800000ns, VDD,
+ 827248.900000ns, VSS,
+ 827368.900000ns, VSS,
+ 827369.000000ns, VDD,
+ 827609.100000ns, VDD,
+ 827609.200000ns, VSS,
+ 827849.300000ns, VSS,
+ 827849.400000ns, VDD,
+ 827969.400000ns, VDD,
+ 827969.500000ns, VSS,
+ 828089.500000ns, VSS,
+ 828089.600000ns, VDD,
+ 828569.900000ns, VDD,
+ 828570.000000ns, VSS,
+ 828810.100000ns, VSS,
+ 828810.200000ns, VDD,
+ 829170.400000ns, VDD,
+ 829170.500000ns, VSS,
+ 829770.900000ns, VSS,
+ 829771.000000ns, VDD,
+ 829891.000000ns, VDD,
+ 829891.100000ns, VSS,
+ 830131.200000ns, VSS,
+ 830131.300000ns, VDD,
+ 830251.300000ns, VDD,
+ 830251.400000ns, VSS,
+ 830371.400000ns, VSS,
+ 830371.500000ns, VDD,
+ 830611.600000ns, VDD,
+ 830611.700000ns, VSS,
+ 830971.900000ns, VSS,
+ 830972.000000ns, VDD,
+ 831092.000000ns, VDD,
+ 831092.100000ns, VSS,
+ 831212.100000ns, VSS,
+ 831212.200000ns, VDD,
+ 831332.200000ns, VDD,
+ 831332.300000ns, VSS,
+ 831812.600000ns, VSS,
+ 831812.700000ns, VDD,
+ 833133.700000ns, VDD,
+ 833133.800000ns, VSS,
+ 833494.000000ns, VSS,
+ 833494.100000ns, VDD,
+ 833854.300000ns, VDD,
+ 833854.400000ns, VSS,
+ 834815.100000ns, VSS,
+ 834815.200000ns, VDD,
+ 835415.600000ns, VDD,
+ 835415.700000ns, VSS,
+ 836376.400000ns, VSS,
+ 836376.500000ns, VDD,
+ 837097.000000ns, VDD,
+ 837097.100000ns, VSS,
+ 837457.300000ns, VSS,
+ 837457.400000ns, VDD,
+ 837697.500000ns, VDD,
+ 837697.600000ns, VSS,
+ 837937.700000ns, VSS,
+ 837937.800000ns, VDD,
+ 838298.000000ns, VDD,
+ 838298.100000ns, VSS,
+ 838418.100000ns, VSS,
+ 838418.200000ns, VDD,
+ 838778.400000ns, VDD,
+ 838778.500000ns, VSS,
+ 839739.200000ns, VSS,
+ 839739.300000ns, VDD,
+ 839979.400000ns, VDD,
+ 839979.500000ns, VSS,
+ 840099.500000ns, VSS,
+ 840099.600000ns, VDD,
+ 840579.900000ns, VDD,
+ 840580.000000ns, VSS,
+ 840940.200000ns, VSS,
+ 840940.300000ns, VDD,
+ 841540.700000ns, VDD,
+ 841540.800000ns, VSS,
+ 842261.300000ns, VSS,
+ 842261.400000ns, VDD,
+ 842381.400000ns, VDD,
+ 842381.500000ns, VSS,
+ 842981.900000ns, VSS,
+ 842982.000000ns, VDD,
+ 843222.100000ns, VDD,
+ 843222.200000ns, VSS,
+ 843342.200000ns, VSS,
+ 843342.300000ns, VDD,
+ 843462.300000ns, VDD,
+ 843462.400000ns, VSS,
+ 843582.400000ns, VSS,
+ 843582.500000ns, VDD,
+ 844062.800000ns, VDD,
+ 844062.900000ns, VSS,
+ 844423.100000ns, VSS,
+ 844423.200000ns, VDD,
+ 844663.300000ns, VDD,
+ 844663.400000ns, VSS,
+ 845744.200000ns, VSS,
+ 845744.300000ns, VDD,
+ 846104.500000ns, VDD,
+ 846104.600000ns, VSS,
+ 846464.800000ns, VSS,
+ 846464.900000ns, VDD,
+ 847425.600000ns, VDD,
+ 847425.700000ns, VSS,
+ 848146.200000ns, VSS,
+ 848146.300000ns, VDD,
+ 848626.600000ns, VDD,
+ 848626.700000ns, VSS,
+ 848746.700000ns, VSS,
+ 848746.800000ns, VDD,
+ 849107.000000ns, VDD,
+ 849107.100000ns, VSS,
+ 849227.100000ns, VSS,
+ 849227.200000ns, VDD,
+ 849587.400000ns, VDD,
+ 849587.500000ns, VSS,
+ 849707.500000ns, VSS,
+ 849707.600000ns, VDD,
+ 849947.700000ns, VDD,
+ 849947.800000ns, VSS,
+ 850067.800000ns, VSS,
+ 850067.900000ns, VDD,
+ 850308.000000ns, VDD,
+ 850308.100000ns, VSS,
+ 850548.200000ns, VSS,
+ 850548.300000ns, VDD,
+ 850668.300000ns, VDD,
+ 850668.400000ns, VSS,
+ 850788.400000ns, VSS,
+ 850788.500000ns, VDD,
+ 851268.800000ns, VDD,
+ 851268.900000ns, VSS,
+ 851629.100000ns, VSS,
+ 851629.200000ns, VDD,
+ 851989.400000ns, VDD,
+ 851989.500000ns, VSS,
+ 852589.900000ns, VSS,
+ 852590.000000ns, VDD,
+ 852830.100000ns, VDD,
+ 852830.200000ns, VSS,
+ 853190.400000ns, VSS,
+ 853190.500000ns, VDD,
+ 853790.900000ns, VDD,
+ 853791.000000ns, VSS,
+ 854031.100000ns, VSS,
+ 854031.200000ns, VDD,
+ 854511.500000ns, VDD,
+ 854511.600000ns, VSS,
+ 854631.600000ns, VSS,
+ 854631.700000ns, VDD,
+ 854991.900000ns, VDD,
+ 854992.000000ns, VSS,
+ 855112.000000ns, VSS,
+ 855112.100000ns, VDD,
+ 855592.400000ns, VDD,
+ 855592.500000ns, VSS,
+ 855712.500000ns, VSS,
+ 855712.600000ns, VDD,
+ 855952.700000ns, VDD,
+ 855952.800000ns, VSS,
+ 856072.800000ns, VSS,
+ 856072.900000ns, VDD,
+ 856673.300000ns, VDD,
+ 856673.400000ns, VSS,
+ 857153.700000ns, VSS,
+ 857153.800000ns, VDD,
+ 857273.800000ns, VDD,
+ 857273.900000ns, VSS,
+ 857754.200000ns, VSS,
+ 857754.300000ns, VDD,
+ 858234.600000ns, VDD,
+ 858234.700000ns, VSS,
+ 858354.700000ns, VSS,
+ 858354.800000ns, VDD,
+ 858594.900000ns, VDD,
+ 858595.000000ns, VSS,
+ 858835.100000ns, VSS,
+ 858835.200000ns, VDD,
+ 859075.300000ns, VDD,
+ 859075.400000ns, VSS,
+ 860156.200000ns, VSS,
+ 860156.300000ns, VDD,
+ 860276.300000ns, VDD,
+ 860276.400000ns, VSS,
+ 860396.400000ns, VSS,
+ 860396.500000ns, VDD,
+ 860996.900000ns, VDD,
+ 860997.000000ns, VSS,
+ 861117.000000ns, VSS,
+ 861117.100000ns, VDD,
+ 861717.500000ns, VDD,
+ 861717.600000ns, VSS,
+ 861837.600000ns, VSS,
+ 861837.700000ns, VDD,
+ 862438.100000ns, VDD,
+ 862438.200000ns, VSS,
+ 863639.100000ns, VSS,
+ 863639.200000ns, VDD,
+ 864119.500000ns, VDD,
+ 864119.600000ns, VSS,
+ 864359.700000ns, VSS,
+ 864359.800000ns, VDD,
+ 865440.600000ns, VDD,
+ 865440.700000ns, VSS,
+ 865800.900000ns, VSS,
+ 865801.000000ns, VDD,
+ 866641.600000ns, VDD,
+ 866641.700000ns, VSS,
+ 866881.800000ns, VSS,
+ 866881.900000ns, VDD,
+ 867001.900000ns, VDD,
+ 867002.000000ns, VSS,
+ 867362.200000ns, VSS,
+ 867362.300000ns, VDD,
+ 867602.400000ns, VDD,
+ 867602.500000ns, VSS,
+ 868443.100000ns, VSS,
+ 868443.200000ns, VDD,
+ 868683.300000ns, VDD,
+ 868683.400000ns, VSS,
+ 869043.600000ns, VSS,
+ 869043.700000ns, VDD,
+ 869644.100000ns, VDD,
+ 869644.200000ns, VSS,
+ 870004.400000ns, VSS,
+ 870004.500000ns, VDD,
+ 870244.600000ns, VDD,
+ 870244.700000ns, VSS,
+ 870364.700000ns, VSS,
+ 870364.800000ns, VDD,
+ 871085.300000ns, VDD,
+ 871085.400000ns, VSS,
+ 871445.600000ns, VSS,
+ 871445.700000ns, VDD,
+ 871805.900000ns, VDD,
+ 871806.000000ns, VSS,
+ 872646.600000ns, VSS,
+ 872646.700000ns, VDD,
+ 872886.800000ns, VDD,
+ 872886.900000ns, VSS,
+ 873247.100000ns, VSS,
+ 873247.200000ns, VDD,
+ 873487.300000ns, VDD,
+ 873487.400000ns, VSS,
+ 874087.800000ns, VSS,
+ 874087.900000ns, VDD,
+ 874568.200000ns, VDD,
+ 874568.300000ns, VSS,
+ 874808.400000ns, VSS,
+ 874808.500000ns, VDD,
+ 875288.800000ns, VDD,
+ 875288.900000ns, VSS,
+ 875649.100000ns, VSS,
+ 875649.200000ns, VDD,
+ 877210.400000ns, VDD,
+ 877210.500000ns, VSS,
+ 877690.800000ns, VSS,
+ 877690.900000ns, VDD,
+ 877810.900000ns, VDD,
+ 877811.000000ns, VSS,
+ 878171.200000ns, VSS,
+ 878171.300000ns, VDD,
+ 878291.300000ns, VDD,
+ 878291.400000ns, VSS,
+ 878651.600000ns, VSS,
+ 878651.700000ns, VDD,
+ 878891.800000ns, VDD,
+ 878891.900000ns, VSS,
+ 879011.900000ns, VSS,
+ 879012.000000ns, VDD,
+ 879372.200000ns, VDD,
+ 879372.300000ns, VSS,
+ 879492.300000ns, VSS,
+ 879492.400000ns, VDD,
+ 879612.400000ns, VDD,
+ 879612.500000ns, VSS,
+ 879732.500000ns, VSS,
+ 879732.600000ns, VDD,
+ 882735.000000ns, VDD,
+ 882735.100000ns, VSS,
+ 883335.500000ns, VSS,
+ 883335.600000ns, VDD,
+ 883815.900000ns, VDD,
+ 883816.000000ns, VSS,
+ 884176.200000ns, VSS,
+ 884176.300000ns, VDD,
+ 884416.400000ns, VDD,
+ 884416.500000ns, VSS,
+ 884896.800000ns, VSS,
+ 884896.900000ns, VDD,
+ 885137.000000ns, VDD,
+ 885137.100000ns, VSS,
+ 885977.700000ns, VSS,
+ 885977.800000ns, VDD,
+ 886578.200000ns, VDD,
+ 886578.300000ns, VSS,
+ 886698.300000ns, VSS,
+ 886698.400000ns, VDD,
+ 887779.200000ns, VDD,
+ 887779.300000ns, VSS,
+ 888379.700000ns, VSS,
+ 888379.800000ns, VDD,
+ 888619.900000ns, VDD,
+ 888620.000000ns, VSS,
+ 888740.000000ns, VSS,
+ 888740.100000ns, VDD,
+ 888980.200000ns, VDD,
+ 888980.300000ns, VSS,
+ 889820.900000ns, VSS,
+ 889821.000000ns, VDD,
+ 890061.100000ns, VDD,
+ 890061.200000ns, VSS,
+ 890181.200000ns, VSS,
+ 890181.300000ns, VDD,
+ 890301.300000ns, VDD,
+ 890301.400000ns, VSS,
+ 890661.600000ns, VSS,
+ 890661.700000ns, VDD,
+ 890781.700000ns, VDD,
+ 890781.800000ns, VSS,
+ 891382.200000ns, VSS,
+ 891382.300000ns, VDD,
+ 892102.800000ns, VDD,
+ 892102.900000ns, VSS,
+ 892343.000000ns, VSS,
+ 892343.100000ns, VDD,
+ 892823.400000ns, VDD,
+ 892823.500000ns, VSS,
+ 892943.500000ns, VSS,
+ 892943.600000ns, VDD,
+ 893183.700000ns, VDD,
+ 893183.800000ns, VSS,
+ 894504.800000ns, VSS,
+ 894504.900000ns, VDD,
+ 894985.200000ns, VDD,
+ 894985.300000ns, VSS,
+ 895825.900000ns, VSS,
+ 895826.000000ns, VDD,
+ 896066.100000ns, VDD,
+ 896066.200000ns, VSS,
+ 896546.500000ns, VSS,
+ 896546.600000ns, VDD,
+ 896786.700000ns, VDD,
+ 896786.800000ns, VSS,
+ 897026.900000ns, VSS,
+ 897027.000000ns, VDD,
+ 897267.100000ns, VDD,
+ 897267.200000ns, VSS,
+ 898227.900000ns, VSS,
+ 898228.000000ns, VDD,
+ 898468.100000ns, VDD,
+ 898468.200000ns, VSS,
+ 898588.200000ns, VSS,
+ 898588.300000ns, VDD,
+ 899068.600000ns, VDD,
+ 899068.700000ns, VSS,
+ 899188.700000ns, VSS,
+ 899188.800000ns, VDD,
+ 900389.700000ns, VDD,
+ 900389.800000ns, VSS,
+ 900870.100000ns, VSS,
+ 900870.200000ns, VDD,
+ 901230.400000ns, VDD,
+ 901230.500000ns, VSS,
+ 901350.500000ns, VSS,
+ 901350.600000ns, VDD,
+ 902071.100000ns, VDD,
+ 902071.200000ns, VSS,
+ 902311.300000ns, VSS,
+ 902311.400000ns, VDD,
+ 902551.500000ns, VDD,
+ 902551.600000ns, VSS,
+ 903512.300000ns, VSS,
+ 903512.400000ns, VDD,
+ 904833.400000ns, VDD,
+ 904833.500000ns, VSS,
+ 904953.500000ns, VSS,
+ 904953.600000ns, VDD,
+ 905433.900000ns, VDD,
+ 905434.000000ns, VSS,
+ 905794.200000ns, VSS,
+ 905794.300000ns, VDD,
+ 905914.300000ns, VDD,
+ 905914.400000ns, VSS,
+ 906514.800000ns, VSS,
+ 906514.900000ns, VDD,
+ 906995.200000ns, VDD,
+ 906995.300000ns, VSS,
+ 907355.500000ns, VSS,
+ 907355.600000ns, VDD,
+ 907595.700000ns, VDD,
+ 907595.800000ns, VSS,
+ 907715.800000ns, VSS,
+ 907715.900000ns, VDD,
+ 907956.000000ns, VDD,
+ 907956.100000ns, VSS,
+ 908316.300000ns, VSS,
+ 908316.400000ns, VDD,
+ 908436.400000ns, VDD,
+ 908436.500000ns, VSS,
+ 908556.500000ns, VSS,
+ 908556.600000ns, VDD,
+ 908796.700000ns, VDD,
+ 908796.800000ns, VSS,
+ 908916.800000ns, VSS,
+ 908916.900000ns, VDD,
+ 909157.000000ns, VDD,
+ 909157.100000ns, VSS,
+ 909517.300000ns, VSS,
+ 909517.400000ns, VDD,
+ 909637.400000ns, VDD,
+ 909637.500000ns, VSS,
+ 910598.200000ns, VSS,
+ 910598.300000ns, VDD,
+ 910838.400000ns, VDD,
+ 910838.500000ns, VSS,
+ 910958.500000ns, VSS,
+ 910958.600000ns, VDD,
+ 911198.700000ns, VDD,
+ 911198.800000ns, VSS,
+ 911559.000000ns, VSS,
+ 911559.100000ns, VDD,
+ 911799.200000ns, VDD,
+ 911799.300000ns, VSS,
+ 913000.200000ns, VSS,
+ 913000.300000ns, VDD,
+ 913240.400000ns, VDD,
+ 913240.500000ns, VSS,
+ 913600.700000ns, VSS,
+ 913600.800000ns, VDD,
+ 913720.800000ns, VDD,
+ 913720.900000ns, VSS,
+ 913840.900000ns, VSS,
+ 913841.000000ns, VDD,
+ 914441.400000ns, VDD,
+ 914441.500000ns, VSS,
+ 914801.700000ns, VSS,
+ 914801.800000ns, VDD,
+ 915162.000000ns, VDD,
+ 915162.100000ns, VSS,
+ 915642.400000ns, VSS,
+ 915642.500000ns, VDD,
+ 916122.800000ns, VDD,
+ 916122.900000ns, VSS,
+ 916242.900000ns, VSS,
+ 916243.000000ns, VDD,
+ 917083.600000ns, VDD,
+ 917083.700000ns, VSS,
+ 917443.900000ns, VSS,
+ 917444.000000ns, VDD,
+ 917564.000000ns, VDD,
+ 917564.100000ns, VSS,
+ 917924.300000ns, VSS,
+ 917924.400000ns, VDD,
+ 918164.500000ns, VDD,
+ 918164.600000ns, VSS,
+ 918284.600000ns, VSS,
+ 918284.700000ns, VDD,
+ 918524.800000ns, VDD,
+ 918524.900000ns, VSS,
+ 918765.000000ns, VSS,
+ 918765.100000ns, VDD,
+ 919005.200000ns, VDD,
+ 919005.300000ns, VSS,
+ 919245.400000ns, VSS,
+ 919245.500000ns, VDD,
+ 919845.900000ns, VDD,
+ 919846.000000ns, VSS,
+ 921287.100000ns, VSS,
+ 921287.200000ns, VDD,
+ 921407.200000ns, VDD,
+ 921407.300000ns, VSS,
+ 921767.500000ns, VSS,
+ 921767.600000ns, VDD,
+ 922127.800000ns, VDD,
+ 922127.900000ns, VSS,
+ 922368.000000ns, VSS,
+ 922368.100000ns, VDD,
+ 922608.200000ns, VDD,
+ 922608.300000ns, VSS,
+ 923448.900000ns, VSS,
+ 923449.000000ns, VDD,
+ 923929.300000ns, VDD,
+ 923929.400000ns, VSS,
+ 924770.000000ns, VSS,
+ 924770.100000ns, VDD,
+ 925010.200000ns, VDD,
+ 925010.300000ns, VSS,
+ 925370.500000ns, VSS,
+ 925370.600000ns, VDD,
+ 925971.000000ns, VDD,
+ 925971.100000ns, VSS,
+ 926091.100000ns, VSS,
+ 926091.200000ns, VDD,
+ 926691.600000ns, VDD,
+ 926691.700000ns, VSS,
+ 926811.700000ns, VSS,
+ 926811.800000ns, VDD,
+ 927051.900000ns, VDD,
+ 927052.000000ns, VSS,
+ 927412.200000ns, VSS,
+ 927412.300000ns, VDD,
+ 927532.300000ns, VDD,
+ 927532.400000ns, VSS,
+ 928012.700000ns, VSS,
+ 928012.800000ns, VDD,
+ 928132.800000ns, VDD,
+ 928132.900000ns, VSS,
+ 928252.900000ns, VSS,
+ 928253.000000ns, VDD,
+ 928733.300000ns, VDD,
+ 928733.400000ns, VSS,
+ 928973.500000ns, VSS,
+ 928973.600000ns, VDD,
+ 929213.700000ns, VDD,
+ 929213.800000ns, VSS,
+ 929333.800000ns, VSS,
+ 929333.900000ns, VDD,
+ 929453.900000ns, VDD,
+ 929454.000000ns, VSS,
+ 929934.300000ns, VSS,
+ 929934.400000ns, VDD,
+ 930294.600000ns, VDD,
+ 930294.700000ns, VSS,
+ 930775.000000ns, VSS,
+ 930775.100000ns, VDD,
+ 931255.400000ns, VDD,
+ 931255.500000ns, VSS,
+ 931495.600000ns, VSS,
+ 931495.700000ns, VDD,
+ 932816.700000ns, VDD,
+ 932816.800000ns, VSS,
+ 933537.300000ns, VSS,
+ 933537.400000ns, VDD,
+ 934498.100000ns, VDD,
+ 934498.200000ns, VSS,
+ 934618.200000ns, VSS,
+ 934618.300000ns, VDD,
+ 935338.800000ns, VDD,
+ 935338.900000ns, VSS,
+ 935819.200000ns, VSS,
+ 935819.300000ns, VDD,
+ 935939.300000ns, VDD,
+ 935939.400000ns, VSS,
+ 936539.800000ns, VSS,
+ 936539.900000ns, VDD,
+ 937020.200000ns, VDD,
+ 937020.300000ns, VSS,
+ 937140.300000ns, VSS,
+ 937140.400000ns, VDD,
+ 937500.600000ns, VDD,
+ 937500.700000ns, VSS,
+ 938341.300000ns, VSS,
+ 938341.400000ns, VDD,
+ 938461.400000ns, VDD,
+ 938461.500000ns, VSS,
+ 938941.800000ns, VSS,
+ 938941.900000ns, VDD,
+ 939422.200000ns, VDD,
+ 939422.300000ns, VSS,
+ 939542.300000ns, VSS,
+ 939542.400000ns, VDD,
+ 940022.700000ns, VDD,
+ 940022.800000ns, VSS,
+ 940262.900000ns, VSS,
+ 940263.000000ns, VDD,
+ 940503.100000ns, VDD,
+ 940503.200000ns, VSS,
+ 941223.700000ns, VSS,
+ 941223.800000ns, VDD,
+ 941704.100000ns, VDD,
+ 941704.200000ns, VSS,
+ 941824.200000ns, VSS,
+ 941824.300000ns, VDD,
+ 942664.900000ns, VDD,
+ 942665.000000ns, VSS,
+ 943745.800000ns, VSS,
+ 943745.900000ns, VDD,
+ 944106.100000ns, VDD,
+ 944106.200000ns, VSS,
+ 944226.200000ns, VSS,
+ 944226.300000ns, VDD,
+ 944586.500000ns, VDD,
+ 944586.600000ns, VSS,
+ 944706.600000ns, VSS,
+ 944706.700000ns, VDD,
+ 944946.800000ns, VDD,
+ 944946.900000ns, VSS,
+ 945187.000000ns, VSS,
+ 945187.100000ns, VDD,
+ 945667.400000ns, VDD,
+ 945667.500000ns, VSS,
+ 945787.500000ns, VSS,
+ 945787.600000ns, VDD,
+ 946628.200000ns, VDD,
+ 946628.300000ns, VSS,
+ 947228.700000ns, VSS,
+ 947228.800000ns, VDD,
+ 947468.900000ns, VDD,
+ 947469.000000ns, VSS,
+ 947589.000000ns, VSS,
+ 947589.100000ns, VDD,
+ 947829.200000ns, VDD,
+ 947829.300000ns, VSS,
+ 948189.500000ns, VSS,
+ 948189.600000ns, VDD,
+ 948309.600000ns, VDD,
+ 948309.700000ns, VSS,
+ 948790.000000ns, VSS,
+ 948790.100000ns, VDD,
+ 949390.500000ns, VDD,
+ 949390.600000ns, VSS,
+ 950591.500000ns, VSS,
+ 950591.600000ns, VDD,
+ 950711.600000ns, VDD,
+ 950711.700000ns, VSS,
+ 950951.800000ns, VSS,
+ 950951.900000ns, VDD,
+ 952032.700000ns, VDD,
+ 952032.800000ns, VSS,
+ 953353.800000ns, VSS,
+ 953353.900000ns, VDD,
+ 954074.400000ns, VDD,
+ 954074.500000ns, VSS,
+ 954314.600000ns, VSS,
+ 954314.700000ns, VDD,
+ 954434.700000ns, VDD,
+ 954434.800000ns, VSS,
+ 954795.000000ns, VSS,
+ 954795.100000ns, VDD,
+ 954915.100000ns, VDD,
+ 954915.200000ns, VSS,
+ 955035.200000ns, VSS,
+ 955035.300000ns, VDD,
+ 955515.600000ns, VDD,
+ 955515.700000ns, VSS,
+ 956116.100000ns, VSS,
+ 956116.200000ns, VDD,
+ 956596.500000ns, VDD,
+ 956596.600000ns, VSS,
+ 956716.600000ns, VSS,
+ 956716.700000ns, VDD,
+ 957076.900000ns, VDD,
+ 957077.000000ns, VSS,
+ 957197.000000ns, VSS,
+ 957197.100000ns, VDD,
+ 957917.600000ns, VDD,
+ 957917.700000ns, VSS,
+ 958037.700000ns, VSS,
+ 958037.800000ns, VDD,
+ 958398.000000ns, VDD,
+ 958398.100000ns, VSS,
+ 958518.100000ns, VSS,
+ 958518.200000ns, VDD,
+ 958998.500000ns, VDD,
+ 958998.600000ns, VSS,
+ 959238.700000ns, VSS,
+ 959238.800000ns, VDD,
+ 959719.100000ns, VDD,
+ 959719.200000ns, VSS,
+ 960079.400000ns, VSS,
+ 960079.500000ns, VDD,
+ 960559.800000ns, VDD,
+ 960559.900000ns, VSS,
+ 960800.000000ns, VSS,
+ 960800.100000ns, VDD,
+ 960920.100000ns, VDD,
+ 960920.200000ns, VSS,
+ 961280.400000ns, VSS,
+ 961280.500000ns, VDD,
+ 961400.500000ns, VDD,
+ 961400.600000ns, VSS,
+ 961880.900000ns, VSS,
+ 961881.000000ns, VDD,
+ 962121.100000ns, VDD,
+ 962121.200000ns, VSS,
+ 962481.400000ns, VSS,
+ 962481.500000ns, VDD,
+ 962601.500000ns, VDD,
+ 962601.600000ns, VSS,
+ 962721.600000ns, VSS,
+ 962721.700000ns, VDD,
+ 963802.500000ns, VDD,
+ 963802.600000ns, VSS,
+ 964523.100000ns, VSS,
+ 964523.200000ns, VDD,
+ 964763.300000ns, VDD,
+ 964763.400000ns, VSS,
+ 965003.500000ns, VSS,
+ 965003.600000ns, VDD,
+ 965243.700000ns, VDD,
+ 965243.800000ns, VSS,
+ 965483.900000ns, VSS,
+ 965484.000000ns, VDD,
+ 966564.800000ns, VDD,
+ 966564.900000ns, VSS,
+ 966684.900000ns, VSS,
+ 966685.000000ns, VDD,
+ 966805.000000ns, VDD,
+ 966805.100000ns, VSS,
+ 967045.200000ns, VSS,
+ 967045.300000ns, VDD,
+ 967645.700000ns, VDD,
+ 967645.800000ns, VSS,
+ 967765.800000ns, VSS,
+ 967765.900000ns, VDD,
+ 968366.300000ns, VDD,
+ 968366.400000ns, VSS,
+ 968606.500000ns, VSS,
+ 968606.600000ns, VDD,
+ 968966.800000ns, VDD,
+ 968966.900000ns, VSS,
+ 969207.000000ns, VSS,
+ 969207.100000ns, VDD,
+ 969327.100000ns, VDD,
+ 969327.200000ns, VSS,
+ 969687.400000ns, VSS,
+ 969687.500000ns, VDD,
+ 969927.600000ns, VDD,
+ 969927.700000ns, VSS,
+ 970648.200000ns, VSS,
+ 970648.300000ns, VDD,
+ 970768.300000ns, VDD,
+ 970768.400000ns, VSS,
+ 971128.600000ns, VSS,
+ 971128.700000ns, VDD,
+ 971248.700000ns, VDD,
+ 971248.800000ns, VSS,
+ 971368.800000ns, VSS,
+ 971368.900000ns, VDD,
+ 971729.100000ns, VDD,
+ 971729.200000ns, VSS,
+ 971969.300000ns, VSS,
+ 971969.400000ns, VDD,
+ 972089.400000ns, VDD,
+ 972089.500000ns, VSS,
+ 972209.500000ns, VSS,
+ 972209.600000ns, VDD,
+ 972449.700000ns, VDD,
+ 972449.800000ns, VSS,
+ 972810.000000ns, VSS,
+ 972810.100000ns, VDD,
+ 973650.700000ns, VDD,
+ 973650.800000ns, VSS,
+ 974251.200000ns, VSS,
+ 974251.300000ns, VDD,
+ 974611.500000ns, VDD,
+ 974611.600000ns, VSS,
+ 976292.900000ns, VSS,
+ 976293.000000ns, VDD,
+ 976773.300000ns, VDD,
+ 976773.400000ns, VSS,
+ 977133.600000ns, VSS,
+ 977133.700000ns, VDD,
+ 977373.800000ns, VDD,
+ 977373.900000ns, VSS,
+ 977493.900000ns, VSS,
+ 977494.000000ns, VDD,
+ 977854.200000ns, VDD,
+ 977854.300000ns, VSS,
+ 978694.900000ns, VSS,
+ 978695.000000ns, VDD,
+ 979415.500000ns, VDD,
+ 979415.600000ns, VSS,
+ 979775.800000ns, VSS,
+ 979775.900000ns, VDD,
+ 979895.900000ns, VDD,
+ 979896.000000ns, VSS,
+ 980256.200000ns, VSS,
+ 980256.300000ns, VDD,
+ 980376.300000ns, VDD,
+ 980376.400000ns, VSS,
+ 980736.600000ns, VSS,
+ 980736.700000ns, VDD,
+ 983258.700000ns, VDD,
+ 983258.800000ns, VSS,
+ 983619.000000ns, VSS,
+ 983619.100000ns, VDD,
+ 984099.400000ns, VDD,
+ 984099.500000ns, VSS,
+ 984820.000000ns, VSS,
+ 984820.100000ns, VDD,
+ 985780.800000ns, VDD,
+ 985780.900000ns, VSS,
+ 985900.900000ns, VSS,
+ 985901.000000ns, VDD,
+ 986381.300000ns, VDD,
+ 986381.400000ns, VSS,
+ 986501.400000ns, VSS,
+ 986501.500000ns, VDD,
+ 986981.800000ns, VDD,
+ 986981.900000ns, VSS,
+ 987222.000000ns, VSS,
+ 987222.100000ns, VDD,
+ 987702.400000ns, VDD,
+ 987702.500000ns, VSS,
+ 989143.600000ns, VSS,
+ 989143.700000ns, VDD,
+ 989624.000000ns, VDD,
+ 989624.100000ns, VSS,
+ 989744.100000ns, VSS,
+ 989744.200000ns, VDD,
+ 989984.300000ns, VDD,
+ 989984.400000ns, VSS,
+ 990104.400000ns, VSS,
+ 990104.500000ns, VDD,
+ 990825.000000ns, VDD,
+ 990825.100000ns, VSS,
+ 991425.500000ns, VSS,
+ 991425.600000ns, VDD,
+ 991665.700000ns, VDD,
+ 991665.800000ns, VSS,
+ 992146.100000ns, VSS,
+ 992146.200000ns, VDD,
+ 992386.300000ns, VDD,
+ 992386.400000ns, VSS,
+ 992746.600000ns, VSS,
+ 992746.700000ns, VDD,
+ 993347.100000ns, VDD,
+ 993347.200000ns, VSS,
+ 993707.400000ns, VSS,
+ 993707.500000ns, VDD,
+ 993827.500000ns, VDD,
+ 993827.600000ns, VSS,
+ 993947.600000ns, VSS,
+ 993947.700000ns, VDD,
+ 994067.700000ns, VDD,
+ 994067.800000ns, VSS,
+ 994668.200000ns, VSS,
+ 994668.300000ns, VDD,
+ 994908.400000ns, VDD,
+ 994908.500000ns, VSS,
+ 995749.100000ns, VSS,
+ 995749.200000ns, VDD,
+ 996349.600000ns, VDD,
+ 996349.700000ns, VSS,
+ 996589.800000ns, VSS,
+ 996589.900000ns, VDD,
+ 996709.900000ns, VDD,
+ 996710.000000ns, VSS,
+ 997190.300000ns, VSS,
+ 997190.400000ns, VDD,
+ 997430.500000ns, VDD,
+ 997430.600000ns, VSS,
+ 997550.600000ns, VSS,
+ 997550.700000ns, VDD,
+ 997670.700000ns, VDD,
+ 997670.800000ns, VSS,
+ 997790.800000ns, VSS,
+ 997790.900000ns, VDD,
+ 998151.100000ns, VDD,
+ 998151.200000ns, VSS,
+ 998271.200000ns, VSS,
+ 998271.300000ns, VDD,
+ 998511.400000ns, VDD,
+ 998511.500000ns, VSS,
+ 999832.500000ns, VSS,
+ 999832.600000ns, VDD,
+ 1000312.900000ns, VDD,
+ 1000313.000000ns, VSS,
+ 1000913.400000ns, VSS,
+ 1000913.500000ns, VDD,
+ 1001153.600000ns, VDD,
+ 1001153.700000ns, VSS,
+ 1001273.700000ns, VSS,
+ 1001273.800000ns, VDD,
+ 1001754.100000ns, VDD,
+ 1001754.200000ns, VSS,
+ 1002114.400000ns, VSS,
+ 1002114.500000ns, VDD,
+ 1002714.900000ns, VDD,
+ 1002715.000000ns, VSS,
+ 1002955.100000ns, VSS,
+ 1002955.200000ns, VDD,
+ 1003435.500000ns, VDD,
+ 1003435.600000ns, VSS,
+ 1003555.600000ns, VSS,
+ 1003555.700000ns, VDD,
+ 1004036.000000ns, VDD,
+ 1004036.100000ns, VSS,
+ 1004756.600000ns, VSS,
+ 1004756.700000ns, VDD,
+ 1005237.000000ns, VDD,
+ 1005237.100000ns, VSS,
+ 1005357.100000ns, VSS,
+ 1005357.200000ns, VDD,
+ 1005597.300000ns, VDD,
+ 1005597.400000ns, VSS,
+ 1005957.600000ns, VSS,
+ 1005957.700000ns, VDD,
+ 1006678.200000ns, VDD,
+ 1006678.300000ns, VSS,
+ 1007038.500000ns, VSS,
+ 1007038.600000ns, VDD,
+ 1007278.700000ns, VDD,
+ 1007278.800000ns, VSS,
+ 1007879.200000ns, VSS,
+ 1007879.300000ns, VDD,
+ 1007999.300000ns, VDD,
+ 1007999.400000ns, VSS,
+ 1008479.700000ns, VSS,
+ 1008479.800000ns, VDD,
+ 1009200.300000ns, VDD,
+ 1009200.400000ns, VSS,
+ 1009680.700000ns, VSS,
+ 1009680.800000ns, VDD,
+ 1010401.300000ns, VDD,
+ 1010401.400000ns, VSS,
+ 1010641.500000ns, VSS,
+ 1010641.600000ns, VDD,
+ 1011121.900000ns, VDD,
+ 1011122.000000ns, VSS,
+ 1011242.000000ns, VSS,
+ 1011242.100000ns, VDD,
+ 1011722.400000ns, VDD,
+ 1011722.500000ns, VSS,
+ 1012202.800000ns, VSS,
+ 1012202.900000ns, VDD,
+ 1012322.900000ns, VDD,
+ 1012323.000000ns, VSS,
+ 1012803.300000ns, VSS,
+ 1012803.400000ns, VDD,
+ 1012923.400000ns, VDD,
+ 1012923.500000ns, VSS,
+ 1013283.700000ns, VSS,
+ 1013283.800000ns, VDD,
+ 1013403.800000ns, VDD,
+ 1013403.900000ns, VSS,
+ 1013523.900000ns, VSS,
+ 1013524.000000ns, VDD,
+ 1013644.000000ns, VDD,
+ 1013644.100000ns, VSS,
+ 1013764.100000ns, VSS,
+ 1013764.200000ns, VDD,
+ 1014484.700000ns, VDD,
+ 1014484.800000ns, VSS,
+ 1014845.000000ns, VSS,
+ 1014845.100000ns, VDD,
+ 1015085.200000ns, VDD,
+ 1015085.300000ns, VSS,
+ 1015325.400000ns, VSS,
+ 1015325.500000ns, VDD,
+ 1015565.600000ns, VDD,
+ 1015565.700000ns, VSS,
+ 1016166.100000ns, VSS,
+ 1016166.200000ns, VDD,
+ 1016286.200000ns, VDD,
+ 1016286.300000ns, VSS,
+ 1016526.400000ns, VSS,
+ 1016526.500000ns, VDD,
+ 1016766.600000ns, VDD,
+ 1016766.700000ns, VSS,
+ 1016886.700000ns, VSS,
+ 1016886.800000ns, VDD,
+ 1017126.900000ns, VDD,
+ 1017127.000000ns, VSS,
+ 1017247.000000ns, VSS,
+ 1017247.100000ns, VDD,
+ 1018207.800000ns, VDD,
+ 1018207.900000ns, VSS,
+ 1018448.000000ns, VSS,
+ 1018448.100000ns, VDD,
+ 1018808.300000ns, VDD,
+ 1018808.400000ns, VSS,
+ 1018928.400000ns, VSS,
+ 1018928.500000ns, VDD,
+ 1019408.800000ns, VDD,
+ 1019408.900000ns, VSS,
+ 1019528.900000ns, VSS,
+ 1019529.000000ns, VDD,
+ 1019769.100000ns, VDD,
+ 1019769.200000ns, VSS,
+ 1020129.400000ns, VSS,
+ 1020129.500000ns, VDD,
+ 1020369.600000ns, VDD,
+ 1020369.700000ns, VSS,
+ 1021450.500000ns, VSS,
+ 1021450.600000ns, VDD,
+ 1021690.700000ns, VDD,
+ 1021690.800000ns, VSS,
+ 1022171.100000ns, VSS,
+ 1022171.200000ns, VDD,
+ 1022291.200000ns, VDD,
+ 1022291.300000ns, VSS,
+ 1022411.300000ns, VSS,
+ 1022411.400000ns, VDD,
+ 1022531.400000ns, VDD,
+ 1022531.500000ns, VSS,
+ 1022651.500000ns, VSS,
+ 1022651.600000ns, VDD,
+ 1023011.800000ns, VDD,
+ 1023011.900000ns, VSS,
+ 1023372.100000ns, VSS,
+ 1023372.200000ns, VDD,
+ 1023612.300000ns, VDD,
+ 1023612.400000ns, VSS,
+ 1023852.500000ns, VSS,
+ 1023852.600000ns, VDD,
+ 1024092.700000ns, VDD,
+ 1024092.800000ns, VSS,
+ 1024332.900000ns, VSS,
+ 1024333.000000ns, VDD,
+ 1025293.700000ns, VDD,
+ 1025293.800000ns, VSS,
+ 1026254.500000ns, VSS,
+ 1026254.600000ns, VDD,
+ 1026975.100000ns, VDD,
+ 1026975.200000ns, VSS,
+ 1027215.300000ns, VSS,
+ 1027215.400000ns, VDD,
+ 1027335.400000ns, VDD,
+ 1027335.500000ns, VSS,
+ 1027695.700000ns, VSS,
+ 1027695.800000ns, VDD,
+ 1027935.900000ns, VDD,
+ 1027936.000000ns, VSS,
+ 1028056.000000ns, VSS,
+ 1028056.100000ns, VDD,
+ 1028296.200000ns, VDD,
+ 1028296.300000ns, VSS,
+ 1028656.500000ns, VSS,
+ 1028656.600000ns, VDD,
+ 1028896.700000ns, VDD,
+ 1028896.800000ns, VSS,
+ 1029136.900000ns, VSS,
+ 1029137.000000ns, VDD,
+ 1029857.500000ns, VDD,
+ 1029857.600000ns, VSS,
+ 1029977.600000ns, VSS,
+ 1029977.700000ns, VDD,
+ 1030698.200000ns, VDD,
+ 1030698.300000ns, VSS,
+ 1030818.300000ns, VSS,
+ 1030818.400000ns, VDD,
+ 1031178.600000ns, VDD,
+ 1031178.700000ns, VSS,
+ 1032259.500000ns, VSS,
+ 1032259.600000ns, VDD,
+ 1032499.700000ns, VDD,
+ 1032499.800000ns, VSS,
+ 1032619.800000ns, VSS,
+ 1032619.900000ns, VDD,
+ 1032860.000000ns, VDD,
+ 1032860.100000ns, VSS,
+ 1032980.100000ns, VSS,
+ 1032980.200000ns, VDD,
+ 1033700.700000ns, VDD,
+ 1033700.800000ns, VSS,
+ 1034061.000000ns, VSS,
+ 1034061.100000ns, VDD,
+ 1034421.300000ns, VDD,
+ 1034421.400000ns, VSS,
+ 1034541.400000ns, VSS,
+ 1034541.500000ns, VDD,
+ 1034781.600000ns, VDD,
+ 1034781.700000ns, VSS,
+ 1035021.800000ns, VSS,
+ 1035021.900000ns, VDD,
+ 1035141.900000ns, VDD,
+ 1035142.000000ns, VSS,
+ 1035262.000000ns, VSS,
+ 1035262.100000ns, VDD,
+ 1035862.500000ns, VDD,
+ 1035862.600000ns, VSS,
+ 1036102.700000ns, VSS,
+ 1036102.800000ns, VDD,
+ 1036222.800000ns, VDD,
+ 1036222.900000ns, VSS,
+ 1036583.100000ns, VSS,
+ 1036583.200000ns, VDD,
+ 1036823.300000ns, VDD,
+ 1036823.400000ns, VSS,
+ 1037183.600000ns, VSS,
+ 1037183.700000ns, VDD,
+ 1037664.000000ns, VDD,
+ 1037664.100000ns, VSS,
+ 1038504.700000ns, VSS,
+ 1038504.800000ns, VDD,
+ 1038744.900000ns, VDD,
+ 1038745.000000ns, VSS,
+ 1039225.300000ns, VSS,
+ 1039225.400000ns, VDD,
+ 1039345.400000ns, VDD,
+ 1039345.500000ns, VSS,
+ 1040546.400000ns, VSS,
+ 1040546.500000ns, VDD,
+ 1040786.600000ns, VDD,
+ 1040786.700000ns, VSS,
+ 1041026.800000ns, VSS,
+ 1041026.900000ns, VDD,
+ 1041267.000000ns, VDD,
+ 1041267.100000ns, VSS,
+ 1042227.800000ns, VSS,
+ 1042227.900000ns, VDD,
+ 1042828.300000ns, VDD,
+ 1042828.400000ns, VSS,
+ 1043188.600000ns, VSS,
+ 1043188.700000ns, VDD,
+ 1043428.800000ns, VDD,
+ 1043428.900000ns, VSS,
+ 1043909.200000ns, VSS,
+ 1043909.300000ns, VDD,
+ 1044389.600000ns, VDD,
+ 1044389.700000ns, VSS,
+ 1044509.700000ns, VSS,
+ 1044509.800000ns, VDD,
+ 1045470.500000ns, VDD,
+ 1045470.600000ns, VSS,
+ 1045830.800000ns, VSS,
+ 1045830.900000ns, VDD,
+ 1046191.100000ns, VDD,
+ 1046191.200000ns, VSS,
+ 1047031.800000ns, VSS,
+ 1047031.900000ns, VDD,
+ 1047392.100000ns, VDD,
+ 1047392.200000ns, VSS,
+ 1047512.200000ns, VSS,
+ 1047512.300000ns, VDD,
+ 1047752.400000ns, VDD,
+ 1047752.500000ns, VSS,
+ 1047872.500000ns, VSS,
+ 1047872.600000ns, VDD,
+ 1048232.800000ns, VDD,
+ 1048232.900000ns, VSS,
+ 1048593.100000ns, VSS,
+ 1048593.200000ns, VDD,
+ 1049193.600000ns, VDD,
+ 1049193.700000ns, VSS,
+ 1049433.800000ns, VSS,
+ 1049433.900000ns, VDD,
+ 1049674.000000ns, VDD,
+ 1049674.100000ns, VSS,
+ 1050034.300000ns, VSS,
+ 1050034.400000ns, VDD,
+ 1050154.400000ns, VDD,
+ 1050154.500000ns, VSS,
+ 1050754.900000ns, VSS,
+ 1050755.000000ns, VDD,
+ 1051115.200000ns, VDD,
+ 1051115.300000ns, VSS,
+ 1051235.300000ns, VSS,
+ 1051235.400000ns, VDD,
+ 1051955.900000ns, VDD,
+ 1051956.000000ns, VSS,
+ 1052556.400000ns, VSS,
+ 1052556.500000ns, VDD,
+ 1052796.600000ns, VDD,
+ 1052796.700000ns, VSS,
+ 1052916.700000ns, VSS,
+ 1052916.800000ns, VDD,
+ 1053277.000000ns, VDD,
+ 1053277.100000ns, VSS,
+ 1053757.400000ns, VSS,
+ 1053757.500000ns, VDD,
+ 1054598.100000ns, VDD,
+ 1054598.200000ns, VSS,
+ 1054958.400000ns, VSS,
+ 1054958.500000ns, VDD,
+ 1055198.600000ns, VDD,
+ 1055198.700000ns, VSS,
+ 1055438.800000ns, VSS,
+ 1055438.900000ns, VDD,
+ 1055799.100000ns, VDD,
+ 1055799.200000ns, VSS,
+ 1056399.600000ns, VSS,
+ 1056399.700000ns, VDD,
+ 1056519.700000ns, VDD,
+ 1056519.800000ns, VSS,
+ 1056880.000000ns, VSS,
+ 1056880.100000ns, VDD,
+ 1057000.100000ns, VDD,
+ 1057000.200000ns, VSS,
+ 1057840.800000ns, VSS,
+ 1057840.900000ns, VDD,
+ 1060242.800000ns, VDD,
+ 1060242.900000ns, VSS,
+ 1060362.900000ns, VSS,
+ 1060363.000000ns, VDD,
+ 1060723.200000ns, VDD,
+ 1060723.300000ns, VSS,
+ 1061083.500000ns, VSS,
+ 1061083.600000ns, VDD,
+ 1061443.800000ns, VDD,
+ 1061443.900000ns, VSS,
+ 1062164.400000ns, VSS,
+ 1062164.500000ns, VDD,
+ 1062284.500000ns, VDD,
+ 1062284.600000ns, VSS,
+ 1062644.800000ns, VSS,
+ 1062644.900000ns, VDD,
+ 1062764.900000ns, VDD,
+ 1062765.000000ns, VSS,
+ 1063005.100000ns, VSS,
+ 1063005.200000ns, VDD,
+ 1063125.200000ns, VDD,
+ 1063125.300000ns, VSS,
+ 1063485.500000ns, VSS,
+ 1063485.600000ns, VDD,
+ 1063725.700000ns, VDD,
+ 1063725.800000ns, VSS,
+ 1063845.800000ns, VSS,
+ 1063845.900000ns, VDD,
+ 1064326.200000ns, VDD,
+ 1064326.300000ns, VSS,
+ 1064806.600000ns, VSS,
+ 1064806.700000ns, VDD,
+ 1065046.800000ns, VDD,
+ 1065046.900000ns, VSS,
+ 1065287.000000ns, VSS,
+ 1065287.100000ns, VDD,
+ 1065527.200000ns, VDD,
+ 1065527.300000ns, VSS,
+ 1067088.500000ns, VSS,
+ 1067088.600000ns, VDD,
+ 1067328.700000ns, VDD,
+ 1067328.800000ns, VSS,
+ 1067448.800000ns, VSS,
+ 1067448.900000ns, VDD,
+ 1068169.400000ns, VDD,
+ 1068169.500000ns, VSS,
+ 1068769.900000ns, VSS,
+ 1068770.000000ns, VDD,
+ 1069010.100000ns, VDD,
+ 1069010.200000ns, VSS,
+ 1069250.300000ns, VSS,
+ 1069250.400000ns, VDD,
+ 1069370.400000ns, VDD,
+ 1069370.500000ns, VSS,
+ 1070091.000000ns, VSS,
+ 1070091.100000ns, VDD,
+ 1070451.300000ns, VDD,
+ 1070451.400000ns, VSS,
+ 1070571.400000ns, VSS,
+ 1070571.500000ns, VDD,
+ 1071171.900000ns, VDD,
+ 1071172.000000ns, VSS,
+ 1071292.000000ns, VSS,
+ 1071292.100000ns, VDD,
+ 1071772.400000ns, VDD,
+ 1071772.500000ns, VSS,
+ 1072132.700000ns, VSS,
+ 1072132.800000ns, VDD,
+ 1072853.300000ns, VDD,
+ 1072853.400000ns, VSS,
+ 1072973.400000ns, VSS,
+ 1072973.500000ns, VDD,
+ 1073333.700000ns, VDD,
+ 1073333.800000ns, VSS,
+ 1073814.100000ns, VSS,
+ 1073814.200000ns, VDD,
+ 1074054.300000ns, VDD,
+ 1074054.400000ns, VSS,
+ 1074654.800000ns, VSS,
+ 1074654.900000ns, VDD,
+ 1075135.200000ns, VDD,
+ 1075135.300000ns, VSS,
+ 1075615.600000ns, VSS,
+ 1075615.700000ns, VDD,
+ 1075735.700000ns, VDD,
+ 1075735.800000ns, VSS,
+ 1076456.300000ns, VSS,
+ 1076456.400000ns, VDD,
+ 1076696.500000ns, VDD,
+ 1076696.600000ns, VSS,
+ 1076936.700000ns, VSS,
+ 1076936.800000ns, VDD,
+ 1077176.900000ns, VDD,
+ 1077177.000000ns, VSS,
+ 1078377.900000ns, VSS,
+ 1078378.000000ns, VDD,
+ 1078738.200000ns, VDD,
+ 1078738.300000ns, VSS,
+ 1079338.700000ns, VSS,
+ 1079338.800000ns, VDD,
+ 1079939.200000ns, VDD,
+ 1079939.300000ns, VSS,
+ 1081020.100000ns, VSS,
+ 1081020.200000ns, VDD,
+ 1081140.200000ns, VDD,
+ 1081140.300000ns, VSS,
+ 1081260.300000ns, VSS,
+ 1081260.400000ns, VDD,
+ 1081500.500000ns, VDD,
+ 1081500.600000ns, VSS,
+ 1081740.700000ns, VSS,
+ 1081740.800000ns, VDD,
+ 1081980.900000ns, VDD,
+ 1081981.000000ns, VSS,
+ 1082101.000000ns, VSS,
+ 1082101.100000ns, VDD,
+ 1082701.500000ns, VDD,
+ 1082701.600000ns, VSS,
+ 1083302.000000ns, VSS,
+ 1083302.100000ns, VDD,
+ 1083422.100000ns, VDD,
+ 1083422.200000ns, VSS,
+ 1084262.800000ns, VSS,
+ 1084262.900000ns, VDD,
+ 1084382.900000ns, VDD,
+ 1084383.000000ns, VSS,
+ 1084743.200000ns, VSS,
+ 1084743.300000ns, VDD,
+ 1084983.400000ns, VDD,
+ 1084983.500000ns, VSS,
+ 1085103.500000ns, VSS,
+ 1085103.600000ns, VDD,
+ 1085704.000000ns, VDD,
+ 1085704.100000ns, VSS,
+ 1085824.100000ns, VSS,
+ 1085824.200000ns, VDD,
+ 1087145.200000ns, VDD,
+ 1087145.300000ns, VSS,
+ 1087505.500000ns, VSS,
+ 1087505.600000ns, VDD,
+ 1087745.700000ns, VDD,
+ 1087745.800000ns, VSS,
+ 1087865.800000ns, VSS,
+ 1087865.900000ns, VDD,
+ 1088106.000000ns, VDD,
+ 1088106.100000ns, VSS,
+ 1088226.100000ns, VSS,
+ 1088226.200000ns, VDD,
+ 1088466.300000ns, VDD,
+ 1088466.400000ns, VSS,
+ 1089307.000000ns, VSS,
+ 1089307.100000ns, VDD,
+ 1090027.600000ns, VDD,
+ 1090027.700000ns, VSS,
+ 1090147.700000ns, VSS,
+ 1090147.800000ns, VDD,
+ 1090508.000000ns, VDD,
+ 1090508.100000ns, VSS,
+ 1090988.400000ns, VSS,
+ 1090988.500000ns, VDD,
+ 1091709.000000ns, VDD,
+ 1091709.100000ns, VSS,
+ 1091829.100000ns, VSS,
+ 1091829.200000ns, VDD,
+ 1092429.600000ns, VDD,
+ 1092429.700000ns, VSS,
+ 1092549.700000ns, VSS,
+ 1092549.800000ns, VDD,
+ 1093150.200000ns, VDD,
+ 1093150.300000ns, VSS,
+ 1093270.300000ns, VSS,
+ 1093270.400000ns, VDD,
+ 1093510.500000ns, VDD,
+ 1093510.600000ns, VSS,
+ 1093870.800000ns, VSS,
+ 1093870.900000ns, VDD,
+ 1094111.000000ns, VDD,
+ 1094111.100000ns, VSS,
+ 1094351.200000ns, VSS,
+ 1094351.300000ns, VDD,
+ 1094831.600000ns, VDD,
+ 1094831.700000ns, VSS,
+ 1094951.700000ns, VSS,
+ 1094951.800000ns, VDD,
+ 1095432.100000ns, VDD,
+ 1095432.200000ns, VSS,
+ 1096152.700000ns, VSS,
+ 1096152.800000ns, VDD,
+ 1096513.000000ns, VDD,
+ 1096513.100000ns, VSS,
+ 1096873.300000ns, VSS,
+ 1096873.400000ns, VDD,
+ 1097834.100000ns, VDD,
+ 1097834.200000ns, VSS,
+ 1098074.300000ns, VSS,
+ 1098074.400000ns, VDD,
+ 1098194.400000ns, VDD,
+ 1098194.500000ns, VSS,
+ 1098434.600000ns, VSS,
+ 1098434.700000ns, VDD,
+ 1099275.300000ns, VDD,
+ 1099275.400000ns, VSS,
+ 1099635.600000ns, VSS,
+ 1099635.700000ns, VDD,
+ 1099755.700000ns, VDD,
+ 1099755.800000ns, VSS,
+ 1099995.900000ns, VSS,
+ 1099996.000000ns, VDD,
+ 1100116.000000ns, VDD,
+ 1100116.100000ns, VSS,
+ 1100476.300000ns, VSS,
+ 1100476.400000ns, VDD,
+ 1100596.400000ns, VDD,
+ 1100596.500000ns, VSS,
+ 1100836.600000ns, VSS,
+ 1100836.700000ns, VDD,
+ 1100956.700000ns, VDD,
+ 1100956.800000ns, VSS,
+ 1101076.800000ns, VSS,
+ 1101076.900000ns, VDD,
+ 1101677.300000ns, VDD,
+ 1101677.400000ns, VSS,
+ 1101797.400000ns, VSS,
+ 1101797.500000ns, VDD,
+ 1102037.600000ns, VDD,
+ 1102037.700000ns, VSS,
+ 1102397.900000ns, VSS,
+ 1102398.000000ns, VDD,
+ 1102518.000000ns, VDD,
+ 1102518.100000ns, VSS,
+ 1102638.100000ns, VSS,
+ 1102638.200000ns, VDD,
+ 1102878.300000ns, VDD,
+ 1102878.400000ns, VSS,
+ 1102998.400000ns, VSS,
+ 1102998.500000ns, VDD,
+ 1103719.000000ns, VDD,
+ 1103719.100000ns, VSS,
+ 1104319.500000ns, VSS,
+ 1104319.600000ns, VDD,
+ 1105280.300000ns, VDD,
+ 1105280.400000ns, VSS,
+ 1105400.400000ns, VSS,
+ 1105400.500000ns, VDD,
+ 1105640.600000ns, VDD,
+ 1105640.700000ns, VSS,
+ 1106000.900000ns, VSS,
+ 1106001.000000ns, VDD,
+ 1106121.000000ns, VDD,
+ 1106121.100000ns, VSS,
+ 1106841.600000ns, VSS,
+ 1106841.700000ns, VDD,
+ 1107081.800000ns, VDD,
+ 1107081.900000ns, VSS,
+ 1107201.900000ns, VSS,
+ 1107202.000000ns, VDD,
+ 1107802.400000ns, VDD,
+ 1107802.500000ns, VSS,
+ 1107922.500000ns, VSS,
+ 1107922.600000ns, VDD,
+ 1108282.800000ns, VDD,
+ 1108282.900000ns, VSS,
+ 1108402.900000ns, VSS,
+ 1108403.000000ns, VDD,
+ 1109123.500000ns, VDD,
+ 1109123.600000ns, VSS,
+ 1109243.600000ns, VSS,
+ 1109243.700000ns, VDD,
+ 1109483.800000ns, VDD,
+ 1109483.900000ns, VSS,
+ 1109844.100000ns, VSS,
+ 1109844.200000ns, VDD,
+ 1109964.200000ns, VDD,
+ 1109964.300000ns, VSS,
+ 1110084.300000ns, VSS,
+ 1110084.400000ns, VDD,
+ 1110564.700000ns, VDD,
+ 1110564.800000ns, VSS,
+ 1110804.900000ns, VSS,
+ 1110805.000000ns, VDD,
+ 1111285.300000ns, VDD,
+ 1111285.400000ns, VSS,
+ 1112246.100000ns, VSS,
+ 1112246.200000ns, VDD,
+ 1112486.300000ns, VDD,
+ 1112486.400000ns, VSS,
+ 1112846.600000ns, VSS,
+ 1112846.700000ns, VDD,
+ 1113567.200000ns, VDD,
+ 1113567.300000ns, VSS,
+ 1113927.500000ns, VSS,
+ 1113927.600000ns, VDD,
+ 1114648.100000ns, VDD,
+ 1114648.200000ns, VSS,
+ 1114768.200000ns, VSS,
+ 1114768.300000ns, VDD,
+ 1115128.500000ns, VDD,
+ 1115128.600000ns, VSS,
+ 1115248.600000ns, VSS,
+ 1115248.700000ns, VDD,
+ 1115729.000000ns, VDD,
+ 1115729.100000ns, VSS,
+ 1116329.500000ns, VSS,
+ 1116329.600000ns, VDD,
+ 1116689.800000ns, VDD,
+ 1116689.900000ns, VSS,
+ 1117290.300000ns, VSS,
+ 1117290.400000ns, VDD,
+ 1117530.500000ns, VDD,
+ 1117530.600000ns, VSS,
+ 1118491.300000ns, VSS,
+ 1118491.400000ns, VDD,
+ 1118851.600000ns, VDD,
+ 1118851.700000ns, VSS,
+ 1119572.200000ns, VSS,
+ 1119572.300000ns, VDD,
+ 1120052.600000ns, VDD,
+ 1120052.700000ns, VSS,
+ 1120773.200000ns, VSS,
+ 1120773.300000ns, VDD,
+ 1121373.700000ns, VDD,
+ 1121373.800000ns, VSS,
+ 1121493.800000ns, VSS,
+ 1121493.900000ns, VDD,
+ 1122094.300000ns, VDD,
+ 1122094.400000ns, VSS,
+ 1123055.100000ns, VSS,
+ 1123055.200000ns, VDD,
+ 1123655.600000ns, VDD,
+ 1123655.700000ns, VSS,
+ 1124136.000000ns, VSS,
+ 1124136.100000ns, VDD,
+ 1124256.100000ns, VDD,
+ 1124256.200000ns, VSS,
+ 1124856.600000ns, VSS,
+ 1124856.700000ns, VDD,
+ 1125337.000000ns, VDD,
+ 1125337.100000ns, VSS,
+ 1125457.100000ns, VSS,
+ 1125457.200000ns, VDD,
+ 1125697.300000ns, VDD,
+ 1125697.400000ns, VSS,
+ 1125937.500000ns, VSS,
+ 1125937.600000ns, VDD,
+ 1126778.200000ns, VDD,
+ 1126778.300000ns, VSS,
+ 1126898.300000ns, VSS,
+ 1126898.400000ns, VDD,
+ 1127859.100000ns, VDD,
+ 1127859.200000ns, VSS,
+ 1127979.200000ns, VSS,
+ 1127979.300000ns, VDD,
+ 1128219.400000ns, VDD,
+ 1128219.500000ns, VSS,
+ 1128339.500000ns, VSS,
+ 1128339.600000ns, VDD,
+ 1128819.900000ns, VDD,
+ 1128820.000000ns, VSS,
+ 1128940.000000ns, VSS,
+ 1128940.100000ns, VDD,
+ 1129180.200000ns, VDD,
+ 1129180.300000ns, VSS,
+ 1129420.400000ns, VSS,
+ 1129420.500000ns, VDD,
+ 1129540.500000ns, VDD,
+ 1129540.600000ns, VSS,
+ 1129660.600000ns, VSS,
+ 1129660.700000ns, VDD,
+ 1130261.100000ns, VDD,
+ 1130261.200000ns, VSS,
+ 1130621.400000ns, VSS,
+ 1130621.500000ns, VDD,
+ 1130741.500000ns, VDD,
+ 1130741.600000ns, VSS,
+ 1131221.900000ns, VSS,
+ 1131222.000000ns, VDD,
+ 1131342.000000ns, VDD,
+ 1131342.100000ns, VSS,
+ 1132062.600000ns, VSS,
+ 1132062.700000ns, VDD,
+ 1132543.000000ns, VDD,
+ 1132543.100000ns, VSS,
+ 1132663.100000ns, VSS,
+ 1132663.200000ns, VDD,
+ 1133143.500000ns, VDD,
+ 1133143.600000ns, VSS,
+ 1133383.700000ns, VSS,
+ 1133383.800000ns, VDD,
+ 1133623.900000ns, VDD,
+ 1133624.000000ns, VSS,
+ 1133984.200000ns, VSS,
+ 1133984.300000ns, VDD,
+ 1134104.300000ns, VDD,
+ 1134104.400000ns, VSS,
+ 1134464.600000ns, VSS,
+ 1134464.700000ns, VDD,
+ 1135185.200000ns, VDD,
+ 1135185.300000ns, VSS,
+ 1135305.300000ns, VSS,
+ 1135305.400000ns, VDD,
+ 1135905.800000ns, VDD,
+ 1135905.900000ns, VSS,
+ 1136386.200000ns, VSS,
+ 1136386.300000ns, VDD,
+ 1136866.600000ns, VDD,
+ 1136866.700000ns, VSS,
+ 1137347.000000ns, VSS,
+ 1137347.100000ns, VDD,
+ 1137467.100000ns, VDD,
+ 1137467.200000ns, VSS,
+ 1137827.400000ns, VSS,
+ 1137827.500000ns, VDD,
+ 1138788.200000ns, VDD,
+ 1138788.300000ns, VSS,
+ 1139148.500000ns, VSS,
+ 1139148.600000ns, VDD,
+ 1139388.700000ns, VDD,
+ 1139388.800000ns, VSS,
+ 1139749.000000ns, VSS,
+ 1139749.100000ns, VDD,
+ 1141310.300000ns, VDD,
+ 1141310.400000ns, VSS,
+ 1142151.000000ns, VSS,
+ 1142151.100000ns, VDD,
+ 1142631.400000ns, VDD,
+ 1142631.500000ns, VSS,
+ 1142991.700000ns, VSS,
+ 1142991.800000ns, VDD,
+ 1143111.800000ns, VDD,
+ 1143111.900000ns, VSS,
+ 1143352.000000ns, VSS,
+ 1143352.100000ns, VDD,
+ 1143472.100000ns, VDD,
+ 1143472.200000ns, VSS,
+ 1143712.300000ns, VSS,
+ 1143712.400000ns, VDD,
+ 1144913.300000ns, VDD,
+ 1144913.400000ns, VSS,
+ 1145033.400000ns, VSS,
+ 1145033.500000ns, VDD,
+ 1145273.600000ns, VDD,
+ 1145273.700000ns, VSS,
+ 1145513.800000ns, VSS,
+ 1145513.900000ns, VDD,
+ 1145874.100000ns, VDD,
+ 1145874.200000ns, VSS,
+ 1145994.200000ns, VSS,
+ 1145994.300000ns, VDD,
+ 1146594.700000ns, VDD,
+ 1146594.800000ns, VSS,
+ 1146955.000000ns, VSS,
+ 1146955.100000ns, VDD,
+ 1147075.100000ns, VDD,
+ 1147075.200000ns, VSS,
+ 1147915.800000ns, VSS,
+ 1147915.900000ns, VDD,
+ 1148276.100000ns, VDD,
+ 1148276.200000ns, VSS,
+ 1148756.500000ns, VSS,
+ 1148756.600000ns, VDD,
+ 1148996.700000ns, VDD,
+ 1148996.800000ns, VSS,
+ 1149597.200000ns, VSS,
+ 1149597.300000ns, VDD,
+ 1149837.400000ns, VDD,
+ 1149837.500000ns, VSS,
+ 1149957.500000ns, VSS,
+ 1149957.600000ns, VDD,
+ 1150317.800000ns, VDD,
+ 1150317.900000ns, VSS,
+ 1150798.200000ns, VSS,
+ 1150798.300000ns, VDD,
+ 1150918.300000ns, VDD,
+ 1150918.400000ns, VSS,
+ 1151278.600000ns, VSS,
+ 1151278.700000ns, VDD,
+ 1152239.400000ns, VDD,
+ 1152239.500000ns, VSS,
+ 1152359.500000ns, VSS,
+ 1152359.600000ns, VDD,
+ 1152839.900000ns, VDD,
+ 1152840.000000ns, VSS,
+ 1153200.200000ns, VSS,
+ 1153200.300000ns, VDD,
+ 1153800.700000ns, VDD,
+ 1153800.800000ns, VSS,
+ 1154161.000000ns, VSS,
+ 1154161.100000ns, VDD,
+ 1154401.200000ns, VDD,
+ 1154401.300000ns, VSS,
+ 1154881.600000ns, VSS,
+ 1154881.700000ns, VDD,
+ 1155241.900000ns, VDD,
+ 1155242.000000ns, VSS,
+ 1155602.200000ns, VSS,
+ 1155602.300000ns, VDD,
+ 1156082.600000ns, VDD,
+ 1156082.700000ns, VSS,
+ 1156202.700000ns, VSS,
+ 1156202.800000ns, VDD,
+ 1156442.900000ns, VDD,
+ 1156443.000000ns, VSS,
+ 1156683.100000ns, VSS,
+ 1156683.200000ns, VDD,
+ 1157523.800000ns, VDD,
+ 1157523.900000ns, VSS,
+ 1157884.100000ns, VSS,
+ 1157884.200000ns, VDD,
+ 1158124.300000ns, VDD,
+ 1158124.400000ns, VSS,
+ 1158244.400000ns, VSS,
+ 1158244.500000ns, VDD,
+ 1158484.600000ns, VDD,
+ 1158484.700000ns, VSS,
+ 1158604.700000ns, VSS,
+ 1158604.800000ns, VDD,
+ 1159205.200000ns, VDD,
+ 1159205.300000ns, VSS,
+ 1159685.600000ns, VSS,
+ 1159685.700000ns, VDD,
+ 1160045.900000ns, VDD,
+ 1160046.000000ns, VSS,
+ 1160166.000000ns, VSS,
+ 1160166.100000ns, VDD,
+ 1160526.300000ns, VDD,
+ 1160526.400000ns, VSS,
+ 1161367.000000ns, VSS,
+ 1161367.100000ns, VDD,
+ 1161847.400000ns, VDD,
+ 1161847.500000ns, VSS,
+ 1162447.900000ns, VSS,
+ 1162448.000000ns, VDD,
+ 1162808.200000ns, VDD,
+ 1162808.300000ns, VSS,
+ 1163769.000000ns, VSS,
+ 1163769.100000ns, VDD,
+ 1164369.500000ns, VDD,
+ 1164369.600000ns, VSS,
+ 1164489.600000ns, VSS,
+ 1164489.700000ns, VDD,
+ 1165210.200000ns, VDD,
+ 1165210.300000ns, VSS,
+ 1165450.400000ns, VSS,
+ 1165450.500000ns, VDD,
+ 1166291.100000ns, VDD,
+ 1166291.200000ns, VSS,
+ 1166411.200000ns, VSS,
+ 1166411.300000ns, VDD,
+ 1166891.600000ns, VDD,
+ 1166891.700000ns, VSS,
+ 1167251.900000ns, VSS,
+ 1167252.000000ns, VDD,
+ 1167492.100000ns, VDD,
+ 1167492.200000ns, VSS,
+ 1167612.200000ns, VSS,
+ 1167612.300000ns, VDD,
+ 1167852.400000ns, VDD,
+ 1167852.500000ns, VSS,
+ 1168092.600000ns, VSS,
+ 1168092.700000ns, VDD,
+ 1168332.800000ns, VDD,
+ 1168332.900000ns, VSS,
+ 1168933.300000ns, VSS,
+ 1168933.400000ns, VDD,
+ 1169533.800000ns, VDD,
+ 1169533.900000ns, VSS,
+ 1169894.100000ns, VSS,
+ 1169894.200000ns, VDD,
+ 1170134.300000ns, VDD,
+ 1170134.400000ns, VSS,
+ 1170374.500000ns, VSS,
+ 1170374.600000ns, VDD,
+ 1170494.600000ns, VDD,
+ 1170494.700000ns, VSS,
+ 1170854.900000ns, VSS,
+ 1170855.000000ns, VDD,
+ 1171095.100000ns, VDD,
+ 1171095.200000ns, VSS,
+ 1172176.000000ns, VSS,
+ 1172176.100000ns, VDD,
+ 1172416.200000ns, VDD,
+ 1172416.300000ns, VSS,
+ 1172776.500000ns, VSS,
+ 1172776.600000ns, VDD,
+ 1173377.000000ns, VDD,
+ 1173377.100000ns, VSS,
+ 1173497.100000ns, VSS,
+ 1173497.200000ns, VDD,
+ 1173737.300000ns, VDD,
+ 1173737.400000ns, VSS,
+ 1173857.400000ns, VSS,
+ 1173857.500000ns, VDD,
+ 1174217.700000ns, VDD,
+ 1174217.800000ns, VSS,
+ 1174578.000000ns, VSS,
+ 1174578.100000ns, VDD,
+ 1174818.200000ns, VDD,
+ 1174818.300000ns, VSS,
+ 1174938.300000ns, VSS,
+ 1174938.400000ns, VDD,
+ 1175178.500000ns, VDD,
+ 1175178.600000ns, VSS,
+ 1175538.800000ns, VSS,
+ 1175538.900000ns, VDD,
+ 1175779.000000ns, VDD,
+ 1175779.100000ns, VSS,
+ 1175899.100000ns, VSS,
+ 1175899.200000ns, VDD,
+ 1176019.200000ns, VDD,
+ 1176019.300000ns, VSS,
+ 1176139.300000ns, VSS,
+ 1176139.400000ns, VDD,
+ 1177340.300000ns, VDD,
+ 1177340.400000ns, VSS,
+ 1177460.400000ns, VSS,
+ 1177460.500000ns, VDD,
+ 1178421.200000ns, VDD,
+ 1178421.300000ns, VSS,
+ 1178541.300000ns, VSS,
+ 1178541.400000ns, VDD,
+ 1178901.600000ns, VDD,
+ 1178901.700000ns, VSS,
+ 1179021.700000ns, VSS,
+ 1179021.800000ns, VDD,
+ 1179502.100000ns, VDD,
+ 1179502.200000ns, VSS,
+ 1179622.200000ns, VSS,
+ 1179622.300000ns, VDD,
+ 1179982.500000ns, VDD,
+ 1179982.600000ns, VSS,
+ 1180102.600000ns, VSS,
+ 1180102.700000ns, VDD,
+ 1180462.900000ns, VDD,
+ 1180463.000000ns, VSS,
+ 1180583.000000ns, VSS,
+ 1180583.100000ns, VDD,
+ 1181423.700000ns, VDD,
+ 1181423.800000ns, VSS,
+ 1182384.500000ns, VSS,
+ 1182384.600000ns, VDD,
+ 1182504.600000ns, VDD,
+ 1182504.700000ns, VSS,
+ 1182864.900000ns, VSS,
+ 1182865.000000ns, VDD,
+ 1183105.100000ns, VDD,
+ 1183105.200000ns, VSS,
+ 1183465.400000ns, VSS,
+ 1183465.500000ns, VDD,
+ 1183705.600000ns, VDD,
+ 1183705.700000ns, VSS,
+ 1184306.100000ns, VSS,
+ 1184306.200000ns, VDD,
+ 1184666.400000ns, VDD,
+ 1184666.500000ns, VSS,
+ 1184786.500000ns, VSS,
+ 1184786.600000ns, VDD,
+ 1185747.300000ns, VDD,
+ 1185747.400000ns, VSS,
+ 1186107.600000ns, VSS,
+ 1186107.700000ns, VDD,
+ 1186347.800000ns, VDD,
+ 1186347.900000ns, VSS,
+ 1186467.900000ns, VSS,
+ 1186468.000000ns, VDD,
+ 1186708.100000ns, VDD,
+ 1186708.200000ns, VSS,
+ 1186948.300000ns, VSS,
+ 1186948.400000ns, VDD,
+ 1187188.500000ns, VDD,
+ 1187188.600000ns, VSS,
+ 1187428.700000ns, VSS,
+ 1187428.800000ns, VDD,
+ 1187789.000000ns, VDD,
+ 1187789.100000ns, VSS,
+ 1187909.100000ns, VSS,
+ 1187909.200000ns, VDD,
+ 1188389.500000ns, VDD,
+ 1188389.600000ns, VSS,
+ 1190191.000000ns, VSS,
+ 1190191.100000ns, VDD,
+ 1190431.200000ns, VDD,
+ 1190431.300000ns, VSS,
+ 1191151.800000ns, VSS,
+ 1191151.900000ns, VDD,
+ 1191512.100000ns, VDD,
+ 1191512.200000ns, VSS,
+ 1191872.400000ns, VSS,
+ 1191872.500000ns, VDD,
+ 1192352.800000ns, VDD,
+ 1192352.900000ns, VSS,
+ 1192472.900000ns, VSS,
+ 1192473.000000ns, VDD,
+ 1192833.200000ns, VDD,
+ 1192833.300000ns, VSS,
+ 1192953.300000ns, VSS,
+ 1192953.400000ns, VDD,
+ 1193193.500000ns, VDD,
+ 1193193.600000ns, VSS,
+ 1193553.800000ns, VSS,
+ 1193553.900000ns, VDD,
+ 1194154.300000ns, VDD,
+ 1194154.400000ns, VSS,
+ 1194274.400000ns, VSS,
+ 1194274.500000ns, VDD,
+ 1194995.000000ns, VDD,
+ 1194995.100000ns, VSS,
+ 1195595.500000ns, VSS,
+ 1195595.600000ns, VDD,
+ 1195955.800000ns, VDD,
+ 1195955.900000ns, VSS,
+ 1196316.100000ns, VSS,
+ 1196316.200000ns, VDD,
+ 1196436.200000ns, VDD,
+ 1196436.300000ns, VSS,
+ 1196796.500000ns, VSS,
+ 1196796.600000ns, VDD,
+ 1197397.000000ns, VDD,
+ 1197397.100000ns, VSS,
+ 1197517.100000ns, VSS,
+ 1197517.200000ns, VDD,
+ 1197877.400000ns, VDD,
+ 1197877.500000ns, VSS,
+ 1197997.500000ns, VSS,
+ 1197997.600000ns, VDD,
+ 1198237.700000ns, VDD,
+ 1198237.800000ns, VSS,
+ 1198718.100000ns, VSS,
+ 1198718.200000ns, VDD,
+ 1199558.800000ns, VDD,
+ 1199558.900000ns, VSS,
+ 1200159.300000ns, VSS,
+ 1200159.400000ns, VDD,
+ 1200399.500000ns, VDD,
+ 1200399.600000ns, VSS,
+ 1200879.900000ns, VSS,
+ 1200880.000000ns, VDD,
+ 1201480.400000ns, VDD,
+ 1201480.500000ns, VSS,
+ 1201600.500000ns, VSS,
+ 1201600.600000ns, VDD,
+ 1202201.000000ns, VDD,
+ 1202201.100000ns, VSS,
+ 1202321.100000ns, VSS,
+ 1202321.200000ns, VDD,
+ 1202561.300000ns, VDD,
+ 1202561.400000ns, VSS,
+ 1202681.400000ns, VSS,
+ 1202681.500000ns, VDD,
+ 1203882.400000ns, VDD,
+ 1203882.500000ns, VSS,
+ 1204122.600000ns, VSS,
+ 1204122.700000ns, VDD,
+ 1204723.100000ns, VDD,
+ 1204723.200000ns, VSS,
+ 1205563.800000ns, VSS,
+ 1205563.900000ns, VDD,
+ 1205683.900000ns, VDD,
+ 1205684.000000ns, VSS,
+ 1206044.200000ns, VSS,
+ 1206044.300000ns, VDD,
+ 1206284.400000ns, VDD,
+ 1206284.500000ns, VSS,
+ 1206764.800000ns, VSS,
+ 1206764.900000ns, VDD,
+ 1207125.100000ns, VDD,
+ 1207125.200000ns, VSS,
+ 1207485.400000ns, VSS,
+ 1207485.500000ns, VDD,
+ 1208806.500000ns, VDD,
+ 1208806.600000ns, VSS,
+ 1208926.600000ns, VSS,
+ 1208926.700000ns, VDD,
+ 1209286.900000ns, VDD,
+ 1209287.000000ns, VSS,
+ 1209407.000000ns, VSS,
+ 1209407.100000ns, VDD,
+ 1209527.100000ns, VDD,
+ 1209527.200000ns, VSS,
+ 1210007.500000ns, VSS,
+ 1210007.600000ns, VDD,
+ 1210608.000000ns, VDD,
+ 1210608.100000ns, VSS,
+ 1211208.500000ns, VSS,
+ 1211208.600000ns, VDD,
+ 1211568.800000ns, VDD,
+ 1211568.900000ns, VSS,
+ 1211688.900000ns, VSS,
+ 1211689.000000ns, VDD,
+ 1211929.100000ns, VDD,
+ 1211929.200000ns, VSS,
+ 1212169.300000ns, VSS,
+ 1212169.400000ns, VDD,
+ 1213970.800000ns, VDD,
+ 1213970.900000ns, VSS,
+ 1214211.000000ns, VSS,
+ 1214211.100000ns, VDD,
+ 1214331.100000ns, VDD,
+ 1214331.200000ns, VSS,
+ 1214691.400000ns, VSS,
+ 1214691.500000ns, VDD,
+ 1214811.500000ns, VDD,
+ 1214811.600000ns, VSS,
+ 1215291.900000ns, VSS,
+ 1215292.000000ns, VDD,
+ 1215532.100000ns, VDD,
+ 1215532.200000ns, VSS,
+ 1215652.200000ns, VSS,
+ 1215652.300000ns, VDD,
+ 1216132.600000ns, VDD,
+ 1216132.700000ns, VSS,
+ 1216492.900000ns, VSS,
+ 1216493.000000ns, VDD,
+ 1216733.100000ns, VDD,
+ 1216733.200000ns, VSS,
+ 1216853.200000ns, VSS,
+ 1216853.300000ns, VDD,
+ 1217093.400000ns, VDD,
+ 1217093.500000ns, VSS,
+ 1217453.700000ns, VSS,
+ 1217453.800000ns, VDD,
+ 1217573.800000ns, VDD,
+ 1217573.900000ns, VSS,
+ 1217693.900000ns, VSS,
+ 1217694.000000ns, VDD,
+ 1217934.100000ns, VDD,
+ 1217934.200000ns, VSS,
+ 1218294.400000ns, VSS,
+ 1218294.500000ns, VDD,
+ 1218774.800000ns, VDD,
+ 1218774.900000ns, VSS,
+ 1219735.600000ns, VSS,
+ 1219735.700000ns, VDD,
+ 1220336.100000ns, VDD,
+ 1220336.200000ns, VSS,
+ 1220456.200000ns, VSS,
+ 1220456.300000ns, VDD,
+ 1220816.500000ns, VDD,
+ 1220816.600000ns, VSS,
+ 1221056.700000ns, VSS,
+ 1221056.800000ns, VDD,
+ 1221777.300000ns, VDD,
+ 1221777.400000ns, VSS,
+ 1222257.700000ns, VSS,
+ 1222257.800000ns, VDD,
+ 1222377.800000ns, VDD,
+ 1222377.900000ns, VSS,
+ 1222858.200000ns, VSS,
+ 1222858.300000ns, VDD,
+ 1223098.400000ns, VDD,
+ 1223098.500000ns, VSS,
+ 1223458.700000ns, VSS,
+ 1223458.800000ns, VDD,
+ 1223578.800000ns, VDD,
+ 1223578.900000ns, VSS,
+ 1224779.800000ns, VSS,
+ 1224779.900000ns, VDD,
+ 1224899.900000ns, VDD,
+ 1224900.000000ns, VSS,
+ 1225380.300000ns, VSS,
+ 1225380.400000ns, VDD,
+ 1225860.700000ns, VDD,
+ 1225860.800000ns, VSS,
+ 1225980.800000ns, VSS,
+ 1225980.900000ns, VDD,
+ 1226341.100000ns, VDD,
+ 1226341.200000ns, VSS,
+ 1226581.300000ns, VSS,
+ 1226581.400000ns, VDD,
+ 1226821.500000ns, VDD,
+ 1226821.600000ns, VSS,
+ 1227061.700000ns, VSS,
+ 1227061.800000ns, VDD,
+ 1227422.000000ns, VDD,
+ 1227422.100000ns, VSS,
+ 1227782.300000ns, VSS,
+ 1227782.400000ns, VDD,
+ 1228142.600000ns, VDD,
+ 1228142.700000ns, VSS,
+ 1228262.700000ns, VSS,
+ 1228262.800000ns, VDD,
+ 1228502.900000ns, VDD,
+ 1228503.000000ns, VSS,
+ 1228863.200000ns, VSS,
+ 1228863.300000ns, VDD,
+ 1229343.600000ns, VDD,
+ 1229343.700000ns, VSS,
+ 1230064.200000ns, VSS,
+ 1230064.300000ns, VDD,
+ 1230304.400000ns, VDD,
+ 1230304.500000ns, VSS,
+ 1230664.700000ns, VSS,
+ 1230664.800000ns, VDD,
+ 1230784.800000ns, VDD,
+ 1230784.900000ns, VSS,
+ 1230904.900000ns, VSS,
+ 1230905.000000ns, VDD,
+ 1231265.200000ns, VDD,
+ 1231265.300000ns, VSS,
+ 1231745.600000ns, VSS,
+ 1231745.700000ns, VDD,
+ 1231865.700000ns, VDD,
+ 1231865.800000ns, VSS,
+ 1232346.100000ns, VSS,
+ 1232346.200000ns, VDD,
+ 1232586.300000ns, VDD,
+ 1232586.400000ns, VSS,
+ 1233427.000000ns, VSS,
+ 1233427.100000ns, VDD,
+ 1233667.200000ns, VDD,
+ 1233667.300000ns, VSS,
+ 1233907.400000ns, VSS,
+ 1233907.500000ns, VDD,
+ 1234748.100000ns, VDD,
+ 1234748.200000ns, VSS,
+ 1235588.800000ns, VSS,
+ 1235588.900000ns, VDD,
+ 1235708.900000ns, VDD,
+ 1235709.000000ns, VSS,
+ 1235829.000000ns, VSS,
+ 1235829.100000ns, VDD,
+ 1236669.700000ns, VDD,
+ 1236669.800000ns, VSS,
+ 1238351.100000ns, VSS,
+ 1238351.200000ns, VDD,
+ 1238591.300000ns, VDD,
+ 1238591.400000ns, VSS,
+ 1238951.600000ns, VSS,
+ 1238951.700000ns, VDD,
+ 1239552.100000ns, VDD,
+ 1239552.200000ns, VSS,
+ 1239672.200000ns, VSS,
+ 1239672.300000ns, VDD,
+ 1240032.500000ns, VDD,
+ 1240032.600000ns, VSS,
+ 1240392.800000ns, VSS,
+ 1240392.900000ns, VDD,
+ 1240633.000000ns, VDD,
+ 1240633.100000ns, VSS,
+ 1240993.300000ns, VSS,
+ 1240993.400000ns, VDD,
+ 1241233.500000ns, VDD,
+ 1241233.600000ns, VSS,
+ 1242194.300000ns, VSS,
+ 1242194.400000ns, VDD,
+ 1242794.800000ns, VDD,
+ 1242794.900000ns, VSS,
+ 1242914.900000ns, VSS,
+ 1242915.000000ns, VDD,
+ 1243395.300000ns, VDD,
+ 1243395.400000ns, VSS,
+ 1243635.500000ns, VSS,
+ 1243635.600000ns, VDD,
+ 1243995.800000ns, VDD,
+ 1243995.900000ns, VSS,
+ 1244236.000000ns, VSS,
+ 1244236.100000ns, VDD,
+ 1245076.700000ns, VDD,
+ 1245076.800000ns, VSS,
+ 1245437.000000ns, VSS,
+ 1245437.100000ns, VDD,
+ 1246157.600000ns, VDD,
+ 1246157.700000ns, VSS,
+ 1246878.200000ns, VSS,
+ 1246878.300000ns, VDD,
+ 1247238.500000ns, VDD,
+ 1247238.600000ns, VSS,
+ 1247959.100000ns, VSS,
+ 1247959.200000ns, VDD,
+ 1248439.500000ns, VDD,
+ 1248439.600000ns, VSS,
+ 1249160.100000ns, VSS,
+ 1249160.200000ns, VDD,
+ 1249280.200000ns, VDD,
+ 1249280.300000ns, VSS,
+ 1250241.000000ns, VSS,
+ 1250241.100000ns, VDD,
+ 1250721.400000ns, VDD,
+ 1250721.500000ns, VSS,
+ 1250841.500000ns, VSS,
+ 1250841.600000ns, VDD,
+ 1251201.800000ns, VDD,
+ 1251201.900000ns, VSS,
+ 1251321.900000ns, VSS,
+ 1251322.000000ns, VDD,
+ 1251802.300000ns, VDD,
+ 1251802.400000ns, VSS,
+ 1253243.500000ns, VSS,
+ 1253243.600000ns, VDD,
+ 1253723.900000ns, VDD,
+ 1253724.000000ns, VSS,
+ 1254084.200000ns, VSS,
+ 1254084.300000ns, VDD,
+ 1254204.300000ns, VDD,
+ 1254204.400000ns, VSS,
+ 1254564.600000ns, VSS,
+ 1254564.700000ns, VDD,
+ 1254924.900000ns, VDD,
+ 1254925.000000ns, VSS,
+ 1255165.100000ns, VSS,
+ 1255165.200000ns, VDD,
+ 1255405.300000ns, VDD,
+ 1255405.400000ns, VSS,
+ 1256005.800000ns, VSS,
+ 1256005.900000ns, VDD,
+ 1256366.100000ns, VDD,
+ 1256366.200000ns, VSS,
+ 1256846.500000ns, VSS,
+ 1256846.600000ns, VDD,
+ 1256966.600000ns, VDD,
+ 1256966.700000ns, VSS,
+ 1257687.200000ns, VSS,
+ 1257687.300000ns, VDD,
+ 1258407.800000ns, VDD,
+ 1258407.900000ns, VSS,
+ 1258527.900000ns, VSS,
+ 1258528.000000ns, VDD,
+ 1259488.700000ns, VDD,
+ 1259488.800000ns, VSS,
+ 1259969.100000ns, VSS,
+ 1259969.200000ns, VDD,
+ 1260209.300000ns, VDD,
+ 1260209.400000ns, VSS,
+ 1260689.700000ns, VSS,
+ 1260689.800000ns, VDD,
+ 1260809.800000ns, VDD,
+ 1260809.900000ns, VSS,
+ 1261290.200000ns, VSS,
+ 1261290.300000ns, VDD,
+ 1262251.000000ns, VDD,
+ 1262251.100000ns, VSS,
+ 1262371.100000ns, VSS,
+ 1262371.200000ns, VDD,
+ 1262731.400000ns, VDD,
+ 1262731.500000ns, VSS,
+ 1262851.500000ns, VSS,
+ 1262851.600000ns, VDD,
+ 1264292.700000ns, VDD,
+ 1264292.800000ns, VSS,
+ 1264412.800000ns, VSS,
+ 1264412.900000ns, VDD,
+ 1264773.100000ns, VDD,
+ 1264773.200000ns, VSS,
+ 1264893.200000ns, VSS,
+ 1264893.300000ns, VDD,
+ 1265133.400000ns, VDD,
+ 1265133.500000ns, VSS,
+ 1265373.600000ns, VSS,
+ 1265373.700000ns, VDD,
+ 1265974.100000ns, VDD,
+ 1265974.200000ns, VSS,
+ 1267055.000000ns, VSS,
+ 1267055.100000ns, VDD,
+ 1267415.300000ns, VDD,
+ 1267415.400000ns, VSS,
+ 1267535.400000ns, VSS,
+ 1267535.500000ns, VDD,
+ 1267775.600000ns, VDD,
+ 1267775.700000ns, VSS,
+ 1267895.700000ns, VSS,
+ 1267895.800000ns, VDD,
+ 1268376.100000ns, VDD,
+ 1268376.200000ns, VSS,
+ 1268856.500000ns, VSS,
+ 1268856.600000ns, VDD,
+ 1269096.700000ns, VDD,
+ 1269096.800000ns, VSS,
+ 1270778.100000ns, VSS,
+ 1270778.200000ns, VDD,
+ 1271018.300000ns, VDD,
+ 1271018.400000ns, VSS,
+ 1271378.600000ns, VSS,
+ 1271378.700000ns, VDD,
+ 1271859.000000ns, VDD,
+ 1271859.100000ns, VSS,
+ 1272099.200000ns, VSS,
+ 1272099.300000ns, VDD,
+ 1272219.300000ns, VDD,
+ 1272219.400000ns, VSS,
+ 1272339.400000ns, VSS,
+ 1272339.500000ns, VDD,
+ 1272579.600000ns, VDD,
+ 1272579.700000ns, VSS,
+ 1272699.700000ns, VSS,
+ 1272699.800000ns, VDD,
+ 1273180.100000ns, VDD,
+ 1273180.200000ns, VSS,
+ 1273540.400000ns, VSS,
+ 1273540.500000ns, VDD,
+ 1273900.700000ns, VDD,
+ 1273900.800000ns, VSS,
+ 1274140.900000ns, VSS,
+ 1274141.000000ns, VDD,
+ 1274261.000000ns, VDD,
+ 1274261.100000ns, VSS,
+ 1274741.400000ns, VSS,
+ 1274741.500000ns, VDD,
+ 1275582.100000ns, VDD,
+ 1275582.200000ns, VSS,
+ 1275822.300000ns, VSS,
+ 1275822.400000ns, VDD,
+ 1275942.400000ns, VDD,
+ 1275942.500000ns, VSS,
+ 1276663.000000ns, VSS,
+ 1276663.100000ns, VDD,
+ 1277023.300000ns, VDD,
+ 1277023.400000ns, VSS,
+ 1277143.400000ns, VSS,
+ 1277143.500000ns, VDD,
+ 1277383.600000ns, VDD,
+ 1277383.700000ns, VSS,
+ 1277623.800000ns, VSS,
+ 1277623.900000ns, VDD,
+ 1279185.100000ns, VDD,
+ 1279185.200000ns, VSS,
+ 1279785.600000ns, VSS,
+ 1279785.700000ns, VDD,
+ 1279905.700000ns, VDD,
+ 1279905.800000ns, VSS,
+ 1280025.800000ns, VSS,
+ 1280025.900000ns, VDD,
+ 1280266.000000ns, VDD,
+ 1280266.100000ns, VSS,
+ 1281587.100000ns, VSS,
+ 1281587.200000ns, VDD,
+ 1282547.900000ns, VDD,
+ 1282548.000000ns, VSS,
+ 1282668.000000ns, VSS,
+ 1282668.100000ns, VDD,
+ 1282908.200000ns, VDD,
+ 1282908.300000ns, VSS,
+ 1283268.500000ns, VSS,
+ 1283268.600000ns, VDD,
+ 1283508.700000ns, VDD,
+ 1283508.800000ns, VSS,
+ 1283869.000000ns, VSS,
+ 1283869.100000ns, VDD,
+ 1283989.100000ns, VDD,
+ 1283989.200000ns, VSS,
+ 1284349.400000ns, VSS,
+ 1284349.500000ns, VDD,
+ 1284709.700000ns, VDD,
+ 1284709.800000ns, VSS,
+ 1285070.000000ns, VSS,
+ 1285070.100000ns, VDD,
+ 1285550.400000ns, VDD,
+ 1285550.500000ns, VSS,
+ 1286030.800000ns, VSS,
+ 1286030.900000ns, VDD,
+ 1286391.100000ns, VDD,
+ 1286391.200000ns, VSS,
+ 1286511.200000ns, VSS,
+ 1286511.300000ns, VDD,
+ 1286631.300000ns, VDD,
+ 1286631.400000ns, VSS,
+ 1286751.400000ns, VSS,
+ 1286751.500000ns, VDD,
+ 1287111.700000ns, VDD,
+ 1287111.800000ns, VSS,
+ 1287231.800000ns, VSS,
+ 1287231.900000ns, VDD,
+ 1287952.400000ns, VDD,
+ 1287952.500000ns, VSS,
+ 1288072.500000ns, VSS,
+ 1288072.600000ns, VDD,
+ 1288312.700000ns, VDD,
+ 1288312.800000ns, VSS,
+ 1288432.800000ns, VSS,
+ 1288432.900000ns, VDD,
+ 1288552.900000ns, VDD,
+ 1288553.000000ns, VSS,
+ 1288673.000000ns, VSS,
+ 1288673.100000ns, VDD,
+ 1288913.200000ns, VDD,
+ 1288913.300000ns, VSS,
+ 1289273.500000ns, VSS,
+ 1289273.600000ns, VDD,
+ 1290114.200000ns, VDD,
+ 1290114.300000ns, VSS,
+ 1290714.700000ns, VSS,
+ 1290714.800000ns, VDD,
+ 1290954.900000ns, VDD,
+ 1290955.000000ns, VSS,
+ 1291435.300000ns, VSS,
+ 1291435.400000ns, VDD,
+ 1291795.600000ns, VDD,
+ 1291795.700000ns, VSS,
+ 1292155.900000ns, VSS,
+ 1292156.000000ns, VDD,
+ 1292276.000000ns, VDD,
+ 1292276.100000ns, VSS,
+ 1292396.100000ns, VSS,
+ 1292396.200000ns, VDD,
+ 1292636.300000ns, VDD,
+ 1292636.400000ns, VSS,
+ 1292756.400000ns, VSS,
+ 1292756.500000ns, VDD,
+ 1293356.900000ns, VDD,
+ 1293357.000000ns, VSS,
+ 1294317.700000ns, VSS,
+ 1294317.800000ns, VDD,
+ 1295038.300000ns, VDD,
+ 1295038.400000ns, VSS,
+ 1295158.400000ns, VSS,
+ 1295158.500000ns, VDD,
+ 1296359.400000ns, VDD,
+ 1296359.500000ns, VSS,
+ 1296479.500000ns, VSS,
+ 1296479.600000ns, VDD,
+ 1296719.700000ns, VDD,
+ 1296719.800000ns, VSS,
+ 1297320.200000ns, VSS,
+ 1297320.300000ns, VDD,
+ 1297440.300000ns, VDD,
+ 1297440.400000ns, VSS,
+ 1297800.600000ns, VSS,
+ 1297800.700000ns, VDD,
+ 1297920.700000ns, VDD,
+ 1297920.800000ns, VSS,
+ 1298401.100000ns, VSS,
+ 1298401.200000ns, VDD,
+ 1298521.200000ns, VDD,
+ 1298521.300000ns, VSS,
+ 1299482.000000ns, VSS,
+ 1299482.100000ns, VDD,
+ 1300082.500000ns, VDD,
+ 1300082.600000ns, VSS,
+ 1301884.000000ns, VSS,
+ 1301884.100000ns, VDD,
+ 1302244.300000ns, VDD,
+ 1302244.400000ns, VSS,
+ 1302484.500000ns, VSS,
+ 1302484.600000ns, VDD,
+ 1302844.800000ns, VDD,
+ 1302844.900000ns, VSS,
+ 1302964.900000ns, VSS,
+ 1302965.000000ns, VDD,
+ 1303445.300000ns, VDD,
+ 1303445.400000ns, VSS,
+ 1303565.400000ns, VSS,
+ 1303565.500000ns, VDD,
+ 1303805.600000ns, VDD,
+ 1303805.700000ns, VSS,
+ 1303925.700000ns, VSS,
+ 1303925.800000ns, VDD,
+ 1304406.100000ns, VDD,
+ 1304406.200000ns, VSS,
+ 1304526.200000ns, VSS,
+ 1304526.300000ns, VDD,
+ 1304886.500000ns, VDD,
+ 1304886.600000ns, VSS,
+ 1305727.200000ns, VSS,
+ 1305727.300000ns, VDD,
+ 1305847.300000ns, VDD,
+ 1305847.400000ns, VSS,
+ 1306087.500000ns, VSS,
+ 1306087.600000ns, VDD,
+ 1306207.600000ns, VDD,
+ 1306207.700000ns, VSS,
+ 1307048.300000ns, VSS,
+ 1307048.400000ns, VDD,
+ 1307648.800000ns, VDD,
+ 1307648.900000ns, VSS,
+ 1307768.900000ns, VSS,
+ 1307769.000000ns, VDD,
+ 1308009.100000ns, VDD,
+ 1308009.200000ns, VSS,
+ 1308369.400000ns, VSS,
+ 1308369.500000ns, VDD,
+ 1308849.800000ns, VDD,
+ 1308849.900000ns, VSS,
+ 1308969.900000ns, VSS,
+ 1308970.000000ns, VDD,
+ 1309450.300000ns, VDD,
+ 1309450.400000ns, VSS,
+ 1309570.400000ns, VSS,
+ 1309570.500000ns, VDD,
+ 1309690.500000ns, VDD,
+ 1309690.600000ns, VSS,
+ 1310291.000000ns, VSS,
+ 1310291.100000ns, VDD,
+ 1311011.600000ns, VDD,
+ 1311011.700000ns, VSS,
+ 1311492.000000ns, VSS,
+ 1311492.100000ns, VDD,
+ 1312212.600000ns, VDD,
+ 1312212.700000ns, VSS,
+ 1312332.700000ns, VSS,
+ 1312332.800000ns, VDD,
+ 1312933.200000ns, VDD,
+ 1312933.300000ns, VSS,
+ 1313053.300000ns, VSS,
+ 1313053.400000ns, VDD,
+ 1313773.900000ns, VDD,
+ 1313774.000000ns, VSS,
+ 1313894.000000ns, VSS,
+ 1313894.100000ns, VDD,
+ 1314134.200000ns, VDD,
+ 1314134.300000ns, VSS,
+ 1314494.500000ns, VSS,
+ 1314494.600000ns, VDD,
+ 1314614.600000ns, VDD,
+ 1314614.700000ns, VSS,
+ 1314734.700000ns, VSS,
+ 1314734.800000ns, VDD,
+ 1315095.000000ns, VDD,
+ 1315095.100000ns, VSS,
+ 1315455.300000ns, VSS,
+ 1315455.400000ns, VDD,
+ 1315935.700000ns, VDD,
+ 1315935.800000ns, VSS,
+ 1316055.800000ns, VSS,
+ 1316055.900000ns, VDD,
+ 1317256.800000ns, VDD,
+ 1317256.900000ns, VSS,
+ 1318577.900000ns, VSS,
+ 1318578.000000ns, VDD,
+ 1319178.400000ns, VDD,
+ 1319178.500000ns, VSS,
+ 1320019.100000ns, VSS,
+ 1320019.200000ns, VDD,
+ 1320139.200000ns, VDD,
+ 1320139.300000ns, VSS,
+ 1320859.800000ns, VSS,
+ 1320859.900000ns, VDD,
+ 1321580.400000ns, VDD,
+ 1321580.500000ns, VSS,
+ 1321940.700000ns, VSS,
+ 1321940.800000ns, VDD,
+ 1322901.500000ns, VDD,
+ 1322901.600000ns, VSS,
+ 1323261.800000ns, VSS,
+ 1323261.900000ns, VDD,
+ 1323982.400000ns, VDD,
+ 1323982.500000ns, VSS,
+ 1324462.800000ns, VSS,
+ 1324462.900000ns, VDD,
+ 1325063.300000ns, VDD,
+ 1325063.400000ns, VSS,
+ 1325303.500000ns, VSS,
+ 1325303.600000ns, VDD,
+ 1325663.800000ns, VDD,
+ 1325663.900000ns, VSS,
+ 1325904.000000ns, VSS,
+ 1325904.100000ns, VDD,
+ 1326024.100000ns, VDD,
+ 1326024.200000ns, VSS,
+ 1327225.100000ns, VSS,
+ 1327225.200000ns, VDD,
+ 1327705.500000ns, VDD,
+ 1327705.600000ns, VSS,
+ 1328185.900000ns, VSS,
+ 1328186.000000ns, VDD,
+ 1328666.300000ns, VDD,
+ 1328666.400000ns, VSS,
+ 1329987.400000ns, VSS,
+ 1329987.500000ns, VDD,
+ 1330227.600000ns, VDD,
+ 1330227.700000ns, VSS,
+ 1330467.800000ns, VSS,
+ 1330467.900000ns, VDD,
+ 1330828.100000ns, VDD,
+ 1330828.200000ns, VSS,
+ 1331428.600000ns, VSS,
+ 1331428.700000ns, VDD,
+ 1331548.700000ns, VDD,
+ 1331548.800000ns, VSS,
+ 1331909.000000ns, VSS,
+ 1331909.100000ns, VDD,
+ 1332269.300000ns, VDD,
+ 1332269.400000ns, VSS,
+ 1332509.500000ns, VSS,
+ 1332509.600000ns, VDD,
+ 1333110.000000ns, VDD,
+ 1333110.100000ns, VSS,
+ 1333710.500000ns, VSS,
+ 1333710.600000ns, VDD,
+ 1334190.900000ns, VDD,
+ 1334191.000000ns, VSS,
+ 1334311.000000ns, VSS,
+ 1334311.100000ns, VDD,
+ 1334551.200000ns, VDD,
+ 1334551.300000ns, VSS,
+ 1334911.500000ns, VSS,
+ 1334911.600000ns, VDD,
+ 1335031.600000ns, VDD,
+ 1335031.700000ns, VSS,
+ 1335271.800000ns, VSS,
+ 1335271.900000ns, VDD,
+ 1336352.700000ns, VDD,
+ 1336352.800000ns, VSS,
+ 1337313.500000ns, VSS,
+ 1337313.600000ns, VDD,
+ 1337553.700000ns, VDD,
+ 1337553.800000ns, VSS,
+ 1337673.800000ns, VSS,
+ 1337673.900000ns, VDD,
+ 1338034.100000ns, VDD,
+ 1338034.200000ns, VSS,
+ 1338634.600000ns, VSS,
+ 1338634.700000ns, VDD,
+ 1339235.100000ns, VDD,
+ 1339235.200000ns, VSS,
+ 1339475.300000ns, VSS,
+ 1339475.400000ns, VDD,
+ 1339595.400000ns, VDD,
+ 1339595.500000ns, VSS,
+ 1340195.900000ns, VSS,
+ 1340196.000000ns, VDD,
+ 1340436.100000ns, VDD,
+ 1340436.200000ns, VSS,
+ 1340556.200000ns, VSS,
+ 1340556.300000ns, VDD,
+ 1340796.400000ns, VDD,
+ 1340796.500000ns, VSS,
+ 1342117.500000ns, VSS,
+ 1342117.600000ns, VDD,
+ 1342357.700000ns, VDD,
+ 1342357.800000ns, VSS,
+ 1342718.000000ns, VSS,
+ 1342718.100000ns, VDD,
+ 1342838.100000ns, VDD,
+ 1342838.200000ns, VSS,
+ 1343678.800000ns, VSS,
+ 1343678.900000ns, VDD,
+ 1344159.200000ns, VDD,
+ 1344159.300000ns, VSS,
+ 1344519.500000ns, VSS,
+ 1344519.600000ns, VDD,
+ 1344879.800000ns, VDD,
+ 1344879.900000ns, VSS,
+ 1344999.900000ns, VSS,
+ 1345000.000000ns, VDD,
+ 1345360.200000ns, VDD,
+ 1345360.300000ns, VSS,
+ 1345480.300000ns, VSS,
+ 1345480.400000ns, VDD,
+ 1345960.700000ns, VDD,
+ 1345960.800000ns, VSS,
+ 1346441.100000ns, VSS,
+ 1346441.200000ns, VDD,
+ 1347522.000000ns, VDD,
+ 1347522.100000ns, VSS,
+ 1347762.200000ns, VSS,
+ 1347762.300000ns, VDD,
+ 1348362.700000ns, VDD,
+ 1348362.800000ns, VSS,
+ 1349203.400000ns, VSS,
+ 1349203.500000ns, VDD,
+ 1349443.600000ns, VDD,
+ 1349443.700000ns, VSS,
+ 1349563.700000ns, VSS,
+ 1349563.800000ns, VDD,
+ 1349924.000000ns, VDD,
+ 1349924.100000ns, VSS,
+ 1350044.100000ns, VSS,
+ 1350044.200000ns, VDD,
+ 1350284.300000ns, VDD,
+ 1350284.400000ns, VSS,
+ 1350404.400000ns, VSS,
+ 1350404.500000ns, VDD,
+ 1350764.700000ns, VDD,
+ 1350764.800000ns, VSS,
+ 1351125.000000ns, VSS,
+ 1351125.100000ns, VDD,
+ 1351365.200000ns, VDD,
+ 1351365.300000ns, VSS,
+ 1351605.400000ns, VSS,
+ 1351605.500000ns, VDD,
+ 1351965.700000ns, VDD,
+ 1351965.800000ns, VSS,
+ 1352326.000000ns, VSS,
+ 1352326.100000ns, VDD,
+ 1353406.900000ns, VDD,
+ 1353407.000000ns, VSS,
+ 1353887.300000ns, VSS,
+ 1353887.400000ns, VDD,
+ 1354367.700000ns, VDD,
+ 1354367.800000ns, VSS,
+ 1354487.800000ns, VSS,
+ 1354487.900000ns, VDD,
+ 1354728.000000ns, VDD,
+ 1354728.100000ns, VSS,
+ 1355929.000000ns, VSS,
+ 1355929.100000ns, VDD,
+ 1356049.100000ns, VDD,
+ 1356049.200000ns, VSS,
+ 1356409.400000ns, VSS,
+ 1356409.500000ns, VDD,
+ 1356889.800000ns, VDD,
+ 1356889.900000ns, VSS,
+ 1357250.100000ns, VSS,
+ 1357250.200000ns, VDD,
+ 1357490.300000ns, VDD,
+ 1357490.400000ns, VSS,
+ 1357610.400000ns, VSS,
+ 1357610.500000ns, VDD,
+ 1358331.000000ns, VDD,
+ 1358331.100000ns, VSS,
+ 1358451.100000ns, VSS,
+ 1358451.200000ns, VDD,
+ 1359051.600000ns, VDD,
+ 1359051.700000ns, VSS,
+ 1359411.900000ns, VSS,
+ 1359412.000000ns, VDD,
+ 1359532.000000ns, VDD,
+ 1359532.100000ns, VSS,
+ 1359652.100000ns, VSS,
+ 1359652.200000ns, VDD,
+ 1359892.300000ns, VDD,
+ 1359892.400000ns, VSS,
+ 1360132.500000ns, VSS,
+ 1360132.600000ns, VDD,
+ 1360252.600000ns, VDD,
+ 1360252.700000ns, VSS,
+ 1361333.500000ns, VSS,
+ 1361333.600000ns, VDD,
+ 1361693.800000ns, VDD,
+ 1361693.900000ns, VSS,
+ 1361813.900000ns, VSS,
+ 1361814.000000ns, VDD,
+ 1362174.200000ns, VDD,
+ 1362174.300000ns, VSS,
+ 1362294.300000ns, VSS,
+ 1362294.400000ns, VDD,
+ 1362534.500000ns, VDD,
+ 1362534.600000ns, VSS,
+ 1362894.800000ns, VSS,
+ 1362894.900000ns, VDD,
+ 1363375.200000ns, VDD,
+ 1363375.300000ns, VSS,
+ 1363735.500000ns, VSS,
+ 1363735.600000ns, VDD,
+ 1363975.700000ns, VDD,
+ 1363975.800000ns, VSS,
+ 1364456.100000ns, VSS,
+ 1364456.200000ns, VDD,
+ 1364696.300000ns, VDD,
+ 1364696.400000ns, VSS,
+ 1364816.400000ns, VSS,
+ 1364816.500000ns, VDD,
+ 1365176.700000ns, VDD,
+ 1365176.800000ns, VSS,
+ 1365296.800000ns, VSS,
+ 1365296.900000ns, VDD,
+ 1366017.400000ns, VDD,
+ 1366017.500000ns, VSS,
+ 1366257.600000ns, VSS,
+ 1366257.700000ns, VDD,
+ 1366738.000000ns, VDD,
+ 1366738.100000ns, VSS,
+ 1367098.300000ns, VSS,
+ 1367098.400000ns, VDD,
+ 1367578.700000ns, VDD,
+ 1367578.800000ns, VSS,
+ 1367818.900000ns, VSS,
+ 1367819.000000ns, VDD,
+ 1368419.400000ns, VDD,
+ 1368419.500000ns, VSS,
+ 1368539.500000ns, VSS,
+ 1368539.600000ns, VDD,
+ 1369140.000000ns, VDD,
+ 1369140.100000ns, VSS,
+ 1369620.400000ns, VSS,
+ 1369620.500000ns, VDD,
+ 1369740.500000ns, VDD,
+ 1369740.600000ns, VSS,
+ 1370100.800000ns, VSS,
+ 1370100.900000ns, VDD,
+ 1370581.200000ns, VDD,
+ 1370581.300000ns, VSS,
+ 1370701.300000ns, VSS,
+ 1370701.400000ns, VDD,
+ 1370821.400000ns, VDD,
+ 1370821.500000ns, VSS,
+ 1370941.500000ns, VSS,
+ 1370941.600000ns, VDD,
+ 1371421.900000ns, VDD,
+ 1371422.000000ns, VSS,
+ 1371782.200000ns, VSS,
+ 1371782.300000ns, VDD,
+ 1372142.500000ns, VDD,
+ 1372142.600000ns, VSS,
+ 1372863.100000ns, VSS,
+ 1372863.200000ns, VDD,
+ 1372983.200000ns, VDD,
+ 1372983.300000ns, VSS,
+ 1373463.600000ns, VSS,
+ 1373463.700000ns, VDD,
+ 1374304.300000ns, VDD,
+ 1374304.400000ns, VSS,
+ 1374424.400000ns, VSS,
+ 1374424.500000ns, VDD,
+ 1374904.800000ns, VDD,
+ 1374904.900000ns, VSS,
+ 1375505.300000ns, VSS,
+ 1375505.400000ns, VDD,
+ 1375985.700000ns, VDD,
+ 1375985.800000ns, VSS,
+ 1376586.200000ns, VSS,
+ 1376586.300000ns, VDD,
+ 1376706.300000ns, VDD,
+ 1376706.400000ns, VSS,
+ 1377186.700000ns, VSS,
+ 1377186.800000ns, VDD,
+ 1377426.900000ns, VDD,
+ 1377427.000000ns, VSS,
+ 1377787.200000ns, VSS,
+ 1377787.300000ns, VDD,
+ 1378027.400000ns, VDD,
+ 1378027.500000ns, VSS,
+ 1378387.700000ns, VSS,
+ 1378387.800000ns, VDD,
+ 1379708.800000ns, VDD,
+ 1379708.900000ns, VSS,
+ 1380069.100000ns, VSS,
+ 1380069.200000ns, VDD,
+ 1380549.500000ns, VDD,
+ 1380549.600000ns, VSS,
+ 1380789.700000ns, VSS,
+ 1380789.800000ns, VDD,
+ 1380909.800000ns, VDD,
+ 1380909.900000ns, VSS,
+ 1381390.200000ns, VSS,
+ 1381390.300000ns, VDD,
+ 1381630.400000ns, VDD,
+ 1381630.500000ns, VSS,
+ 1381990.700000ns, VSS,
+ 1381990.800000ns, VDD,
+ 1382351.000000ns, VDD,
+ 1382351.100000ns, VSS,
+ 1382471.100000ns, VSS,
+ 1382471.200000ns, VDD,
+ 1382831.400000ns, VDD,
+ 1382831.500000ns, VSS,
+ 1382951.500000ns, VSS,
+ 1382951.600000ns, VDD,
+ 1383431.900000ns, VDD,
+ 1383432.000000ns, VSS,
+ 1384032.400000ns, VSS,
+ 1384032.500000ns, VDD,
+ 1384152.500000ns, VDD,
+ 1384152.600000ns, VSS,
+ 1384272.600000ns, VSS,
+ 1384272.700000ns, VDD,
+ 1384993.200000ns, VDD,
+ 1384993.300000ns, VSS,
+ 1385233.400000ns, VSS,
+ 1385233.500000ns, VDD,
+ 1385353.500000ns, VDD,
+ 1385353.600000ns, VSS,
+ 1385833.900000ns, VSS,
+ 1385834.000000ns, VDD,
+ 1386074.100000ns, VDD,
+ 1386074.200000ns, VSS,
+ 1386434.400000ns, VSS,
+ 1386434.500000ns, VDD,
+ 1386554.500000ns, VDD,
+ 1386554.600000ns, VSS,
+ 1387635.400000ns, VSS,
+ 1387635.500000ns, VDD,
+ 1388235.900000ns, VDD,
+ 1388236.000000ns, VSS,
+ 1388356.000000ns, VSS,
+ 1388356.100000ns, VDD,
+ 1388716.300000ns, VDD,
+ 1388716.400000ns, VSS,
+ 1389196.700000ns, VSS,
+ 1389196.800000ns, VDD,
+ 1389917.300000ns, VDD,
+ 1389917.400000ns, VSS,
+ 1390758.000000ns, VSS,
+ 1390758.100000ns, VDD,
+ 1390998.200000ns, VDD,
+ 1390998.300000ns, VSS,
+ 1391238.400000ns, VSS,
+ 1391238.500000ns, VDD,
+ 1391358.500000ns, VDD,
+ 1391358.600000ns, VSS,
+ 1391718.800000ns, VSS,
+ 1391718.900000ns, VDD,
+ 1391959.000000ns, VDD,
+ 1391959.100000ns, VSS,
+ 1392439.400000ns, VSS,
+ 1392439.500000ns, VDD,
+ 1392679.600000ns, VDD,
+ 1392679.700000ns, VSS,
+ 1392919.800000ns, VSS,
+ 1392919.900000ns, VDD,
+ 1393160.000000ns, VDD,
+ 1393160.100000ns, VSS,
+ 1393400.200000ns, VSS,
+ 1393400.300000ns, VDD,
+ 1393520.300000ns, VDD,
+ 1393520.400000ns, VSS,
+ 1393880.600000ns, VSS,
+ 1393880.700000ns, VDD,
+ 1394961.500000ns, VDD,
+ 1394961.600000ns, VSS,
+ 1396522.800000ns, VSS,
+ 1396522.900000ns, VDD,
+ 1396763.000000ns, VDD,
+ 1396763.100000ns, VSS,
+ 1397003.200000ns, VSS,
+ 1397003.300000ns, VDD,
+ 1397243.400000ns, VDD,
+ 1397243.500000ns, VSS,
+ 1398684.600000ns, VSS,
+ 1398684.700000ns, VDD,
+ 1399285.100000ns, VDD,
+ 1399285.200000ns, VSS,
+ 1399765.500000ns, VSS,
+ 1399765.600000ns, VDD,
+ 1400366.000000ns, VDD,
+ 1400366.100000ns, VSS,
+ 1400846.400000ns, VSS,
+ 1400846.500000ns, VDD,
+ 1401927.300000ns, VDD,
+ 1401927.400000ns, VSS,
+ 1402167.500000ns, VSS,
+ 1402167.600000ns, VDD,
+ 1403728.800000ns, VDD,
+ 1403728.900000ns, VSS,
+ 1403969.000000ns, VSS,
+ 1403969.100000ns, VDD,
+ 1404209.200000ns, VDD,
+ 1404209.300000ns, VSS,
+ 1404689.600000ns, VSS,
+ 1404689.700000ns, VDD,
+ 1404929.800000ns, VDD,
+ 1404929.900000ns, VSS,
+ 1405290.100000ns, VSS,
+ 1405290.200000ns, VDD,
+ 1405650.400000ns, VDD,
+ 1405650.500000ns, VSS,
+ 1405770.500000ns, VSS,
+ 1405770.600000ns, VDD,
+ 1406250.900000ns, VDD,
+ 1406251.000000ns, VSS,
+ 1406371.000000ns, VSS,
+ 1406371.100000ns, VDD,
+ 1406731.300000ns, VDD,
+ 1406731.400000ns, VSS,
+ 1407211.700000ns, VSS,
+ 1407211.800000ns, VDD,
+ 1407451.900000ns, VDD,
+ 1407452.000000ns, VSS,
+ 1408052.400000ns, VSS,
+ 1408052.500000ns, VDD,
+ 1408893.100000ns, VDD,
+ 1408893.200000ns, VSS,
+ 1409013.200000ns, VSS,
+ 1409013.300000ns, VDD,
+ 1409253.400000ns, VDD,
+ 1409253.500000ns, VSS,
+ 1409613.700000ns, VSS,
+ 1409613.800000ns, VDD,
+ 1410214.200000ns, VDD,
+ 1410214.300000ns, VSS,
+ 1410934.800000ns, VSS,
+ 1410934.900000ns, VDD,
+ 1411175.000000ns, VDD,
+ 1411175.100000ns, VSS,
+ 1411535.300000ns, VSS,
+ 1411535.400000ns, VDD,
+ 1411655.400000ns, VDD,
+ 1411655.500000ns, VSS,
+ 1411895.600000ns, VSS,
+ 1411895.700000ns, VDD,
+ 1412135.800000ns, VDD,
+ 1412135.900000ns, VSS,
+ 1412496.100000ns, VSS,
+ 1412496.200000ns, VDD,
+ 1412616.200000ns, VDD,
+ 1412616.300000ns, VSS,
+ 1413577.000000ns, VSS,
+ 1413577.100000ns, VDD,
+ 1414898.100000ns, VDD,
+ 1414898.200000ns, VSS,
+ 1415258.400000ns, VSS,
+ 1415258.500000ns, VDD,
+ 1415858.900000ns, VDD,
+ 1415859.000000ns, VSS,
+ 1416219.200000ns, VSS,
+ 1416219.300000ns, VDD,
+ 1416339.300000ns, VDD,
+ 1416339.400000ns, VSS,
+ 1416699.600000ns, VSS,
+ 1416699.700000ns, VDD,
+ 1416939.800000ns, VDD,
+ 1416939.900000ns, VSS,
+ 1417059.900000ns, VSS,
+ 1417060.000000ns, VDD,
+ 1417900.600000ns, VDD,
+ 1417900.700000ns, VSS,
+ 1418621.200000ns, VSS,
+ 1418621.300000ns, VDD,
+ 1419101.600000ns, VDD,
+ 1419101.700000ns, VSS,
+ 1419461.900000ns, VSS,
+ 1419462.000000ns, VDD,
+ 1419582.000000ns, VDD,
+ 1419582.100000ns, VSS,
+ 1420422.700000ns, VSS,
+ 1420422.800000ns, VDD,
+ 1420783.000000ns, VDD,
+ 1420783.100000ns, VSS,
+ 1421143.300000ns, VSS,
+ 1421143.400000ns, VDD,
+ 1422224.200000ns, VDD,
+ 1422224.300000ns, VSS,
+ 1422464.400000ns, VSS,
+ 1422464.500000ns, VDD,
+ 1422584.500000ns, VDD,
+ 1422584.600000ns, VSS,
+ 1422824.700000ns, VSS,
+ 1422824.800000ns, VDD,
+ 1422944.800000ns, VDD,
+ 1422944.900000ns, VSS,
+ 1423545.300000ns, VSS,
+ 1423545.400000ns, VDD,
+ 1423785.500000ns, VDD,
+ 1423785.600000ns, VSS,
+ 1424025.700000ns, VSS,
+ 1424025.800000ns, VDD,
+ 1424145.800000ns, VDD,
+ 1424145.900000ns, VSS,
+ 1424506.100000ns, VSS,
+ 1424506.200000ns, VDD,
+ 1424626.200000ns, VDD,
+ 1424626.300000ns, VSS,
+ 1425106.600000ns, VSS,
+ 1425106.700000ns, VDD,
+ 1425947.300000ns, VDD,
+ 1425947.400000ns, VSS,
+ 1426067.400000ns, VSS,
+ 1426067.500000ns, VDD,
+ 1426307.600000ns, VDD,
+ 1426307.700000ns, VSS,
+ 1427748.800000ns, VSS,
+ 1427748.900000ns, VDD,
+ 1427989.000000ns, VDD,
+ 1427989.100000ns, VSS,
+ 1428109.100000ns, VSS,
+ 1428109.200000ns, VDD,
+ 1428229.200000ns, VDD,
+ 1428229.300000ns, VSS,
+ 1428949.800000ns, VSS,
+ 1428949.900000ns, VDD,
+ 1429069.900000ns, VDD,
+ 1429070.000000ns, VSS,
+ 1429790.500000ns, VSS,
+ 1429790.600000ns, VDD,
+ 1430030.700000ns, VDD,
+ 1430030.800000ns, VSS,
+ 1430270.900000ns, VSS,
+ 1430271.000000ns, VDD,
+ 1430991.500000ns, VDD,
+ 1430991.600000ns, VSS,
+ 1431111.600000ns, VSS,
+ 1431111.700000ns, VDD,
+ 1431231.700000ns, VDD,
+ 1431231.800000ns, VSS,
+ 1432552.800000ns, VSS,
+ 1432552.900000ns, VDD,
+ 1433273.400000ns, VDD,
+ 1433273.500000ns, VSS,
+ 1433393.500000ns, VSS,
+ 1433393.600000ns, VDD,
+ 1434234.200000ns, VDD,
+ 1434234.300000ns, VSS,
+ 1434354.300000ns, VSS,
+ 1434354.400000ns, VDD,
+ 1434594.500000ns, VDD,
+ 1434594.600000ns, VSS,
+ 1434954.800000ns, VSS,
+ 1434954.900000ns, VDD,
+ 1435195.000000ns, VDD,
+ 1435195.100000ns, VSS,
+ 1435675.400000ns, VSS,
+ 1435675.500000ns, VDD,
+ 1436035.700000ns, VDD,
+ 1436035.800000ns, VSS,
+ 1436275.900000ns, VSS,
+ 1436276.000000ns, VDD,
+ 1437356.800000ns, VDD,
+ 1437356.900000ns, VSS,
+ 1437717.100000ns, VSS,
+ 1437717.200000ns, VDD,
+ 1437957.300000ns, VDD,
+ 1437957.400000ns, VSS,
+ 1438077.400000ns, VSS,
+ 1438077.500000ns, VDD,
+ 1438317.600000ns, VDD,
+ 1438317.700000ns, VSS,
+ 1438437.700000ns, VSS,
+ 1438437.800000ns, VDD,
+ 1438798.000000ns, VDD,
+ 1438798.100000ns, VSS,
+ 1439038.200000ns, VSS,
+ 1439038.300000ns, VDD,
+ 1439158.300000ns, VDD,
+ 1439158.400000ns, VSS,
+ 1439518.600000ns, VSS,
+ 1439518.700000ns, VDD,
+ 1440119.100000ns, VDD,
+ 1440119.200000ns, VSS,
+ 1440359.300000ns, VSS,
+ 1440359.400000ns, VDD,
+ 1440839.700000ns, VDD,
+ 1440839.800000ns, VSS,
+ 1441079.900000ns, VSS,
+ 1441080.000000ns, VDD,
+ 1441320.100000ns, VDD,
+ 1441320.200000ns, VSS,
+ 1441440.200000ns, VSS,
+ 1441440.300000ns, VDD,
+ 1441560.300000ns, VDD,
+ 1441560.400000ns, VSS,
+ 1441680.400000ns, VSS,
+ 1441680.500000ns, VDD,
+ 1442280.900000ns, VDD,
+ 1442281.000000ns, VSS,
+ 1442401.000000ns, VSS,
+ 1442401.100000ns, VDD,
+ 1442641.200000ns, VDD,
+ 1442641.300000ns, VSS,
+ 1442761.300000ns, VSS,
+ 1442761.400000ns, VDD,
+ 1443001.500000ns, VDD,
+ 1443001.600000ns, VSS,
+ 1443481.900000ns, VSS,
+ 1443482.000000ns, VDD,
+ 1444082.400000ns, VDD,
+ 1444082.500000ns, VSS,
+ 1444322.600000ns, VSS,
+ 1444322.700000ns, VDD,
+ 1444923.100000ns, VDD,
+ 1444923.200000ns, VSS,
+ 1445043.200000ns, VSS,
+ 1445043.300000ns, VDD,
+ 1445403.500000ns, VDD,
+ 1445403.600000ns, VSS,
+ 1445523.600000ns, VSS,
+ 1445523.700000ns, VDD,
+ 1446364.300000ns, VDD,
+ 1446364.400000ns, VSS,
+ 1446484.400000ns, VSS,
+ 1446484.500000ns, VDD,
+ 1446844.700000ns, VDD,
+ 1446844.800000ns, VSS,
+ 1446964.800000ns, VSS,
+ 1446964.900000ns, VDD,
+ 1447205.000000ns, VDD,
+ 1447205.100000ns, VSS,
+ 1447325.100000ns, VSS,
+ 1447325.200000ns, VDD,
+ 1447565.300000ns, VDD,
+ 1447565.400000ns, VSS,
+ 1447925.600000ns, VSS,
+ 1447925.700000ns, VDD,
+ 1448045.700000ns, VDD,
+ 1448045.800000ns, VSS,
+ 1448646.200000ns, VSS,
+ 1448646.300000ns, VDD,
+ 1448886.400000ns, VDD,
+ 1448886.500000ns, VSS,
+ 1449006.500000ns, VSS,
+ 1449006.600000ns, VDD,
+ 1449126.600000ns, VDD,
+ 1449126.700000ns, VSS,
+ 1449366.800000ns, VSS,
+ 1449366.900000ns, VDD,
+ 1449847.200000ns, VDD,
+ 1449847.300000ns, VSS,
+ 1449967.300000ns, VSS,
+ 1449967.400000ns, VDD,
+ 1450447.700000ns, VDD,
+ 1450447.800000ns, VSS,
+ 1451648.700000ns, VSS,
+ 1451648.800000ns, VDD,
+ 1452129.100000ns, VDD,
+ 1452129.200000ns, VSS,
+ 1452489.400000ns, VSS,
+ 1452489.500000ns, VDD,
+ 1453330.100000ns, VDD,
+ 1453330.200000ns, VSS,
+ 1453690.400000ns, VSS,
+ 1453690.500000ns, VDD,
+ 1453810.500000ns, VDD,
+ 1453810.600000ns, VSS,
+ 1454531.100000ns, VSS,
+ 1454531.200000ns, VDD,
+ 1455011.500000ns, VDD,
+ 1455011.600000ns, VSS,
+ 1455251.700000ns, VSS,
+ 1455251.800000ns, VDD,
+ 1455371.800000ns, VDD,
+ 1455371.900000ns, VSS,
+ 1455491.900000ns, VSS,
+ 1455492.000000ns, VDD,
+ 1455612.000000ns, VDD,
+ 1455612.100000ns, VSS,
+ 1455732.100000ns, VSS,
+ 1455732.200000ns, VDD,
+ 1456212.500000ns, VDD,
+ 1456212.600000ns, VSS,
+ 1456332.600000ns, VSS,
+ 1456332.700000ns, VDD,
+ 1456572.800000ns, VDD,
+ 1456572.900000ns, VSS,
+ 1456692.900000ns, VSS,
+ 1456693.000000ns, VDD,
+ 1456933.100000ns, VDD,
+ 1456933.200000ns, VSS,
+ 1457053.200000ns, VSS,
+ 1457053.300000ns, VDD,
+ 1457413.500000ns, VDD,
+ 1457413.600000ns, VSS,
+ 1458254.200000ns, VSS,
+ 1458254.300000ns, VDD,
+ 1458374.300000ns, VDD,
+ 1458374.400000ns, VSS,
+ 1458614.500000ns, VSS,
+ 1458614.600000ns, VDD,
+ 1458734.600000ns, VDD,
+ 1458734.700000ns, VSS,
+ 1459335.100000ns, VSS,
+ 1459335.200000ns, VDD,
+ 1459695.400000ns, VDD,
+ 1459695.500000ns, VSS,
+ 1460175.800000ns, VSS,
+ 1460175.900000ns, VDD,
+ 1460295.900000ns, VDD,
+ 1460296.000000ns, VSS,
+ 1460536.100000ns, VSS,
+ 1460536.200000ns, VDD,
+ 1460656.200000ns, VDD,
+ 1460656.300000ns, VSS,
+ 1461256.700000ns, VSS,
+ 1461256.800000ns, VDD,
+ 1461977.300000ns, VDD,
+ 1461977.400000ns, VSS,
+ 1462457.700000ns, VSS,
+ 1462457.800000ns, VDD,
+ 1462938.100000ns, VDD,
+ 1462938.200000ns, VSS,
+ 1463298.400000ns, VSS,
+ 1463298.500000ns, VDD,
+ 1464139.100000ns, VDD,
+ 1464139.200000ns, VSS,
+ 1464259.200000ns, VSS,
+ 1464259.300000ns, VDD,
+ 1465220.000000ns, VDD,
+ 1465220.100000ns, VSS,
+ 1465700.400000ns, VSS,
+ 1465700.500000ns, VDD,
+ 1466060.700000ns, VDD,
+ 1466060.800000ns, VSS,
+ 1466180.800000ns, VSS,
+ 1466180.900000ns, VDD,
+ 1466661.200000ns, VDD,
+ 1466661.300000ns, VSS,
+ 1466781.300000ns, VSS,
+ 1466781.400000ns, VDD,
+ 1467261.700000ns, VDD,
+ 1467261.800000ns, VSS,
+ 1468462.700000ns, VSS,
+ 1468462.800000ns, VDD,
+ 1468582.800000ns, VDD,
+ 1468582.900000ns, VSS,
+ 1469183.300000ns, VSS,
+ 1469183.400000ns, VDD,
+ 1469303.400000ns, VDD,
+ 1469303.500000ns, VSS,
+ 1469423.500000ns, VSS,
+ 1469423.600000ns, VDD,
+ 1469663.700000ns, VDD,
+ 1469663.800000ns, VSS,
+ 1469783.800000ns, VSS,
+ 1469783.900000ns, VDD,
+ 1470144.100000ns, VDD,
+ 1470144.200000ns, VSS,
+ 1470744.600000ns, VSS,
+ 1470744.700000ns, VDD,
+ 1471225.000000ns, VDD,
+ 1471225.100000ns, VSS,
+ 1471345.100000ns, VSS,
+ 1471345.200000ns, VDD,
+ 1471465.200000ns, VDD,
+ 1471465.300000ns, VSS,
+ 1471705.400000ns, VSS,
+ 1471705.500000ns, VDD,
+ 1471825.500000ns, VDD,
+ 1471825.600000ns, VSS,
+ 1472426.000000ns, VSS,
+ 1472426.100000ns, VDD,
+ 1473146.600000ns, VDD,
+ 1473146.700000ns, VSS,
+ 1474707.900000ns, VSS,
+ 1474708.000000ns, VDD,
+ 1474828.000000ns, VDD,
+ 1474828.100000ns, VSS,
+ 1475308.400000ns, VSS,
+ 1475308.500000ns, VDD,
+ 1475668.700000ns, VDD,
+ 1475668.800000ns, VSS,
+ 1476269.200000ns, VSS,
+ 1476269.300000ns, VDD,
+ 1476509.400000ns, VDD,
+ 1476509.500000ns, VSS,
+ 1476749.600000ns, VSS,
+ 1476749.700000ns, VDD,
+ 1476989.800000ns, VDD,
+ 1476989.900000ns, VSS,
+ 1477350.100000ns, VSS,
+ 1477350.200000ns, VDD,
+ 1477590.300000ns, VDD,
+ 1477590.400000ns, VSS,
+ 1478070.700000ns, VSS,
+ 1478070.800000ns, VDD,
+ 1478310.900000ns, VDD,
+ 1478311.000000ns, VSS,
+ 1478911.400000ns, VSS,
+ 1478911.500000ns, VDD,
+ 1479391.800000ns, VDD,
+ 1479391.900000ns, VSS,
+ 1479511.900000ns, VSS,
+ 1479512.000000ns, VDD,
+ 1479992.300000ns, VDD,
+ 1479992.400000ns, VSS,
+ 1480592.800000ns, VSS,
+ 1480592.900000ns, VDD,
+ 1481073.200000ns, VDD,
+ 1481073.300000ns, VSS,
+ 1481913.900000ns, VSS,
+ 1481914.000000ns, VDD,
+ 1482394.300000ns, VDD,
+ 1482394.400000ns, VSS,
+ 1482754.600000ns, VSS,
+ 1482754.700000ns, VDD,
+ 1483235.000000ns, VDD,
+ 1483235.100000ns, VSS,
+ 1483475.200000ns, VSS,
+ 1483475.300000ns, VDD,
+ 1483955.600000ns, VDD,
+ 1483955.700000ns, VSS,
+ 1484075.700000ns, VSS,
+ 1484075.800000ns, VDD,
+ 1484315.900000ns, VDD,
+ 1484316.000000ns, VSS,
+ 1484556.100000ns, VSS,
+ 1484556.200000ns, VDD,
+ 1484796.300000ns, VDD,
+ 1484796.400000ns, VSS,
+ 1485036.500000ns, VSS,
+ 1485036.600000ns, VDD,
+ 1485156.600000ns, VDD,
+ 1485156.700000ns, VSS,
+ 1485276.700000ns, VSS,
+ 1485276.800000ns, VDD,
+ 1485997.300000ns, VDD,
+ 1485997.400000ns, VSS,
+ 1486357.600000ns, VSS,
+ 1486357.700000ns, VDD,
+ 1486597.800000ns, VDD,
+ 1486597.900000ns, VSS,
+ 1486958.100000ns, VSS,
+ 1486958.200000ns, VDD,
+ 1487798.800000ns, VDD,
+ 1487798.900000ns, VSS,
+ 1488279.200000ns, VSS,
+ 1488279.300000ns, VDD,
+ 1488879.700000ns, VDD,
+ 1488879.800000ns, VSS,
+ 1489119.900000ns, VSS,
+ 1489120.000000ns, VDD,
+ 1489360.100000ns, VDD,
+ 1489360.200000ns, VSS,
+ 1489720.400000ns, VSS,
+ 1489720.500000ns, VDD,
+ 1489840.500000ns, VDD,
+ 1489840.600000ns, VSS,
+ 1489960.600000ns, VSS,
+ 1489960.700000ns, VDD,
+ 1490441.000000ns, VDD,
+ 1490441.100000ns, VSS,
+ 1490921.400000ns, VSS,
+ 1490921.500000ns, VDD,
+ 1491041.500000ns, VDD,
+ 1491041.600000ns, VSS,
+ 1491161.600000ns, VSS,
+ 1491161.700000ns, VDD,
+ 1491762.100000ns, VDD,
+ 1491762.200000ns, VSS,
+ 1491882.200000ns, VSS,
+ 1491882.300000ns, VDD,
+ 1492843.000000ns, VDD,
+ 1492843.100000ns, VSS,
+ 1492963.100000ns, VSS,
+ 1492963.200000ns, VDD,
+ 1493323.400000ns, VDD,
+ 1493323.500000ns, VSS,
+ 1493683.700000ns, VSS,
+ 1493683.800000ns, VDD,
+ 1493923.900000ns, VDD,
+ 1493924.000000ns, VSS,
+ 1494164.100000ns, VSS,
+ 1494164.200000ns, VDD,
+ 1494404.300000ns, VDD,
+ 1494404.400000ns, VSS,
+ 1495124.900000ns, VSS,
+ 1495125.000000ns, VDD,
+ 1495365.100000ns, VDD,
+ 1495365.200000ns, VSS,
+ 1495965.600000ns, VSS,
+ 1495965.700000ns, VDD,
+ 1496325.900000ns, VDD,
+ 1496326.000000ns, VSS,
+ 1496926.400000ns, VSS,
+ 1496926.500000ns, VDD,
+ 1498007.300000ns, VDD,
+ 1498007.400000ns, VSS,
+ 1499088.200000ns, VSS,
+ 1499088.300000ns, VDD,
+ 1499568.600000ns, VDD,
+ 1499568.700000ns, VSS,
+ 1500169.100000ns, VSS,
+ 1500169.200000ns, VDD,
+ 1500889.700000ns, VDD,
+ 1500889.800000ns, VSS,
+ 1501250.000000ns, VSS,
+ 1501250.100000ns, VDD,
+ 1501850.500000ns, VDD,
+ 1501850.600000ns, VSS,
+ 1501970.600000ns, VSS,
+ 1501970.700000ns, VDD,
+ 1502330.900000ns, VDD,
+ 1502331.000000ns, VSS,
+ 1502571.100000ns, VSS,
+ 1502571.200000ns, VDD,
+ 1503051.500000ns, VDD,
+ 1503051.600000ns, VSS,
+ 1503411.800000ns, VSS,
+ 1503411.900000ns, VDD,
+ 1504252.500000ns, VDD,
+ 1504252.600000ns, VSS,
+ 1504372.600000ns, VSS,
+ 1504372.700000ns, VDD,
+ 1505693.700000ns, VDD,
+ 1505693.800000ns, VSS,
+ 1506534.400000ns, VSS,
+ 1506534.500000ns, VDD,
+ 1506894.700000ns, VDD,
+ 1506894.800000ns, VSS,
+ 1507495.200000ns, VSS,
+ 1507495.300000ns, VDD,
+ 1508095.700000ns, VDD,
+ 1508095.800000ns, VSS,
+ 1508936.400000ns, VSS,
+ 1508936.500000ns, VDD,
+ 1510377.600000ns, VDD,
+ 1510377.700000ns, VSS,
+ 1510737.900000ns, VSS,
+ 1510738.000000ns, VDD,
+ 1511218.300000ns, VDD,
+ 1511218.400000ns, VSS,
+ 1511698.700000ns, VSS,
+ 1511698.800000ns, VDD,
+ 1511938.900000ns, VDD,
+ 1511939.000000ns, VSS,
+ 1512299.200000ns, VSS,
+ 1512299.300000ns, VDD,
+ 1512419.300000ns, VDD,
+ 1512419.400000ns, VSS,
+ 1513019.800000ns, VSS,
+ 1513019.900000ns, VDD,
+ 1514100.700000ns, VDD,
+ 1514100.800000ns, VSS,
+ 1514220.800000ns, VSS,
+ 1514220.900000ns, VDD,
+ 1514340.900000ns, VDD,
+ 1514341.000000ns, VSS,
+ 1514461.000000ns, VSS,
+ 1514461.100000ns, VDD,
+ 1514581.100000ns, VDD,
+ 1514581.200000ns, VSS,
+ 1515902.200000ns, VSS,
+ 1515902.300000ns, VDD,
+ 1516742.900000ns, VDD,
+ 1516743.000000ns, VSS,
+ 1516863.000000ns, VSS,
+ 1516863.100000ns, VDD,
+ 1517463.500000ns, VDD,
+ 1517463.600000ns, VSS,
+ 1519745.400000ns, VSS,
+ 1519745.500000ns, VDD,
+ 1519865.500000ns, VDD,
+ 1519865.600000ns, VSS,
+ 1520466.000000ns, VSS,
+ 1520466.100000ns, VDD,
+ 1520706.200000ns, VDD,
+ 1520706.300000ns, VSS,
+ 1521306.700000ns, VSS,
+ 1521306.800000ns, VDD,
+ 1522147.400000ns, VDD,
+ 1522147.500000ns, VSS,
+ 1522387.600000ns, VSS,
+ 1522387.700000ns, VDD,
+ 1523108.200000ns, VDD,
+ 1523108.300000ns, VSS,
+ 1523348.400000ns, VSS,
+ 1523348.500000ns, VDD,
+ 1523708.700000ns, VDD,
+ 1523708.800000ns, VSS,
+ 1523828.800000ns, VSS,
+ 1523828.900000ns, VDD,
+ 1524669.500000ns, VDD,
+ 1524669.600000ns, VSS,
+ 1524789.600000ns, VSS,
+ 1524789.700000ns, VDD,
+ 1525029.800000ns, VDD,
+ 1525029.900000ns, VSS,
+ 1525750.400000ns, VSS,
+ 1525750.500000ns, VDD,
+ 1526350.900000ns, VDD,
+ 1526351.000000ns, VSS,
+ 1526471.000000ns, VSS,
+ 1526471.100000ns, VDD,
+ 1526831.300000ns, VDD,
+ 1526831.400000ns, VSS,
+ 1526951.400000ns, VSS,
+ 1526951.500000ns, VDD,
+ 1527311.700000ns, VDD,
+ 1527311.800000ns, VSS,
+ 1527672.000000ns, VSS,
+ 1527672.100000ns, VDD,
+ 1527792.100000ns, VDD,
+ 1527792.200000ns, VSS,
+ 1528392.600000ns, VSS,
+ 1528392.700000ns, VDD,
+ 1529353.400000ns, VDD,
+ 1529353.500000ns, VSS,
+ 1529713.700000ns, VSS,
+ 1529713.800000ns, VDD,
+ 1530434.300000ns, VDD,
+ 1530434.400000ns, VSS,
+ 1530674.500000ns, VSS,
+ 1530674.600000ns, VDD,
+ 1530794.600000ns, VDD,
+ 1530794.700000ns, VSS,
+ 1531515.200000ns, VSS,
+ 1531515.300000ns, VDD,
+ 1531755.400000ns, VDD,
+ 1531755.500000ns, VSS,
+ 1531875.500000ns, VSS,
+ 1531875.600000ns, VDD,
+ 1532115.700000ns, VDD,
+ 1532115.800000ns, VSS,
+ 1532476.000000ns, VSS,
+ 1532476.100000ns, VDD,
+ 1532596.100000ns, VDD,
+ 1532596.200000ns, VSS,
+ 1532836.300000ns, VSS,
+ 1532836.400000ns, VDD,
+ 1533316.700000ns, VDD,
+ 1533316.800000ns, VSS,
+ 1533677.000000ns, VSS,
+ 1533677.100000ns, VDD,
+ 1534037.300000ns, VDD,
+ 1534037.400000ns, VSS,
+ 1534157.400000ns, VSS,
+ 1534157.500000ns, VDD,
+ 1534397.600000ns, VDD,
+ 1534397.700000ns, VSS,
+ 1534757.900000ns, VSS,
+ 1534758.000000ns, VDD,
+ 1535238.300000ns, VDD,
+ 1535238.400000ns, VSS,
+ 1535718.700000ns, VSS,
+ 1535718.800000ns, VDD,
+ 1535838.800000ns, VDD,
+ 1535838.900000ns, VSS,
+ 1536079.000000ns, VSS,
+ 1536079.100000ns, VDD,
+ 1536199.100000ns, VDD,
+ 1536199.200000ns, VSS,
+ 1537280.000000ns, VSS,
+ 1537280.100000ns, VDD,
+ 1537520.200000ns, VDD,
+ 1537520.300000ns, VSS,
+ 1537880.500000ns, VSS,
+ 1537880.600000ns, VDD,
+ 1538120.700000ns, VDD,
+ 1538120.800000ns, VSS,
+ 1538961.400000ns, VSS,
+ 1538961.500000ns, VDD,
+ 1539441.800000ns, VDD,
+ 1539441.900000ns, VSS,
+ 1540162.400000ns, VSS,
+ 1540162.500000ns, VDD,
+ 1540762.900000ns, VDD,
+ 1540763.000000ns, VSS,
+ 1541123.200000ns, VSS,
+ 1541123.300000ns, VDD,
+ 1541363.400000ns, VDD,
+ 1541363.500000ns, VSS,
+ 1541483.500000ns, VSS,
+ 1541483.600000ns, VDD,
+ 1541843.800000ns, VDD,
+ 1541843.900000ns, VSS,
+ 1542204.100000ns, VSS,
+ 1542204.200000ns, VDD,
+ 1542324.200000ns, VDD,
+ 1542324.300000ns, VSS,
+ 1542684.500000ns, VSS,
+ 1542684.600000ns, VDD,
+ 1543044.800000ns, VDD,
+ 1543044.900000ns, VSS,
+ 1543645.300000ns, VSS,
+ 1543645.400000ns, VDD,
+ 1543765.400000ns, VDD,
+ 1543765.500000ns, VSS,
+ 1544245.800000ns, VSS,
+ 1544245.900000ns, VDD,
+ 1544726.200000ns, VDD,
+ 1544726.300000ns, VSS,
+ 1544846.300000ns, VSS,
+ 1544846.400000ns, VDD,
+ 1545326.700000ns, VDD,
+ 1545326.800000ns, VSS,
+ 1545446.800000ns, VSS,
+ 1545446.900000ns, VDD,
+ 1545807.100000ns, VDD,
+ 1545807.200000ns, VSS,
+ 1545927.200000ns, VSS,
+ 1545927.300000ns, VDD,
+ 1546167.400000ns, VDD,
+ 1546167.500000ns, VSS,
+ 1546407.600000ns, VSS,
+ 1546407.700000ns, VDD,
+ 1546647.800000ns, VDD,
+ 1546647.900000ns, VSS,
+ 1546767.900000ns, VSS,
+ 1546768.000000ns, VDD,
+ 1547248.300000ns, VDD,
+ 1547248.400000ns, VSS,
+ 1548209.100000ns, VSS,
+ 1548209.200000ns, VDD,
+ 1548329.200000ns, VDD,
+ 1548329.300000ns, VSS,
+ 1548689.500000ns, VSS,
+ 1548689.600000ns, VDD,
+ 1548809.600000ns, VDD,
+ 1548809.700000ns, VSS,
+ 1549049.800000ns, VSS,
+ 1549049.900000ns, VDD,
+ 1549290.000000ns, VDD,
+ 1549290.100000ns, VSS,
+ 1549410.100000ns, VSS,
+ 1549410.200000ns, VDD,
+ 1549650.300000ns, VDD,
+ 1549650.400000ns, VSS,
+ 1549770.400000ns, VSS,
+ 1549770.500000ns, VDD
+)}


RD in_D 0 1.0
BD in_D 0 V={table(time,
+ 0.100000ns, VSS,
+ 240.200000ns, VSS,
+ 240.300000ns, VDD,
+ 1441.200000ns, VDD,
+ 1441.300000ns, VSS,
+ 1921.600000ns, VSS,
+ 1921.700000ns, VDD,
+ 2161.800000ns, VDD,
+ 2161.900000ns, VSS,
+ 2281.900000ns, VSS,
+ 2282.000000ns, VDD,
+ 2402.000000ns, VDD,
+ 2402.100000ns, VSS,
+ 2882.400000ns, VSS,
+ 2882.500000ns, VDD,
+ 4563.800000ns, VDD,
+ 4563.900000ns, VSS,
+ 4924.100000ns, VSS,
+ 4924.200000ns, VDD,
+ 6125.100000ns, VDD,
+ 6125.200000ns, VSS,
+ 6605.500000ns, VSS,
+ 6605.600000ns, VDD,
+ 6845.700000ns, VDD,
+ 6845.800000ns, VSS,
+ 7085.900000ns, VSS,
+ 7086.000000ns, VDD,
+ 7206.000000ns, VDD,
+ 7206.100000ns, VSS,
+ 7926.600000ns, VSS,
+ 7926.700000ns, VDD,
+ 9247.700000ns, VDD,
+ 9247.800000ns, VSS,
+ 9728.100000ns, VSS,
+ 9728.200000ns, VDD,
+ 10088.400000ns, VDD,
+ 10088.500000ns, VSS,
+ 10929.100000ns, VSS,
+ 10929.200000ns, VDD,
+ 12130.100000ns, VDD,
+ 12130.200000ns, VSS,
+ 12850.700000ns, VSS,
+ 12850.800000ns, VDD,
+ 13090.900000ns, VDD,
+ 13091.000000ns, VSS,
+ 13451.200000ns, VSS,
+ 13451.300000ns, VDD,
+ 14051.700000ns, VDD,
+ 14051.800000ns, VSS,
+ 14171.800000ns, VSS,
+ 14171.900000ns, VDD,
+ 15613.000000ns, VDD,
+ 15613.100000ns, VSS,
+ 16093.400000ns, VSS,
+ 16093.500000ns, VDD,
+ 16573.800000ns, VDD,
+ 16573.900000ns, VSS,
+ 17054.200000ns, VSS,
+ 17054.300000ns, VDD,
+ 18015.000000ns, VDD,
+ 18015.100000ns, VSS,
+ 18495.400000ns, VSS,
+ 18495.500000ns, VDD,
+ 18855.700000ns, VDD,
+ 18855.800000ns, VSS,
+ 19816.500000ns, VSS,
+ 19816.600000ns, VDD,
+ 20657.200000ns, VDD,
+ 20657.300000ns, VSS,
+ 20897.400000ns, VSS,
+ 20897.500000ns, VDD,
+ 21017.500000ns, VDD,
+ 21017.600000ns, VSS,
+ 21137.600000ns, VSS,
+ 21137.700000ns, VDD,
+ 21377.800000ns, VDD,
+ 21377.900000ns, VSS,
+ 21858.200000ns, VSS,
+ 21858.300000ns, VDD,
+ 21978.300000ns, VDD,
+ 21978.400000ns, VSS,
+ 23059.200000ns, VSS,
+ 23059.300000ns, VDD,
+ 23179.300000ns, VDD,
+ 23179.400000ns, VSS,
+ 23299.400000ns, VSS,
+ 23299.500000ns, VDD,
+ 23779.800000ns, VDD,
+ 23779.900000ns, VSS,
+ 24740.600000ns, VSS,
+ 24740.700000ns, VDD,
+ 24980.800000ns, VDD,
+ 24980.900000ns, VSS,
+ 25100.900000ns, VSS,
+ 25101.000000ns, VDD,
+ 25701.400000ns, VDD,
+ 25701.500000ns, VSS,
+ 26422.000000ns, VSS,
+ 26422.100000ns, VDD,
+ 28343.600000ns, VDD,
+ 28343.700000ns, VSS,
+ 30505.400000ns, VSS,
+ 30505.500000ns, VDD,
+ 30985.800000ns, VDD,
+ 30985.900000ns, VSS,
+ 31226.000000ns, VSS,
+ 31226.100000ns, VDD,
+ 31466.200000ns, VDD,
+ 31466.300000ns, VSS,
+ 32547.100000ns, VSS,
+ 32547.200000ns, VDD,
+ 33387.800000ns, VDD,
+ 33387.900000ns, VSS,
+ 34829.000000ns, VSS,
+ 34829.100000ns, VDD,
+ 35429.500000ns, VDD,
+ 35429.600000ns, VSS,
+ 36390.300000ns, VSS,
+ 36390.400000ns, VDD,
+ 37351.100000ns, VDD,
+ 37351.200000ns, VSS,
+ 37471.200000ns, VSS,
+ 37471.300000ns, VDD,
+ 37951.600000ns, VDD,
+ 37951.700000ns, VSS,
+ 38792.300000ns, VSS,
+ 38792.400000ns, VDD,
+ 40113.400000ns, VDD,
+ 40113.500000ns, VSS,
+ 40593.800000ns, VSS,
+ 40593.900000ns, VDD,
+ 41074.200000ns, VDD,
+ 41074.300000ns, VSS,
+ 41434.500000ns, VSS,
+ 41434.600000ns, VDD,
+ 41914.900000ns, VDD,
+ 41915.000000ns, VSS,
+ 42515.400000ns, VSS,
+ 42515.500000ns, VDD,
+ 42995.800000ns, VDD,
+ 42995.900000ns, VSS,
+ 43476.200000ns, VSS,
+ 43476.300000ns, VDD,
+ 44076.700000ns, VDD,
+ 44076.800000ns, VSS,
+ 44797.300000ns, VSS,
+ 44797.400000ns, VDD,
+ 45037.500000ns, VDD,
+ 45037.600000ns, VSS,
+ 45397.800000ns, VSS,
+ 45397.900000ns, VDD,
+ 45638.000000ns, VDD,
+ 45638.100000ns, VSS,
+ 45758.100000ns, VSS,
+ 45758.200000ns, VDD,
+ 46238.500000ns, VDD,
+ 46238.600000ns, VSS,
+ 46478.700000ns, VSS,
+ 46478.800000ns, VDD,
+ 47319.400000ns, VDD,
+ 47319.500000ns, VSS,
+ 48400.300000ns, VSS,
+ 48400.400000ns, VDD,
+ 48640.500000ns, VDD,
+ 48640.600000ns, VSS,
+ 49120.900000ns, VSS,
+ 49121.000000ns, VDD,
+ 50081.700000ns, VDD,
+ 50081.800000ns, VSS,
+ 51522.900000ns, VSS,
+ 51523.000000ns, VDD,
+ 51643.000000ns, VDD,
+ 51643.100000ns, VSS,
+ 52123.400000ns, VSS,
+ 52123.500000ns, VDD,
+ 53324.400000ns, VDD,
+ 53324.500000ns, VSS,
+ 54645.500000ns, VSS,
+ 54645.600000ns, VDD,
+ 56326.900000ns, VDD,
+ 56327.000000ns, VSS,
+ 56447.000000ns, VSS,
+ 56447.100000ns, VDD,
+ 56567.100000ns, VDD,
+ 56567.200000ns, VSS,
+ 57047.500000ns, VSS,
+ 57047.600000ns, VDD,
+ 57527.900000ns, VDD,
+ 57528.000000ns, VSS,
+ 57768.100000ns, VSS,
+ 57768.200000ns, VDD,
+ 58728.900000ns, VDD,
+ 58729.000000ns, VSS,
+ 58969.100000ns, VSS,
+ 58969.200000ns, VDD,
+ 59089.200000ns, VDD,
+ 59089.300000ns, VSS,
+ 59689.700000ns, VSS,
+ 59689.800000ns, VDD,
+ 60290.200000ns, VDD,
+ 60290.300000ns, VSS,
+ 60650.500000ns, VSS,
+ 60650.600000ns, VDD,
+ 61130.900000ns, VDD,
+ 61131.000000ns, VSS,
+ 62091.700000ns, VSS,
+ 62091.800000ns, VDD,
+ 62572.100000ns, VDD,
+ 62572.200000ns, VSS,
+ 63893.200000ns, VSS,
+ 63893.300000ns, VDD,
+ 64613.800000ns, VDD,
+ 64613.900000ns, VSS,
+ 64854.000000ns, VSS,
+ 64854.100000ns, VDD,
+ 65574.600000ns, VDD,
+ 65574.700000ns, VSS,
+ 65934.900000ns, VSS,
+ 65935.000000ns, VDD,
+ 66295.200000ns, VDD,
+ 66295.300000ns, VSS,
+ 66655.500000ns, VSS,
+ 66655.600000ns, VDD,
+ 68096.700000ns, VDD,
+ 68096.800000ns, VSS,
+ 69898.200000ns, VSS,
+ 69898.300000ns, VDD,
+ 70498.700000ns, VDD,
+ 70498.800000ns, VSS,
+ 70979.100000ns, VSS,
+ 70979.200000ns, VDD,
+ 72060.000000ns, VDD,
+ 72060.100000ns, VSS,
+ 72540.400000ns, VSS,
+ 72540.500000ns, VDD,
+ 72900.700000ns, VDD,
+ 72900.800000ns, VSS,
+ 73020.800000ns, VSS,
+ 73020.900000ns, VDD,
+ 73140.900000ns, VDD,
+ 73141.000000ns, VSS,
+ 73861.500000ns, VSS,
+ 73861.600000ns, VDD,
+ 74942.400000ns, VDD,
+ 74942.500000ns, VSS,
+ 75302.700000ns, VSS,
+ 75302.800000ns, VDD,
+ 75663.000000ns, VDD,
+ 75663.100000ns, VSS,
+ 76383.600000ns, VSS,
+ 76383.700000ns, VDD,
+ 76503.700000ns, VDD,
+ 76503.800000ns, VSS,
+ 77104.200000ns, VSS,
+ 77104.300000ns, VDD,
+ 79986.600000ns, VDD,
+ 79986.700000ns, VSS,
+ 80346.900000ns, VSS,
+ 80347.000000ns, VDD,
+ 80467.000000ns, VDD,
+ 80467.100000ns, VSS,
+ 80587.100000ns, VSS,
+ 80587.200000ns, VDD,
+ 81908.200000ns, VDD,
+ 81908.300000ns, VSS,
+ 82748.900000ns, VSS,
+ 82749.000000ns, VDD,
+ 82989.100000ns, VDD,
+ 82989.200000ns, VSS,
+ 83469.500000ns, VSS,
+ 83469.600000ns, VDD,
+ 83949.900000ns, VDD,
+ 83950.000000ns, VSS,
+ 84790.600000ns, VSS,
+ 84790.700000ns, VDD,
+ 84910.700000ns, VDD,
+ 84910.800000ns, VSS,
+ 85030.800000ns, VSS,
+ 85030.900000ns, VDD,
+ 86832.300000ns, VDD,
+ 86832.400000ns, VSS,
+ 87192.600000ns, VSS,
+ 87192.700000ns, VDD,
+ 87793.100000ns, VDD,
+ 87793.200000ns, VSS,
+ 88033.300000ns, VSS,
+ 88033.400000ns, VDD,
+ 88513.700000ns, VDD,
+ 88513.800000ns, VSS,
+ 88753.900000ns, VSS,
+ 88754.000000ns, VDD,
+ 89474.500000ns, VDD,
+ 89474.600000ns, VSS,
+ 90195.100000ns, VSS,
+ 90195.200000ns, VDD,
+ 91876.500000ns, VDD,
+ 91876.600000ns, VSS,
+ 93557.900000ns, VSS,
+ 93558.000000ns, VDD,
+ 95719.700000ns, VDD,
+ 95719.800000ns, VSS,
+ 96920.700000ns, VSS,
+ 96920.800000ns, VDD,
+ 99082.500000ns, VDD,
+ 99082.600000ns, VSS,
+ 100163.400000ns, VSS,
+ 100163.500000ns, VDD,
+ 101844.800000ns, VDD,
+ 101844.900000ns, VSS,
+ 102445.300000ns, VSS,
+ 102445.400000ns, VDD,
+ 103286.000000ns, VDD,
+ 103286.100000ns, VSS,
+ 103646.300000ns, VSS,
+ 103646.400000ns, VDD,
+ 103886.500000ns, VDD,
+ 103886.600000ns, VSS,
+ 104006.600000ns, VSS,
+ 104006.700000ns, VDD,
+ 104246.800000ns, VDD,
+ 104246.900000ns, VSS,
+ 105928.200000ns, VSS,
+ 105928.300000ns, VDD,
+ 106168.400000ns, VDD,
+ 106168.500000ns, VSS,
+ 106288.500000ns, VSS,
+ 106288.600000ns, VDD,
+ 106768.900000ns, VDD,
+ 106769.000000ns, VSS,
+ 106889.000000ns, VSS,
+ 106889.100000ns, VDD,
+ 107249.300000ns, VDD,
+ 107249.400000ns, VSS,
+ 107369.400000ns, VSS,
+ 107369.500000ns, VDD,
+ 107489.500000ns, VDD,
+ 107489.600000ns, VSS,
+ 107729.700000ns, VSS,
+ 107729.800000ns, VDD,
+ 107849.800000ns, VDD,
+ 107849.900000ns, VSS,
+ 109050.800000ns, VSS,
+ 109050.900000ns, VDD,
+ 109411.100000ns, VDD,
+ 109411.200000ns, VSS,
+ 110732.200000ns, VSS,
+ 110732.300000ns, VDD,
+ 111092.500000ns, VDD,
+ 111092.600000ns, VSS,
+ 112053.300000ns, VSS,
+ 112053.400000ns, VDD,
+ 112653.800000ns, VDD,
+ 112653.900000ns, VSS,
+ 114575.400000ns, VSS,
+ 114575.500000ns, VDD,
+ 114935.700000ns, VDD,
+ 114935.800000ns, VSS,
+ 115175.900000ns, VSS,
+ 115176.000000ns, VDD,
+ 115536.200000ns, VDD,
+ 115536.300000ns, VSS,
+ 115896.500000ns, VSS,
+ 115896.600000ns, VDD,
+ 116136.700000ns, VDD,
+ 116136.800000ns, VSS,
+ 116857.300000ns, VSS,
+ 116857.400000ns, VDD,
+ 117818.100000ns, VDD,
+ 117818.200000ns, VSS,
+ 118178.400000ns, VSS,
+ 118178.500000ns, VDD,
+ 118899.000000ns, VDD,
+ 118899.100000ns, VSS,
+ 120100.000000ns, VSS,
+ 120100.100000ns, VDD,
+ 120220.100000ns, VDD,
+ 120220.200000ns, VSS,
+ 120340.200000ns, VSS,
+ 120340.300000ns, VDD,
+ 120820.600000ns, VDD,
+ 120820.700000ns, VSS,
+ 121301.000000ns, VSS,
+ 121301.100000ns, VDD,
+ 122021.600000ns, VDD,
+ 122021.700000ns, VSS,
+ 122862.300000ns, VSS,
+ 122862.400000ns, VDD,
+ 123703.000000ns, VDD,
+ 123703.100000ns, VSS,
+ 124183.400000ns, VSS,
+ 124183.500000ns, VDD,
+ 125024.100000ns, VDD,
+ 125024.200000ns, VSS,
+ 125504.500000ns, VSS,
+ 125504.600000ns, VDD,
+ 126345.200000ns, VDD,
+ 126345.300000ns, VSS,
+ 126825.600000ns, VSS,
+ 126825.700000ns, VDD,
+ 127065.800000ns, VDD,
+ 127065.900000ns, VSS,
+ 128627.100000ns, VSS,
+ 128627.200000ns, VDD,
+ 128747.200000ns, VDD,
+ 128747.300000ns, VSS,
+ 128867.300000ns, VSS,
+ 128867.400000ns, VDD,
+ 129227.600000ns, VDD,
+ 129227.700000ns, VSS,
+ 129347.700000ns, VSS,
+ 129347.800000ns, VDD,
+ 130188.400000ns, VDD,
+ 130188.500000ns, VSS,
+ 131149.200000ns, VSS,
+ 131149.300000ns, VDD,
+ 131869.800000ns, VDD,
+ 131869.900000ns, VSS,
+ 132230.100000ns, VSS,
+ 132230.200000ns, VDD,
+ 132470.300000ns, VDD,
+ 132470.400000ns, VSS,
+ 132710.500000ns, VSS,
+ 132710.600000ns, VDD,
+ 133311.000000ns, VDD,
+ 133311.100000ns, VSS,
+ 134271.800000ns, VSS,
+ 134271.900000ns, VDD,
+ 135352.700000ns, VDD,
+ 135352.800000ns, VSS,
+ 136673.800000ns, VSS,
+ 136673.900000ns, VDD,
+ 136793.900000ns, VDD,
+ 136794.000000ns, VSS,
+ 136914.000000ns, VSS,
+ 136914.100000ns, VDD,
+ 137274.300000ns, VDD,
+ 137274.400000ns, VSS,
+ 137514.500000ns, VSS,
+ 137514.600000ns, VDD,
+ 137634.600000ns, VDD,
+ 137634.700000ns, VSS,
+ 138355.200000ns, VSS,
+ 138355.300000ns, VDD,
+ 139195.900000ns, VDD,
+ 139196.000000ns, VSS,
+ 139556.200000ns, VSS,
+ 139556.300000ns, VDD,
+ 140517.000000ns, VDD,
+ 140517.100000ns, VSS,
+ 141597.900000ns, VSS,
+ 141598.000000ns, VDD,
+ 141718.000000ns, VDD,
+ 141718.100000ns, VSS,
+ 143039.100000ns, VSS,
+ 143039.200000ns, VDD,
+ 143279.300000ns, VDD,
+ 143279.400000ns, VSS,
+ 143639.600000ns, VSS,
+ 143639.700000ns, VDD,
+ 143759.700000ns, VDD,
+ 143759.800000ns, VSS,
+ 143879.800000ns, VSS,
+ 143879.900000ns, VDD,
+ 144120.000000ns, VDD,
+ 144120.100000ns, VSS,
+ 145200.900000ns, VSS,
+ 145201.000000ns, VDD,
+ 145801.400000ns, VDD,
+ 145801.500000ns, VSS,
+ 146762.200000ns, VSS,
+ 146762.300000ns, VDD,
+ 147362.700000ns, VDD,
+ 147362.800000ns, VSS,
+ 147843.100000ns, VSS,
+ 147843.200000ns, VDD,
+ 150004.900000ns, VDD,
+ 150005.000000ns, VSS,
+ 151205.900000ns, VSS,
+ 151206.000000ns, VDD,
+ 153728.000000ns, VDD,
+ 153728.100000ns, VSS,
+ 154088.300000ns, VSS,
+ 154088.400000ns, VDD,
+ 154688.800000ns, VDD,
+ 154688.900000ns, VSS,
+ 155049.100000ns, VSS,
+ 155049.200000ns, VDD,
+ 155289.300000ns, VDD,
+ 155289.400000ns, VSS,
+ 155409.400000ns, VSS,
+ 155409.500000ns, VDD,
+ 155529.500000ns, VDD,
+ 155529.600000ns, VSS,
+ 156009.900000ns, VSS,
+ 156010.000000ns, VDD,
+ 156130.000000ns, VDD,
+ 156130.100000ns, VSS,
+ 156250.100000ns, VSS,
+ 156250.200000ns, VDD,
+ 157210.900000ns, VDD,
+ 157211.000000ns, VSS,
+ 157451.100000ns, VSS,
+ 157451.200000ns, VDD,
+ 157691.300000ns, VDD,
+ 157691.400000ns, VSS,
+ 157931.500000ns, VSS,
+ 157931.600000ns, VDD,
+ 158291.800000ns, VDD,
+ 158291.900000ns, VSS,
+ 158652.100000ns, VSS,
+ 158652.200000ns, VDD,
+ 159612.900000ns, VDD,
+ 159613.000000ns, VSS,
+ 159973.200000ns, VSS,
+ 159973.300000ns, VDD,
+ 161174.200000ns, VDD,
+ 161174.300000ns, VSS,
+ 161654.600000ns, VSS,
+ 161654.700000ns, VDD,
+ 162014.900000ns, VDD,
+ 162015.000000ns, VSS,
+ 162975.700000ns, VSS,
+ 162975.800000ns, VDD,
+ 163696.300000ns, VDD,
+ 163696.400000ns, VSS,
+ 165137.500000ns, VSS,
+ 165137.600000ns, VDD,
+ 165497.800000ns, VDD,
+ 165497.900000ns, VSS,
+ 165978.200000ns, VSS,
+ 165978.300000ns, VDD,
+ 166939.000000ns, VDD,
+ 166939.100000ns, VSS,
+ 167779.700000ns, VSS,
+ 167779.800000ns, VDD,
+ 168500.300000ns, VDD,
+ 168500.400000ns, VSS,
+ 170061.600000ns, VSS,
+ 170061.700000ns, VDD,
+ 170542.000000ns, VDD,
+ 170542.100000ns, VSS,
+ 172703.800000ns, VSS,
+ 172703.900000ns, VDD,
+ 173184.200000ns, VDD,
+ 173184.300000ns, VSS,
+ 173664.600000ns, VSS,
+ 173664.700000ns, VDD,
+ 174145.000000ns, VDD,
+ 174145.100000ns, VSS,
+ 174865.600000ns, VSS,
+ 174865.700000ns, VDD,
+ 175225.900000ns, VDD,
+ 175226.000000ns, VSS,
+ 175586.200000ns, VSS,
+ 175586.300000ns, VDD,
+ 175706.300000ns, VDD,
+ 175706.400000ns, VSS,
+ 175826.400000ns, VSS,
+ 175826.500000ns, VDD,
+ 177507.800000ns, VDD,
+ 177507.900000ns, VSS,
+ 177748.000000ns, VSS,
+ 177748.100000ns, VDD,
+ 178348.500000ns, VDD,
+ 178348.600000ns, VSS,
+ 179549.500000ns, VSS,
+ 179549.600000ns, VDD,
+ 179789.700000ns, VDD,
+ 179789.800000ns, VSS,
+ 180029.900000ns, VSS,
+ 180030.000000ns, VDD,
+ 180630.400000ns, VDD,
+ 180630.500000ns, VSS,
+ 181110.800000ns, VSS,
+ 181110.900000ns, VDD,
+ 181711.300000ns, VDD,
+ 181711.400000ns, VSS,
+ 181831.400000ns, VSS,
+ 181831.500000ns, VDD,
+ 186155.000000ns, VDD,
+ 186155.100000ns, VSS,
+ 186395.200000ns, VSS,
+ 186395.300000ns, VDD,
+ 186515.300000ns, VDD,
+ 186515.400000ns, VSS,
+ 186635.400000ns, VSS,
+ 186635.500000ns, VDD,
+ 186995.700000ns, VDD,
+ 186995.800000ns, VSS,
+ 187476.100000ns, VSS,
+ 187476.200000ns, VDD,
+ 189037.400000ns, VDD,
+ 189037.500000ns, VSS,
+ 189397.700000ns, VSS,
+ 189397.800000ns, VDD,
+ 189637.900000ns, VDD,
+ 189638.000000ns, VSS,
+ 190238.400000ns, VSS,
+ 190238.500000ns, VDD,
+ 190959.000000ns, VDD,
+ 190959.100000ns, VSS,
+ 193240.900000ns, VSS,
+ 193241.000000ns, VDD,
+ 193601.200000ns, VDD,
+ 193601.300000ns, VSS,
+ 193721.300000ns, VSS,
+ 193721.400000ns, VDD,
+ 193841.400000ns, VDD,
+ 193841.500000ns, VSS,
+ 194201.700000ns, VSS,
+ 194201.800000ns, VDD,
+ 194802.200000ns, VDD,
+ 194802.300000ns, VSS,
+ 195162.500000ns, VSS,
+ 195162.600000ns, VDD,
+ 198044.900000ns, VDD,
+ 198045.000000ns, VSS,
+ 198165.000000ns, VSS,
+ 198165.100000ns, VDD,
+ 199245.900000ns, VDD,
+ 199246.000000ns, VSS,
+ 199726.300000ns, VSS,
+ 199726.400000ns, VDD,
+ 199846.400000ns, VDD,
+ 199846.500000ns, VSS,
+ 199966.500000ns, VSS,
+ 199966.600000ns, VDD,
+ 201407.700000ns, VDD,
+ 201407.800000ns, VSS,
+ 202368.500000ns, VSS,
+ 202368.600000ns, VDD,
+ 203209.200000ns, VDD,
+ 203209.300000ns, VSS,
+ 203449.400000ns, VSS,
+ 203449.500000ns, VDD,
+ 203689.600000ns, VDD,
+ 203689.700000ns, VSS,
+ 204290.100000ns, VSS,
+ 204290.200000ns, VDD,
+ 204410.200000ns, VDD,
+ 204410.300000ns, VSS,
+ 204530.300000ns, VSS,
+ 204530.400000ns, VDD,
+ 207292.600000ns, VDD,
+ 207292.700000ns, VSS,
+ 209094.100000ns, VSS,
+ 209094.200000ns, VDD,
+ 209814.700000ns, VDD,
+ 209814.800000ns, VSS,
+ 209934.800000ns, VSS,
+ 209934.900000ns, VDD,
+ 210175.000000ns, VDD,
+ 210175.100000ns, VSS,
+ 210655.400000ns, VSS,
+ 210655.500000ns, VDD,
+ 211135.800000ns, VDD,
+ 211135.900000ns, VSS,
+ 211856.400000ns, VSS,
+ 211856.500000ns, VDD,
+ 212577.000000ns, VDD,
+ 212577.100000ns, VSS,
+ 212817.200000ns, VSS,
+ 212817.300000ns, VDD,
+ 213657.900000ns, VDD,
+ 213658.000000ns, VSS,
+ 214138.300000ns, VSS,
+ 214138.400000ns, VDD,
+ 214258.400000ns, VDD,
+ 214258.500000ns, VSS,
+ 214979.000000ns, VSS,
+ 214979.100000ns, VDD,
+ 215579.500000ns, VDD,
+ 215579.600000ns, VSS,
+ 216540.300000ns, VSS,
+ 216540.400000ns, VDD,
+ 216780.500000ns, VDD,
+ 216780.600000ns, VSS,
+ 217501.100000ns, VSS,
+ 217501.200000ns, VDD,
+ 218221.700000ns, VDD,
+ 218221.800000ns, VSS,
+ 218702.100000ns, VSS,
+ 218702.200000ns, VDD,
+ 218942.300000ns, VDD,
+ 218942.400000ns, VSS,
+ 219182.500000ns, VSS,
+ 219182.600000ns, VDD,
+ 219783.000000ns, VDD,
+ 219783.100000ns, VSS,
+ 220143.300000ns, VSS,
+ 220143.400000ns, VDD,
+ 220503.600000ns, VDD,
+ 220503.700000ns, VSS,
+ 220743.800000ns, VSS,
+ 220743.900000ns, VDD,
+ 222185.000000ns, VDD,
+ 222185.100000ns, VSS,
+ 222665.400000ns, VSS,
+ 222665.500000ns, VDD,
+ 222905.600000ns, VDD,
+ 222905.700000ns, VSS,
+ 223025.700000ns, VSS,
+ 223025.800000ns, VDD,
+ 223265.900000ns, VDD,
+ 223266.000000ns, VSS,
+ 223386.000000ns, VSS,
+ 223386.100000ns, VDD,
+ 223746.300000ns, VDD,
+ 223746.400000ns, VSS,
+ 224466.900000ns, VSS,
+ 224467.000000ns, VDD,
+ 225788.000000ns, VDD,
+ 225788.100000ns, VSS,
+ 226148.300000ns, VSS,
+ 226148.400000ns, VDD,
+ 226628.700000ns, VDD,
+ 226628.800000ns, VSS,
+ 227109.100000ns, VSS,
+ 227109.200000ns, VDD,
+ 227709.600000ns, VDD,
+ 227709.700000ns, VSS,
+ 227829.700000ns, VSS,
+ 227829.800000ns, VDD,
+ 227949.800000ns, VDD,
+ 227949.900000ns, VSS,
+ 228310.100000ns, VSS,
+ 228310.200000ns, VDD,
+ 229150.800000ns, VDD,
+ 229150.900000ns, VSS,
+ 230111.600000ns, VSS,
+ 230111.700000ns, VDD,
+ 231072.400000ns, VDD,
+ 231072.500000ns, VSS,
+ 231793.000000ns, VSS,
+ 231793.100000ns, VDD,
+ 231913.100000ns, VDD,
+ 231913.200000ns, VSS,
+ 233714.600000ns, VSS,
+ 233714.700000ns, VDD,
+ 234074.900000ns, VDD,
+ 234075.000000ns, VSS,
+ 234315.100000ns, VSS,
+ 234315.200000ns, VDD,
+ 234795.500000ns, VDD,
+ 234795.600000ns, VSS,
+ 236236.700000ns, VSS,
+ 236236.800000ns, VDD,
+ 236717.100000ns, VDD,
+ 236717.200000ns, VSS,
+ 236837.200000ns, VSS,
+ 236837.300000ns, VDD,
+ 237557.800000ns, VDD,
+ 237557.900000ns, VSS,
+ 238638.700000ns, VSS,
+ 238638.800000ns, VDD,
+ 239359.300000ns, VDD,
+ 239359.400000ns, VSS,
+ 239839.700000ns, VSS,
+ 239839.800000ns, VDD,
+ 240920.600000ns, VDD,
+ 240920.700000ns, VSS,
+ 241761.300000ns, VSS,
+ 241761.400000ns, VDD,
+ 242481.900000ns, VDD,
+ 242482.000000ns, VSS,
+ 243082.400000ns, VSS,
+ 243082.500000ns, VDD,
+ 243562.800000ns, VDD,
+ 243562.900000ns, VSS,
+ 243682.900000ns, VSS,
+ 243683.000000ns, VDD,
+ 243923.100000ns, VDD,
+ 243923.200000ns, VSS,
+ 245604.500000ns, VSS,
+ 245604.600000ns, VDD,
+ 246205.000000ns, VDD,
+ 246205.100000ns, VSS,
+ 246325.100000ns, VSS,
+ 246325.200000ns, VDD,
+ 246805.500000ns, VDD,
+ 246805.600000ns, VSS,
+ 247526.100000ns, VSS,
+ 247526.200000ns, VDD,
+ 248006.500000ns, VDD,
+ 248006.600000ns, VSS,
+ 248126.600000ns, VSS,
+ 248126.700000ns, VDD,
+ 248366.800000ns, VDD,
+ 248366.900000ns, VSS,
+ 248967.300000ns, VSS,
+ 248967.400000ns, VDD,
+ 249687.900000ns, VDD,
+ 249688.000000ns, VSS,
+ 250048.200000ns, VSS,
+ 250048.300000ns, VDD,
+ 250408.500000ns, VDD,
+ 250408.600000ns, VSS,
+ 251009.000000ns, VSS,
+ 251009.100000ns, VDD,
+ 251489.400000ns, VDD,
+ 251489.500000ns, VSS,
+ 251969.800000ns, VSS,
+ 251969.900000ns, VDD,
+ 252810.500000ns, VDD,
+ 252810.600000ns, VSS,
+ 253891.400000ns, VSS,
+ 253891.500000ns, VDD,
+ 254131.600000ns, VDD,
+ 254131.700000ns, VSS,
+ 254732.100000ns, VSS,
+ 254732.200000ns, VDD,
+ 255212.500000ns, VDD,
+ 255212.600000ns, VSS,
+ 255332.600000ns, VSS,
+ 255332.700000ns, VDD,
+ 255813.000000ns, VDD,
+ 255813.100000ns, VSS,
+ 256413.500000ns, VSS,
+ 256413.600000ns, VDD,
+ 256773.800000ns, VDD,
+ 256773.900000ns, VSS,
+ 258094.900000ns, VSS,
+ 258095.000000ns, VDD,
+ 258575.300000ns, VDD,
+ 258575.400000ns, VSS,
+ 258695.400000ns, VSS,
+ 258695.500000ns, VDD,
+ 260136.600000ns, VDD,
+ 260136.700000ns, VSS,
+ 260617.000000ns, VSS,
+ 260617.100000ns, VDD,
+ 260737.100000ns, VDD,
+ 260737.200000ns, VSS,
+ 261097.400000ns, VSS,
+ 261097.500000ns, VDD,
+ 261217.500000ns, VDD,
+ 261217.600000ns, VSS,
+ 261457.700000ns, VSS,
+ 261457.800000ns, VDD,
+ 261938.100000ns, VDD,
+ 261938.200000ns, VSS,
+ 262538.600000ns, VSS,
+ 262538.700000ns, VDD,
+ 263019.000000ns, VDD,
+ 263019.100000ns, VSS,
+ 263619.500000ns, VSS,
+ 263619.600000ns, VDD,
+ 263739.600000ns, VDD,
+ 263739.700000ns, VSS,
+ 264700.400000ns, VSS,
+ 264700.500000ns, VDD,
+ 265060.700000ns, VDD,
+ 265060.800000ns, VSS,
+ 266501.900000ns, VSS,
+ 266502.000000ns, VDD,
+ 266982.300000ns, VDD,
+ 266982.400000ns, VSS,
+ 267342.600000ns, VSS,
+ 267342.700000ns, VDD,
+ 268303.400000ns, VDD,
+ 268303.500000ns, VSS,
+ 269264.200000ns, VSS,
+ 269264.300000ns, VDD,
+ 269864.700000ns, VDD,
+ 269864.800000ns, VSS,
+ 269984.800000ns, VSS,
+ 269984.900000ns, VDD,
+ 270104.900000ns, VDD,
+ 270105.000000ns, VSS,
+ 270225.000000ns, VSS,
+ 270225.100000ns, VDD,
+ 270345.100000ns, VDD,
+ 270345.200000ns, VSS,
+ 273107.400000ns, VSS,
+ 273107.500000ns, VDD,
+ 273828.000000ns, VDD,
+ 273828.100000ns, VSS,
+ 274668.700000ns, VSS,
+ 274668.800000ns, VDD,
+ 274788.800000ns, VDD,
+ 274788.900000ns, VSS,
+ 275149.100000ns, VSS,
+ 275149.200000ns, VDD,
+ 275629.500000ns, VDD,
+ 275629.600000ns, VSS,
+ 277551.100000ns, VSS,
+ 277551.200000ns, VDD,
+ 277911.400000ns, VDD,
+ 277911.500000ns, VSS,
+ 278391.800000ns, VSS,
+ 278391.900000ns, VDD,
+ 281274.200000ns, VDD,
+ 281274.300000ns, VSS,
+ 282355.100000ns, VSS,
+ 282355.200000ns, VDD,
+ 282715.400000ns, VDD,
+ 282715.500000ns, VSS,
+ 283315.900000ns, VSS,
+ 283316.000000ns, VDD,
+ 283436.000000ns, VDD,
+ 283436.100000ns, VSS,
+ 283556.100000ns, VSS,
+ 283556.200000ns, VDD,
+ 284997.300000ns, VDD,
+ 284997.400000ns, VSS,
+ 285597.800000ns, VSS,
+ 285597.900000ns, VDD,
+ 285838.000000ns, VDD,
+ 285838.100000ns, VSS,
+ 286078.200000ns, VSS,
+ 286078.300000ns, VDD,
+ 286198.300000ns, VDD,
+ 286198.400000ns, VSS,
+ 286918.900000ns, VSS,
+ 286919.000000ns, VDD,
+ 287999.800000ns, VDD,
+ 287999.900000ns, VSS,
+ 288240.000000ns, VSS,
+ 288240.100000ns, VDD,
+ 288840.500000ns, VDD,
+ 288840.600000ns, VSS,
+ 289080.700000ns, VSS,
+ 289080.800000ns, VDD,
+ 289801.300000ns, VDD,
+ 289801.400000ns, VSS,
+ 290161.600000ns, VSS,
+ 290161.700000ns, VDD,
+ 290642.000000ns, VDD,
+ 290642.100000ns, VSS,
+ 290762.100000ns, VSS,
+ 290762.200000ns, VDD,
+ 292683.700000ns, VDD,
+ 292683.800000ns, VSS,
+ 294365.100000ns, VSS,
+ 294365.200000ns, VDD,
+ 294965.600000ns, VDD,
+ 294965.700000ns, VSS,
+ 295205.800000ns, VSS,
+ 295205.900000ns, VDD,
+ 298568.600000ns, VDD,
+ 298568.700000ns, VSS,
+ 298808.800000ns, VSS,
+ 298808.900000ns, VDD,
+ 299169.100000ns, VDD,
+ 299169.200000ns, VSS,
+ 299769.600000ns, VSS,
+ 299769.700000ns, VDD,
+ 300250.000000ns, VDD,
+ 300250.100000ns, VSS,
+ 300370.100000ns, VSS,
+ 300370.200000ns, VDD,
+ 300490.200000ns, VDD,
+ 300490.300000ns, VSS,
+ 301330.900000ns, VSS,
+ 301331.000000ns, VDD,
+ 301811.300000ns, VDD,
+ 301811.400000ns, VSS,
+ 302652.000000ns, VSS,
+ 302652.100000ns, VDD,
+ 303612.800000ns, VDD,
+ 303612.900000ns, VSS,
+ 304213.300000ns, VSS,
+ 304213.400000ns, VDD,
+ 306735.400000ns, VDD,
+ 306735.500000ns, VSS,
+ 307215.800000ns, VSS,
+ 307215.900000ns, VDD,
+ 308296.700000ns, VDD,
+ 308296.800000ns, VSS,
+ 308416.800000ns, VSS,
+ 308416.900000ns, VDD,
+ 308897.200000ns, VDD,
+ 308897.300000ns, VSS,
+ 310218.300000ns, VSS,
+ 310218.400000ns, VDD,
+ 311419.300000ns, VDD,
+ 311419.400000ns, VSS,
+ 311779.600000ns, VSS,
+ 311779.700000ns, VDD,
+ 311899.700000ns, VDD,
+ 311899.800000ns, VSS,
+ 312019.800000ns, VSS,
+ 312019.900000ns, VDD,
+ 312740.400000ns, VDD,
+ 312740.500000ns, VSS,
+ 314061.500000ns, VSS,
+ 314061.600000ns, VDD,
+ 314782.100000ns, VDD,
+ 314782.200000ns, VSS,
+ 315142.400000ns, VSS,
+ 315142.500000ns, VDD,
+ 315622.800000ns, VDD,
+ 315622.900000ns, VSS,
+ 315863.000000ns, VSS,
+ 315863.100000ns, VDD,
+ 316583.600000ns, VDD,
+ 316583.700000ns, VSS,
+ 316823.800000ns, VSS,
+ 316823.900000ns, VDD,
+ 317064.000000ns, VDD,
+ 317064.100000ns, VSS,
+ 317544.400000ns, VSS,
+ 317544.500000ns, VDD,
+ 318745.400000ns, VDD,
+ 318745.500000ns, VSS,
+ 319706.200000ns, VSS,
+ 319706.300000ns, VDD,
+ 321627.800000ns, VDD,
+ 321627.900000ns, VSS,
+ 323429.300000ns, VSS,
+ 323429.400000ns, VDD,
+ 324390.100000ns, VDD,
+ 324390.200000ns, VSS,
+ 324990.600000ns, VSS,
+ 324990.700000ns, VDD,
+ 325110.700000ns, VDD,
+ 325110.800000ns, VSS,
+ 326311.700000ns, VSS,
+ 326311.800000ns, VDD,
+ 326431.800000ns, VDD,
+ 326431.900000ns, VSS,
+ 329794.600000ns, VSS,
+ 329794.700000ns, VDD,
+ 330034.800000ns, VDD,
+ 330034.900000ns, VSS,
+ 331235.800000ns, VSS,
+ 331235.900000ns, VDD,
+ 331956.400000ns, VDD,
+ 331956.500000ns, VSS,
+ 332076.500000ns, VSS,
+ 332076.600000ns, VDD,
+ 332556.900000ns, VDD,
+ 332557.000000ns, VSS,
+ 333998.100000ns, VSS,
+ 333998.200000ns, VDD,
+ 334718.700000ns, VDD,
+ 334718.800000ns, VSS,
+ 335199.100000ns, VSS,
+ 335199.200000ns, VDD,
+ 335679.500000ns, VDD,
+ 335679.600000ns, VSS,
+ 336039.800000ns, VSS,
+ 336039.900000ns, VDD,
+ 336159.900000ns, VDD,
+ 336160.000000ns, VSS,
+ 336880.500000ns, VSS,
+ 336880.600000ns, VDD,
+ 337000.600000ns, VDD,
+ 337000.700000ns, VSS,
+ 337360.900000ns, VSS,
+ 337361.000000ns, VDD,
+ 338441.800000ns, VDD,
+ 338441.900000ns, VSS,
+ 338802.100000ns, VSS,
+ 338802.200000ns, VDD,
+ 338922.200000ns, VDD,
+ 338922.300000ns, VSS,
+ 339762.900000ns, VSS,
+ 339763.000000ns, VDD,
+ 340243.300000ns, VDD,
+ 340243.400000ns, VSS,
+ 340363.400000ns, VSS,
+ 340363.500000ns, VDD,
+ 340483.500000ns, VDD,
+ 340483.600000ns, VSS,
+ 340843.800000ns, VSS,
+ 340843.900000ns, VDD,
+ 341684.500000ns, VDD,
+ 341684.600000ns, VSS,
+ 342044.800000ns, VSS,
+ 342044.900000ns, VDD,
+ 342164.900000ns, VDD,
+ 342165.000000ns, VSS,
+ 342285.000000ns, VSS,
+ 342285.100000ns, VDD,
+ 343125.700000ns, VDD,
+ 343125.800000ns, VSS,
+ 343245.800000ns, VSS,
+ 343245.900000ns, VDD,
+ 343606.100000ns, VDD,
+ 343606.200000ns, VSS,
+ 344687.000000ns, VSS,
+ 344687.100000ns, VDD,
+ 345167.400000ns, VDD,
+ 345167.500000ns, VSS,
+ 345287.500000ns, VSS,
+ 345287.600000ns, VDD,
+ 345407.600000ns, VDD,
+ 345407.700000ns, VSS,
+ 346128.200000ns, VSS,
+ 346128.300000ns, VDD,
+ 347329.200000ns, VDD,
+ 347329.300000ns, VSS,
+ 347689.500000ns, VSS,
+ 347689.600000ns, VDD,
+ 347809.600000ns, VDD,
+ 347809.700000ns, VSS,
+ 348049.800000ns, VSS,
+ 348049.900000ns, VDD,
+ 348410.100000ns, VDD,
+ 348410.200000ns, VSS,
+ 349250.800000ns, VSS,
+ 349250.900000ns, VDD,
+ 349851.300000ns, VDD,
+ 349851.400000ns, VSS,
+ 350331.700000ns, VSS,
+ 350331.800000ns, VDD,
+ 350812.100000ns, VDD,
+ 350812.200000ns, VSS,
+ 351172.400000ns, VSS,
+ 351172.500000ns, VDD,
+ 352013.100000ns, VDD,
+ 352013.200000ns, VSS,
+ 352373.400000ns, VSS,
+ 352373.500000ns, VDD,
+ 353934.700000ns, VDD,
+ 353934.800000ns, VSS,
+ 355255.800000ns, VSS,
+ 355255.900000ns, VDD,
+ 355496.000000ns, VDD,
+ 355496.100000ns, VSS,
+ 355616.100000ns, VSS,
+ 355616.200000ns, VDD,
+ 355736.200000ns, VDD,
+ 355736.300000ns, VSS,
+ 358018.100000ns, VSS,
+ 358018.200000ns, VDD,
+ 359099.000000ns, VDD,
+ 359099.100000ns, VSS,
+ 359339.200000ns, VSS,
+ 359339.300000ns, VDD,
+ 359819.600000ns, VDD,
+ 359819.700000ns, VSS,
+ 360300.000000ns, VSS,
+ 360300.100000ns, VDD,
+ 360780.400000ns, VDD,
+ 360780.500000ns, VSS,
+ 360900.500000ns, VSS,
+ 360900.600000ns, VDD,
+ 361020.600000ns, VDD,
+ 361020.700000ns, VSS,
+ 362822.100000ns, VSS,
+ 362822.200000ns, VDD,
+ 363422.600000ns, VDD,
+ 363422.700000ns, VSS,
+ 363662.800000ns, VSS,
+ 363662.900000ns, VDD,
+ 364023.100000ns, VDD,
+ 364023.200000ns, VSS,
+ 364263.300000ns, VSS,
+ 364263.400000ns, VDD,
+ 364623.600000ns, VDD,
+ 364623.700000ns, VSS,
+ 364743.700000ns, VSS,
+ 364743.800000ns, VDD,
+ 365584.400000ns, VDD,
+ 365584.500000ns, VSS,
+ 366184.900000ns, VSS,
+ 366185.000000ns, VDD,
+ 367746.200000ns, VDD,
+ 367746.300000ns, VSS,
+ 368226.600000ns, VSS,
+ 368226.700000ns, VDD,
+ 368466.800000ns, VDD,
+ 368466.900000ns, VSS,
+ 369067.300000ns, VSS,
+ 369067.400000ns, VDD,
+ 369667.800000ns, VDD,
+ 369667.900000ns, VSS,
+ 372670.300000ns, VSS,
+ 372670.400000ns, VDD,
+ 373270.800000ns, VDD,
+ 373270.900000ns, VSS,
+ 373390.900000ns, VSS,
+ 373391.000000ns, VDD,
+ 373631.100000ns, VDD,
+ 373631.200000ns, VSS,
+ 373751.200000ns, VSS,
+ 373751.300000ns, VDD,
+ 375192.400000ns, VDD,
+ 375192.500000ns, VSS,
+ 376513.500000ns, VSS,
+ 376513.600000ns, VDD,
+ 376993.900000ns, VDD,
+ 376994.000000ns, VSS,
+ 377114.000000ns, VSS,
+ 377114.100000ns, VDD,
+ 377234.100000ns, VDD,
+ 377234.200000ns, VSS,
+ 377834.600000ns, VSS,
+ 377834.700000ns, VDD,
+ 378074.800000ns, VDD,
+ 378074.900000ns, VSS,
+ 378194.900000ns, VSS,
+ 378195.000000ns, VDD,
+ 378555.200000ns, VDD,
+ 378555.300000ns, VSS,
+ 378675.300000ns, VSS,
+ 378675.400000ns, VDD,
+ 379275.800000ns, VDD,
+ 379275.900000ns, VSS,
+ 379756.200000ns, VSS,
+ 379756.300000ns, VDD,
+ 379876.300000ns, VDD,
+ 379876.400000ns, VSS,
+ 379996.400000ns, VSS,
+ 379996.500000ns, VDD,
+ 380717.000000ns, VDD,
+ 380717.100000ns, VSS,
+ 382398.400000ns, VSS,
+ 382398.500000ns, VDD,
+ 384320.000000ns, VDD,
+ 384320.100000ns, VSS,
+ 384680.300000ns, VSS,
+ 384680.400000ns, VDD,
+ 385040.600000ns, VDD,
+ 385040.700000ns, VSS,
+ 385641.100000ns, VSS,
+ 385641.200000ns, VDD,
+ 386241.600000ns, VDD,
+ 386241.700000ns, VSS,
+ 387082.300000ns, VSS,
+ 387082.400000ns, VDD,
+ 388043.100000ns, VDD,
+ 388043.200000ns, VSS,
+ 388283.300000ns, VSS,
+ 388283.400000ns, VDD,
+ 389364.200000ns, VDD,
+ 389364.300000ns, VSS,
+ 390084.800000ns, VSS,
+ 390084.900000ns, VDD,
+ 390204.900000ns, VDD,
+ 390205.000000ns, VSS,
+ 390805.400000ns, VSS,
+ 390805.500000ns, VDD,
+ 391405.900000ns, VDD,
+ 391406.000000ns, VSS,
+ 392126.500000ns, VSS,
+ 392126.600000ns, VDD,
+ 392246.600000ns, VDD,
+ 392246.700000ns, VSS,
+ 392486.800000ns, VSS,
+ 392486.900000ns, VDD,
+ 392967.200000ns, VDD,
+ 392967.300000ns, VSS,
+ 393327.500000ns, VSS,
+ 393327.600000ns, VDD,
+ 393567.700000ns, VDD,
+ 393567.800000ns, VSS,
+ 393807.900000ns, VSS,
+ 393808.000000ns, VDD,
+ 394888.800000ns, VDD,
+ 394888.900000ns, VSS,
+ 395729.500000ns, VSS,
+ 395729.600000ns, VDD,
+ 396810.400000ns, VDD,
+ 396810.500000ns, VSS,
+ 397290.800000ns, VSS,
+ 397290.900000ns, VDD,
+ 398611.900000ns, VDD,
+ 398612.000000ns, VSS,
+ 400053.100000ns, VSS,
+ 400053.200000ns, VDD,
+ 401494.300000ns, VDD,
+ 401494.400000ns, VSS,
+ 401854.600000ns, VSS,
+ 401854.700000ns, VDD,
+ 402214.900000ns, VDD,
+ 402215.000000ns, VSS,
+ 402335.000000ns, VSS,
+ 402335.100000ns, VDD,
+ 402455.100000ns, VDD,
+ 402455.200000ns, VSS,
+ 402695.300000ns, VSS,
+ 402695.400000ns, VDD,
+ 403415.900000ns, VDD,
+ 403416.000000ns, VSS,
+ 404016.400000ns, VSS,
+ 404016.500000ns, VDD,
+ 404857.100000ns, VDD,
+ 404857.200000ns, VSS,
+ 406178.200000ns, VSS,
+ 406178.300000ns, VDD,
+ 406418.400000ns, VDD,
+ 406418.500000ns, VSS,
+ 407859.600000ns, VSS,
+ 407859.700000ns, VDD,
+ 408340.000000ns, VDD,
+ 408340.100000ns, VSS,
+ 408460.100000ns, VSS,
+ 408460.200000ns, VDD,
+ 409541.000000ns, VDD,
+ 409541.100000ns, VSS,
+ 410021.400000ns, VSS,
+ 410021.500000ns, VDD,
+ 410381.700000ns, VDD,
+ 410381.800000ns, VSS,
+ 410862.100000ns, VSS,
+ 410862.200000ns, VDD,
+ 411342.500000ns, VDD,
+ 411342.600000ns, VSS,
+ 411822.900000ns, VSS,
+ 411823.000000ns, VDD,
+ 412303.300000ns, VDD,
+ 412303.400000ns, VSS,
+ 413744.500000ns, VSS,
+ 413744.600000ns, VDD,
+ 414705.300000ns, VDD,
+ 414705.400000ns, VSS,
+ 415185.700000ns, VSS,
+ 415185.800000ns, VDD,
+ 415666.100000ns, VDD,
+ 415666.200000ns, VSS,
+ 416867.100000ns, VSS,
+ 416867.200000ns, VDD,
+ 419509.300000ns, VDD,
+ 419509.400000ns, VSS,
+ 420229.900000ns, VSS,
+ 420230.000000ns, VDD,
+ 420470.100000ns, VDD,
+ 420470.200000ns, VSS,
+ 420710.300000ns, VSS,
+ 420710.400000ns, VDD,
+ 421190.700000ns, VDD,
+ 421190.800000ns, VSS,
+ 421551.000000ns, VSS,
+ 421551.100000ns, VDD,
+ 422271.600000ns, VDD,
+ 422271.700000ns, VSS,
+ 422752.000000ns, VSS,
+ 422752.100000ns, VDD,
+ 422872.100000ns, VDD,
+ 422872.200000ns, VSS,
+ 423953.000000ns, VSS,
+ 423953.100000ns, VDD,
+ 426595.200000ns, VDD,
+ 426595.300000ns, VSS,
+ 428276.600000ns, VSS,
+ 428276.700000ns, VDD,
+ 428877.100000ns, VDD,
+ 428877.200000ns, VSS,
+ 428997.200000ns, VSS,
+ 428997.300000ns, VDD,
+ 429117.300000ns, VDD,
+ 429117.400000ns, VSS,
+ 429717.800000ns, VSS,
+ 429717.900000ns, VDD,
+ 430198.200000ns, VDD,
+ 430198.300000ns, VSS,
+ 430438.400000ns, VSS,
+ 430438.500000ns, VDD,
+ 432840.400000ns, VDD,
+ 432840.500000ns, VSS,
+ 433320.800000ns, VSS,
+ 433320.900000ns, VDD,
+ 436083.100000ns, VDD,
+ 436083.200000ns, VSS,
+ 436203.200000ns, VSS,
+ 436203.300000ns, VDD,
+ 437524.300000ns, VDD,
+ 437524.400000ns, VSS,
+ 437644.400000ns, VSS,
+ 437644.500000ns, VDD,
+ 438244.900000ns, VDD,
+ 438245.000000ns, VSS,
+ 438485.100000ns, VSS,
+ 438485.200000ns, VDD,
+ 438605.200000ns, VDD,
+ 438605.300000ns, VSS,
+ 438845.400000ns, VSS,
+ 438845.500000ns, VDD,
+ 438965.500000ns, VDD,
+ 438965.600000ns, VSS,
+ 439926.300000ns, VSS,
+ 439926.400000ns, VDD,
+ 441247.400000ns, VDD,
+ 441247.500000ns, VSS,
+ 441367.500000ns, VSS,
+ 441367.600000ns, VDD,
+ 441487.600000ns, VDD,
+ 441487.700000ns, VSS,
+ 441727.800000ns, VSS,
+ 441727.900000ns, VDD,
+ 442568.500000ns, VDD,
+ 442568.600000ns, VSS,
+ 442808.700000ns, VSS,
+ 442808.800000ns, VDD,
+ 443289.100000ns, VDD,
+ 443289.200000ns, VSS,
+ 443649.400000ns, VSS,
+ 443649.500000ns, VDD,
+ 443769.500000ns, VDD,
+ 443769.600000ns, VSS,
+ 444129.800000ns, VSS,
+ 444129.900000ns, VDD,
+ 445691.100000ns, VDD,
+ 445691.200000ns, VSS,
+ 445931.300000ns, VSS,
+ 445931.400000ns, VDD,
+ 446892.100000ns, VDD,
+ 446892.200000ns, VSS,
+ 447852.900000ns, VSS,
+ 447853.000000ns, VDD,
+ 448093.100000ns, VDD,
+ 448093.200000ns, VSS,
+ 448213.200000ns, VSS,
+ 448213.300000ns, VDD,
+ 448333.300000ns, VDD,
+ 448333.400000ns, VSS,
+ 449174.000000ns, VSS,
+ 449174.100000ns, VDD,
+ 449294.100000ns, VDD,
+ 449294.200000ns, VSS,
+ 449894.600000ns, VSS,
+ 449894.700000ns, VDD,
+ 450254.900000ns, VDD,
+ 450255.000000ns, VSS,
+ 451936.300000ns, VSS,
+ 451936.400000ns, VDD,
+ 452296.600000ns, VDD,
+ 452296.700000ns, VSS,
+ 453377.500000ns, VSS,
+ 453377.600000ns, VDD,
+ 453737.800000ns, VDD,
+ 453737.900000ns, VSS,
+ 453978.000000ns, VSS,
+ 453978.100000ns, VDD,
+ 454338.300000ns, VDD,
+ 454338.400000ns, VSS,
+ 454458.400000ns, VSS,
+ 454458.500000ns, VDD,
+ 455058.900000ns, VDD,
+ 455059.000000ns, VSS,
+ 455419.200000ns, VSS,
+ 455419.300000ns, VDD,
+ 455539.300000ns, VDD,
+ 455539.400000ns, VSS,
+ 455659.400000ns, VSS,
+ 455659.500000ns, VDD,
+ 456019.700000ns, VDD,
+ 456019.800000ns, VSS,
+ 456139.800000ns, VSS,
+ 456139.900000ns, VDD,
+ 458541.800000ns, VDD,
+ 458541.900000ns, VSS,
+ 458902.100000ns, VSS,
+ 458902.200000ns, VDD,
+ 459622.700000ns, VDD,
+ 459622.800000ns, VSS,
+ 460463.400000ns, VSS,
+ 460463.500000ns, VDD,
+ 461063.900000ns, VDD,
+ 461064.000000ns, VSS,
+ 462144.800000ns, VSS,
+ 462144.900000ns, VDD,
+ 462625.200000ns, VDD,
+ 462625.300000ns, VSS,
+ 463586.000000ns, VSS,
+ 463586.100000ns, VDD,
+ 463946.300000ns, VDD,
+ 463946.400000ns, VSS,
+ 464546.800000ns, VSS,
+ 464546.900000ns, VDD,
+ 465627.700000ns, VDD,
+ 465627.800000ns, VSS,
+ 465867.900000ns, VSS,
+ 465868.000000ns, VDD,
+ 466468.400000ns, VDD,
+ 466468.500000ns, VSS,
+ 466708.600000ns, VSS,
+ 466708.700000ns, VDD,
+ 466948.800000ns, VDD,
+ 466948.900000ns, VSS,
+ 468029.700000ns, VSS,
+ 468029.800000ns, VDD,
+ 468269.900000ns, VDD,
+ 468270.000000ns, VSS,
+ 468510.100000ns, VSS,
+ 468510.200000ns, VDD,
+ 470431.700000ns, VDD,
+ 470431.800000ns, VSS,
+ 470912.100000ns, VSS,
+ 470912.200000ns, VDD,
+ 471392.500000ns, VDD,
+ 471392.600000ns, VSS,
+ 472113.100000ns, VSS,
+ 472113.200000ns, VDD,
+ 472473.400000ns, VDD,
+ 472473.500000ns, VSS,
+ 473434.200000ns, VSS,
+ 473434.300000ns, VDD,
+ 473554.300000ns, VDD,
+ 473554.400000ns, VSS,
+ 474154.800000ns, VSS,
+ 474154.900000ns, VDD,
+ 475235.700000ns, VDD,
+ 475235.800000ns, VSS,
+ 475716.100000ns, VSS,
+ 475716.200000ns, VDD,
+ 477757.800000ns, VDD,
+ 477757.900000ns, VSS,
+ 478358.300000ns, VSS,
+ 478358.400000ns, VDD,
+ 478958.800000ns, VDD,
+ 478958.900000ns, VSS,
+ 480760.300000ns, VSS,
+ 480760.400000ns, VDD,
+ 482081.400000ns, VDD,
+ 482081.500000ns, VSS,
+ 482321.600000ns, VSS,
+ 482321.700000ns, VDD,
+ 482441.700000ns, VDD,
+ 482441.800000ns, VSS,
+ 483402.500000ns, VSS,
+ 483402.600000ns, VDD,
+ 484363.300000ns, VDD,
+ 484363.400000ns, VSS,
+ 484723.600000ns, VSS,
+ 484723.700000ns, VDD,
+ 484843.700000ns, VDD,
+ 484843.800000ns, VSS,
+ 485684.400000ns, VSS,
+ 485684.500000ns, VDD,
+ 486284.900000ns, VDD,
+ 486285.000000ns, VSS,
+ 487005.500000ns, VSS,
+ 487005.600000ns, VDD,
+ 487125.600000ns, VDD,
+ 487125.700000ns, VSS,
+ 489047.200000ns, VSS,
+ 489047.300000ns, VDD,
+ 489527.600000ns, VDD,
+ 489527.700000ns, VSS,
+ 490368.300000ns, VSS,
+ 490368.400000ns, VDD,
+ 491449.200000ns, VDD,
+ 491449.300000ns, VSS,
+ 491809.500000ns, VSS,
+ 491809.600000ns, VDD,
+ 492289.900000ns, VDD,
+ 492290.000000ns, VSS,
+ 492650.200000ns, VSS,
+ 492650.300000ns, VDD,
+ 493010.500000ns, VDD,
+ 493010.600000ns, VSS,
+ 495532.600000ns, VSS,
+ 495532.700000ns, VDD,
+ 496133.100000ns, VDD,
+ 496133.200000ns, VSS,
+ 496613.500000ns, VSS,
+ 496613.600000ns, VDD,
+ 497214.000000ns, VDD,
+ 497214.100000ns, VSS,
+ 497574.300000ns, VSS,
+ 497574.400000ns, VDD,
+ 498294.900000ns, VDD,
+ 498295.000000ns, VSS,
+ 498535.100000ns, VSS,
+ 498535.200000ns, VDD,
+ 499736.100000ns, VDD,
+ 499736.200000ns, VSS,
+ 500096.400000ns, VSS,
+ 500096.500000ns, VDD,
+ 502018.000000ns, VDD,
+ 502018.100000ns, VSS,
+ 503579.300000ns, VSS,
+ 503579.400000ns, VDD,
+ 505861.200000ns, VDD,
+ 505861.300000ns, VSS,
+ 506221.500000ns, VSS,
+ 506221.600000ns, VDD,
+ 506581.800000ns, VDD,
+ 506581.900000ns, VSS,
+ 508023.000000ns, VSS,
+ 508023.100000ns, VDD,
+ 508143.100000ns, VDD,
+ 508143.200000ns, VSS,
+ 508503.400000ns, VSS,
+ 508503.500000ns, VDD,
+ 509224.000000ns, VDD,
+ 509224.100000ns, VSS,
+ 509704.400000ns, VSS,
+ 509704.500000ns, VDD,
+ 509944.600000ns, VDD,
+ 509944.700000ns, VSS,
+ 510785.300000ns, VSS,
+ 510785.400000ns, VDD,
+ 511986.300000ns, VDD,
+ 511986.400000ns, VSS,
+ 513187.300000ns, VSS,
+ 513187.400000ns, VDD,
+ 513547.600000ns, VDD,
+ 513547.700000ns, VSS,
+ 513907.900000ns, VSS,
+ 513908.000000ns, VDD,
+ 514628.500000ns, VDD,
+ 514628.600000ns, VSS,
+ 514868.700000ns, VSS,
+ 514868.800000ns, VDD,
+ 515829.500000ns, VDD,
+ 515829.600000ns, VSS,
+ 516309.900000ns, VSS,
+ 516310.000000ns, VDD,
+ 516790.300000ns, VDD,
+ 516790.400000ns, VSS,
+ 517270.700000ns, VSS,
+ 517270.800000ns, VDD,
+ 517510.900000ns, VDD,
+ 517511.000000ns, VSS,
+ 517631.000000ns, VSS,
+ 517631.100000ns, VDD,
+ 518111.400000ns, VDD,
+ 518111.500000ns, VSS,
+ 518711.900000ns, VSS,
+ 518712.000000ns, VDD,
+ 518952.100000ns, VDD,
+ 518952.200000ns, VSS,
+ 519192.300000ns, VSS,
+ 519192.400000ns, VDD,
+ 519432.500000ns, VDD,
+ 519432.600000ns, VSS,
+ 519792.800000ns, VSS,
+ 519792.900000ns, VDD,
+ 520153.100000ns, VDD,
+ 520153.200000ns, VSS,
+ 520273.200000ns, VSS,
+ 520273.300000ns, VDD,
+ 520753.600000ns, VDD,
+ 520753.700000ns, VSS,
+ 520993.800000ns, VSS,
+ 520993.900000ns, VDD,
+ 521234.000000ns, VDD,
+ 521234.100000ns, VSS,
+ 521954.600000ns, VSS,
+ 521954.700000ns, VDD,
+ 522435.000000ns, VDD,
+ 522435.100000ns, VSS,
+ 522915.400000ns, VSS,
+ 522915.500000ns, VDD,
+ 525077.200000ns, VDD,
+ 525077.300000ns, VSS,
+ 525317.400000ns, VSS,
+ 525317.500000ns, VDD,
+ 527359.100000ns, VDD,
+ 527359.200000ns, VSS,
+ 527479.200000ns, VSS,
+ 527479.300000ns, VDD,
+ 528440.000000ns, VDD,
+ 528440.100000ns, VSS,
+ 528560.100000ns, VSS,
+ 528560.200000ns, VDD,
+ 528680.200000ns, VDD,
+ 528680.300000ns, VSS,
+ 528800.300000ns, VSS,
+ 528800.400000ns, VDD,
+ 529400.800000ns, VDD,
+ 529400.900000ns, VSS,
+ 530121.400000ns, VSS,
+ 530121.500000ns, VDD,
+ 531082.200000ns, VDD,
+ 531082.300000ns, VSS,
+ 531922.900000ns, VSS,
+ 531923.000000ns, VDD,
+ 532043.000000ns, VDD,
+ 532043.100000ns, VSS,
+ 532643.500000ns, VSS,
+ 532643.600000ns, VDD,
+ 533123.900000ns, VDD,
+ 533124.000000ns, VSS,
+ 534925.400000ns, VSS,
+ 534925.500000ns, VDD,
+ 535285.700000ns, VDD,
+ 535285.800000ns, VSS,
+ 536126.400000ns, VSS,
+ 536126.500000ns, VDD,
+ 536366.600000ns, VDD,
+ 536366.700000ns, VSS,
+ 536486.700000ns, VSS,
+ 536486.800000ns, VDD,
+ 536967.100000ns, VDD,
+ 536967.200000ns, VSS,
+ 537207.300000ns, VSS,
+ 537207.400000ns, VDD,
+ 537327.400000ns, VDD,
+ 537327.500000ns, VSS,
+ 538288.200000ns, VSS,
+ 538288.300000ns, VDD,
+ 538648.500000ns, VDD,
+ 538648.600000ns, VSS,
+ 539609.300000ns, VSS,
+ 539609.400000ns, VDD,
+ 539969.600000ns, VDD,
+ 539969.700000ns, VSS,
+ 541891.200000ns, VSS,
+ 541891.300000ns, VDD,
+ 542611.800000ns, VDD,
+ 542611.900000ns, VSS,
+ 543092.200000ns, VSS,
+ 543092.300000ns, VDD,
+ 543212.300000ns, VDD,
+ 543212.400000ns, VSS,
+ 544293.200000ns, VSS,
+ 544293.300000ns, VDD,
+ 546935.400000ns, VDD,
+ 546935.500000ns, VSS,
+ 548016.300000ns, VSS,
+ 548016.400000ns, VDD,
+ 549337.400000ns, VDD,
+ 549337.500000ns, VSS,
+ 549817.800000ns, VSS,
+ 549817.900000ns, VDD,
+ 550418.300000ns, VDD,
+ 550418.400000ns, VSS,
+ 550658.500000ns, VSS,
+ 550658.600000ns, VDD,
+ 551379.100000ns, VDD,
+ 551379.200000ns, VSS,
+ 551499.200000ns, VSS,
+ 551499.300000ns, VDD,
+ 552820.300000ns, VDD,
+ 552820.400000ns, VSS,
+ 553420.800000ns, VSS,
+ 553420.900000ns, VDD,
+ 554862.000000ns, VDD,
+ 554862.100000ns, VSS,
+ 555462.500000ns, VSS,
+ 555462.600000ns, VDD,
+ 556063.000000ns, VDD,
+ 556063.100000ns, VSS,
+ 556183.100000ns, VSS,
+ 556183.200000ns, VDD,
+ 556783.600000ns, VDD,
+ 556783.700000ns, VSS,
+ 557143.900000ns, VSS,
+ 557144.000000ns, VDD,
+ 557384.100000ns, VDD,
+ 557384.200000ns, VSS,
+ 557504.200000ns, VSS,
+ 557504.300000ns, VDD,
+ 557624.300000ns, VDD,
+ 557624.400000ns, VSS,
+ 558224.800000ns, VSS,
+ 558224.900000ns, VDD,
+ 558585.100000ns, VDD,
+ 558585.200000ns, VSS,
+ 558825.300000ns, VSS,
+ 558825.400000ns, VDD,
+ 559065.500000ns, VDD,
+ 559065.600000ns, VSS,
+ 560626.800000ns, VSS,
+ 560626.900000ns, VDD,
+ 561467.500000ns, VDD,
+ 561467.600000ns, VSS,
+ 562188.100000ns, VSS,
+ 562188.200000ns, VDD,
+ 562548.400000ns, VDD,
+ 562548.500000ns, VSS,
+ 562908.700000ns, VSS,
+ 562908.800000ns, VDD,
+ 563028.800000ns, VDD,
+ 563028.900000ns, VSS,
+ 565310.700000ns, VSS,
+ 565310.800000ns, VDD,
+ 566511.700000ns, VDD,
+ 566511.800000ns, VSS,
+ 566872.000000ns, VSS,
+ 566872.100000ns, VDD,
+ 568193.100000ns, VDD,
+ 568193.200000ns, VSS,
+ 568433.300000ns, VSS,
+ 568433.400000ns, VDD,
+ 569754.400000ns, VDD,
+ 569754.500000ns, VSS,
+ 570114.700000ns, VSS,
+ 570114.800000ns, VDD,
+ 570595.100000ns, VDD,
+ 570595.200000ns, VSS,
+ 570835.300000ns, VSS,
+ 570835.400000ns, VDD,
+ 571195.600000ns, VDD,
+ 571195.700000ns, VSS,
+ 572756.900000ns, VSS,
+ 572757.000000ns, VDD,
+ 572877.000000ns, VDD,
+ 572877.100000ns, VSS,
+ 573117.200000ns, VSS,
+ 573117.300000ns, VDD,
+ 573237.300000ns, VDD,
+ 573237.400000ns, VSS,
+ 573597.600000ns, VSS,
+ 573597.700000ns, VDD,
+ 573717.700000ns, VDD,
+ 573717.800000ns, VSS,
+ 573957.900000ns, VSS,
+ 573958.000000ns, VDD,
+ 574078.000000ns, VDD,
+ 574078.100000ns, VSS,
+ 574918.700000ns, VSS,
+ 574918.800000ns, VDD,
+ 575158.900000ns, VDD,
+ 575159.000000ns, VSS,
+ 575399.100000ns, VSS,
+ 575399.200000ns, VDD,
+ 575519.200000ns, VDD,
+ 575519.300000ns, VSS,
+ 575759.400000ns, VSS,
+ 575759.500000ns, VDD,
+ 576239.800000ns, VDD,
+ 576239.900000ns, VSS,
+ 576720.200000ns, VSS,
+ 576720.300000ns, VDD,
+ 577681.000000ns, VDD,
+ 577681.100000ns, VSS,
+ 578281.500000ns, VSS,
+ 578281.600000ns, VDD,
+ 578882.000000ns, VDD,
+ 578882.100000ns, VSS,
+ 579722.700000ns, VSS,
+ 579722.800000ns, VDD,
+ 579842.800000ns, VDD,
+ 579842.900000ns, VSS,
+ 580803.600000ns, VSS,
+ 580803.700000ns, VDD,
+ 582124.700000ns, VDD,
+ 582124.800000ns, VSS,
+ 582845.300000ns, VSS,
+ 582845.400000ns, VDD,
+ 583085.500000ns, VDD,
+ 583085.600000ns, VSS,
+ 584286.500000ns, VSS,
+ 584286.600000ns, VDD,
+ 585247.300000ns, VDD,
+ 585247.400000ns, VSS,
+ 585367.400000ns, VSS,
+ 585367.500000ns, VDD,
+ 585847.800000ns, VDD,
+ 585847.900000ns, VSS,
+ 586208.100000ns, VSS,
+ 586208.200000ns, VDD,
+ 587529.200000ns, VDD,
+ 587529.300000ns, VSS,
+ 587769.400000ns, VSS,
+ 587769.500000ns, VDD,
+ 588490.000000ns, VDD,
+ 588490.100000ns, VSS,
+ 589090.500000ns, VSS,
+ 589090.600000ns, VDD,
+ 589691.000000ns, VDD,
+ 589691.100000ns, VSS,
+ 590171.400000ns, VSS,
+ 590171.500000ns, VDD,
+ 590771.900000ns, VDD,
+ 590772.000000ns, VSS,
+ 591612.600000ns, VSS,
+ 591612.700000ns, VDD,
+ 592093.000000ns, VDD,
+ 592093.100000ns, VSS,
+ 593053.800000ns, VSS,
+ 593053.900000ns, VDD,
+ 593534.200000ns, VDD,
+ 593534.300000ns, VSS,
+ 594254.800000ns, VSS,
+ 594254.900000ns, VDD,
+ 594374.900000ns, VDD,
+ 594375.000000ns, VSS,
+ 594855.300000ns, VSS,
+ 594855.400000ns, VDD,
+ 595095.500000ns, VDD,
+ 595095.600000ns, VSS,
+ 595335.700000ns, VSS,
+ 595335.800000ns, VDD,
+ 595575.900000ns, VDD,
+ 595576.000000ns, VSS,
+ 595696.000000ns, VSS,
+ 595696.100000ns, VDD,
+ 595936.200000ns, VDD,
+ 595936.300000ns, VSS,
+ 596776.900000ns, VSS,
+ 596777.000000ns, VDD,
+ 598578.400000ns, VDD,
+ 598578.500000ns, VSS,
+ 599779.400000ns, VSS,
+ 599779.500000ns, VDD,
+ 600259.800000ns, VDD,
+ 600259.900000ns, VSS,
+ 600500.000000ns, VSS,
+ 600500.100000ns, VDD,
+ 601340.700000ns, VDD,
+ 601340.800000ns, VSS,
+ 601460.800000ns, VSS,
+ 601460.900000ns, VDD,
+ 601580.900000ns, VDD,
+ 601581.000000ns, VSS,
+ 602781.900000ns, VSS,
+ 602782.000000ns, VDD,
+ 603262.300000ns, VDD,
+ 603262.400000ns, VSS,
+ 603502.500000ns, VSS,
+ 603502.600000ns, VDD,
+ 603742.700000ns, VDD,
+ 603742.800000ns, VSS,
+ 604103.000000ns, VSS,
+ 604103.100000ns, VDD,
+ 604343.200000ns, VDD,
+ 604343.300000ns, VSS,
+ 604583.400000ns, VSS,
+ 604583.500000ns, VDD,
+ 605304.000000ns, VDD,
+ 605304.100000ns, VSS,
+ 605784.400000ns, VSS,
+ 605784.500000ns, VDD,
+ 606384.900000ns, VDD,
+ 606385.000000ns, VSS,
+ 606505.000000ns, VSS,
+ 606505.100000ns, VDD,
+ 606625.100000ns, VDD,
+ 606625.200000ns, VSS,
+ 607225.600000ns, VSS,
+ 607225.700000ns, VDD,
+ 607465.800000ns, VDD,
+ 607465.900000ns, VSS,
+ 607585.900000ns, VSS,
+ 607586.000000ns, VDD,
+ 607826.100000ns, VDD,
+ 607826.200000ns, VSS,
+ 607946.200000ns, VSS,
+ 607946.300000ns, VDD,
+ 608306.500000ns, VDD,
+ 608306.600000ns, VSS,
+ 608786.900000ns, VSS,
+ 608787.000000ns, VDD,
+ 609507.500000ns, VDD,
+ 609507.600000ns, VSS,
+ 609987.900000ns, VSS,
+ 609988.000000ns, VDD,
+ 610348.200000ns, VDD,
+ 610348.300000ns, VSS,
+ 612750.200000ns, VSS,
+ 612750.300000ns, VDD,
+ 613951.200000ns, VDD,
+ 613951.300000ns, VSS,
+ 614671.800000ns, VSS,
+ 614671.900000ns, VDD,
+ 614912.000000ns, VDD,
+ 614912.100000ns, VSS,
+ 615752.700000ns, VSS,
+ 615752.800000ns, VDD,
+ 615992.900000ns, VDD,
+ 615993.000000ns, VSS,
+ 616233.100000ns, VSS,
+ 616233.200000ns, VDD,
+ 616353.200000ns, VDD,
+ 616353.300000ns, VSS,
+ 616473.300000ns, VSS,
+ 616473.400000ns, VDD,
+ 617554.200000ns, VDD,
+ 617554.300000ns, VSS,
+ 618034.600000ns, VSS,
+ 618034.700000ns, VDD,
+ 619355.700000ns, VDD,
+ 619355.800000ns, VSS,
+ 619475.800000ns, VSS,
+ 619475.900000ns, VDD,
+ 620556.700000ns, VDD,
+ 620556.800000ns, VSS,
+ 621277.300000ns, VSS,
+ 621277.400000ns, VDD,
+ 622118.000000ns, VDD,
+ 622118.100000ns, VSS,
+ 622358.200000ns, VSS,
+ 622358.300000ns, VDD,
+ 622958.700000ns, VDD,
+ 622958.800000ns, VSS,
+ 623319.000000ns, VSS,
+ 623319.100000ns, VDD,
+ 623679.300000ns, VDD,
+ 623679.400000ns, VSS,
+ 624039.600000ns, VSS,
+ 624039.700000ns, VDD,
+ 624279.800000ns, VDD,
+ 624279.900000ns, VSS,
+ 625120.500000ns, VSS,
+ 625120.600000ns, VDD,
+ 626201.400000ns, VDD,
+ 626201.500000ns, VSS,
+ 626681.800000ns, VSS,
+ 626681.900000ns, VDD,
+ 626801.900000ns, VDD,
+ 626802.000000ns, VSS,
+ 627882.800000ns, VSS,
+ 627882.900000ns, VDD,
+ 628843.600000ns, VDD,
+ 628843.700000ns, VSS,
+ 628963.700000ns, VSS,
+ 628963.800000ns, VDD,
+ 629444.100000ns, VDD,
+ 629444.200000ns, VSS,
+ 629564.200000ns, VSS,
+ 629564.300000ns, VDD,
+ 629684.300000ns, VDD,
+ 629684.400000ns, VSS,
+ 629924.500000ns, VSS,
+ 629924.600000ns, VDD,
+ 630885.300000ns, VDD,
+ 630885.400000ns, VSS,
+ 631125.500000ns, VSS,
+ 631125.600000ns, VDD,
+ 631846.100000ns, VDD,
+ 631846.200000ns, VSS,
+ 632806.900000ns, VSS,
+ 632807.000000ns, VDD,
+ 633167.200000ns, VDD,
+ 633167.300000ns, VSS,
+ 633767.700000ns, VSS,
+ 633767.800000ns, VDD,
+ 633887.800000ns, VDD,
+ 633887.900000ns, VSS,
+ 634368.200000ns, VSS,
+ 634368.300000ns, VDD,
+ 634968.700000ns, VDD,
+ 634968.800000ns, VSS,
+ 635929.500000ns, VSS,
+ 635929.600000ns, VDD,
+ 636049.600000ns, VDD,
+ 636049.700000ns, VSS,
+ 637490.800000ns, VSS,
+ 637490.900000ns, VDD,
+ 637731.000000ns, VDD,
+ 637731.100000ns, VSS,
+ 637971.200000ns, VSS,
+ 637971.300000ns, VDD,
+ 638451.600000ns, VDD,
+ 638451.700000ns, VSS,
+ 638811.900000ns, VSS,
+ 638812.000000ns, VDD,
+ 639412.400000ns, VDD,
+ 639412.500000ns, VSS,
+ 639892.800000ns, VSS,
+ 639892.900000ns, VDD,
+ 640253.100000ns, VDD,
+ 640253.200000ns, VSS,
+ 641454.100000ns, VSS,
+ 641454.200000ns, VDD,
+ 642895.300000ns, VDD,
+ 642895.400000ns, VSS,
+ 643495.800000ns, VSS,
+ 643495.900000ns, VDD,
+ 644456.600000ns, VDD,
+ 644456.700000ns, VSS,
+ 644816.900000ns, VSS,
+ 644817.000000ns, VDD,
+ 645297.300000ns, VDD,
+ 645297.400000ns, VSS,
+ 645417.400000ns, VSS,
+ 645417.500000ns, VDD,
+ 645777.700000ns, VDD,
+ 645777.800000ns, VSS,
+ 645897.800000ns, VSS,
+ 645897.900000ns, VDD,
+ 646978.700000ns, VDD,
+ 646978.800000ns, VSS,
+ 647218.900000ns, VSS,
+ 647219.000000ns, VDD,
+ 647819.400000ns, VDD,
+ 647819.500000ns, VSS,
+ 647939.500000ns, VSS,
+ 647939.600000ns, VDD,
+ 648059.600000ns, VDD,
+ 648059.700000ns, VSS,
+ 648419.900000ns, VSS,
+ 648420.000000ns, VDD,
+ 649260.600000ns, VDD,
+ 649260.700000ns, VSS,
+ 649620.900000ns, VSS,
+ 649621.000000ns, VDD,
+ 649741.000000ns, VDD,
+ 649741.100000ns, VSS,
+ 649981.200000ns, VSS,
+ 649981.300000ns, VDD,
+ 650101.300000ns, VDD,
+ 650101.400000ns, VSS,
+ 650701.800000ns, VSS,
+ 650701.900000ns, VDD,
+ 651662.600000ns, VDD,
+ 651662.700000ns, VSS,
+ 651782.700000ns, VSS,
+ 651782.800000ns, VDD,
+ 652263.100000ns, VDD,
+ 652263.200000ns, VSS,
+ 652623.400000ns, VSS,
+ 652623.500000ns, VDD,
+ 653103.800000ns, VDD,
+ 653103.900000ns, VSS,
+ 653704.300000ns, VSS,
+ 653704.400000ns, VDD,
+ 654304.800000ns, VDD,
+ 654304.900000ns, VSS,
+ 655385.700000ns, VSS,
+ 655385.800000ns, VDD,
+ 655625.900000ns, VDD,
+ 655626.000000ns, VSS,
+ 655746.000000ns, VSS,
+ 655746.100000ns, VDD,
+ 656947.000000ns, VDD,
+ 656947.100000ns, VSS,
+ 657187.200000ns, VSS,
+ 657187.300000ns, VDD,
+ 657547.500000ns, VDD,
+ 657547.600000ns, VSS,
+ 657787.700000ns, VSS,
+ 657787.800000ns, VDD,
+ 658268.100000ns, VDD,
+ 658268.200000ns, VSS,
+ 658628.400000ns, VSS,
+ 658628.500000ns, VDD,
+ 659349.000000ns, VDD,
+ 659349.100000ns, VSS,
+ 659829.400000ns, VSS,
+ 659829.500000ns, VDD,
+ 660189.700000ns, VDD,
+ 660189.800000ns, VSS,
+ 660670.100000ns, VSS,
+ 660670.200000ns, VDD,
+ 660910.300000ns, VDD,
+ 660910.400000ns, VSS,
+ 661030.400000ns, VSS,
+ 661030.500000ns, VDD,
+ 661751.000000ns, VDD,
+ 661751.100000ns, VSS,
+ 661991.200000ns, VSS,
+ 661991.300000ns, VDD,
+ 662711.800000ns, VDD,
+ 662711.900000ns, VSS,
+ 663912.800000ns, VSS,
+ 663912.900000ns, VDD,
+ 664032.900000ns, VDD,
+ 664033.000000ns, VSS,
+ 665954.500000ns, VSS,
+ 665954.600000ns, VDD,
+ 666314.800000ns, VDD,
+ 666314.900000ns, VSS,
+ 666675.100000ns, VSS,
+ 666675.200000ns, VDD,
+ 668476.600000ns, VDD,
+ 668476.700000ns, VSS,
+ 668596.700000ns, VSS,
+ 668596.800000ns, VDD,
+ 668716.800000ns, VDD,
+ 668716.900000ns, VSS,
+ 669917.800000ns, VSS,
+ 669917.900000ns, VDD,
+ 670037.900000ns, VDD,
+ 670038.000000ns, VSS,
+ 670518.300000ns, VSS,
+ 670518.400000ns, VDD,
+ 671599.200000ns, VDD,
+ 671599.300000ns, VSS,
+ 673761.000000ns, VSS,
+ 673761.100000ns, VDD,
+ 674001.200000ns, VDD,
+ 674001.300000ns, VSS,
+ 674121.300000ns, VSS,
+ 674121.400000ns, VDD,
+ 674241.400000ns, VDD,
+ 674241.500000ns, VSS,
+ 674721.800000ns, VSS,
+ 674721.900000ns, VDD,
+ 674841.900000ns, VDD,
+ 674842.000000ns, VSS,
+ 675322.300000ns, VSS,
+ 675322.400000ns, VDD,
+ 675682.600000ns, VDD,
+ 675682.700000ns, VSS,
+ 676643.400000ns, VSS,
+ 676643.500000ns, VDD,
+ 677364.000000ns, VDD,
+ 677364.100000ns, VSS,
+ 679766.000000ns, VSS,
+ 679766.100000ns, VDD,
+ 680486.600000ns, VDD,
+ 680486.700000ns, VSS,
+ 680846.900000ns, VSS,
+ 680847.000000ns, VDD,
+ 683609.200000ns, VDD,
+ 683609.300000ns, VSS,
+ 684690.100000ns, VSS,
+ 684690.200000ns, VDD,
+ 685530.800000ns, VDD,
+ 685530.900000ns, VSS,
+ 686731.800000ns, VSS,
+ 686731.900000ns, VDD,
+ 687332.300000ns, VDD,
+ 687332.400000ns, VSS,
+ 688413.200000ns, VSS,
+ 688413.300000ns, VDD,
+ 688533.300000ns, VDD,
+ 688533.400000ns, VSS,
+ 689013.700000ns, VSS,
+ 689013.800000ns, VDD,
+ 689374.000000ns, VDD,
+ 689374.100000ns, VSS,
+ 690214.700000ns, VSS,
+ 690214.800000ns, VDD,
+ 690454.900000ns, VDD,
+ 690455.000000ns, VSS,
+ 690815.200000ns, VSS,
+ 690815.300000ns, VDD,
+ 691415.700000ns, VDD,
+ 691415.800000ns, VSS,
+ 691776.000000ns, VSS,
+ 691776.100000ns, VDD,
+ 692256.400000ns, VDD,
+ 692256.500000ns, VSS,
+ 692736.800000ns, VSS,
+ 692736.900000ns, VDD,
+ 693457.400000ns, VDD,
+ 693457.500000ns, VSS,
+ 694418.200000ns, VSS,
+ 694418.300000ns, VDD,
+ 696219.700000ns, VDD,
+ 696219.800000ns, VSS,
+ 697781.000000ns, VSS,
+ 697781.100000ns, VDD,
+ 698261.400000ns, VDD,
+ 698261.500000ns, VSS,
+ 698982.000000ns, VSS,
+ 698982.100000ns, VDD,
+ 699342.300000ns, VDD,
+ 699342.400000ns, VSS,
+ 700783.500000ns, VSS,
+ 700783.600000ns, VDD,
+ 701023.700000ns, VDD,
+ 701023.800000ns, VSS,
+ 702464.900000ns, VSS,
+ 702465.000000ns, VDD,
+ 703065.400000ns, VDD,
+ 703065.500000ns, VSS,
+ 703185.500000ns, VSS,
+ 703185.600000ns, VDD,
+ 705107.100000ns, VDD,
+ 705107.200000ns, VSS,
+ 705347.300000ns, VSS,
+ 705347.400000ns, VDD,
+ 705467.400000ns, VDD,
+ 705467.500000ns, VSS,
+ 706548.300000ns, VSS,
+ 706548.400000ns, VDD,
+ 707148.800000ns, VDD,
+ 707148.900000ns, VSS,
+ 707509.100000ns, VSS,
+ 707509.200000ns, VDD,
+ 707989.500000ns, VDD,
+ 707989.600000ns, VSS,
+ 708830.200000ns, VSS,
+ 708830.300000ns, VDD,
+ 709070.400000ns, VDD,
+ 709070.500000ns, VSS,
+ 709550.800000ns, VSS,
+ 709550.900000ns, VDD,
+ 711112.100000ns, VDD,
+ 711112.200000ns, VSS,
+ 712072.900000ns, VSS,
+ 712073.000000ns, VDD,
+ 712553.300000ns, VDD,
+ 712553.400000ns, VSS,
+ 712673.400000ns, VSS,
+ 712673.500000ns, VDD,
+ 712913.600000ns, VDD,
+ 712913.700000ns, VSS,
+ 713153.800000ns, VSS,
+ 713153.900000ns, VDD,
+ 713634.200000ns, VDD,
+ 713634.300000ns, VSS,
+ 714595.000000ns, VSS,
+ 714595.100000ns, VDD,
+ 714715.100000ns, VDD,
+ 714715.200000ns, VSS,
+ 714955.300000ns, VSS,
+ 714955.400000ns, VDD,
+ 715435.700000ns, VDD,
+ 715435.800000ns, VSS,
+ 715916.100000ns, VSS,
+ 715916.200000ns, VDD,
+ 716156.300000ns, VDD,
+ 716156.400000ns, VSS,
+ 716276.400000ns, VSS,
+ 716276.500000ns, VDD,
+ 716636.700000ns, VDD,
+ 716636.800000ns, VSS,
+ 717117.100000ns, VSS,
+ 717117.200000ns, VDD,
+ 718558.300000ns, VDD,
+ 718558.400000ns, VSS,
+ 719278.900000ns, VSS,
+ 719279.000000ns, VDD,
+ 720359.800000ns, VDD,
+ 720359.900000ns, VSS,
+ 720600.000000ns, VSS,
+ 720600.100000ns, VDD,
+ 720960.300000ns, VDD,
+ 720960.400000ns, VSS,
+ 722041.200000ns, VSS,
+ 722041.300000ns, VDD,
+ 722521.600000ns, VDD,
+ 722521.700000ns, VSS,
+ 724443.200000ns, VSS,
+ 724443.300000ns, VDD,
+ 726364.800000ns, VDD,
+ 726364.900000ns, VSS,
+ 727325.600000ns, VSS,
+ 727325.700000ns, VDD,
+ 728646.700000ns, VDD,
+ 728646.800000ns, VSS,
+ 729007.000000ns, VSS,
+ 729007.100000ns, VDD,
+ 729727.600000ns, VDD,
+ 729727.700000ns, VSS,
+ 729967.800000ns, VSS,
+ 729967.900000ns, VDD,
+ 730328.100000ns, VDD,
+ 730328.200000ns, VSS,
+ 730448.200000ns, VSS,
+ 730448.300000ns, VDD,
+ 730568.300000ns, VDD,
+ 730568.400000ns, VSS,
+ 733690.900000ns, VSS,
+ 733691.000000ns, VDD,
+ 734411.500000ns, VDD,
+ 734411.600000ns, VSS,
+ 735972.800000ns, VSS,
+ 735972.900000ns, VDD,
+ 736573.300000ns, VDD,
+ 736573.400000ns, VSS,
+ 738134.600000ns, VSS,
+ 738134.700000ns, VDD,
+ 738735.100000ns, VDD,
+ 738735.200000ns, VSS,
+ 738855.200000ns, VSS,
+ 738855.300000ns, VDD,
+ 739095.400000ns, VDD,
+ 739095.500000ns, VSS,
+ 739816.000000ns, VSS,
+ 739816.100000ns, VDD,
+ 740056.200000ns, VDD,
+ 740056.300000ns, VSS,
+ 740176.300000ns, VSS,
+ 740176.400000ns, VDD,
+ 740776.800000ns, VDD,
+ 740776.900000ns, VSS,
+ 741737.600000ns, VSS,
+ 741737.700000ns, VDD,
+ 743178.800000ns, VDD,
+ 743178.900000ns, VSS,
+ 743659.200000ns, VSS,
+ 743659.300000ns, VDD,
+ 744019.500000ns, VDD,
+ 744019.600000ns, VSS,
+ 744620.000000ns, VSS,
+ 744620.100000ns, VDD,
+ 745340.600000ns, VDD,
+ 745340.700000ns, VSS,
+ 746781.800000ns, VSS,
+ 746781.900000ns, VDD,
+ 748583.300000ns, VDD,
+ 748583.400000ns, VSS,
+ 748943.600000ns, VSS,
+ 748943.700000ns, VDD,
+ 749303.900000ns, VDD,
+ 749304.000000ns, VSS,
+ 749664.200000ns, VSS,
+ 749664.300000ns, VDD,
+ 749784.300000ns, VDD,
+ 749784.400000ns, VSS,
+ 750264.700000ns, VSS,
+ 750264.800000ns, VDD,
+ 751345.600000ns, VDD,
+ 751345.700000ns, VSS,
+ 752186.300000ns, VSS,
+ 752186.400000ns, VDD,
+ 752426.500000ns, VDD,
+ 752426.600000ns, VSS,
+ 752906.900000ns, VSS,
+ 752907.000000ns, VDD,
+ 753147.100000ns, VDD,
+ 753147.200000ns, VSS,
+ 753267.200000ns, VSS,
+ 753267.300000ns, VDD,
+ 754828.500000ns, VDD,
+ 754828.600000ns, VSS,
+ 755068.700000ns, VSS,
+ 755068.800000ns, VDD,
+ 755308.900000ns, VDD,
+ 755309.000000ns, VSS,
+ 756029.500000ns, VSS,
+ 756029.600000ns, VDD,
+ 756389.800000ns, VDD,
+ 756389.900000ns, VSS,
+ 756750.100000ns, VSS,
+ 756750.200000ns, VDD,
+ 756990.300000ns, VDD,
+ 756990.400000ns, VSS,
+ 758071.200000ns, VSS,
+ 758071.300000ns, VDD,
+ 760953.600000ns, VDD,
+ 760953.700000ns, VSS,
+ 761434.000000ns, VSS,
+ 761434.100000ns, VDD,
+ 762635.000000ns, VDD,
+ 762635.100000ns, VSS,
+ 762995.300000ns, VSS,
+ 762995.400000ns, VDD,
+ 763355.600000ns, VDD,
+ 763355.700000ns, VSS,
+ 764436.500000ns, VSS,
+ 764436.600000ns, VDD,
+ 765277.200000ns, VDD,
+ 765277.300000ns, VSS,
+ 765877.700000ns, VSS,
+ 765877.800000ns, VDD,
+ 768279.700000ns, VDD,
+ 768279.800000ns, VSS,
+ 768760.100000ns, VSS,
+ 768760.200000ns, VDD,
+ 769600.800000ns, VDD,
+ 769600.900000ns, VSS,
+ 769841.000000ns, VSS,
+ 769841.100000ns, VDD,
+ 770081.200000ns, VDD,
+ 770081.300000ns, VSS,
+ 770561.600000ns, VSS,
+ 770561.700000ns, VDD,
+ 770681.700000ns, VDD,
+ 770681.800000ns, VSS,
+ 770801.800000ns, VSS,
+ 770801.900000ns, VDD,
+ 771282.200000ns, VDD,
+ 771282.300000ns, VSS,
+ 772723.400000ns, VSS,
+ 772723.500000ns, VDD,
+ 773083.700000ns, VDD,
+ 773083.800000ns, VSS,
+ 773203.800000ns, VSS,
+ 773203.900000ns, VDD,
+ 773684.200000ns, VDD,
+ 773684.300000ns, VSS,
+ 774164.600000ns, VSS,
+ 774164.700000ns, VDD,
+ 777887.700000ns, VDD,
+ 777887.800000ns, VSS,
+ 778248.000000ns, VSS,
+ 778248.100000ns, VDD,
+ 778488.200000ns, VDD,
+ 778488.300000ns, VSS,
+ 779689.200000ns, VSS,
+ 779689.300000ns, VDD,
+ 782571.600000ns, VDD,
+ 782571.700000ns, VSS,
+ 782811.800000ns, VSS,
+ 782811.900000ns, VDD,
+ 783292.200000ns, VDD,
+ 783292.300000ns, VSS,
+ 783892.700000ns, VSS,
+ 783892.800000ns, VDD,
+ 784012.800000ns, VDD,
+ 784012.900000ns, VSS,
+ 786895.200000ns, VSS,
+ 786895.300000ns, VDD,
+ 788696.700000ns, VDD,
+ 788696.800000ns, VSS,
+ 789417.300000ns, VSS,
+ 789417.400000ns, VDD,
+ 790017.800000ns, VDD,
+ 790017.900000ns, VSS,
+ 790378.100000ns, VSS,
+ 790378.200000ns, VDD,
+ 790498.200000ns, VDD,
+ 790498.300000ns, VSS,
+ 790618.300000ns, VSS,
+ 790618.400000ns, VDD,
+ 792059.500000ns, VDD,
+ 792059.600000ns, VSS,
+ 792299.700000ns, VSS,
+ 792299.800000ns, VDD,
+ 792900.200000ns, VDD,
+ 792900.300000ns, VSS,
+ 793500.700000ns, VSS,
+ 793500.800000ns, VDD,
+ 793861.000000ns, VDD,
+ 793861.100000ns, VSS,
+ 794941.900000ns, VSS,
+ 794942.000000ns, VDD,
+ 795062.000000ns, VDD,
+ 795062.100000ns, VSS,
+ 795782.600000ns, VSS,
+ 795782.700000ns, VDD,
+ 796142.900000ns, VDD,
+ 796143.000000ns, VSS,
+ 796863.500000ns, VSS,
+ 796863.600000ns, VDD,
+ 797584.100000ns, VDD,
+ 797584.200000ns, VSS,
+ 798304.700000ns, VSS,
+ 798304.800000ns, VDD,
+ 798905.200000ns, VDD,
+ 798905.300000ns, VSS,
+ 800226.300000ns, VSS,
+ 800226.400000ns, VDD,
+ 800706.700000ns, VDD,
+ 800706.800000ns, VSS,
+ 800826.800000ns, VSS,
+ 800826.900000ns, VDD,
+ 801547.400000ns, VDD,
+ 801547.500000ns, VSS,
+ 801667.500000ns, VSS,
+ 801667.600000ns, VDD,
+ 801787.600000ns, VDD,
+ 801787.700000ns, VSS,
+ 802268.000000ns, VSS,
+ 802268.100000ns, VDD,
+ 802388.100000ns, VDD,
+ 802388.200000ns, VSS,
+ 802988.600000ns, VSS,
+ 802988.700000ns, VDD,
+ 803829.300000ns, VDD,
+ 803829.400000ns, VSS,
+ 804189.600000ns, VSS,
+ 804189.700000ns, VDD,
+ 804309.700000ns, VDD,
+ 804309.800000ns, VSS,
+ 804790.100000ns, VSS,
+ 804790.200000ns, VDD,
+ 805150.400000ns, VDD,
+ 805150.500000ns, VSS,
+ 805270.500000ns, VSS,
+ 805270.600000ns, VDD,
+ 805750.900000ns, VDD,
+ 805751.000000ns, VSS,
+ 806231.300000ns, VSS,
+ 806231.400000ns, VDD,
+ 806711.700000ns, VDD,
+ 806711.800000ns, VSS,
+ 806831.800000ns, VSS,
+ 806831.900000ns, VDD,
+ 807432.300000ns, VDD,
+ 807432.400000ns, VSS,
+ 808393.100000ns, VSS,
+ 808393.200000ns, VDD,
+ 808873.500000ns, VDD,
+ 808873.600000ns, VSS,
+ 809714.200000ns, VSS,
+ 809714.300000ns, VDD,
+ 810915.200000ns, VDD,
+ 810915.300000ns, VSS,
+ 813197.100000ns, VSS,
+ 813197.200000ns, VDD,
+ 814157.900000ns, VDD,
+ 814158.000000ns, VSS,
+ 814758.400000ns, VSS,
+ 814758.500000ns, VDD,
+ 814878.500000ns, VDD,
+ 814878.600000ns, VSS,
+ 815959.400000ns, VSS,
+ 815959.500000ns, VDD,
+ 816079.500000ns, VDD,
+ 816079.600000ns, VSS,
+ 817160.400000ns, VSS,
+ 817160.500000ns, VDD,
+ 817881.000000ns, VDD,
+ 817881.100000ns, VSS,
+ 818721.700000ns, VSS,
+ 818721.800000ns, VDD,
+ 819562.400000ns, VDD,
+ 819562.500000ns, VSS,
+ 820042.800000ns, VSS,
+ 820042.900000ns, VDD,
+ 820523.200000ns, VDD,
+ 820523.300000ns, VSS,
+ 821123.700000ns, VSS,
+ 821123.800000ns, VDD,
+ 821724.200000ns, VDD,
+ 821724.300000ns, VSS,
+ 823165.400000ns, VSS,
+ 823165.500000ns, VDD,
+ 823886.000000ns, VDD,
+ 823886.100000ns, VSS,
+ 824126.200000ns, VSS,
+ 824126.300000ns, VDD,
+ 824486.500000ns, VDD,
+ 824486.600000ns, VSS,
+ 825207.100000ns, VSS,
+ 825207.200000ns, VDD,
+ 825807.600000ns, VDD,
+ 825807.700000ns, VSS,
+ 826528.200000ns, VSS,
+ 826528.300000ns, VDD,
+ 827969.400000ns, VDD,
+ 827969.500000ns, VSS,
+ 829170.400000ns, VSS,
+ 829170.500000ns, VDD,
+ 829770.900000ns, VDD,
+ 829771.000000ns, VSS,
+ 831212.100000ns, VSS,
+ 831212.200000ns, VDD,
+ 831692.500000ns, VDD,
+ 831692.600000ns, VSS,
+ 831812.600000ns, VSS,
+ 831812.700000ns, VDD,
+ 833734.200000ns, VDD,
+ 833734.300000ns, VSS,
+ 834454.800000ns, VSS,
+ 834454.900000ns, VDD,
+ 835775.900000ns, VDD,
+ 835776.000000ns, VSS,
+ 835896.000000ns, VSS,
+ 835896.100000ns, VDD,
+ 838057.800000ns, VDD,
+ 838057.900000ns, VSS,
+ 838298.000000ns, VSS,
+ 838298.100000ns, VDD,
+ 838538.200000ns, VDD,
+ 838538.300000ns, VSS,
+ 838658.300000ns, VSS,
+ 838658.400000ns, VDD,
+ 838778.400000ns, VDD,
+ 838778.500000ns, VSS,
+ 839499.000000ns, VSS,
+ 839499.100000ns, VDD,
+ 839739.200000ns, VDD,
+ 839739.300000ns, VSS,
+ 840459.800000ns, VSS,
+ 840459.900000ns, VDD,
+ 840820.100000ns, VDD,
+ 840820.200000ns, VSS,
+ 841540.700000ns, VSS,
+ 841540.800000ns, VDD,
+ 841780.900000ns, VDD,
+ 841781.000000ns, VSS,
+ 842861.800000ns, VSS,
+ 842861.900000ns, VDD,
+ 843462.300000ns, VDD,
+ 843462.400000ns, VSS,
+ 844182.900000ns, VSS,
+ 844183.000000ns, VDD,
+ 844543.200000ns, VDD,
+ 844543.300000ns, VSS,
+ 844663.300000ns, VSS,
+ 844663.400000ns, VDD,
+ 844903.500000ns, VDD,
+ 844903.600000ns, VSS,
+ 845023.600000ns, VSS,
+ 845023.700000ns, VDD,
+ 846825.100000ns, VDD,
+ 846825.200000ns, VSS,
+ 846945.200000ns, VSS,
+ 846945.300000ns, VDD,
+ 847185.400000ns, VDD,
+ 847185.500000ns, VSS,
+ 847305.500000ns, VSS,
+ 847305.600000ns, VDD,
+ 848146.200000ns, VDD,
+ 848146.300000ns, VSS,
+ 848626.600000ns, VSS,
+ 848626.700000ns, VDD,
+ 849587.400000ns, VDD,
+ 849587.500000ns, VSS,
+ 849827.600000ns, VSS,
+ 849827.700000ns, VDD,
+ 850187.900000ns, VDD,
+ 850188.000000ns, VSS,
+ 852229.600000ns, VSS,
+ 852229.700000ns, VDD,
+ 853550.700000ns, VDD,
+ 853550.800000ns, VSS,
+ 853911.000000ns, VSS,
+ 853911.100000ns, VDD,
+ 854991.900000ns, VDD,
+ 854992.000000ns, VSS,
+ 855952.700000ns, VSS,
+ 855952.800000ns, VDD,
+ 857153.700000ns, VDD,
+ 857153.800000ns, VSS,
+ 859195.400000ns, VSS,
+ 859195.500000ns, VDD,
+ 859675.800000ns, VDD,
+ 859675.900000ns, VSS,
+ 861237.100000ns, VSS,
+ 861237.200000ns, VDD,
+ 861357.200000ns, VDD,
+ 861357.300000ns, VSS,
+ 861957.700000ns, VSS,
+ 861957.800000ns, VDD,
+ 863759.200000ns, VDD,
+ 863759.300000ns, VSS,
+ 864239.600000ns, VSS,
+ 864239.700000ns, VDD,
+ 864960.200000ns, VDD,
+ 864960.300000ns, VSS,
+ 865200.400000ns, VSS,
+ 865200.500000ns, VDD,
+ 865440.600000ns, VDD,
+ 865440.700000ns, VSS,
+ 865560.700000ns, VSS,
+ 865560.800000ns, VDD,
+ 866881.800000ns, VDD,
+ 866881.900000ns, VSS,
+ 867362.200000ns, VSS,
+ 867362.300000ns, VDD,
+ 867602.400000ns, VDD,
+ 867602.500000ns, VSS,
+ 868563.200000ns, VSS,
+ 868563.300000ns, VDD,
+ 869764.200000ns, VDD,
+ 869764.300000ns, VSS,
+ 870965.200000ns, VSS,
+ 870965.300000ns, VDD,
+ 872046.100000ns, VDD,
+ 872046.200000ns, VSS,
+ 872286.300000ns, VSS,
+ 872286.400000ns, VDD,
+ 872406.400000ns, VDD,
+ 872406.500000ns, VSS,
+ 872526.500000ns, VSS,
+ 872526.600000ns, VDD,
+ 872886.800000ns, VDD,
+ 872886.900000ns, VSS,
+ 873487.300000ns, VSS,
+ 873487.400000ns, VDD,
+ 874688.300000ns, VDD,
+ 874688.400000ns, VSS,
+ 875408.900000ns, VSS,
+ 875409.000000ns, VDD,
+ 875529.000000ns, VDD,
+ 875529.100000ns, VSS,
+ 876249.600000ns, VSS,
+ 876249.700000ns, VDD,
+ 877090.300000ns, VDD,
+ 877090.400000ns, VSS,
+ 879132.000000ns, VSS,
+ 879132.100000ns, VDD,
+ 880693.300000ns, VDD,
+ 880693.400000ns, VSS,
+ 880933.500000ns, VSS,
+ 880933.600000ns, VDD,
+ 881173.700000ns, VDD,
+ 881173.800000ns, VSS,
+ 881413.900000ns, VSS,
+ 881414.000000ns, VDD,
+ 881534.000000ns, VDD,
+ 881534.100000ns, VSS,
+ 881894.300000ns, VSS,
+ 881894.400000ns, VDD,
+ 882134.500000ns, VDD,
+ 882134.600000ns, VSS,
+ 882735.000000ns, VSS,
+ 882735.100000ns, VDD,
+ 883695.800000ns, VDD,
+ 883695.900000ns, VSS,
+ 884776.700000ns, VSS,
+ 884776.800000ns, VDD,
+ 885257.100000ns, VDD,
+ 885257.200000ns, VSS,
+ 885377.200000ns, VSS,
+ 885377.300000ns, VDD,
+ 885857.600000ns, VDD,
+ 885857.700000ns, VSS,
+ 886578.200000ns, VSS,
+ 886578.300000ns, VDD,
+ 887058.600000ns, VDD,
+ 887058.700000ns, VSS,
+ 887418.900000ns, VSS,
+ 887419.000000ns, VDD,
+ 887539.000000ns, VDD,
+ 887539.100000ns, VSS,
+ 888139.500000ns, VSS,
+ 888139.600000ns, VDD,
+ 888259.600000ns, VDD,
+ 888259.700000ns, VSS,
+ 889580.700000ns, VSS,
+ 889580.800000ns, VDD,
+ 889941.000000ns, VDD,
+ 889941.100000ns, VSS,
+ 890061.100000ns, VSS,
+ 890061.200000ns, VDD,
+ 890661.600000ns, VDD,
+ 890661.700000ns, VSS,
+ 891382.200000ns, VSS,
+ 891382.300000ns, VDD,
+ 892343.000000ns, VDD,
+ 892343.100000ns, VSS,
+ 892823.400000ns, VSS,
+ 892823.500000ns, VDD,
+ 894985.200000ns, VDD,
+ 894985.300000ns, VSS,
+ 896066.100000ns, VSS,
+ 896066.200000ns, VDD,
+ 897867.600000ns, VDD,
+ 897867.700000ns, VSS,
+ 898468.100000ns, VSS,
+ 898468.200000ns, VDD,
+ 898948.500000ns, VDD,
+ 898948.600000ns, VSS,
+ 903031.900000ns, VSS,
+ 903032.000000ns, VDD,
+ 903512.300000ns, VDD,
+ 903512.400000ns, VSS,
+ 904593.200000ns, VSS,
+ 904593.300000ns, VDD,
+ 905794.200000ns, VDD,
+ 905794.300000ns, VSS,
+ 906274.600000ns, VSS,
+ 906274.700000ns, VDD,
+ 906394.700000ns, VDD,
+ 906394.800000ns, VSS,
+ 906755.000000ns, VSS,
+ 906755.100000ns, VDD,
+ 907475.600000ns, VDD,
+ 907475.700000ns, VSS,
+ 907595.700000ns, VSS,
+ 907595.800000ns, VDD,
+ 908796.700000ns, VDD,
+ 908796.800000ns, VSS,
+ 909757.500000ns, VSS,
+ 909757.600000ns, VDD,
+ 910237.900000ns, VDD,
+ 910238.000000ns, VSS,
+ 910718.300000ns, VSS,
+ 910718.400000ns, VDD,
+ 911679.100000ns, VDD,
+ 911679.200000ns, VSS,
+ 912159.500000ns, VSS,
+ 912159.600000ns, VDD,
+ 912279.600000ns, VDD,
+ 912279.700000ns, VSS,
+ 912399.700000ns, VSS,
+ 912399.800000ns, VDD,
+ 912639.900000ns, VDD,
+ 912640.000000ns, VSS,
+ 912880.100000ns, VSS,
+ 912880.200000ns, VDD,
+ 914321.300000ns, VDD,
+ 914321.400000ns, VSS,
+ 914561.500000ns, VSS,
+ 914561.600000ns, VDD,
+ 915162.000000ns, VDD,
+ 915162.100000ns, VSS,
+ 916122.800000ns, VSS,
+ 916122.900000ns, VDD,
+ 917443.900000ns, VDD,
+ 917444.000000ns, VSS,
+ 918164.500000ns, VSS,
+ 918164.600000ns, VDD,
+ 919605.700000ns, VDD,
+ 919605.800000ns, VSS,
+ 919966.000000ns, VSS,
+ 919966.100000ns, VDD,
+ 920326.300000ns, VDD,
+ 920326.400000ns, VSS,
+ 920446.400000ns, VSS,
+ 920446.500000ns, VDD,
+ 920806.700000ns, VDD,
+ 920806.800000ns, VSS,
+ 921287.100000ns, VSS,
+ 921287.200000ns, VDD,
+ 921887.600000ns, VDD,
+ 921887.700000ns, VSS,
+ 922007.700000ns, VSS,
+ 922007.800000ns, VDD,
+ 923208.700000ns, VDD,
+ 923208.800000ns, VSS,
+ 923328.800000ns, VSS,
+ 923328.900000ns, VDD,
+ 923448.900000ns, VDD,
+ 923449.000000ns, VSS,
+ 923809.200000ns, VSS,
+ 923809.300000ns, VDD,
+ 924049.400000ns, VDD,
+ 924049.500000ns, VSS,
+ 924169.500000ns, VSS,
+ 924169.600000ns, VDD,
+ 925010.200000ns, VDD,
+ 925010.300000ns, VSS,
+ 925370.500000ns, VSS,
+ 925370.600000ns, VDD,
+ 925971.000000ns, VDD,
+ 925971.100000ns, VSS,
+ 926451.400000ns, VSS,
+ 926451.500000ns, VDD,
+ 926571.500000ns, VDD,
+ 926571.600000ns, VSS,
+ 927412.200000ns, VSS,
+ 927412.300000ns, VDD,
+ 928132.800000ns, VDD,
+ 928132.900000ns, VSS,
+ 929093.600000ns, VSS,
+ 929093.700000ns, VDD,
+ 929694.100000ns, VDD,
+ 929694.200000ns, VSS,
+ 929814.200000ns, VSS,
+ 929814.300000ns, VDD,
+ 929934.300000ns, VDD,
+ 929934.400000ns, VSS,
+ 930054.400000ns, VSS,
+ 930054.500000ns, VDD,
+ 930174.500000ns, VDD,
+ 930174.600000ns, VSS,
+ 930775.000000ns, VSS,
+ 930775.100000ns, VDD,
+ 931495.600000ns, VDD,
+ 931495.700000ns, VSS,
+ 931976.000000ns, VSS,
+ 931976.100000ns, VDD,
+ 932336.300000ns, VDD,
+ 932336.400000ns, VSS,
+ 933297.100000ns, VSS,
+ 933297.200000ns, VDD,
+ 933537.300000ns, VDD,
+ 933537.400000ns, VSS,
+ 935338.800000ns, VSS,
+ 935338.900000ns, VDD,
+ 935819.200000ns, VDD,
+ 935819.300000ns, VSS,
+ 937020.200000ns, VSS,
+ 937020.300000ns, VDD,
+ 937260.400000ns, VDD,
+ 937260.500000ns, VSS,
+ 937380.500000ns, VSS,
+ 937380.600000ns, VDD,
+ 937860.900000ns, VDD,
+ 937861.000000ns, VSS,
+ 939422.200000ns, VSS,
+ 939422.300000ns, VDD,
+ 940022.700000ns, VDD,
+ 940022.800000ns, VSS,
+ 940863.400000ns, VSS,
+ 940863.500000ns, VDD,
+ 940983.500000ns, VDD,
+ 940983.600000ns, VSS,
+ 941704.100000ns, VSS,
+ 941704.200000ns, VDD,
+ 942664.900000ns, VDD,
+ 942665.000000ns, VSS,
+ 942905.100000ns, VSS,
+ 942905.200000ns, VDD,
+ 943745.800000ns, VDD,
+ 943745.900000ns, VSS,
+ 944586.500000ns, VSS,
+ 944586.600000ns, VDD,
+ 945187.000000ns, VDD,
+ 945187.100000ns, VSS,
+ 945427.200000ns, VSS,
+ 945427.300000ns, VDD,
+ 945547.300000ns, VDD,
+ 945547.400000ns, VSS,
+ 946388.000000ns, VSS,
+ 946388.100000ns, VDD,
+ 947108.600000ns, VDD,
+ 947108.700000ns, VSS,
+ 947468.900000ns, VSS,
+ 947469.000000ns, VDD,
+ 948309.600000ns, VDD,
+ 948309.700000ns, VSS,
+ 948669.900000ns, VSS,
+ 948670.000000ns, VDD,
+ 949390.500000ns, VDD,
+ 949390.600000ns, VSS,
+ 949870.900000ns, VSS,
+ 949871.000000ns, VDD,
+ 950231.200000ns, VDD,
+ 950231.300000ns, VSS,
+ 950471.400000ns, VSS,
+ 950471.500000ns, VDD,
+ 950951.800000ns, VDD,
+ 950951.900000ns, VSS,
+ 952993.500000ns, VSS,
+ 952993.600000ns, VDD,
+ 953113.600000ns, VDD,
+ 953113.700000ns, VSS,
+ 953954.300000ns, VSS,
+ 953954.400000ns, VDD,
+ 954314.600000ns, VDD,
+ 954314.700000ns, VSS,
+ 957917.600000ns, VSS,
+ 957917.700000ns, VDD,
+ 958398.000000ns, VDD,
+ 958398.100000ns, VSS,
+ 958878.400000ns, VSS,
+ 958878.500000ns, VDD,
+ 958998.500000ns, VDD,
+ 958998.600000ns, VSS,
+ 959599.000000ns, VSS,
+ 959599.100000ns, VDD,
+ 960439.700000ns, VDD,
+ 960439.800000ns, VSS,
+ 960920.100000ns, VSS,
+ 960920.200000ns, VDD,
+ 961520.600000ns, VDD,
+ 961520.700000ns, VSS,
+ 961640.700000ns, VSS,
+ 961640.800000ns, VDD,
+ 962721.600000ns, VDD,
+ 962721.700000ns, VSS,
+ 963802.500000ns, VSS,
+ 963802.600000ns, VDD,
+ 966684.900000ns, VDD,
+ 966685.000000ns, VSS,
+ 967045.200000ns, VSS,
+ 967045.300000ns, VDD,
+ 967525.600000ns, VDD,
+ 967525.700000ns, VSS,
+ 968126.100000ns, VSS,
+ 968126.200000ns, VDD,
+ 968246.200000ns, VDD,
+ 968246.300000ns, VSS,
+ 969086.900000ns, VSS,
+ 969087.000000ns, VDD,
+ 969207.000000ns, VDD,
+ 969207.100000ns, VSS,
+ 969927.600000ns, VSS,
+ 969927.700000ns, VDD,
+ 970287.900000ns, VDD,
+ 970288.000000ns, VSS,
+ 970648.200000ns, VSS,
+ 970648.300000ns, VDD,
+ 970888.400000ns, VDD,
+ 970888.500000ns, VSS,
+ 971008.500000ns, VSS,
+ 971008.600000ns, VDD,
+ 971488.900000ns, VDD,
+ 971489.000000ns, VSS,
+ 971729.100000ns, VSS,
+ 971729.200000ns, VDD,
+ 972329.600000ns, VDD,
+ 972329.700000ns, VSS,
+ 973170.300000ns, VSS,
+ 973170.400000ns, VDD,
+ 973650.700000ns, VDD,
+ 973650.800000ns, VSS,
+ 974131.100000ns, VSS,
+ 974131.200000ns, VDD,
+ 976773.300000ns, VDD,
+ 976773.400000ns, VSS,
+ 978214.500000ns, VSS,
+ 978214.600000ns, VDD,
+ 978574.800000ns, VDD,
+ 978574.900000ns, VSS,
+ 980736.600000ns, VSS,
+ 980736.700000ns, VDD,
+ 981096.900000ns, VDD,
+ 981097.000000ns, VSS,
+ 981337.100000ns, VSS,
+ 981337.200000ns, VDD,
+ 981457.200000ns, VDD,
+ 981457.300000ns, VSS,
+ 982297.900000ns, VSS,
+ 982298.000000ns, VDD,
+ 983258.700000ns, VDD,
+ 983258.800000ns, VSS,
+ 984219.500000ns, VSS,
+ 984219.600000ns, VDD,
+ 985780.800000ns, VDD,
+ 985780.900000ns, VSS,
+ 986381.300000ns, VSS,
+ 986381.400000ns, VDD,
+ 987462.200000ns, VDD,
+ 987462.300000ns, VSS,
+ 987702.400000ns, VSS,
+ 987702.500000ns, VDD,
+ 988423.000000ns, VDD,
+ 988423.100000ns, VSS,
+ 988543.100000ns, VSS,
+ 988543.200000ns, VDD,
+ 988903.400000ns, VDD,
+ 988903.500000ns, VSS,
+ 989023.500000ns, VSS,
+ 989023.600000ns, VDD,
+ 989143.600000ns, VDD,
+ 989143.700000ns, VSS,
+ 989984.300000ns, VSS,
+ 989984.400000ns, VDD,
+ 990704.900000ns, VDD,
+ 990705.000000ns, VSS,
+ 991425.500000ns, VSS,
+ 991425.600000ns, VDD,
+ 991545.600000ns, VDD,
+ 991545.700000ns, VSS,
+ 991665.700000ns, VSS,
+ 991665.800000ns, VDD,
+ 992146.100000ns, VDD,
+ 992146.200000ns, VSS,
+ 992746.600000ns, VSS,
+ 992746.700000ns, VDD,
+ 993467.200000ns, VDD,
+ 993467.300000ns, VSS,
+ 993587.300000ns, VSS,
+ 993587.400000ns, VDD,
+ 995148.600000ns, VDD,
+ 995148.700000ns, VSS,
+ 995629.000000ns, VSS,
+ 995629.100000ns, VDD,
+ 996109.400000ns, VDD,
+ 996109.500000ns, VSS,
+ 996229.500000ns, VSS,
+ 996229.600000ns, VDD,
+ 996349.600000ns, VDD,
+ 996349.700000ns, VSS,
+ 996589.800000ns, VSS,
+ 996589.900000ns, VDD,
+ 996830.000000ns, VDD,
+ 996830.100000ns, VSS,
+ 996950.100000ns, VSS,
+ 996950.200000ns, VDD,
+ 997910.900000ns, VDD,
+ 997911.000000ns, VSS,
+ 998751.600000ns, VSS,
+ 998751.700000ns, VDD,
+ 999232.000000ns, VDD,
+ 999232.100000ns, VSS,
+ 999472.200000ns, VSS,
+ 999472.300000ns, VDD,
+ 999712.400000ns, VDD,
+ 999712.500000ns, VSS,
+ 999832.500000ns, VSS,
+ 999832.600000ns, VDD,
+ 1000433.000000ns, VDD,
+ 1000433.100000ns, VSS,
+ 1001273.700000ns, VSS,
+ 1001273.800000ns, VDD,
+ 1001754.100000ns, VDD,
+ 1001754.200000ns, VSS,
+ 1002955.100000ns, VSS,
+ 1002955.200000ns, VDD,
+ 1003195.300000ns, VDD,
+ 1003195.400000ns, VSS,
+ 1003915.900000ns, VSS,
+ 1003916.000000ns, VDD,
+ 1004396.300000ns, VDD,
+ 1004396.400000ns, VSS,
+ 1004516.400000ns, VSS,
+ 1004516.500000ns, VDD,
+ 1004636.500000ns, VDD,
+ 1004636.600000ns, VSS,
+ 1005116.900000ns, VSS,
+ 1005117.000000ns, VDD,
+ 1005237.000000ns, VDD,
+ 1005237.100000ns, VSS,
+ 1006678.200000ns, VSS,
+ 1006678.300000ns, VDD,
+ 1007398.800000ns, VDD,
+ 1007398.900000ns, VSS,
+ 1008359.600000ns, VSS,
+ 1008359.700000ns, VDD,
+ 1008840.000000ns, VDD,
+ 1008840.100000ns, VSS,
+ 1008960.100000ns, VSS,
+ 1008960.200000ns, VDD,
+ 1009320.400000ns, VDD,
+ 1009320.500000ns, VSS,
+ 1009440.500000ns, VSS,
+ 1009440.600000ns, VDD,
+ 1010281.200000ns, VDD,
+ 1010281.300000ns, VSS,
+ 1010881.700000ns, VSS,
+ 1010881.800000ns, VDD,
+ 1011121.900000ns, VDD,
+ 1011122.000000ns, VSS,
+ 1011602.300000ns, VSS,
+ 1011602.400000ns, VDD,
+ 1013283.700000ns, VDD,
+ 1013283.800000ns, VSS,
+ 1014604.800000ns, VSS,
+ 1014604.900000ns, VDD,
+ 1014724.900000ns, VDD,
+ 1014725.000000ns, VSS,
+ 1016766.600000ns, VSS,
+ 1016766.700000ns, VDD,
+ 1018087.700000ns, VDD,
+ 1018087.800000ns, VSS,
+ 1018327.900000ns, VSS,
+ 1018328.000000ns, VDD,
+ 1018808.300000ns, VDD,
+ 1018808.400000ns, VSS,
+ 1020249.500000ns, VSS,
+ 1020249.600000ns, VDD,
+ 1020970.100000ns, VDD,
+ 1020970.200000ns, VSS,
+ 1021090.200000ns, VSS,
+ 1021090.300000ns, VDD,
+ 1021210.300000ns, VDD,
+ 1021210.400000ns, VSS,
+ 1021690.700000ns, VSS,
+ 1021690.800000ns, VDD,
+ 1023011.800000ns, VDD,
+ 1023011.900000ns, VSS,
+ 1023732.400000ns, VSS,
+ 1023732.500000ns, VDD,
+ 1024453.000000ns, VDD,
+ 1024453.100000ns, VSS,
+ 1027095.200000ns, VSS,
+ 1027095.300000ns, VDD,
+ 1027335.400000ns, VDD,
+ 1027335.500000ns, VSS,
+ 1027935.900000ns, VSS,
+ 1027936.000000ns, VDD,
+ 1029016.800000ns, VDD,
+ 1029016.900000ns, VSS,
+ 1029497.200000ns, VSS,
+ 1029497.300000ns, VDD,
+ 1029857.500000ns, VDD,
+ 1029857.600000ns, VSS,
+ 1030458.000000ns, VSS,
+ 1030458.100000ns, VDD,
+ 1031058.500000ns, VDD,
+ 1031058.600000ns, VSS,
+ 1032379.600000ns, VSS,
+ 1032379.700000ns, VDD,
+ 1032860.000000ns, VDD,
+ 1032860.100000ns, VSS,
+ 1033340.400000ns, VSS,
+ 1033340.500000ns, VDD,
+ 1033460.500000ns, VDD,
+ 1033460.600000ns, VSS,
+ 1033580.600000ns, VSS,
+ 1033580.700000ns, VDD,
+ 1035141.900000ns, VDD,
+ 1035142.000000ns, VSS,
+ 1035622.300000ns, VSS,
+ 1035622.400000ns, VDD,
+ 1035742.400000ns, VDD,
+ 1035742.500000ns, VSS,
+ 1035982.600000ns, VSS,
+ 1035982.700000ns, VDD,
+ 1036102.700000ns, VDD,
+ 1036102.800000ns, VSS,
+ 1036463.000000ns, VSS,
+ 1036463.100000ns, VDD,
+ 1037423.800000ns, VDD,
+ 1037423.900000ns, VSS,
+ 1037664.000000ns, VSS,
+ 1037664.100000ns, VDD,
+ 1038865.000000ns, VDD,
+ 1038865.100000ns, VSS,
+ 1039105.200000ns, VSS,
+ 1039105.300000ns, VDD,
+ 1039225.300000ns, VDD,
+ 1039225.400000ns, VSS,
+ 1039705.700000ns, VSS,
+ 1039705.800000ns, VDD,
+ 1039825.800000ns, VDD,
+ 1039825.900000ns, VSS,
+ 1041867.500000ns, VSS,
+ 1041867.600000ns, VDD,
+ 1042107.700000ns, VDD,
+ 1042107.800000ns, VSS,
+ 1042588.100000ns, VSS,
+ 1042588.200000ns, VDD,
+ 1042708.200000ns, VDD,
+ 1042708.300000ns, VSS,
+ 1042828.300000ns, VSS,
+ 1042828.400000ns, VDD,
+ 1042948.400000ns, VDD,
+ 1042948.500000ns, VSS,
+ 1044389.600000ns, VSS,
+ 1044389.700000ns, VDD,
+ 1044990.100000ns, VDD,
+ 1044990.200000ns, VSS,
+ 1045350.400000ns, VSS,
+ 1045350.500000ns, VDD,
+ 1046191.100000ns, VDD,
+ 1046191.200000ns, VSS,
+ 1047031.800000ns, VSS,
+ 1047031.900000ns, VDD,
+ 1047872.500000ns, VDD,
+ 1047872.600000ns, VSS,
+ 1048112.700000ns, VSS,
+ 1048112.800000ns, VDD,
+ 1048352.900000ns, VDD,
+ 1048353.000000ns, VSS,
+ 1049193.600000ns, VSS,
+ 1049193.700000ns, VDD,
+ 1051115.200000ns, VDD,
+ 1051115.300000ns, VSS,
+ 1053277.000000ns, VSS,
+ 1053277.100000ns, VDD,
+ 1054478.000000ns, VDD,
+ 1054478.100000ns, VSS,
+ 1055318.700000ns, VSS,
+ 1055318.800000ns, VDD,
+ 1055679.000000ns, VDD,
+ 1055679.100000ns, VSS,
+ 1056399.600000ns, VSS,
+ 1056399.700000ns, VDD,
+ 1056639.800000ns, VDD,
+ 1056639.900000ns, VSS,
+ 1056759.900000ns, VSS,
+ 1056760.000000ns, VDD,
+ 1058681.500000ns, VDD,
+ 1058681.600000ns, VSS,
+ 1059762.400000ns, VSS,
+ 1059762.500000ns, VDD,
+ 1060242.800000ns, VDD,
+ 1060242.900000ns, VSS,
+ 1060963.400000ns, VSS,
+ 1060963.500000ns, VDD,
+ 1061323.700000ns, VDD,
+ 1061323.800000ns, VSS,
+ 1062644.800000ns, VSS,
+ 1062644.900000ns, VDD,
+ 1063965.900000ns, VDD,
+ 1063966.000000ns, VSS,
+ 1064086.000000ns, VSS,
+ 1064086.100000ns, VDD,
+ 1064686.500000ns, VDD,
+ 1064686.600000ns, VSS,
+ 1065887.500000ns, VSS,
+ 1065887.600000ns, VDD,
+ 1066488.000000ns, VDD,
+ 1066488.100000ns, VSS,
+ 1067088.500000ns, VSS,
+ 1067088.600000ns, VDD,
+ 1067809.100000ns, VDD,
+ 1067809.200000ns, VSS,
+ 1067929.200000ns, VSS,
+ 1067929.300000ns, VDD,
+ 1068049.300000ns, VDD,
+ 1068049.400000ns, VSS,
+ 1068529.700000ns, VSS,
+ 1068529.800000ns, VDD,
+ 1069490.500000ns, VDD,
+ 1069490.600000ns, VSS,
+ 1069610.600000ns, VSS,
+ 1069610.700000ns, VDD,
+ 1069730.700000ns, VDD,
+ 1069730.800000ns, VSS,
+ 1071171.900000ns, VSS,
+ 1071172.000000ns, VDD,
+ 1071412.100000ns, VDD,
+ 1071412.200000ns, VSS,
+ 1071532.200000ns, VSS,
+ 1071532.300000ns, VDD,
+ 1071652.300000ns, VDD,
+ 1071652.400000ns, VSS,
+ 1073333.700000ns, VSS,
+ 1073333.800000ns, VDD,
+ 1074054.300000ns, VDD,
+ 1074054.400000ns, VSS,
+ 1074294.500000ns, VSS,
+ 1074294.600000ns, VDD,
+ 1075015.100000ns, VDD,
+ 1075015.200000ns, VSS,
+ 1075135.200000ns, VSS,
+ 1075135.300000ns, VDD,
+ 1075615.600000ns, VDD,
+ 1075615.700000ns, VSS,
+ 1076336.200000ns, VSS,
+ 1076336.300000ns, VDD,
+ 1077537.200000ns, VDD,
+ 1077537.300000ns, VSS,
+ 1078377.900000ns, VSS,
+ 1078378.000000ns, VDD,
+ 1079338.700000ns, VDD,
+ 1079338.800000ns, VSS,
+ 1080419.600000ns, VSS,
+ 1080419.700000ns, VDD,
+ 1080659.800000ns, VDD,
+ 1080659.900000ns, VSS,
+ 1081620.600000ns, VSS,
+ 1081620.700000ns, VDD,
+ 1081980.900000ns, VDD,
+ 1081981.000000ns, VSS,
+ 1082341.200000ns, VSS,
+ 1082341.300000ns, VDD,
+ 1082581.400000ns, VDD,
+ 1082581.500000ns, VSS,
+ 1083302.000000ns, VSS,
+ 1083302.100000ns, VDD,
+ 1083662.300000ns, VDD,
+ 1083662.400000ns, VSS,
+ 1084262.800000ns, VSS,
+ 1084262.900000ns, VDD,
+ 1085463.800000ns, VDD,
+ 1085463.900000ns, VSS,
+ 1085583.900000ns, VSS,
+ 1085584.000000ns, VDD,
+ 1086905.000000ns, VDD,
+ 1086905.100000ns, VSS,
+ 1087025.100000ns, VSS,
+ 1087025.200000ns, VDD,
+ 1087865.800000ns, VDD,
+ 1087865.900000ns, VSS,
+ 1089307.000000ns, VSS,
+ 1089307.100000ns, VDD,
+ 1090027.600000ns, VDD,
+ 1090027.700000ns, VSS,
+ 1090988.400000ns, VSS,
+ 1090988.500000ns, VDD,
+ 1091228.600000ns, VDD,
+ 1091228.700000ns, VSS,
+ 1091468.800000ns, VSS,
+ 1091468.900000ns, VDD,
+ 1092429.600000ns, VDD,
+ 1092429.700000ns, VSS,
+ 1093150.200000ns, VSS,
+ 1093150.300000ns, VDD,
+ 1093630.600000ns, VDD,
+ 1093630.700000ns, VSS,
+ 1093990.900000ns, VSS,
+ 1093991.000000ns, VDD,
+ 1094231.100000ns, VDD,
+ 1094231.200000ns, VSS,
+ 1094351.200000ns, VSS,
+ 1094351.300000ns, VDD,
+ 1095552.200000ns, VDD,
+ 1095552.300000ns, VSS,
+ 1095912.500000ns, VSS,
+ 1095912.600000ns, VDD,
+ 1096032.600000ns, VDD,
+ 1096032.700000ns, VSS,
+ 1096392.900000ns, VSS,
+ 1096393.000000ns, VDD,
+ 1097473.800000ns, VDD,
+ 1097473.900000ns, VSS,
+ 1098434.600000ns, VSS,
+ 1098434.700000ns, VDD,
+ 1098674.800000ns, VDD,
+ 1098674.900000ns, VSS,
+ 1099155.200000ns, VSS,
+ 1099155.300000ns, VDD,
+ 1099635.600000ns, VDD,
+ 1099635.700000ns, VSS,
+ 1099995.900000ns, VSS,
+ 1099996.000000ns, VDD,
+ 1100476.300000ns, VDD,
+ 1100476.400000ns, VSS,
+ 1100836.600000ns, VSS,
+ 1100836.700000ns, VDD,
+ 1101196.900000ns, VDD,
+ 1101197.000000ns, VSS,
+ 1103118.500000ns, VSS,
+ 1103118.600000ns, VDD,
+ 1103598.900000ns, VDD,
+ 1103599.000000ns, VSS,
+ 1104079.300000ns, VSS,
+ 1104079.400000ns, VDD,
+ 1104799.900000ns, VDD,
+ 1104800.000000ns, VSS,
+ 1106241.100000ns, VSS,
+ 1106241.200000ns, VDD,
+ 1106961.700000ns, VDD,
+ 1106961.800000ns, VSS,
+ 1107322.000000ns, VSS,
+ 1107322.100000ns, VDD,
+ 1108282.800000ns, VDD,
+ 1108282.900000ns, VSS,
+ 1109123.500000ns, VSS,
+ 1109123.600000ns, VDD,
+ 1109603.900000ns, VDD,
+ 1109604.000000ns, VSS,
+ 1110925.000000ns, VSS,
+ 1110925.100000ns, VDD,
+ 1111645.600000ns, VDD,
+ 1111645.700000ns, VSS,
+ 1113086.800000ns, VSS,
+ 1113086.900000ns, VDD,
+ 1114648.100000ns, VDD,
+ 1114648.200000ns, VSS,
+ 1115128.500000ns, VSS,
+ 1115128.600000ns, VDD,
+ 1115608.900000ns, VDD,
+ 1115609.000000ns, VSS,
+ 1115729.000000ns, VSS,
+ 1115729.100000ns, VDD,
+ 1116689.800000ns, VDD,
+ 1116689.900000ns, VSS,
+ 1116930.000000ns, VSS,
+ 1116930.100000ns, VDD,
+ 1117170.200000ns, VDD,
+ 1117170.300000ns, VSS,
+ 1118010.900000ns, VSS,
+ 1118011.000000ns, VDD,
+ 1118851.600000ns, VDD,
+ 1118851.700000ns, VSS,
+ 1119211.900000ns, VSS,
+ 1119212.000000ns, VDD,
+ 1120052.600000ns, VDD,
+ 1120052.700000ns, VSS,
+ 1120653.100000ns, VSS,
+ 1120653.200000ns, VDD,
+ 1121373.700000ns, VDD,
+ 1121373.800000ns, VSS,
+ 1121613.900000ns, VSS,
+ 1121614.000000ns, VDD,
+ 1121734.000000ns, VDD,
+ 1121734.100000ns, VSS,
+ 1122574.700000ns, VSS,
+ 1122574.800000ns, VDD,
+ 1123415.400000ns, VDD,
+ 1123415.500000ns, VSS,
+ 1123535.500000ns, VSS,
+ 1123535.600000ns, VDD,
+ 1123655.600000ns, VDD,
+ 1123655.700000ns, VSS,
+ 1125337.000000ns, VSS,
+ 1125337.100000ns, VDD,
+ 1126658.100000ns, VDD,
+ 1126658.200000ns, VSS,
+ 1127258.600000ns, VSS,
+ 1127258.700000ns, VDD,
+ 1127618.900000ns, VDD,
+ 1127619.000000ns, VSS,
+ 1127739.000000ns, VSS,
+ 1127739.100000ns, VDD,
+ 1127859.100000ns, VDD,
+ 1127859.200000ns, VSS,
+ 1128219.400000ns, VSS,
+ 1128219.500000ns, VDD,
+ 1128819.900000ns, VDD,
+ 1128820.000000ns, VSS,
+ 1130020.900000ns, VSS,
+ 1130021.000000ns, VDD,
+ 1130621.400000ns, VDD,
+ 1130621.500000ns, VSS,
+ 1131221.900000ns, VSS,
+ 1131222.000000ns, VDD,
+ 1131702.300000ns, VDD,
+ 1131702.400000ns, VSS,
+ 1131822.400000ns, VSS,
+ 1131822.500000ns, VDD,
+ 1133503.800000ns, VDD,
+ 1133503.900000ns, VSS,
+ 1134464.600000ns, VSS,
+ 1134464.700000ns, VDD,
+ 1134584.700000ns, VDD,
+ 1134584.800000ns, VSS,
+ 1135305.300000ns, VSS,
+ 1135305.400000ns, VDD,
+ 1136866.600000ns, VDD,
+ 1136866.700000ns, VSS,
+ 1137347.000000ns, VSS,
+ 1137347.100000ns, VDD,
+ 1137827.400000ns, VDD,
+ 1137827.500000ns, VSS,
+ 1138788.200000ns, VSS,
+ 1138788.300000ns, VDD,
+ 1138908.300000ns, VDD,
+ 1138908.400000ns, VSS,
+ 1141310.300000ns, VSS,
+ 1141310.400000ns, VDD,
+ 1142751.500000ns, VDD,
+ 1142751.600000ns, VSS,
+ 1142991.700000ns, VSS,
+ 1142991.800000ns, VDD,
+ 1143231.900000ns, VDD,
+ 1143232.000000ns, VSS,
+ 1143352.000000ns, VSS,
+ 1143352.100000ns, VDD,
+ 1144192.700000ns, VDD,
+ 1144192.800000ns, VSS,
+ 1144432.900000ns, VSS,
+ 1144433.000000ns, VDD,
+ 1145994.200000ns, VDD,
+ 1145994.300000ns, VSS,
+ 1147555.500000ns, VSS,
+ 1147555.600000ns, VDD,
+ 1148156.000000ns, VDD,
+ 1148156.100000ns, VSS,
+ 1148636.400000ns, VSS,
+ 1148636.500000ns, VDD,
+ 1149357.000000ns, VDD,
+ 1149357.100000ns, VSS,
+ 1149717.300000ns, VSS,
+ 1149717.400000ns, VDD,
+ 1149837.400000ns, VDD,
+ 1149837.500000ns, VSS,
+ 1150317.800000ns, VSS,
+ 1150317.900000ns, VDD,
+ 1150798.200000ns, VDD,
+ 1150798.300000ns, VSS,
+ 1151158.500000ns, VSS,
+ 1151158.600000ns, VDD,
+ 1151759.000000ns, VDD,
+ 1151759.100000ns, VSS,
+ 1152960.000000ns, VSS,
+ 1152960.100000ns, VDD,
+ 1153320.300000ns, VDD,
+ 1153320.400000ns, VSS,
+ 1153440.400000ns, VSS,
+ 1153440.500000ns, VDD,
+ 1154521.300000ns, VDD,
+ 1154521.400000ns, VSS,
+ 1154761.500000ns, VSS,
+ 1154761.600000ns, VDD,
+ 1155241.900000ns, VDD,
+ 1155242.000000ns, VSS,
+ 1155602.200000ns, VSS,
+ 1155602.300000ns, VDD,
+ 1157283.600000ns, VDD,
+ 1157283.700000ns, VSS,
+ 1157403.700000ns, VSS,
+ 1157403.800000ns, VDD,
+ 1157643.900000ns, VDD,
+ 1157644.000000ns, VSS,
+ 1158124.300000ns, VSS,
+ 1158124.400000ns, VDD,
+ 1159085.100000ns, VDD,
+ 1159085.200000ns, VSS,
+ 1159445.400000ns, VSS,
+ 1159445.500000ns, VDD,
+ 1159685.600000ns, VDD,
+ 1159685.700000ns, VSS,
+ 1161847.400000ns, VSS,
+ 1161847.500000ns, VDD,
+ 1162808.200000ns, VDD,
+ 1162808.300000ns, VSS,
+ 1163288.600000ns, VSS,
+ 1163288.700000ns, VDD,
+ 1164369.500000ns, VDD,
+ 1164369.600000ns, VSS,
+ 1165090.100000ns, VSS,
+ 1165090.200000ns, VDD,
+ 1165570.500000ns, VDD,
+ 1165570.600000ns, VSS,
+ 1165690.600000ns, VSS,
+ 1165690.700000ns, VDD,
+ 1166771.500000ns, VDD,
+ 1166771.600000ns, VSS,
+ 1167251.900000ns, VSS,
+ 1167252.000000ns, VDD,
+ 1167852.400000ns, VDD,
+ 1167852.500000ns, VSS,
+ 1168332.800000ns, VSS,
+ 1168332.900000ns, VDD,
+ 1170134.300000ns, VDD,
+ 1170134.400000ns, VSS,
+ 1170374.500000ns, VSS,
+ 1170374.600000ns, VDD,
+ 1171095.100000ns, VDD,
+ 1171095.200000ns, VSS,
+ 1171575.500000ns, VSS,
+ 1171575.600000ns, VDD,
+ 1171815.700000ns, VDD,
+ 1171815.800000ns, VSS,
+ 1172536.300000ns, VSS,
+ 1172536.400000ns, VDD,
+ 1172896.600000ns, VDD,
+ 1172896.700000ns, VSS,
+ 1173737.300000ns, VSS,
+ 1173737.400000ns, VDD,
+ 1174097.600000ns, VDD,
+ 1174097.700000ns, VSS,
+ 1174578.000000ns, VSS,
+ 1174578.100000ns, VDD,
+ 1175418.700000ns, VDD,
+ 1175418.800000ns, VSS,
+ 1176019.200000ns, VSS,
+ 1176019.300000ns, VDD,
+ 1177340.300000ns, VDD,
+ 1177340.400000ns, VSS,
+ 1178901.600000ns, VSS,
+ 1178901.700000ns, VDD,
+ 1180462.900000ns, VDD,
+ 1180463.000000ns, VSS,
+ 1180823.200000ns, VSS,
+ 1180823.300000ns, VDD,
+ 1181303.600000ns, VDD,
+ 1181303.700000ns, VSS,
+ 1181784.000000ns, VSS,
+ 1181784.100000ns, VDD,
+ 1181904.100000ns, VDD,
+ 1181904.200000ns, VSS,
+ 1183225.200000ns, VSS,
+ 1183225.300000ns, VDD,
+ 1183705.600000ns, VDD,
+ 1183705.700000ns, VSS,
+ 1184426.200000ns, VSS,
+ 1184426.300000ns, VDD,
+ 1184666.400000ns, VDD,
+ 1184666.500000ns, VSS,
+ 1185146.800000ns, VSS,
+ 1185146.900000ns, VDD,
+ 1185747.300000ns, VDD,
+ 1185747.400000ns, VSS,
+ 1186347.800000ns, VSS,
+ 1186347.900000ns, VDD,
+ 1187308.600000ns, VDD,
+ 1187308.700000ns, VSS,
+ 1187789.000000ns, VSS,
+ 1187789.100000ns, VDD,
+ 1189830.700000ns, VDD,
+ 1189830.800000ns, VSS,
+ 1190551.300000ns, VSS,
+ 1190551.400000ns, VDD,
+ 1191512.100000ns, VDD,
+ 1191512.200000ns, VSS,
+ 1191752.300000ns, VSS,
+ 1191752.400000ns, VDD,
+ 1193673.900000ns, VDD,
+ 1193674.000000ns, VSS,
+ 1193794.000000ns, VSS,
+ 1193794.100000ns, VDD,
+ 1194034.200000ns, VDD,
+ 1194034.300000ns, VSS,
+ 1194154.300000ns, VSS,
+ 1194154.400000ns, VDD,
+ 1194514.600000ns, VDD,
+ 1194514.700000ns, VSS,
+ 1194995.000000ns, VSS,
+ 1194995.100000ns, VDD,
+ 1195235.200000ns, VDD,
+ 1195235.300000ns, VSS,
+ 1195355.300000ns, VSS,
+ 1195355.400000ns, VDD,
+ 1195475.400000ns, VDD,
+ 1195475.500000ns, VSS,
+ 1196316.100000ns, VSS,
+ 1196316.200000ns, VDD,
+ 1197877.400000ns, VDD,
+ 1197877.500000ns, VSS,
+ 1198357.800000ns, VSS,
+ 1198357.900000ns, VDD,
+ 1198718.100000ns, VDD,
+ 1198718.200000ns, VSS,
+ 1198958.300000ns, VSS,
+ 1198958.400000ns, VDD,
+ 1199198.500000ns, VDD,
+ 1199198.600000ns, VSS,
+ 1200639.700000ns, VSS,
+ 1200639.800000ns, VDD,
+ 1200759.800000ns, VDD,
+ 1200759.900000ns, VSS,
+ 1201240.200000ns, VSS,
+ 1201240.300000ns, VDD,
+ 1201360.300000ns, VDD,
+ 1201360.400000ns, VSS,
+ 1202201.000000ns, VSS,
+ 1202201.100000ns, VDD,
+ 1202561.300000ns, VDD,
+ 1202561.400000ns, VSS,
+ 1202801.500000ns, VSS,
+ 1202801.600000ns, VDD,
+ 1203041.700000ns, VDD,
+ 1203041.800000ns, VSS,
+ 1203402.000000ns, VSS,
+ 1203402.100000ns, VDD,
+ 1204122.600000ns, VDD,
+ 1204122.700000ns, VSS,
+ 1204603.000000ns, VSS,
+ 1204603.100000ns, VDD,
+ 1205083.400000ns, VDD,
+ 1205083.500000ns, VSS,
+ 1206044.200000ns, VSS,
+ 1206044.300000ns, VDD,
+ 1207125.100000ns, VDD,
+ 1207125.200000ns, VSS,
+ 1207965.800000ns, VSS,
+ 1207965.900000ns, VDD,
+ 1208806.500000ns, VDD,
+ 1208806.600000ns, VSS,
+ 1212169.300000ns, VSS,
+ 1212169.400000ns, VDD,
+ 1212409.500000ns, VDD,
+ 1212409.600000ns, VSS,
+ 1213370.300000ns, VSS,
+ 1213370.400000ns, VDD,
+ 1214811.500000ns, VDD,
+ 1214811.600000ns, VSS,
+ 1215772.300000ns, VSS,
+ 1215772.400000ns, VDD,
+ 1216132.600000ns, VDD,
+ 1216132.700000ns, VSS,
+ 1216492.900000ns, VSS,
+ 1216493.000000ns, VDD,
+ 1216613.000000ns, VDD,
+ 1216613.100000ns, VSS,
+ 1216733.100000ns, VSS,
+ 1216733.200000ns, VDD,
+ 1218054.200000ns, VDD,
+ 1218054.300000ns, VSS,
+ 1218174.300000ns, VSS,
+ 1218174.400000ns, VDD,
+ 1218294.400000ns, VDD,
+ 1218294.500000ns, VSS,
+ 1218534.600000ns, VSS,
+ 1218534.700000ns, VDD,
+ 1219495.400000ns, VDD,
+ 1219495.500000ns, VSS,
+ 1220336.100000ns, VSS,
+ 1220336.200000ns, VDD,
+ 1220816.500000ns, VDD,
+ 1220816.600000ns, VSS,
+ 1221056.700000ns, VSS,
+ 1221056.800000ns, VDD,
+ 1221657.200000ns, VDD,
+ 1221657.300000ns, VSS,
+ 1222497.900000ns, VSS,
+ 1222498.000000ns, VDD,
+ 1222618.000000ns, VDD,
+ 1222618.100000ns, VSS,
+ 1223218.500000ns, VSS,
+ 1223218.600000ns, VDD,
+ 1223939.100000ns, VDD,
+ 1223939.200000ns, VSS,
+ 1225260.200000ns, VSS,
+ 1225260.300000ns, VDD,
+ 1225740.600000ns, VDD,
+ 1225740.700000ns, VSS,
+ 1225860.700000ns, VSS,
+ 1225860.800000ns, VDD,
+ 1226341.100000ns, VDD,
+ 1226341.200000ns, VSS,
+ 1226461.200000ns, VSS,
+ 1226461.300000ns, VDD,
+ 1226821.500000ns, VDD,
+ 1226821.600000ns, VSS,
+ 1227061.700000ns, VSS,
+ 1227061.800000ns, VDD,
+ 1228743.100000ns, VDD,
+ 1228743.200000ns, VSS,
+ 1231265.200000ns, VSS,
+ 1231265.300000ns, VDD,
+ 1232826.500000ns, VDD,
+ 1232826.600000ns, VSS,
+ 1233306.900000ns, VSS,
+ 1233307.000000ns, VDD,
+ 1234387.800000ns, VDD,
+ 1234387.900000ns, VSS,
+ 1234748.100000ns, VSS,
+ 1234748.200000ns, VDD,
+ 1237270.200000ns, VDD,
+ 1237270.300000ns, VSS,
+ 1237990.800000ns, VSS,
+ 1237990.900000ns, VDD,
+ 1238231.000000ns, VDD,
+ 1238231.100000ns, VSS,
+ 1239912.400000ns, VSS,
+ 1239912.500000ns, VDD,
+ 1240272.700000ns, VDD,
+ 1240272.800000ns, VSS,
+ 1241473.700000ns, VSS,
+ 1241473.800000ns, VDD,
+ 1241954.100000ns, VDD,
+ 1241954.200000ns, VSS,
+ 1242314.400000ns, VSS,
+ 1242314.500000ns, VDD,
+ 1244115.900000ns, VDD,
+ 1244116.000000ns, VSS,
+ 1244236.000000ns, VSS,
+ 1244236.100000ns, VDD,
+ 1244476.200000ns, VDD,
+ 1244476.300000ns, VSS,
+ 1244716.400000ns, VSS,
+ 1244716.500000ns, VDD,
+ 1245557.100000ns, VDD,
+ 1245557.200000ns, VSS,
+ 1246037.500000ns, VSS,
+ 1246037.600000ns, VDD,
+ 1246517.900000ns, VDD,
+ 1246518.000000ns, VSS,
+ 1246638.000000ns, VSS,
+ 1246638.100000ns, VDD,
+ 1246758.100000ns, VDD,
+ 1246758.200000ns, VSS,
+ 1246998.300000ns, VSS,
+ 1246998.400000ns, VDD,
+ 1247238.500000ns, VDD,
+ 1247238.600000ns, VSS,
+ 1248559.600000ns, VSS,
+ 1248559.700000ns, VDD,
+ 1250120.900000ns, VDD,
+ 1250121.000000ns, VSS,
+ 1250601.300000ns, VSS,
+ 1250601.400000ns, VDD,
+ 1250721.400000ns, VDD,
+ 1250721.500000ns, VSS,
+ 1251201.800000ns, VSS,
+ 1251201.900000ns, VDD,
+ 1251682.200000ns, VDD,
+ 1251682.300000ns, VSS,
+ 1252522.900000ns, VSS,
+ 1252523.000000ns, VDD,
+ 1252643.000000ns, VDD,
+ 1252643.100000ns, VSS,
+ 1252883.200000ns, VSS,
+ 1252883.300000ns, VDD,
+ 1253603.800000ns, VDD,
+ 1253603.900000ns, VSS,
+ 1253723.900000ns, VSS,
+ 1253724.000000ns, VDD,
+ 1254324.400000ns, VDD,
+ 1254324.500000ns, VSS,
+ 1254444.500000ns, VSS,
+ 1254444.600000ns, VDD,
+ 1254684.700000ns, VDD,
+ 1254684.800000ns, VSS,
+ 1254924.900000ns, VSS,
+ 1254925.000000ns, VDD,
+ 1255645.500000ns, VDD,
+ 1255645.600000ns, VSS,
+ 1256846.500000ns, VSS,
+ 1256846.600000ns, VDD,
+ 1257807.300000ns, VDD,
+ 1257807.400000ns, VSS,
+ 1258407.800000ns, VSS,
+ 1258407.900000ns, VDD,
+ 1259008.300000ns, VDD,
+ 1259008.400000ns, VSS,
+ 1259488.700000ns, VSS,
+ 1259488.800000ns, VDD,
+ 1259849.000000ns, VDD,
+ 1259849.100000ns, VSS,
+ 1259969.100000ns, VSS,
+ 1259969.200000ns, VDD,
+ 1260689.700000ns, VDD,
+ 1260689.800000ns, VSS,
+ 1260929.900000ns, VSS,
+ 1260930.000000ns, VDD,
+ 1261050.000000ns, VDD,
+ 1261050.100000ns, VSS,
+ 1261170.100000ns, VSS,
+ 1261170.200000ns, VDD,
+ 1262251.000000ns, VDD,
+ 1262251.100000ns, VSS,
+ 1264773.100000ns, VSS,
+ 1264773.200000ns, VDD,
+ 1265013.300000ns, VDD,
+ 1265013.400000ns, VSS,
+ 1265133.400000ns, VSS,
+ 1265133.500000ns, VDD,
+ 1265373.600000ns, VDD,
+ 1265373.700000ns, VSS,
+ 1268256.000000ns, VSS,
+ 1268256.100000ns, VDD,
+ 1269697.200000ns, VDD,
+ 1269697.300000ns, VSS,
+ 1272219.300000ns, VSS,
+ 1272219.400000ns, VDD,
+ 1273420.300000ns, VDD,
+ 1273420.400000ns, VSS,
+ 1273780.600000ns, VSS,
+ 1273780.700000ns, VDD,
+ 1274140.900000ns, VDD,
+ 1274141.000000ns, VSS,
+ 1274861.500000ns, VSS,
+ 1274861.600000ns, VDD,
+ 1275101.700000ns, VDD,
+ 1275101.800000ns, VSS,
+ 1275221.800000ns, VSS,
+ 1275221.900000ns, VDD,
+ 1275462.000000ns, VDD,
+ 1275462.100000ns, VSS,
+ 1275582.100000ns, VSS,
+ 1275582.200000ns, VDD,
+ 1276302.700000ns, VDD,
+ 1276302.800000ns, VSS,
+ 1276422.800000ns, VSS,
+ 1276422.900000ns, VDD,
+ 1277023.300000ns, VDD,
+ 1277023.400000ns, VSS,
+ 1278104.200000ns, VSS,
+ 1278104.300000ns, VDD,
+ 1278584.600000ns, VDD,
+ 1278584.700000ns, VSS,
+ 1280386.100000ns, VSS,
+ 1280386.200000ns, VDD,
+ 1280506.200000ns, VDD,
+ 1280506.300000ns, VSS,
+ 1280986.600000ns, VSS,
+ 1280986.700000ns, VDD,
+ 1281346.900000ns, VDD,
+ 1281347.000000ns, VSS,
+ 1281467.000000ns, VSS,
+ 1281467.100000ns, VDD,
+ 1283508.700000ns, VDD,
+ 1283508.800000ns, VSS,
+ 1283989.100000ns, VSS,
+ 1283989.200000ns, VDD,
+ 1285430.300000ns, VDD,
+ 1285430.400000ns, VSS,
+ 1286271.000000ns, VSS,
+ 1286271.100000ns, VDD,
+ 1286631.300000ns, VDD,
+ 1286631.400000ns, VSS,
+ 1287351.900000ns, VSS,
+ 1287352.000000ns, VDD,
+ 1287472.000000ns, VDD,
+ 1287472.100000ns, VSS,
+ 1287592.100000ns, VSS,
+ 1287592.200000ns, VDD,
+ 1289393.600000ns, VDD,
+ 1289393.700000ns, VSS,
+ 1289994.100000ns, VSS,
+ 1289994.200000ns, VDD,
+ 1290354.400000ns, VDD,
+ 1290354.500000ns, VSS,
+ 1291795.600000ns, VSS,
+ 1291795.700000ns, VDD,
+ 1292876.500000ns, VDD,
+ 1292876.600000ns, VSS,
+ 1293356.900000ns, VSS,
+ 1293357.000000ns, VDD,
+ 1294077.500000ns, VDD,
+ 1294077.600000ns, VSS,
+ 1294317.700000ns, VSS,
+ 1294317.800000ns, VDD,
+ 1294557.900000ns, VDD,
+ 1294558.000000ns, VSS,
+ 1295038.300000ns, VSS,
+ 1295038.400000ns, VDD,
+ 1295758.900000ns, VDD,
+ 1295759.000000ns, VSS,
+ 1296119.200000ns, VSS,
+ 1296119.300000ns, VDD,
+ 1296239.300000ns, VDD,
+ 1296239.400000ns, VSS,
+ 1297320.200000ns, VSS,
+ 1297320.300000ns, VDD,
+ 1297800.600000ns, VDD,
+ 1297800.700000ns, VSS,
+ 1298401.100000ns, VSS,
+ 1298401.200000ns, VDD,
+ 1300082.500000ns, VDD,
+ 1300082.600000ns, VSS,
+ 1300803.100000ns, VSS,
+ 1300803.200000ns, VDD,
+ 1300923.200000ns, VDD,
+ 1300923.300000ns, VSS,
+ 1301523.700000ns, VSS,
+ 1301523.800000ns, VDD,
+ 1302124.200000ns, VDD,
+ 1302124.300000ns, VSS,
+ 1302244.300000ns, VSS,
+ 1302244.400000ns, VDD,
+ 1302844.800000ns, VDD,
+ 1302844.900000ns, VSS,
+ 1303685.500000ns, VSS,
+ 1303685.600000ns, VDD,
+ 1303805.600000ns, VDD,
+ 1303805.700000ns, VSS,
+ 1304406.100000ns, VSS,
+ 1304406.200000ns, VDD,
+ 1304646.300000ns, VDD,
+ 1304646.400000ns, VSS,
+ 1304766.400000ns, VSS,
+ 1304766.500000ns, VDD,
+ 1304886.500000ns, VDD,
+ 1304886.600000ns, VSS,
+ 1305727.200000ns, VSS,
+ 1305727.300000ns, VDD,
+ 1306087.500000ns, VDD,
+ 1306087.600000ns, VSS,
+ 1306688.000000ns, VSS,
+ 1306688.100000ns, VDD,
+ 1306928.200000ns, VDD,
+ 1306928.300000ns, VSS,
+ 1308969.900000ns, VSS,
+ 1308970.000000ns, VDD,
+ 1309570.400000ns, VDD,
+ 1309570.500000ns, VSS,
+ 1310170.900000ns, VSS,
+ 1310171.000000ns, VDD,
+ 1310291.000000ns, VDD,
+ 1310291.100000ns, VSS,
+ 1310891.500000ns, VSS,
+ 1310891.600000ns, VDD,
+ 1311612.100000ns, VDD,
+ 1311612.200000ns, VSS,
+ 1311732.200000ns, VSS,
+ 1311732.300000ns, VDD,
+ 1312212.600000ns, VDD,
+ 1312212.700000ns, VSS,
+ 1312933.200000ns, VSS,
+ 1312933.300000ns, VDD,
+ 1313413.600000ns, VDD,
+ 1313413.700000ns, VSS,
+ 1313773.900000ns, VSS,
+ 1313774.000000ns, VDD,
+ 1314254.300000ns, VDD,
+ 1314254.400000ns, VSS,
+ 1314614.600000ns, VSS,
+ 1314614.700000ns, VDD,
+ 1314974.900000ns, VDD,
+ 1314975.000000ns, VSS,
+ 1315455.300000ns, VSS,
+ 1315455.400000ns, VDD,
+ 1315695.500000ns, VDD,
+ 1315695.600000ns, VSS,
+ 1315815.600000ns, VSS,
+ 1315815.700000ns, VDD,
+ 1315935.700000ns, VDD,
+ 1315935.800000ns, VSS,
+ 1316175.900000ns, VSS,
+ 1316176.000000ns, VDD,
+ 1317857.300000ns, VDD,
+ 1317857.400000ns, VSS,
+ 1318938.200000ns, VSS,
+ 1318938.300000ns, VDD,
+ 1319418.600000ns, VDD,
+ 1319418.700000ns, VSS,
+ 1320019.100000ns, VSS,
+ 1320019.200000ns, VDD,
+ 1320499.500000ns, VDD,
+ 1320499.600000ns, VSS,
+ 1320979.900000ns, VSS,
+ 1320980.000000ns, VDD,
+ 1321100.000000ns, VDD,
+ 1321100.100000ns, VSS,
+ 1321700.500000ns, VSS,
+ 1321700.600000ns, VDD,
+ 1322421.100000ns, VDD,
+ 1322421.200000ns, VSS,
+ 1322901.500000ns, VSS,
+ 1322901.600000ns, VDD,
+ 1323381.900000ns, VDD,
+ 1323382.000000ns, VSS,
+ 1323862.300000ns, VSS,
+ 1323862.400000ns, VDD,
+ 1324462.800000ns, VDD,
+ 1324462.900000ns, VSS,
+ 1324823.100000ns, VSS,
+ 1324823.200000ns, VDD,
+ 1325303.500000ns, VDD,
+ 1325303.600000ns, VSS,
+ 1325543.700000ns, VSS,
+ 1325543.800000ns, VDD,
+ 1325904.000000ns, VDD,
+ 1325904.100000ns, VSS,
+ 1326504.500000ns, VSS,
+ 1326504.600000ns, VDD,
+ 1327105.000000ns, VDD,
+ 1327105.100000ns, VSS,
+ 1327345.200000ns, VSS,
+ 1327345.300000ns, VDD,
+ 1328185.900000ns, VDD,
+ 1328186.000000ns, VSS,
+ 1328546.200000ns, VSS,
+ 1328546.300000ns, VDD,
+ 1329987.400000ns, VDD,
+ 1329987.500000ns, VSS,
+ 1330227.600000ns, VSS,
+ 1330227.700000ns, VDD,
+ 1330467.800000ns, VDD,
+ 1330467.900000ns, VSS,
+ 1332629.600000ns, VSS,
+ 1332629.700000ns, VDD,
+ 1333230.100000ns, VDD,
+ 1333230.200000ns, VSS,
+ 1333350.200000ns, VSS,
+ 1333350.300000ns, VDD,
+ 1333710.500000ns, VDD,
+ 1333710.600000ns, VSS,
+ 1334190.900000ns, VSS,
+ 1334191.000000ns, VDD,
+ 1334671.300000ns, VDD,
+ 1334671.400000ns, VSS,
+ 1335031.600000ns, VSS,
+ 1335031.700000ns, VDD,
+ 1335752.200000ns, VDD,
+ 1335752.300000ns, VSS,
+ 1336953.200000ns, VSS,
+ 1336953.300000ns, VDD,
+ 1337193.400000ns, VDD,
+ 1337193.500000ns, VSS,
+ 1337553.700000ns, VSS,
+ 1337553.800000ns, VDD,
+ 1339115.000000ns, VDD,
+ 1339115.100000ns, VSS,
+ 1340316.000000ns, VSS,
+ 1340316.100000ns, VDD,
+ 1340796.400000ns, VDD,
+ 1340796.500000ns, VSS,
+ 1341276.800000ns, VSS,
+ 1341276.900000ns, VDD,
+ 1342718.000000ns, VDD,
+ 1342718.100000ns, VSS,
+ 1343318.500000ns, VSS,
+ 1343318.600000ns, VDD,
+ 1343558.700000ns, VDD,
+ 1343558.800000ns, VSS,
+ 1344039.100000ns, VSS,
+ 1344039.200000ns, VDD,
+ 1344879.800000ns, VDD,
+ 1344879.900000ns, VSS,
+ 1345360.200000ns, VSS,
+ 1345360.300000ns, VDD,
+ 1346080.800000ns, VDD,
+ 1346080.900000ns, VSS,
+ 1346200.900000ns, VSS,
+ 1346201.000000ns, VDD,
+ 1347041.600000ns, VDD,
+ 1347041.700000ns, VSS,
+ 1347762.200000ns, VSS,
+ 1347762.300000ns, VDD,
+ 1348242.600000ns, VDD,
+ 1348242.700000ns, VSS,
+ 1348602.900000ns, VSS,
+ 1348603.000000ns, VDD,
+ 1348963.200000ns, VDD,
+ 1348963.300000ns, VSS,
+ 1349083.300000ns, VSS,
+ 1349083.400000ns, VDD,
+ 1349683.800000ns, VDD,
+ 1349683.900000ns, VSS,
+ 1350044.100000ns, VSS,
+ 1350044.200000ns, VDD,
+ 1350284.300000ns, VDD,
+ 1350284.400000ns, VSS,
+ 1351004.900000ns, VSS,
+ 1351005.000000ns, VDD,
+ 1351965.700000ns, VDD,
+ 1351965.800000ns, VSS,
+ 1353166.700000ns, VSS,
+ 1353166.800000ns, VDD,
+ 1353406.900000ns, VDD,
+ 1353407.000000ns, VSS,
+ 1354848.100000ns, VSS,
+ 1354848.200000ns, VDD,
+ 1354968.200000ns, VDD,
+ 1354968.300000ns, VSS,
+ 1355328.500000ns, VSS,
+ 1355328.600000ns, VDD,
+ 1355929.000000ns, VDD,
+ 1355929.100000ns, VSS,
+ 1356289.300000ns, VSS,
+ 1356289.400000ns, VDD,
+ 1356769.700000ns, VDD,
+ 1356769.800000ns, VSS,
+ 1356889.800000ns, VSS,
+ 1356889.900000ns, VDD,
+ 1357490.300000ns, VDD,
+ 1357490.400000ns, VSS,
+ 1357970.700000ns, VSS,
+ 1357970.800000ns, VDD,
+ 1358811.400000ns, VDD,
+ 1358811.500000ns, VSS,
+ 1358931.500000ns, VSS,
+ 1358931.600000ns, VDD,
+ 1359051.600000ns, VDD,
+ 1359051.700000ns, VSS,
+ 1359532.000000ns, VSS,
+ 1359532.100000ns, VDD,
+ 1360252.600000ns, VDD,
+ 1360252.700000ns, VSS,
+ 1360733.000000ns, VSS,
+ 1360733.100000ns, VDD,
+ 1361213.400000ns, VDD,
+ 1361213.500000ns, VSS,
+ 1361693.800000ns, VSS,
+ 1361693.900000ns, VDD,
+ 1362174.200000ns, VDD,
+ 1362174.300000ns, VSS,
+ 1362534.500000ns, VSS,
+ 1362534.600000ns, VDD,
+ 1362894.800000ns, VDD,
+ 1362894.900000ns, VSS,
+ 1363255.100000ns, VSS,
+ 1363255.200000ns, VDD,
+ 1363855.600000ns, VDD,
+ 1363855.700000ns, VSS,
+ 1363975.700000ns, VSS,
+ 1363975.800000ns, VDD,
+ 1364936.500000ns, VDD,
+ 1364936.600000ns, VSS,
+ 1365056.600000ns, VSS,
+ 1365056.700000ns, VDD,
+ 1365176.700000ns, VDD,
+ 1365176.800000ns, VSS,
+ 1365537.000000ns, VSS,
+ 1365537.100000ns, VDD,
+ 1366257.600000ns, VDD,
+ 1366257.700000ns, VSS,
+ 1366978.200000ns, VSS,
+ 1366978.300000ns, VDD,
+ 1367698.800000ns, VDD,
+ 1367698.900000ns, VSS,
+ 1370821.400000ns, VSS,
+ 1370821.500000ns, VDD,
+ 1372142.500000ns, VDD,
+ 1372142.600000ns, VSS,
+ 1373463.600000ns, VSS,
+ 1373463.700000ns, VDD,
+ 1373823.900000ns, VDD,
+ 1373824.000000ns, VSS,
+ 1374304.300000ns, VSS,
+ 1374304.400000ns, VDD,
+ 1374904.800000ns, VDD,
+ 1374904.900000ns, VSS,
+ 1375985.700000ns, VSS,
+ 1375985.800000ns, VDD,
+ 1376225.900000ns, VDD,
+ 1376226.000000ns, VSS,
+ 1376706.300000ns, VSS,
+ 1376706.400000ns, VDD,
+ 1377186.700000ns, VDD,
+ 1377186.800000ns, VSS,
+ 1377667.100000ns, VSS,
+ 1377667.200000ns, VDD,
+ 1378147.500000ns, VDD,
+ 1378147.600000ns, VSS,
+ 1378507.800000ns, VSS,
+ 1378507.900000ns, VDD,
+ 1378627.900000ns, VDD,
+ 1378628.000000ns, VSS,
+ 1379108.300000ns, VSS,
+ 1379108.400000ns, VDD,
+ 1379708.800000ns, VDD,
+ 1379708.900000ns, VSS,
+ 1380429.400000ns, VSS,
+ 1380429.500000ns, VDD,
+ 1382351.000000ns, VDD,
+ 1382351.100000ns, VSS,
+ 1383071.600000ns, VSS,
+ 1383071.700000ns, VDD,
+ 1383672.100000ns, VDD,
+ 1383672.200000ns, VSS,
+ 1385233.400000ns, VSS,
+ 1385233.500000ns, VDD,
+ 1386554.500000ns, VDD,
+ 1386554.600000ns, VSS,
+ 1387875.600000ns, VSS,
+ 1387875.700000ns, VDD,
+ 1388235.900000ns, VDD,
+ 1388236.000000ns, VSS,
+ 1389677.100000ns, VSS,
+ 1389677.200000ns, VDD,
+ 1390157.500000ns, VDD,
+ 1390157.600000ns, VSS,
+ 1390758.000000ns, VSS,
+ 1390758.100000ns, VDD,
+ 1392919.800000ns, VDD,
+ 1392919.900000ns, VSS,
+ 1393039.900000ns, VSS,
+ 1393040.000000ns, VDD,
+ 1393280.100000ns, VDD,
+ 1393280.200000ns, VSS,
+ 1393880.600000ns, VSS,
+ 1393880.700000ns, VDD,
+ 1394240.900000ns, VDD,
+ 1394241.000000ns, VSS,
+ 1395441.900000ns, VSS,
+ 1395442.000000ns, VDD,
+ 1395802.200000ns, VDD,
+ 1395802.300000ns, VSS,
+ 1396883.100000ns, VSS,
+ 1396883.200000ns, VDD,
+ 1397003.200000ns, VDD,
+ 1397003.300000ns, VSS,
+ 1397723.800000ns, VSS,
+ 1397723.900000ns, VDD,
+ 1397843.900000ns, VDD,
+ 1397844.000000ns, VSS,
+ 1398084.100000ns, VSS,
+ 1398084.200000ns, VDD,
+ 1398204.200000ns, VDD,
+ 1398204.300000ns, VSS,
+ 1398324.300000ns, VSS,
+ 1398324.400000ns, VDD,
+ 1398924.800000ns, VDD,
+ 1398924.900000ns, VSS,
+ 1399044.900000ns, VSS,
+ 1399045.000000ns, VDD,
+ 1399165.000000ns, VDD,
+ 1399165.100000ns, VSS,
+ 1399765.500000ns, VSS,
+ 1399765.600000ns, VDD,
+ 1400005.700000ns, VDD,
+ 1400005.800000ns, VSS,
+ 1400726.300000ns, VSS,
+ 1400726.400000ns, VDD,
+ 1400966.500000ns, VDD,
+ 1400966.600000ns, VSS,
+ 1401086.600000ns, VSS,
+ 1401086.700000ns, VDD,
+ 1402647.900000ns, VDD,
+ 1402648.000000ns, VSS,
+ 1403848.900000ns, VSS,
+ 1403849.000000ns, VDD,
+ 1405170.000000ns, VDD,
+ 1405170.100000ns, VSS,
+ 1406250.900000ns, VSS,
+ 1406251.000000ns, VDD,
+ 1406731.300000ns, VDD,
+ 1406731.400000ns, VSS,
+ 1407211.700000ns, VSS,
+ 1407211.800000ns, VDD,
+ 1407331.800000ns, VDD,
+ 1407331.900000ns, VSS,
+ 1407812.200000ns, VSS,
+ 1407812.300000ns, VDD,
+ 1407932.300000ns, VDD,
+ 1407932.400000ns, VSS,
+ 1408652.900000ns, VSS,
+ 1408653.000000ns, VDD,
+ 1408773.000000ns, VDD,
+ 1408773.100000ns, VSS,
+ 1408893.100000ns, VSS,
+ 1408893.200000ns, VDD,
+ 1409613.700000ns, VDD,
+ 1409613.800000ns, VSS,
+ 1410574.500000ns, VSS,
+ 1410574.600000ns, VDD,
+ 1410694.600000ns, VDD,
+ 1410694.700000ns, VSS,
+ 1410814.700000ns, VSS,
+ 1410814.800000ns, VDD,
+ 1411775.500000ns, VDD,
+ 1411775.600000ns, VSS,
+ 1414417.700000ns, VSS,
+ 1414417.800000ns, VDD,
+ 1414537.800000ns, VDD,
+ 1414537.900000ns, VSS,
+ 1415858.900000ns, VSS,
+ 1415859.000000ns, VDD,
+ 1416819.700000ns, VDD,
+ 1416819.800000ns, VSS,
+ 1416939.800000ns, VSS,
+ 1416939.900000ns, VDD,
+ 1417420.200000ns, VDD,
+ 1417420.300000ns, VSS,
+ 1418140.800000ns, VSS,
+ 1418140.900000ns, VDD,
+ 1421263.400000ns, VDD,
+ 1421263.500000ns, VSS,
+ 1421383.500000ns, VSS,
+ 1421383.600000ns, VDD,
+ 1421503.600000ns, VDD,
+ 1421503.700000ns, VSS,
+ 1422824.700000ns, VSS,
+ 1422824.800000ns, VDD,
+ 1423064.900000ns, VDD,
+ 1423065.000000ns, VSS,
+ 1424265.900000ns, VSS,
+ 1424266.000000ns, VDD,
+ 1424386.000000ns, VDD,
+ 1424386.100000ns, VSS,
+ 1425106.600000ns, VSS,
+ 1425106.700000ns, VDD,
+ 1425587.000000ns, VDD,
+ 1425587.100000ns, VSS,
+ 1427268.400000ns, VSS,
+ 1427268.500000ns, VDD,
+ 1427628.700000ns, VDD,
+ 1427628.800000ns, VSS,
+ 1428589.500000ns, VSS,
+ 1428589.600000ns, VDD,
+ 1428709.600000ns, VDD,
+ 1428709.700000ns, VSS,
+ 1429190.000000ns, VSS,
+ 1429190.100000ns, VDD,
+ 1430150.800000ns, VDD,
+ 1430150.900000ns, VSS,
+ 1430391.000000ns, VSS,
+ 1430391.100000ns, VDD,
+ 1430631.200000ns, VDD,
+ 1430631.300000ns, VSS,
+ 1433393.500000ns, VSS,
+ 1433393.600000ns, VDD,
+ 1433633.700000ns, VDD,
+ 1433633.800000ns, VSS,
+ 1433873.900000ns, VSS,
+ 1433874.000000ns, VDD,
+ 1434114.100000ns, VDD,
+ 1434114.200000ns, VSS,
+ 1434714.600000ns, VSS,
+ 1434714.700000ns, VDD,
+ 1435555.300000ns, VDD,
+ 1435555.400000ns, VSS,
+ 1435675.400000ns, VSS,
+ 1435675.500000ns, VDD,
+ 1435915.600000ns, VDD,
+ 1435915.700000ns, VSS,
+ 1436275.900000ns, VSS,
+ 1436276.000000ns, VDD,
+ 1436756.300000ns, VDD,
+ 1436756.400000ns, VSS,
+ 1437837.200000ns, VSS,
+ 1437837.300000ns, VDD,
+ 1437957.300000ns, VDD,
+ 1437957.400000ns, VSS,
+ 1438317.600000ns, VSS,
+ 1438317.700000ns, VDD,
+ 1439038.200000ns, VDD,
+ 1439038.300000ns, VSS,
+ 1439518.600000ns, VSS,
+ 1439518.700000ns, VDD,
+ 1439999.000000ns, VDD,
+ 1439999.100000ns, VSS,
+ 1440239.200000ns, VSS,
+ 1440239.300000ns, VDD,
+ 1440959.800000ns, VDD,
+ 1440959.900000ns, VSS,
+ 1441200.000000ns, VSS,
+ 1441200.100000ns, VDD,
+ 1442040.700000ns, VDD,
+ 1442040.800000ns, VSS,
+ 1442160.800000ns, VSS,
+ 1442160.900000ns, VDD,
+ 1442881.400000ns, VDD,
+ 1442881.500000ns, VSS,
+ 1443241.700000ns, VSS,
+ 1443241.800000ns, VDD,
+ 1444082.400000ns, VDD,
+ 1444082.500000ns, VSS,
+ 1444322.600000ns, VSS,
+ 1444322.700000ns, VDD,
+ 1445403.500000ns, VDD,
+ 1445403.600000ns, VSS,
+ 1446364.300000ns, VSS,
+ 1446364.400000ns, VDD,
+ 1447685.400000ns, VDD,
+ 1447685.500000ns, VSS,
+ 1448165.800000ns, VSS,
+ 1448165.900000ns, VDD,
+ 1450087.400000ns, VDD,
+ 1450087.500000ns, VSS,
+ 1450207.500000ns, VSS,
+ 1450207.600000ns, VDD,
+ 1450327.600000ns, VDD,
+ 1450327.700000ns, VSS,
+ 1451528.600000ns, VSS,
+ 1451528.700000ns, VDD,
+ 1452849.700000ns, VDD,
+ 1452849.800000ns, VSS,
+ 1454170.800000ns, VSS,
+ 1454170.900000ns, VDD,
+ 1454290.900000ns, VDD,
+ 1454291.000000ns, VSS,
+ 1454411.000000ns, VSS,
+ 1454411.100000ns, VDD,
+ 1454771.300000ns, VDD,
+ 1454771.400000ns, VSS,
+ 1455251.700000ns, VSS,
+ 1455251.800000ns, VDD,
+ 1455612.000000ns, VDD,
+ 1455612.100000ns, VSS,
+ 1455972.300000ns, VSS,
+ 1455972.400000ns, VDD,
+ 1456212.500000ns, VDD,
+ 1456212.600000ns, VSS,
+ 1458494.400000ns, VSS,
+ 1458494.500000ns, VDD,
+ 1458614.500000ns, VDD,
+ 1458614.600000ns, VSS,
+ 1460536.100000ns, VSS,
+ 1460536.200000ns, VDD,
+ 1460896.400000ns, VDD,
+ 1460896.500000ns, VSS,
+ 1461857.200000ns, VSS,
+ 1461857.300000ns, VDD,
+ 1462217.500000ns, VDD,
+ 1462217.600000ns, VSS,
+ 1462457.700000ns, VSS,
+ 1462457.800000ns, VDD,
+ 1462697.900000ns, VDD,
+ 1462698.000000ns, VSS,
+ 1462818.000000ns, VSS,
+ 1462818.100000ns, VDD,
+ 1463658.700000ns, VDD,
+ 1463658.800000ns, VSS,
+ 1464019.000000ns, VSS,
+ 1464019.100000ns, VDD,
+ 1464619.500000ns, VDD,
+ 1464619.600000ns, VSS,
+ 1464859.700000ns, VSS,
+ 1464859.800000ns, VDD,
+ 1465099.900000ns, VDD,
+ 1465100.000000ns, VSS,
+ 1466661.200000ns, VSS,
+ 1466661.300000ns, VDD,
+ 1467141.600000ns, VDD,
+ 1467141.700000ns, VSS,
+ 1467742.100000ns, VSS,
+ 1467742.200000ns, VDD,
+ 1467862.200000ns, VDD,
+ 1467862.300000ns, VSS,
+ 1467982.300000ns, VSS,
+ 1467982.400000ns, VDD,
+ 1468222.500000ns, VDD,
+ 1468222.600000ns, VSS,
+ 1469303.400000ns, VSS,
+ 1469303.500000ns, VDD,
+ 1469663.700000ns, VDD,
+ 1469663.800000ns, VSS,
+ 1470024.000000ns, VSS,
+ 1470024.100000ns, VDD,
+ 1470504.400000ns, VDD,
+ 1470504.500000ns, VSS,
+ 1470624.500000ns, VSS,
+ 1470624.600000ns, VDD,
+ 1471225.000000ns, VDD,
+ 1471225.100000ns, VSS,
+ 1471585.300000ns, VSS,
+ 1471585.400000ns, VDD,
+ 1471825.500000ns, VDD,
+ 1471825.600000ns, VSS,
+ 1472426.000000ns, VSS,
+ 1472426.100000ns, VDD,
+ 1473146.600000ns, VDD,
+ 1473146.700000ns, VSS,
+ 1475308.400000ns, VSS,
+ 1475308.500000ns, VDD,
+ 1476269.200000ns, VDD,
+ 1476269.300000ns, VSS,
+ 1476629.500000ns, VSS,
+ 1476629.600000ns, VDD,
+ 1479391.800000ns, VDD,
+ 1479391.900000ns, VSS,
+ 1479632.000000ns, VSS,
+ 1479632.100000ns, VDD,
+ 1479752.100000ns, VDD,
+ 1479752.200000ns, VSS,
+ 1481193.300000ns, VSS,
+ 1481193.400000ns, VDD,
+ 1481313.400000ns, VDD,
+ 1481313.500000ns, VSS,
+ 1481433.500000ns, VSS,
+ 1481433.600000ns, VDD,
+ 1481913.900000ns, VDD,
+ 1481914.000000ns, VSS,
+ 1482394.300000ns, VSS,
+ 1482394.400000ns, VDD,
+ 1482634.500000ns, VDD,
+ 1482634.600000ns, VSS,
+ 1483955.600000ns, VSS,
+ 1483955.700000ns, VDD,
+ 1484436.000000ns, VDD,
+ 1484436.100000ns, VSS,
+ 1485156.600000ns, VSS,
+ 1485156.700000ns, VDD,
+ 1485757.100000ns, VDD,
+ 1485757.200000ns, VSS,
+ 1485877.200000ns, VSS,
+ 1485877.300000ns, VDD,
+ 1485997.300000ns, VDD,
+ 1485997.400000ns, VSS,
+ 1486237.500000ns, VSS,
+ 1486237.600000ns, VDD,
+ 1486597.800000ns, VDD,
+ 1486597.900000ns, VSS,
+ 1487198.300000ns, VSS,
+ 1487198.400000ns, VDD,
+ 1487438.500000ns, VDD,
+ 1487438.600000ns, VSS,
+ 1490561.100000ns, VSS,
+ 1490561.200000ns, VDD,
+ 1491041.500000ns, VDD,
+ 1491041.600000ns, VSS,
+ 1492843.000000ns, VSS,
+ 1492843.100000ns, VDD,
+ 1493083.200000ns, VDD,
+ 1493083.300000ns, VSS,
+ 1493323.400000ns, VSS,
+ 1493323.500000ns, VDD,
+ 1493563.600000ns, VDD,
+ 1493563.700000ns, VSS,
+ 1494524.400000ns, VSS,
+ 1494524.500000ns, VDD,
+ 1495965.600000ns, VDD,
+ 1495965.700000ns, VSS,
+ 1496205.800000ns, VSS,
+ 1496205.900000ns, VDD,
+ 1497526.900000ns, VDD,
+ 1497527.000000ns, VSS,
+ 1498247.500000ns, VSS,
+ 1498247.600000ns, VDD,
+ 1498727.900000ns, VDD,
+ 1498728.000000ns, VSS,
+ 1499688.700000ns, VSS,
+ 1499688.800000ns, VDD,
+ 1500529.400000ns, VDD,
+ 1500529.500000ns, VSS,
+ 1500649.500000ns, VSS,
+ 1500649.600000ns, VDD,
+ 1501250.000000ns, VDD,
+ 1501250.100000ns, VSS,
+ 1502811.300000ns, VSS,
+ 1502811.400000ns, VDD,
+ 1503772.100000ns, VDD,
+ 1503772.200000ns, VSS,
+ 1504492.700000ns, VSS,
+ 1504492.800000ns, VDD,
+ 1506054.000000ns, VDD,
+ 1506054.100000ns, VSS,
+ 1507134.900000ns, VSS,
+ 1507135.000000ns, VDD,
+ 1507255.000000ns, VDD,
+ 1507255.100000ns, VSS,
+ 1508456.000000ns, VSS,
+ 1508456.100000ns, VDD,
+ 1508936.400000ns, VDD,
+ 1508936.500000ns, VSS,
+ 1509416.800000ns, VSS,
+ 1509416.900000ns, VDD,
+ 1509536.900000ns, VDD,
+ 1509537.000000ns, VSS,
+ 1509657.000000ns, VSS,
+ 1509657.100000ns, VDD,
+ 1509897.200000ns, VDD,
+ 1509897.300000ns, VSS,
+ 1510137.400000ns, VSS,
+ 1510137.500000ns, VDD,
+ 1511578.600000ns, VDD,
+ 1511578.700000ns, VSS,
+ 1513380.100000ns, VSS,
+ 1513380.200000ns, VDD,
+ 1513500.200000ns, VDD,
+ 1513500.300000ns, VSS,
+ 1513620.300000ns, VSS,
+ 1513620.400000ns, VDD,
+ 1513980.600000ns, VDD,
+ 1513980.700000ns, VSS,
+ 1514100.700000ns, VSS,
+ 1514100.800000ns, VDD,
+ 1514461.000000ns, VDD,
+ 1514461.100000ns, VSS,
+ 1514941.400000ns, VSS,
+ 1514941.500000ns, VDD,
+ 1515061.500000ns, VDD,
+ 1515061.600000ns, VSS,
+ 1515181.600000ns, VSS,
+ 1515181.700000ns, VDD,
+ 1515301.700000ns, VDD,
+ 1515301.800000ns, VSS,
+ 1515782.100000ns, VSS,
+ 1515782.200000ns, VDD,
+ 1516742.900000ns, VDD,
+ 1516743.000000ns, VSS,
+ 1518424.300000ns, VSS,
+ 1518424.400000ns, VDD,
+ 1518784.600000ns, VDD,
+ 1518784.700000ns, VSS,
+ 1518904.700000ns, VSS,
+ 1518904.800000ns, VDD,
+ 1519745.400000ns, VDD,
+ 1519745.500000ns, VSS,
+ 1521426.800000ns, VSS,
+ 1521426.900000ns, VDD,
+ 1521546.900000ns, VDD,
+ 1521547.000000ns, VSS,
+ 1521667.000000ns, VSS,
+ 1521667.100000ns, VDD,
+ 1522147.400000ns, VDD,
+ 1522147.500000ns, VSS,
+ 1522387.600000ns, VSS,
+ 1522387.700000ns, VDD,
+ 1523348.400000ns, VDD,
+ 1523348.500000ns, VSS,
+ 1523708.700000ns, VSS,
+ 1523708.800000ns, VDD,
+ 1525029.800000ns, VDD,
+ 1525029.900000ns, VSS,
+ 1525630.300000ns, VSS,
+ 1525630.400000ns, VDD,
+ 1526110.700000ns, VDD,
+ 1526110.800000ns, VSS,
+ 1526230.800000ns, VSS,
+ 1526230.900000ns, VDD,
+ 1526350.900000ns, VDD,
+ 1526351.000000ns, VSS,
+ 1527311.700000ns, VSS,
+ 1527311.800000ns, VDD,
+ 1527672.000000ns, VDD,
+ 1527672.100000ns, VSS,
+ 1528272.500000ns, VSS,
+ 1528272.600000ns, VDD,
+ 1528873.000000ns, VDD,
+ 1528873.100000ns, VSS,
+ 1532716.200000ns, VSS,
+ 1532716.300000ns, VDD,
+ 1533196.600000ns, VDD,
+ 1533196.700000ns, VSS,
+ 1533677.000000ns, VSS,
+ 1533677.100000ns, VDD,
+ 1534397.600000ns, VDD,
+ 1534397.700000ns, VSS,
+ 1534637.800000ns, VSS,
+ 1534637.900000ns, VDD,
+ 1535238.300000ns, VDD,
+ 1535238.400000ns, VSS,
+ 1536079.000000ns, VSS,
+ 1536079.100000ns, VDD,
+ 1538721.200000ns, VDD,
+ 1538721.300000ns, VSS,
+ 1538841.300000ns, VSS,
+ 1538841.400000ns, VDD,
+ 1539321.700000ns, VDD,
+ 1539321.800000ns, VSS,
+ 1540042.300000ns, VSS,
+ 1540042.400000ns, VDD,
+ 1540642.800000ns, VDD,
+ 1540642.900000ns, VSS,
+ 1541363.400000ns, VSS,
+ 1541363.500000ns, VDD,
+ 1542324.200000ns, VDD,
+ 1542324.300000ns, VSS,
+ 1542804.600000ns, VSS,
+ 1542804.700000ns, VDD,
+ 1543765.400000ns, VDD,
+ 1543765.500000ns, VSS,
+ 1544486.000000ns, VSS,
+ 1544486.100000ns, VDD,
+ 1545206.600000ns, VDD,
+ 1545206.700000ns, VSS,
+ 1545326.700000ns, VSS,
+ 1545326.800000ns, VDD,
+ 1545807.100000ns, VDD,
+ 1545807.200000ns, VSS,
+ 1546767.900000ns, VSS,
+ 1546768.000000ns, VDD,
+ 1547248.300000ns, VDD,
+ 1547248.400000ns, VSS,
+ 1547728.700000ns, VSS,
+ 1547728.800000ns, VDD,
+ 1548209.100000ns, VDD,
+ 1548209.200000ns, VSS,
+ 1548689.500000ns, VSS,
+ 1548689.600000ns, VDD,
+ 1549290.000000ns, VDD,
+ 1549290.100000ns, VSS,
+ 1549890.500000ns, VSS,
+ 1549890.600000ns, VDD,
+ 1550250.800000ns, VDD,
+ 1550250.900000ns, VSS,
+ 1550370.900000ns, VSS,
+ 1550371.000000ns, VDD
+)}



RSDN in_SDN 0 1.0
BSDN in_SDN 0 V={table(time,
+ 0.100000ns, VSS,
+ 360.300000ns, VSS,
+ 360.400000ns, VDD,
+ 720.600000ns, VDD,
+ 720.700000ns, VSS,
+ 1080.900000ns, VSS,
+ 1081.000000ns, VDD,
+ 1561.300000ns, VDD,
+ 1561.400000ns, VSS,
+ 2522.100000ns, VSS,
+ 2522.200000ns, VDD,
+ 3242.700000ns, VDD,
+ 3242.800000ns, VSS,
+ 3482.900000ns, VSS,
+ 3483.000000ns, VDD,
+ 3843.200000ns, VDD,
+ 3843.300000ns, VSS,
+ 4203.500000ns, VSS,
+ 4203.600000ns, VDD,
+ 5164.300000ns, VDD,
+ 5164.400000ns, VSS,
+ 5284.400000ns, VSS,
+ 5284.500000ns, VDD,
+ 5404.500000ns, VDD,
+ 5404.600000ns, VSS,
+ 5764.800000ns, VSS,
+ 5764.900000ns, VDD,
+ 6725.600000ns, VDD,
+ 6725.700000ns, VSS,
+ 7566.300000ns, VSS,
+ 7566.400000ns, VDD,
+ 8046.700000ns, VDD,
+ 8046.800000ns, VSS,
+ 8767.300000ns, VSS,
+ 8767.400000ns, VDD,
+ 9487.900000ns, VDD,
+ 9488.000000ns, VSS,
+ 9848.200000ns, VSS,
+ 9848.300000ns, VDD,
+ 10809.000000ns, VDD,
+ 10809.100000ns, VSS,
+ 10929.100000ns, VSS,
+ 10929.200000ns, VDD,
+ 11649.700000ns, VDD,
+ 11649.800000ns, VSS,
+ 11889.900000ns, VSS,
+ 11890.000000ns, VDD,
+ 12010.000000ns, VDD,
+ 12010.100000ns, VSS,
+ 12250.200000ns, VSS,
+ 12250.300000ns, VDD,
+ 12490.400000ns, VDD,
+ 12490.500000ns, VSS,
+ 13211.000000ns, VSS,
+ 13211.100000ns, VDD,
+ 13331.100000ns, VDD,
+ 13331.200000ns, VSS,
+ 13451.200000ns, VSS,
+ 13451.300000ns, VDD,
+ 13571.300000ns, VDD,
+ 13571.400000ns, VSS,
+ 14291.900000ns, VSS,
+ 14292.000000ns, VDD,
+ 15613.000000ns, VDD,
+ 15613.100000ns, VSS,
+ 15853.200000ns, VSS,
+ 15853.300000ns, VDD,
+ 15973.300000ns, VDD,
+ 15973.400000ns, VSS,
+ 16213.500000ns, VSS,
+ 16213.600000ns, VDD,
+ 17774.800000ns, VDD,
+ 17774.900000ns, VSS,
+ 17894.900000ns, VSS,
+ 17895.000000ns, VDD,
+ 18975.800000ns, VDD,
+ 18975.900000ns, VSS,
+ 19816.500000ns, VSS,
+ 19816.600000ns, VDD,
+ 19936.600000ns, VDD,
+ 19936.700000ns, VSS,
+ 21257.700000ns, VSS,
+ 21257.800000ns, VDD,
+ 21618.000000ns, VDD,
+ 21618.100000ns, VSS,
+ 22939.100000ns, VSS,
+ 22939.200000ns, VDD,
+ 23539.600000ns, VDD,
+ 23539.700000ns, VSS,
+ 23659.700000ns, VSS,
+ 23659.800000ns, VDD,
+ 24140.100000ns, VDD,
+ 24140.200000ns, VSS,
+ 24260.200000ns, VSS,
+ 24260.300000ns, VDD,
+ 24380.300000ns, VDD,
+ 24380.400000ns, VSS,
+ 24620.500000ns, VSS,
+ 24620.600000ns, VDD,
+ 26061.700000ns, VDD,
+ 26061.800000ns, VSS,
+ 26422.000000ns, VSS,
+ 26422.100000ns, VDD,
+ 26542.100000ns, VDD,
+ 26542.200000ns, VSS,
+ 26902.400000ns, VSS,
+ 26902.500000ns, VDD,
+ 27142.600000ns, VDD,
+ 27142.700000ns, VSS,
+ 27262.700000ns, VSS,
+ 27262.800000ns, VDD,
+ 27623.000000ns, VDD,
+ 27623.100000ns, VSS,
+ 27983.300000ns, VSS,
+ 27983.400000ns, VDD,
+ 28223.500000ns, VDD,
+ 28223.600000ns, VSS,
+ 28343.600000ns, VSS,
+ 28343.700000ns, VDD,
+ 29064.200000ns, VDD,
+ 29064.300000ns, VSS,
+ 29184.300000ns, VSS,
+ 29184.400000ns, VDD,
+ 30385.300000ns, VDD,
+ 30385.400000ns, VSS,
+ 30745.600000ns, VSS,
+ 30745.700000ns, VDD,
+ 30865.700000ns, VDD,
+ 30865.800000ns, VSS,
+ 30985.800000ns, VSS,
+ 30985.900000ns, VDD,
+ 31346.100000ns, VDD,
+ 31346.200000ns, VSS,
+ 31466.200000ns, VSS,
+ 31466.300000ns, VDD,
+ 31706.400000ns, VDD,
+ 31706.500000ns, VSS,
+ 32306.900000ns, VSS,
+ 32307.000000ns, VDD,
+ 32427.000000ns, VDD,
+ 32427.100000ns, VSS,
+ 32787.300000ns, VSS,
+ 32787.400000ns, VDD,
+ 33027.500000ns, VDD,
+ 33027.600000ns, VSS,
+ 33507.900000ns, VSS,
+ 33508.000000ns, VDD,
+ 33748.100000ns, VDD,
+ 33748.200000ns, VSS,
+ 34588.800000ns, VSS,
+ 34588.900000ns, VDD,
+ 35189.300000ns, VDD,
+ 35189.400000ns, VSS,
+ 35309.400000ns, VSS,
+ 35309.500000ns, VDD,
+ 35429.500000ns, VDD,
+ 35429.600000ns, VSS,
+ 35549.600000ns, VSS,
+ 35549.700000ns, VDD,
+ 35909.900000ns, VDD,
+ 35910.000000ns, VSS,
+ 36150.100000ns, VSS,
+ 36150.200000ns, VDD,
+ 36270.200000ns, VDD,
+ 36270.300000ns, VSS,
+ 36390.300000ns, VSS,
+ 36390.400000ns, VDD,
+ 36870.700000ns, VDD,
+ 36870.800000ns, VSS,
+ 36990.800000ns, VSS,
+ 36990.900000ns, VDD,
+ 37110.900000ns, VDD,
+ 37111.000000ns, VSS,
+ 37471.200000ns, VSS,
+ 37471.300000ns, VDD,
+ 38432.000000ns, VDD,
+ 38432.100000ns, VSS,
+ 38792.300000ns, VSS,
+ 38792.400000ns, VDD,
+ 39032.500000ns, VDD,
+ 39032.600000ns, VSS,
+ 39392.800000ns, VSS,
+ 39392.900000ns, VDD,
+ 39512.900000ns, VDD,
+ 39513.000000ns, VSS,
+ 39633.000000ns, VSS,
+ 39633.100000ns, VDD,
+ 39753.100000ns, VDD,
+ 39753.200000ns, VSS,
+ 40113.400000ns, VSS,
+ 40113.500000ns, VDD,
+ 40954.100000ns, VDD,
+ 40954.200000ns, VSS,
+ 41194.300000ns, VSS,
+ 41194.400000ns, VDD,
+ 41314.400000ns, VDD,
+ 41314.500000ns, VSS,
+ 41794.800000ns, VSS,
+ 41794.900000ns, VDD,
+ 42035.000000ns, VDD,
+ 42035.100000ns, VSS,
+ 42275.200000ns, VSS,
+ 42275.300000ns, VDD,
+ 43236.000000ns, VDD,
+ 43236.100000ns, VSS,
+ 43356.100000ns, VSS,
+ 43356.200000ns, VDD,
+ 43956.600000ns, VDD,
+ 43956.700000ns, VSS,
+ 44196.800000ns, VSS,
+ 44196.900000ns, VDD,
+ 44557.100000ns, VDD,
+ 44557.200000ns, VSS,
+ 44677.200000ns, VSS,
+ 44677.300000ns, VDD,
+ 45037.500000ns, VDD,
+ 45037.600000ns, VSS,
+ 45157.600000ns, VSS,
+ 45157.700000ns, VDD,
+ 45397.800000ns, VDD,
+ 45397.900000ns, VSS,
+ 46718.900000ns, VSS,
+ 46719.000000ns, VDD,
+ 47679.700000ns, VDD,
+ 47679.800000ns, VSS,
+ 48040.000000ns, VSS,
+ 48040.100000ns, VDD,
+ 48400.300000ns, VDD,
+ 48400.400000ns, VSS,
+ 48640.500000ns, VSS,
+ 48640.600000ns, VDD,
+ 50081.700000ns, VDD,
+ 50081.800000ns, VSS,
+ 50442.000000ns, VSS,
+ 50442.100000ns, VDD,
+ 50682.200000ns, VDD,
+ 50682.300000ns, VSS,
+ 51042.500000ns, VSS,
+ 51042.600000ns, VDD,
+ 51402.800000ns, VDD,
+ 51402.900000ns, VSS,
+ 51643.000000ns, VSS,
+ 51643.100000ns, VDD,
+ 51763.100000ns, VDD,
+ 51763.200000ns, VSS,
+ 52123.400000ns, VSS,
+ 52123.500000ns, VDD,
+ 52483.700000ns, VDD,
+ 52483.800000ns, VSS,
+ 52603.800000ns, VSS,
+ 52603.900000ns, VDD,
+ 53564.600000ns, VDD,
+ 53564.700000ns, VSS,
+ 54165.100000ns, VSS,
+ 54165.200000ns, VDD,
+ 54285.200000ns, VDD,
+ 54285.300000ns, VSS,
+ 54525.400000ns, VSS,
+ 54525.500000ns, VDD,
+ 55726.400000ns, VDD,
+ 55726.500000ns, VSS,
+ 55846.500000ns, VSS,
+ 55846.600000ns, VDD,
+ 56567.100000ns, VDD,
+ 56567.200000ns, VSS,
+ 56807.300000ns, VSS,
+ 56807.400000ns, VDD,
+ 57047.500000ns, VDD,
+ 57047.600000ns, VSS,
+ 57287.700000ns, VSS,
+ 57287.800000ns, VDD,
+ 57527.900000ns, VDD,
+ 57528.000000ns, VSS,
+ 57648.000000ns, VSS,
+ 57648.100000ns, VDD,
+ 58008.300000ns, VDD,
+ 58008.400000ns, VSS,
+ 58368.600000ns, VSS,
+ 58368.700000ns, VDD,
+ 58728.900000ns, VDD,
+ 58729.000000ns, VSS,
+ 59209.300000ns, VSS,
+ 59209.400000ns, VDD,
+ 59329.400000ns, VDD,
+ 59329.500000ns, VSS,
+ 59809.800000ns, VSS,
+ 59809.900000ns, VDD,
+ 60290.200000ns, VDD,
+ 60290.300000ns, VSS,
+ 60770.600000ns, VSS,
+ 60770.700000ns, VDD,
+ 61130.900000ns, VDD,
+ 61131.000000ns, VSS,
+ 61491.200000ns, VSS,
+ 61491.300000ns, VDD,
+ 61971.600000ns, VDD,
+ 61971.700000ns, VSS,
+ 62932.400000ns, VSS,
+ 62932.500000ns, VDD,
+ 63052.500000ns, VDD,
+ 63052.600000ns, VSS,
+ 63172.600000ns, VSS,
+ 63172.700000ns, VDD,
+ 63532.900000ns, VDD,
+ 63533.000000ns, VSS,
+ 63893.200000ns, VSS,
+ 63893.300000ns, VDD,
+ 64013.300000ns, VDD,
+ 64013.400000ns, VSS,
+ 64373.600000ns, VSS,
+ 64373.700000ns, VDD,
+ 64733.900000ns, VDD,
+ 64734.000000ns, VSS,
+ 64854.000000ns, VSS,
+ 64854.100000ns, VDD,
+ 65214.300000ns, VDD,
+ 65214.400000ns, VSS,
+ 65334.400000ns, VSS,
+ 65334.500000ns, VDD,
+ 65454.500000ns, VDD,
+ 65454.600000ns, VSS,
+ 65934.900000ns, VSS,
+ 65935.000000ns, VDD,
+ 66295.200000ns, VDD,
+ 66295.300000ns, VSS,
+ 67015.800000ns, VSS,
+ 67015.900000ns, VDD,
+ 68096.700000ns, VDD,
+ 68096.800000ns, VSS,
+ 68216.800000ns, VSS,
+ 68216.900000ns, VDD,
+ 68457.000000ns, VDD,
+ 68457.100000ns, VSS,
+ 69057.500000ns, VSS,
+ 69057.600000ns, VDD,
+ 69537.900000ns, VDD,
+ 69538.000000ns, VSS,
+ 69658.000000ns, VSS,
+ 69658.100000ns, VDD,
+ 69778.100000ns, VDD,
+ 69778.200000ns, VSS,
+ 69898.200000ns, VSS,
+ 69898.300000ns, VDD,
+ 70258.500000ns, VDD,
+ 70258.600000ns, VSS,
+ 70378.600000ns, VSS,
+ 70378.700000ns, VDD,
+ 70498.700000ns, VDD,
+ 70498.800000ns, VSS,
+ 70738.900000ns, VSS,
+ 70739.000000ns, VDD,
+ 71339.400000ns, VDD,
+ 71339.500000ns, VSS,
+ 71819.800000ns, VSS,
+ 71819.900000ns, VDD,
+ 71939.900000ns, VDD,
+ 71940.000000ns, VSS,
+ 72060.000000ns, VSS,
+ 72060.100000ns, VDD,
+ 72420.300000ns, VDD,
+ 72420.400000ns, VSS,
+ 72780.600000ns, VSS,
+ 72780.700000ns, VDD,
+ 73140.900000ns, VDD,
+ 73141.000000ns, VSS,
+ 73501.200000ns, VSS,
+ 73501.300000ns, VDD,
+ 74101.700000ns, VDD,
+ 74101.800000ns, VSS,
+ 74341.900000ns, VSS,
+ 74342.000000ns, VDD,
+ 74582.100000ns, VDD,
+ 74582.200000ns, VSS,
+ 74702.200000ns, VSS,
+ 74702.300000ns, VDD,
+ 74822.300000ns, VDD,
+ 74822.400000ns, VSS,
+ 75182.600000ns, VSS,
+ 75182.700000ns, VDD,
+ 75302.700000ns, VDD,
+ 75302.800000ns, VSS,
+ 75422.800000ns, VSS,
+ 75422.900000ns, VDD,
+ 76023.300000ns, VDD,
+ 76023.400000ns, VSS,
+ 76743.900000ns, VSS,
+ 76744.000000ns, VDD,
+ 77104.200000ns, VDD,
+ 77104.300000ns, VSS,
+ 77944.900000ns, VSS,
+ 77945.000000ns, VDD,
+ 79386.100000ns, VDD,
+ 79386.200000ns, VSS,
+ 80106.700000ns, VSS,
+ 80106.800000ns, VDD,
+ 82388.600000ns, VDD,
+ 82388.700000ns, VSS,
+ 82628.800000ns, VSS,
+ 82628.900000ns, VDD,
+ 82748.900000ns, VDD,
+ 82749.000000ns, VSS,
+ 82869.000000ns, VSS,
+ 82869.100000ns, VDD,
+ 83469.500000ns, VDD,
+ 83469.600000ns, VSS,
+ 83589.600000ns, VSS,
+ 83589.700000ns, VDD,
+ 84190.100000ns, VDD,
+ 84190.200000ns, VSS,
+ 84310.200000ns, VSS,
+ 84310.300000ns, VDD,
+ 84790.600000ns, VDD,
+ 84790.700000ns, VSS,
+ 85391.100000ns, VSS,
+ 85391.200000ns, VDD,
+ 85631.300000ns, VDD,
+ 85631.400000ns, VSS,
+ 85871.500000ns, VSS,
+ 85871.600000ns, VDD,
+ 85991.600000ns, VDD,
+ 85991.700000ns, VSS,
+ 86472.000000ns, VSS,
+ 86472.100000ns, VDD,
+ 87432.800000ns, VDD,
+ 87432.900000ns, VSS,
+ 87673.000000ns, VSS,
+ 87673.100000ns, VDD,
+ 88513.700000ns, VDD,
+ 88513.800000ns, VSS,
+ 88633.800000ns, VSS,
+ 88633.900000ns, VDD,
+ 88994.100000ns, VDD,
+ 88994.200000ns, VSS,
+ 89114.200000ns, VSS,
+ 89114.300000ns, VDD,
+ 89474.500000ns, VDD,
+ 89474.600000ns, VSS,
+ 89834.800000ns, VSS,
+ 89834.900000ns, VDD,
+ 90435.300000ns, VDD,
+ 90435.400000ns, VSS,
+ 90795.600000ns, VSS,
+ 90795.700000ns, VDD,
+ 91756.400000ns, VDD,
+ 91756.500000ns, VSS,
+ 91876.500000ns, VSS,
+ 91876.600000ns, VDD,
+ 92116.700000ns, VDD,
+ 92116.800000ns, VSS,
+ 92236.800000ns, VSS,
+ 92236.900000ns, VDD,
+ 92717.200000ns, VDD,
+ 92717.300000ns, VSS,
+ 92957.400000ns, VSS,
+ 92957.500000ns, VDD,
+ 94518.700000ns, VDD,
+ 94518.800000ns, VSS,
+ 94638.800000ns, VSS,
+ 94638.900000ns, VDD,
+ 94758.900000ns, VDD,
+ 94759.000000ns, VSS,
+ 94879.000000ns, VSS,
+ 94879.100000ns, VDD,
+ 96080.000000ns, VDD,
+ 96080.100000ns, VSS,
+ 96800.600000ns, VSS,
+ 96800.700000ns, VDD,
+ 98842.300000ns, VDD,
+ 98842.400000ns, VSS,
+ 98962.400000ns, VSS,
+ 98962.500000ns, VDD,
+ 99202.600000ns, VDD,
+ 99202.700000ns, VSS,
+ 99322.700000ns, VSS,
+ 99322.800000ns, VDD,
+ 99683.000000ns, VDD,
+ 99683.100000ns, VSS,
+ 99803.100000ns, VSS,
+ 99803.200000ns, VDD,
+ 100643.800000ns, VDD,
+ 100643.900000ns, VSS,
+ 100884.000000ns, VSS,
+ 100884.100000ns, VDD,
+ 101484.500000ns, VDD,
+ 101484.600000ns, VSS,
+ 101604.600000ns, VSS,
+ 101604.700000ns, VDD,
+ 101724.700000ns, VDD,
+ 101724.800000ns, VSS,
+ 101844.800000ns, VSS,
+ 101844.900000ns, VDD,
+ 102085.000000ns, VDD,
+ 102085.100000ns, VSS,
+ 102565.400000ns, VSS,
+ 102565.500000ns, VDD,
+ 103165.900000ns, VDD,
+ 103166.000000ns, VSS,
+ 103286.000000ns, VSS,
+ 103286.100000ns, VDD,
+ 103526.200000ns, VDD,
+ 103526.300000ns, VSS,
+ 104126.700000ns, VSS,
+ 104126.800000ns, VDD,
+ 104246.800000ns, VDD,
+ 104246.900000ns, VSS,
+ 104727.200000ns, VSS,
+ 104727.300000ns, VDD,
+ 104967.400000ns, VDD,
+ 104967.500000ns, VSS,
+ 105567.900000ns, VSS,
+ 105568.000000ns, VDD,
+ 106048.300000ns, VDD,
+ 106048.400000ns, VSS,
+ 106288.500000ns, VSS,
+ 106288.600000ns, VDD,
+ 107129.200000ns, VDD,
+ 107129.300000ns, VSS,
+ 107489.500000ns, VSS,
+ 107489.600000ns, VDD,
+ 107609.600000ns, VDD,
+ 107609.700000ns, VSS,
+ 108210.100000ns, VSS,
+ 108210.200000ns, VDD,
+ 108450.300000ns, VDD,
+ 108450.400000ns, VSS,
+ 108570.400000ns, VSS,
+ 108570.500000ns, VDD,
+ 108690.500000ns, VDD,
+ 108690.600000ns, VSS,
+ 108810.600000ns, VSS,
+ 108810.700000ns, VDD,
+ 108930.700000ns, VDD,
+ 108930.800000ns, VSS,
+ 109050.800000ns, VSS,
+ 109050.900000ns, VDD,
+ 109771.400000ns, VDD,
+ 109771.500000ns, VSS,
+ 110011.600000ns, VSS,
+ 110011.700000ns, VDD,
+ 110371.900000ns, VDD,
+ 110372.000000ns, VSS,
+ 110732.200000ns, VSS,
+ 110732.300000ns, VDD,
+ 111092.500000ns, VDD,
+ 111092.600000ns, VSS,
+ 111933.200000ns, VSS,
+ 111933.300000ns, VDD,
+ 112173.400000ns, VDD,
+ 112173.500000ns, VSS,
+ 112413.600000ns, VSS,
+ 112413.700000ns, VDD,
+ 112773.900000ns, VDD,
+ 112774.000000ns, VSS,
+ 113254.300000ns, VSS,
+ 113254.400000ns, VDD,
+ 113614.600000ns, VDD,
+ 113614.700000ns, VSS,
+ 113854.800000ns, VSS,
+ 113854.900000ns, VDD,
+ 113974.900000ns, VDD,
+ 113975.000000ns, VSS,
+ 114335.200000ns, VSS,
+ 114335.300000ns, VDD,
+ 114455.300000ns, VDD,
+ 114455.400000ns, VSS,
+ 114575.400000ns, VSS,
+ 114575.500000ns, VDD,
+ 114695.500000ns, VDD,
+ 114695.600000ns, VSS,
+ 114815.600000ns, VSS,
+ 114815.700000ns, VDD,
+ 114935.700000ns, VDD,
+ 114935.800000ns, VSS,
+ 115536.200000ns, VSS,
+ 115536.300000ns, VDD,
+ 115776.400000ns, VDD,
+ 115776.500000ns, VSS,
+ 116136.700000ns, VSS,
+ 116136.800000ns, VDD,
+ 116376.900000ns, VDD,
+ 116377.000000ns, VSS,
+ 116737.200000ns, VSS,
+ 116737.300000ns, VDD,
+ 117818.100000ns, VDD,
+ 117818.200000ns, VSS,
+ 118058.300000ns, VSS,
+ 118058.400000ns, VDD,
+ 118538.700000ns, VDD,
+ 118538.800000ns, VSS,
+ 118899.000000ns, VSS,
+ 118899.100000ns, VDD,
+ 119019.100000ns, VDD,
+ 119019.200000ns, VSS,
+ 119379.400000ns, VSS,
+ 119379.500000ns, VDD,
+ 119739.700000ns, VDD,
+ 119739.800000ns, VSS,
+ 120700.500000ns, VSS,
+ 120700.600000ns, VDD,
+ 121060.800000ns, VDD,
+ 121060.900000ns, VSS,
+ 121661.300000ns, VSS,
+ 121661.400000ns, VDD,
+ 122021.600000ns, VDD,
+ 122021.700000ns, VSS,
+ 122502.000000ns, VSS,
+ 122502.100000ns, VDD,
+ 122862.300000ns, VDD,
+ 122862.400000ns, VSS,
+ 122982.400000ns, VSS,
+ 122982.500000ns, VDD,
+ 123703.000000ns, VDD,
+ 123703.100000ns, VSS,
+ 124183.400000ns, VSS,
+ 124183.500000ns, VDD,
+ 124663.800000ns, VDD,
+ 124663.900000ns, VSS,
+ 124783.900000ns, VSS,
+ 124784.000000ns, VDD,
+ 125264.300000ns, VDD,
+ 125264.400000ns, VSS,
+ 125984.900000ns, VSS,
+ 125985.000000ns, VDD,
+ 126105.000000ns, VDD,
+ 126105.100000ns, VSS,
+ 126465.300000ns, VSS,
+ 126465.400000ns, VDD,
+ 127426.100000ns, VDD,
+ 127426.200000ns, VSS,
+ 128026.600000ns, VSS,
+ 128026.700000ns, VDD,
+ 128507.000000ns, VDD,
+ 128507.100000ns, VSS,
+ 129587.900000ns, VSS,
+ 129588.000000ns, VDD,
+ 129948.200000ns, VDD,
+ 129948.300000ns, VSS,
+ 130068.300000ns, VSS,
+ 130068.400000ns, VDD,
+ 130188.400000ns, VDD,
+ 130188.500000ns, VSS,
+ 130308.500000ns, VSS,
+ 130308.600000ns, VDD,
+ 130788.900000ns, VDD,
+ 130789.000000ns, VSS,
+ 130909.000000ns, VSS,
+ 130909.100000ns, VDD,
+ 131029.100000ns, VDD,
+ 131029.200000ns, VSS,
+ 131509.500000ns, VSS,
+ 131509.600000ns, VDD,
+ 132110.000000ns, VDD,
+ 132110.100000ns, VSS,
+ 132230.100000ns, VSS,
+ 132230.200000ns, VDD,
+ 132590.400000ns, VDD,
+ 132590.500000ns, VSS,
+ 132710.500000ns, VSS,
+ 132710.600000ns, VDD,
+ 133190.900000ns, VDD,
+ 133191.000000ns, VSS,
+ 133311.000000ns, VSS,
+ 133311.100000ns, VDD,
+ 133431.100000ns, VDD,
+ 133431.200000ns, VSS,
+ 133911.500000ns, VSS,
+ 133911.600000ns, VDD,
+ 134872.300000ns, VDD,
+ 134872.400000ns, VSS,
+ 135232.600000ns, VSS,
+ 135232.700000ns, VDD,
+ 135352.700000ns, VDD,
+ 135352.800000ns, VSS,
+ 135472.800000ns, VSS,
+ 135472.900000ns, VDD,
+ 136193.400000ns, VDD,
+ 136193.500000ns, VSS,
+ 136313.500000ns, VSS,
+ 136313.600000ns, VDD,
+ 136433.600000ns, VDD,
+ 136433.700000ns, VSS,
+ 136553.700000ns, VSS,
+ 136553.800000ns, VDD,
+ 137154.200000ns, VDD,
+ 137154.300000ns, VSS,
+ 137994.900000ns, VSS,
+ 137995.000000ns, VDD,
+ 138355.200000ns, VDD,
+ 138355.300000ns, VSS,
+ 139195.900000ns, VSS,
+ 139196.000000ns, VDD,
+ 139436.100000ns, VDD,
+ 139436.200000ns, VSS,
+ 139556.200000ns, VSS,
+ 139556.300000ns, VDD,
+ 140276.800000ns, VDD,
+ 140276.900000ns, VSS,
+ 140396.900000ns, VSS,
+ 140397.000000ns, VDD,
+ 140877.300000ns, VDD,
+ 140877.400000ns, VSS,
+ 141117.500000ns, VSS,
+ 141117.600000ns, VDD,
+ 141597.900000ns, VDD,
+ 141598.000000ns, VSS,
+ 141838.100000ns, VSS,
+ 141838.200000ns, VDD,
+ 142078.300000ns, VDD,
+ 142078.400000ns, VSS,
+ 142198.400000ns, VSS,
+ 142198.500000ns, VDD,
+ 142678.800000ns, VDD,
+ 142678.900000ns, VSS,
+ 143039.100000ns, VSS,
+ 143039.200000ns, VDD,
+ 143399.400000ns, VDD,
+ 143399.500000ns, VSS,
+ 143879.800000ns, VSS,
+ 143879.900000ns, VDD,
+ 143999.900000ns, VDD,
+ 144000.000000ns, VSS,
+ 144360.200000ns, VSS,
+ 144360.300000ns, VDD,
+ 144840.600000ns, VDD,
+ 144840.700000ns, VSS,
+ 145080.800000ns, VSS,
+ 145080.900000ns, VDD,
+ 145921.500000ns, VDD,
+ 145921.600000ns, VSS,
+ 146161.700000ns, VSS,
+ 146161.800000ns, VDD,
+ 146762.200000ns, VDD,
+ 146762.300000ns, VSS,
+ 146882.300000ns, VSS,
+ 146882.400000ns, VDD,
+ 147482.800000ns, VDD,
+ 147482.900000ns, VSS,
+ 147843.100000ns, VSS,
+ 147843.200000ns, VDD,
+ 148203.400000ns, VDD,
+ 148203.500000ns, VSS,
+ 148443.600000ns, VSS,
+ 148443.700000ns, VDD,
+ 149764.700000ns, VDD,
+ 149764.800000ns, VSS,
+ 150245.100000ns, VSS,
+ 150245.200000ns, VDD,
+ 150365.200000ns, VDD,
+ 150365.300000ns, VSS,
+ 150485.300000ns, VSS,
+ 150485.400000ns, VDD,
+ 150725.500000ns, VDD,
+ 150725.600000ns, VSS,
+ 150845.600000ns, VSS,
+ 150845.700000ns, VDD,
+ 150965.700000ns, VDD,
+ 150965.800000ns, VSS,
+ 151085.800000ns, VSS,
+ 151085.900000ns, VDD,
+ 152046.600000ns, VDD,
+ 152046.700000ns, VSS,
+ 152406.900000ns, VSS,
+ 152407.000000ns, VDD,
+ 153007.400000ns, VDD,
+ 153007.500000ns, VSS,
+ 153367.700000ns, VSS,
+ 153367.800000ns, VDD,
+ 153728.000000ns, VDD,
+ 153728.100000ns, VSS,
+ 154088.300000ns, VSS,
+ 154088.400000ns, VDD,
+ 154328.500000ns, VDD,
+ 154328.600000ns, VSS,
+ 154448.600000ns, VSS,
+ 154448.700000ns, VDD,
+ 154568.700000ns, VDD,
+ 154568.800000ns, VSS,
+ 155049.100000ns, VSS,
+ 155049.200000ns, VDD,
+ 155529.500000ns, VDD,
+ 155529.600000ns, VSS,
+ 156250.100000ns, VSS,
+ 156250.200000ns, VDD,
+ 157210.900000ns, VDD,
+ 157211.000000ns, VSS,
+ 157451.100000ns, VSS,
+ 157451.200000ns, VDD,
+ 158772.200000ns, VDD,
+ 158772.300000ns, VSS,
+ 158892.300000ns, VSS,
+ 158892.400000ns, VDD,
+ 159372.700000ns, VDD,
+ 159372.800000ns, VSS,
+ 159612.900000ns, VSS,
+ 159613.000000ns, VDD,
+ 160333.500000ns, VDD,
+ 160333.600000ns, VSS,
+ 161294.300000ns, VSS,
+ 161294.400000ns, VDD,
+ 163576.200000ns, VDD,
+ 163576.300000ns, VSS,
+ 163696.300000ns, VSS,
+ 163696.400000ns, VDD,
+ 164416.900000ns, VDD,
+ 164417.000000ns, VSS,
+ 164777.200000ns, VSS,
+ 164777.300000ns, VDD,
+ 165137.500000ns, VDD,
+ 165137.600000ns, VSS,
+ 165257.600000ns, VSS,
+ 165257.700000ns, VDD,
+ 165497.800000ns, VDD,
+ 165497.900000ns, VSS,
+ 165617.900000ns, VSS,
+ 165618.000000ns, VDD,
+ 165978.200000ns, VDD,
+ 165978.300000ns, VSS,
+ 166458.600000ns, VSS,
+ 166458.700000ns, VDD,
+ 166818.900000ns, VDD,
+ 166819.000000ns, VSS,
+ 167659.600000ns, VSS,
+ 167659.700000ns, VDD,
+ 167779.700000ns, VDD,
+ 167779.800000ns, VSS,
+ 167899.800000ns, VSS,
+ 167899.900000ns, VDD,
+ 168380.200000ns, VDD,
+ 168380.300000ns, VSS,
+ 168740.500000ns, VSS,
+ 168740.600000ns, VDD,
+ 168860.600000ns, VDD,
+ 168860.700000ns, VSS,
+ 169220.900000ns, VSS,
+ 169221.000000ns, VDD,
+ 169701.300000ns, VDD,
+ 169701.400000ns, VSS,
+ 169941.500000ns, VSS,
+ 169941.600000ns, VDD,
+ 170061.600000ns, VDD,
+ 170061.700000ns, VSS,
+ 170181.700000ns, VSS,
+ 170181.800000ns, VDD,
+ 170902.300000ns, VDD,
+ 170902.400000ns, VSS,
+ 171262.600000ns, VSS,
+ 171262.700000ns, VDD,
+ 172343.500000ns, VDD,
+ 172343.600000ns, VSS,
+ 172703.800000ns, VSS,
+ 172703.900000ns, VDD,
+ 174865.600000ns, VDD,
+ 174865.700000ns, VSS,
+ 175105.800000ns, VSS,
+ 175105.900000ns, VDD,
+ 175466.100000ns, VDD,
+ 175466.200000ns, VSS,
+ 176066.600000ns, VSS,
+ 176066.700000ns, VDD,
+ 176787.200000ns, VDD,
+ 176787.300000ns, VSS,
+ 177027.400000ns, VSS,
+ 177027.500000ns, VDD,
+ 177147.500000ns, VDD,
+ 177147.600000ns, VSS,
+ 177627.900000ns, VSS,
+ 177628.000000ns, VDD,
+ 178468.600000ns, VDD,
+ 178468.700000ns, VSS,
+ 178828.900000ns, VSS,
+ 178829.000000ns, VDD,
+ 179189.200000ns, VDD,
+ 179189.300000ns, VSS,
+ 179549.500000ns, VSS,
+ 179549.600000ns, VDD,
+ 179909.800000ns, VDD,
+ 179909.900000ns, VSS,
+ 180029.900000ns, VSS,
+ 180030.000000ns, VDD,
+ 180870.600000ns, VDD,
+ 180870.700000ns, VSS,
+ 180990.700000ns, VSS,
+ 180990.800000ns, VDD,
+ 181110.800000ns, VDD,
+ 181110.900000ns, VSS,
+ 181230.900000ns, VSS,
+ 181231.000000ns, VDD,
+ 181591.200000ns, VDD,
+ 181591.300000ns, VSS,
+ 181831.400000ns, VSS,
+ 181831.500000ns, VDD,
+ 181951.500000ns, VDD,
+ 181951.600000ns, VSS,
+ 182311.800000ns, VSS,
+ 182311.900000ns, VDD,
+ 182912.300000ns, VDD,
+ 182912.400000ns, VSS,
+ 183032.400000ns, VSS,
+ 183032.500000ns, VDD,
+ 183753.000000ns, VDD,
+ 183753.100000ns, VSS,
+ 183873.100000ns, VSS,
+ 183873.200000ns, VDD,
+ 185314.300000ns, VDD,
+ 185314.400000ns, VSS,
+ 185674.600000ns, VSS,
+ 185674.700000ns, VDD,
+ 185914.800000ns, VDD,
+ 185914.900000ns, VSS,
+ 186155.000000ns, VSS,
+ 186155.100000ns, VDD,
+ 186995.700000ns, VDD,
+ 186995.800000ns, VSS,
+ 187476.100000ns, VSS,
+ 187476.200000ns, VDD,
+ 187956.500000ns, VDD,
+ 187956.600000ns, VSS,
+ 188076.600000ns, VSS,
+ 188076.700000ns, VDD,
+ 189397.700000ns, VDD,
+ 189397.800000ns, VSS,
+ 189517.800000ns, VSS,
+ 189517.900000ns, VDD,
+ 190238.400000ns, VDD,
+ 190238.500000ns, VSS,
+ 191079.100000ns, VSS,
+ 191079.200000ns, VDD,
+ 191199.200000ns, VDD,
+ 191199.300000ns, VSS,
+ 191319.300000ns, VSS,
+ 191319.400000ns, VDD,
+ 191439.400000ns, VDD,
+ 191439.500000ns, VSS,
+ 191799.700000ns, VSS,
+ 191799.800000ns, VDD,
+ 192160.000000ns, VDD,
+ 192160.100000ns, VSS,
+ 192880.600000ns, VSS,
+ 192880.700000ns, VDD,
+ 193120.800000ns, VDD,
+ 193120.900000ns, VSS,
+ 193481.100000ns, VSS,
+ 193481.200000ns, VDD,
+ 193841.400000ns, VDD,
+ 193841.500000ns, VSS,
+ 194081.600000ns, VSS,
+ 194081.700000ns, VDD,
+ 194562.000000ns, VDD,
+ 194562.100000ns, VSS,
+ 194802.200000ns, VSS,
+ 194802.300000ns, VDD,
+ 195042.400000ns, VDD,
+ 195042.500000ns, VSS,
+ 195162.500000ns, VSS,
+ 195162.600000ns, VDD,
+ 195642.900000ns, VDD,
+ 195643.000000ns, VSS,
+ 195883.100000ns, VSS,
+ 195883.200000ns, VDD,
+ 196243.400000ns, VDD,
+ 196243.500000ns, VSS,
+ 196483.600000ns, VSS,
+ 196483.700000ns, VDD,
+ 197204.200000ns, VDD,
+ 197204.300000ns, VSS,
+ 197324.300000ns, VSS,
+ 197324.400000ns, VDD,
+ 197684.600000ns, VDD,
+ 197684.700000ns, VSS,
+ 197924.800000ns, VSS,
+ 197924.900000ns, VDD,
+ 198525.300000ns, VDD,
+ 198525.400000ns, VSS,
+ 198645.400000ns, VSS,
+ 198645.500000ns, VDD,
+ 198885.600000ns, VDD,
+ 198885.700000ns, VSS,
+ 199366.000000ns, VSS,
+ 199366.100000ns, VDD,
+ 199486.100000ns, VDD,
+ 199486.200000ns, VSS,
+ 199966.500000ns, VSS,
+ 199966.600000ns, VDD,
+ 200687.100000ns, VDD,
+ 200687.200000ns, VSS,
+ 200927.300000ns, VSS,
+ 200927.400000ns, VDD,
+ 202128.300000ns, VDD,
+ 202128.400000ns, VSS,
+ 202368.500000ns, VSS,
+ 202368.600000ns, VDD,
+ 202969.000000ns, VDD,
+ 202969.100000ns, VSS,
+ 203089.100000ns, VSS,
+ 203089.200000ns, VDD,
+ 203209.200000ns, VDD,
+ 203209.300000ns, VSS,
+ 203329.300000ns, VSS,
+ 203329.400000ns, VDD,
+ 204530.300000ns, VDD,
+ 204530.400000ns, VSS,
+ 204890.600000ns, VSS,
+ 204890.700000ns, VDD,
+ 205851.400000ns, VDD,
+ 205851.500000ns, VSS,
+ 205971.500000ns, VSS,
+ 205971.600000ns, VDD,
+ 206331.800000ns, VDD,
+ 206331.900000ns, VSS,
+ 206572.000000ns, VSS,
+ 206572.100000ns, VDD,
+ 206932.300000ns, VDD,
+ 206932.400000ns, VSS,
+ 207292.600000ns, VSS,
+ 207292.700000ns, VDD,
+ 207893.100000ns, VDD,
+ 207893.200000ns, VSS,
+ 208013.200000ns, VSS,
+ 208013.300000ns, VDD,
+ 208253.400000ns, VDD,
+ 208253.500000ns, VSS,
+ 208613.700000ns, VSS,
+ 208613.800000ns, VDD,
+ 209454.400000ns, VDD,
+ 209454.500000ns, VSS,
+ 210655.400000ns, VSS,
+ 210655.500000ns, VDD,
+ 210895.600000ns, VDD,
+ 210895.700000ns, VSS,
+ 211015.700000ns, VSS,
+ 211015.800000ns, VDD,
+ 211135.800000ns, VDD,
+ 211135.900000ns, VSS,
+ 211856.400000ns, VSS,
+ 211856.500000ns, VDD,
+ 213297.600000ns, VDD,
+ 213297.700000ns, VSS,
+ 213657.900000ns, VSS,
+ 213658.000000ns, VDD,
+ 214018.200000ns, VDD,
+ 214018.300000ns, VSS,
+ 214378.500000ns, VSS,
+ 214378.600000ns, VDD,
+ 214738.800000ns, VDD,
+ 214738.900000ns, VSS,
+ 214979.000000ns, VSS,
+ 214979.100000ns, VDD,
+ 216420.200000ns, VDD,
+ 216420.300000ns, VSS,
+ 217140.800000ns, VSS,
+ 217140.900000ns, VDD,
+ 217621.200000ns, VDD,
+ 217621.300000ns, VSS,
+ 217741.300000ns, VSS,
+ 217741.400000ns, VDD,
+ 218101.600000ns, VDD,
+ 218101.700000ns, VSS,
+ 218461.900000ns, VSS,
+ 218462.000000ns, VDD,
+ 218582.000000ns, VDD,
+ 218582.100000ns, VSS,
+ 218702.100000ns, VSS,
+ 218702.200000ns, VDD,
+ 219542.800000ns, VDD,
+ 219542.900000ns, VSS,
+ 220023.200000ns, VSS,
+ 220023.300000ns, VDD,
+ 220383.500000ns, VDD,
+ 220383.600000ns, VSS,
+ 220623.700000ns, VSS,
+ 220623.800000ns, VDD,
+ 221344.300000ns, VDD,
+ 221344.400000ns, VSS,
+ 221704.600000ns, VSS,
+ 221704.700000ns, VDD,
+ 222425.200000ns, VDD,
+ 222425.300000ns, VSS,
+ 222545.300000ns, VSS,
+ 222545.400000ns, VDD,
+ 222665.400000ns, VDD,
+ 222665.500000ns, VSS,
+ 223025.700000ns, VSS,
+ 223025.800000ns, VDD,
+ 223145.800000ns, VDD,
+ 223145.900000ns, VSS,
+ 223506.100000ns, VSS,
+ 223506.200000ns, VDD,
+ 224106.600000ns, VDD,
+ 224106.700000ns, VSS,
+ 224466.900000ns, VSS,
+ 224467.000000ns, VDD,
+ 224707.100000ns, VDD,
+ 224707.200000ns, VSS,
+ 224827.200000ns, VSS,
+ 224827.300000ns, VDD,
+ 225307.600000ns, VDD,
+ 225307.700000ns, VSS,
+ 226028.200000ns, VSS,
+ 226028.300000ns, VDD,
+ 226148.300000ns, VDD,
+ 226148.400000ns, VSS,
+ 226268.400000ns, VSS,
+ 226268.500000ns, VDD,
+ 226628.700000ns, VDD,
+ 226628.800000ns, VSS,
+ 227349.300000ns, VSS,
+ 227349.400000ns, VDD,
+ 227469.400000ns, VDD,
+ 227469.500000ns, VSS,
+ 228310.100000ns, VSS,
+ 228310.200000ns, VDD,
+ 229871.400000ns, VDD,
+ 229871.500000ns, VSS,
+ 229991.500000ns, VSS,
+ 229991.600000ns, VDD,
+ 230471.900000ns, VDD,
+ 230472.000000ns, VSS,
+ 230592.000000ns, VSS,
+ 230592.100000ns, VDD,
+ 230952.300000ns, VDD,
+ 230952.400000ns, VSS,
+ 231312.600000ns, VSS,
+ 231312.700000ns, VDD,
+ 232153.300000ns, VDD,
+ 232153.400000ns, VSS,
+ 232753.800000ns, VSS,
+ 232753.900000ns, VDD,
+ 232873.900000ns, VDD,
+ 232874.000000ns, VSS,
+ 232994.000000ns, VSS,
+ 232994.100000ns, VDD,
+ 233714.600000ns, VDD,
+ 233714.700000ns, VSS,
+ 233834.700000ns, VSS,
+ 233834.800000ns, VDD,
+ 234195.000000ns, VDD,
+ 234195.100000ns, VSS,
+ 234555.300000ns, VSS,
+ 234555.400000ns, VDD,
+ 234795.500000ns, VDD,
+ 234795.600000ns, VSS,
+ 234915.600000ns, VSS,
+ 234915.700000ns, VDD,
+ 235155.800000ns, VDD,
+ 235155.900000ns, VSS,
+ 235636.200000ns, VSS,
+ 235636.300000ns, VDD,
+ 236116.600000ns, VDD,
+ 236116.700000ns, VSS,
+ 236597.000000ns, VSS,
+ 236597.100000ns, VDD,
+ 236957.300000ns, VDD,
+ 236957.400000ns, VSS,
+ 237077.400000ns, VSS,
+ 237077.500000ns, VDD,
+ 237197.500000ns, VDD,
+ 237197.600000ns, VSS,
+ 237437.700000ns, VSS,
+ 237437.800000ns, VDD,
+ 237798.000000ns, VDD,
+ 237798.100000ns, VSS,
+ 237918.100000ns, VSS,
+ 237918.200000ns, VDD,
+ 238038.200000ns, VDD,
+ 238038.300000ns, VSS,
+ 238278.400000ns, VSS,
+ 238278.500000ns, VDD,
+ 238398.500000ns, VDD,
+ 238398.600000ns, VSS,
+ 238999.000000ns, VSS,
+ 238999.100000ns, VDD,
+ 239479.400000ns, VDD,
+ 239479.500000ns, VSS,
+ 240320.100000ns, VSS,
+ 240320.200000ns, VDD,
+ 240920.600000ns, VDD,
+ 240920.700000ns, VSS,
+ 241160.800000ns, VSS,
+ 241160.900000ns, VDD,
+ 241280.900000ns, VDD,
+ 241281.000000ns, VSS,
+ 241761.300000ns, VSS,
+ 241761.400000ns, VDD,
+ 242001.500000ns, VDD,
+ 242001.600000ns, VSS,
+ 242241.700000ns, VSS,
+ 242241.800000ns, VDD,
+ 242722.100000ns, VDD,
+ 242722.200000ns, VSS,
+ 242842.200000ns, VSS,
+ 242842.300000ns, VDD,
+ 242962.300000ns, VDD,
+ 242962.400000ns, VSS,
+ 243082.400000ns, VSS,
+ 243082.500000ns, VDD,
+ 244163.300000ns, VDD,
+ 244163.400000ns, VSS,
+ 244283.400000ns, VSS,
+ 244283.500000ns, VDD,
+ 244883.900000ns, VDD,
+ 244884.000000ns, VSS,
+ 245004.000000ns, VSS,
+ 245004.100000ns, VDD,
+ 245964.800000ns, VDD,
+ 245964.900000ns, VSS,
+ 246685.400000ns, VSS,
+ 246685.500000ns, VDD,
+ 247285.900000ns, VDD,
+ 247286.000000ns, VSS,
+ 247406.000000ns, VSS,
+ 247406.100000ns, VDD,
+ 249567.800000ns, VDD,
+ 249567.900000ns, VSS,
+ 249687.900000ns, VSS,
+ 249688.000000ns, VDD,
+ 250048.200000ns, VDD,
+ 250048.300000ns, VSS,
+ 250168.300000ns, VSS,
+ 250168.400000ns, VDD,
+ 250408.500000ns, VDD,
+ 250408.600000ns, VSS,
+ 250768.800000ns, VSS,
+ 250768.900000ns, VDD,
+ 253170.800000ns, VDD,
+ 253170.900000ns, VSS,
+ 253411.000000ns, VSS,
+ 253411.100000ns, VDD,
+ 253891.400000ns, VDD,
+ 253891.500000ns, VSS,
+ 254011.500000ns, VSS,
+ 254011.600000ns, VDD,
+ 254131.600000ns, VDD,
+ 254131.700000ns, VSS,
+ 254491.900000ns, VSS,
+ 254492.000000ns, VDD,
+ 254612.000000ns, VDD,
+ 254612.100000ns, VSS,
+ 254732.100000ns, VSS,
+ 254732.200000ns, VDD,
+ 255452.700000ns, VDD,
+ 255452.800000ns, VSS,
+ 256053.200000ns, VSS,
+ 256053.300000ns, VDD,
+ 256413.500000ns, VDD,
+ 256413.600000ns, VSS,
+ 256653.700000ns, VSS,
+ 256653.800000ns, VDD,
+ 257734.600000ns, VDD,
+ 257734.700000ns, VSS,
+ 257854.700000ns, VSS,
+ 257854.800000ns, VDD,
+ 257974.800000ns, VDD,
+ 257974.900000ns, VSS,
+ 258094.900000ns, VSS,
+ 258095.000000ns, VDD,
+ 258455.200000ns, VDD,
+ 258455.300000ns, VSS,
+ 258575.300000ns, VSS,
+ 258575.400000ns, VDD,
+ 259896.400000ns, VDD,
+ 259896.500000ns, VSS,
+ 260016.500000ns, VSS,
+ 260016.600000ns, VDD,
+ 260496.900000ns, VDD,
+ 260497.000000ns, VSS,
+ 261217.500000ns, VSS,
+ 261217.600000ns, VDD,
+ 261457.700000ns, VDD,
+ 261457.800000ns, VSS,
+ 261577.800000ns, VSS,
+ 261577.900000ns, VDD,
+ 261938.100000ns, VDD,
+ 261938.200000ns, VSS,
+ 262178.300000ns, VSS,
+ 262178.400000ns, VDD,
+ 262658.700000ns, VDD,
+ 262658.800000ns, VSS,
+ 263139.100000ns, VSS,
+ 263139.200000ns, VDD,
+ 263379.300000ns, VDD,
+ 263379.400000ns, VSS,
+ 264220.000000ns, VSS,
+ 264220.100000ns, VDD,
+ 264460.200000ns, VDD,
+ 264460.300000ns, VSS,
+ 264580.300000ns, VSS,
+ 264580.400000ns, VDD,
+ 264700.400000ns, VDD,
+ 264700.500000ns, VSS,
+ 264940.600000ns, VSS,
+ 264940.700000ns, VDD,
+ 265781.300000ns, VDD,
+ 265781.400000ns, VSS,
+ 265901.400000ns, VSS,
+ 265901.500000ns, VDD,
+ 266261.700000ns, VDD,
+ 266261.800000ns, VSS,
+ 266381.800000ns, VSS,
+ 266381.900000ns, VDD,
+ 266742.100000ns, VDD,
+ 266742.200000ns, VSS,
+ 266862.200000ns, VSS,
+ 266862.300000ns, VDD,
+ 267102.400000ns, VDD,
+ 267102.500000ns, VSS,
+ 267342.600000ns, VSS,
+ 267342.700000ns, VDD,
+ 268063.200000ns, VDD,
+ 268063.300000ns, VSS,
+ 268183.300000ns, VSS,
+ 268183.400000ns, VDD,
+ 268783.800000ns, VDD,
+ 268783.900000ns, VSS,
+ 269384.300000ns, VSS,
+ 269384.400000ns, VDD,
+ 270104.900000ns, VDD,
+ 270105.000000ns, VSS,
+ 270345.100000ns, VSS,
+ 270345.200000ns, VDD,
+ 270705.400000ns, VDD,
+ 270705.500000ns, VSS,
+ 271305.900000ns, VSS,
+ 271306.000000ns, VDD,
+ 272026.500000ns, VDD,
+ 272026.600000ns, VSS,
+ 272386.800000ns, VSS,
+ 272386.900000ns, VDD,
+ 272747.100000ns, VDD,
+ 272747.200000ns, VSS,
+ 273107.400000ns, VSS,
+ 273107.500000ns, VDD,
+ 273828.000000ns, VDD,
+ 273828.100000ns, VSS,
+ 274308.400000ns, VSS,
+ 274308.500000ns, VDD,
+ 274548.600000ns, VDD,
+ 274548.700000ns, VSS,
+ 275029.000000ns, VSS,
+ 275029.100000ns, VDD,
+ 275989.800000ns, VDD,
+ 275989.900000ns, VSS,
+ 276830.500000ns, VSS,
+ 276830.600000ns, VDD,
+ 277551.100000ns, VDD,
+ 277551.200000ns, VSS,
+ 277911.400000ns, VSS,
+ 277911.500000ns, VDD,
+ 278031.500000ns, VDD,
+ 278031.600000ns, VSS,
+ 278752.100000ns, VSS,
+ 278752.200000ns, VDD,
+ 280553.600000ns, VDD,
+ 280553.700000ns, VSS,
+ 280673.700000ns, VSS,
+ 280673.800000ns, VDD,
+ 281394.300000ns, VDD,
+ 281394.400000ns, VSS,
+ 281994.800000ns, VSS,
+ 281994.900000ns, VDD,
+ 282595.300000ns, VDD,
+ 282595.400000ns, VSS,
+ 282715.400000ns, VSS,
+ 282715.500000ns, VDD,
+ 282955.600000ns, VDD,
+ 282955.700000ns, VSS,
+ 283075.700000ns, VSS,
+ 283075.800000ns, VDD,
+ 283195.800000ns, VDD,
+ 283195.900000ns, VSS,
+ 283916.400000ns, VSS,
+ 283916.500000ns, VDD,
+ 284156.600000ns, VDD,
+ 284156.700000ns, VSS,
+ 284276.700000ns, VSS,
+ 284276.800000ns, VDD,
+ 284396.800000ns, VDD,
+ 284396.900000ns, VSS,
+ 284516.900000ns, VSS,
+ 284517.000000ns, VDD,
+ 284877.200000ns, VDD,
+ 284877.300000ns, VSS,
+ 285117.400000ns, VSS,
+ 285117.500000ns, VDD,
+ 285717.900000ns, VDD,
+ 285718.000000ns, VSS,
+ 285958.100000ns, VSS,
+ 285958.200000ns, VDD,
+ 286678.700000ns, VDD,
+ 286678.800000ns, VSS,
+ 286918.900000ns, VSS,
+ 286919.000000ns, VDD,
+ 287279.200000ns, VDD,
+ 287279.300000ns, VSS,
+ 287639.500000ns, VSS,
+ 287639.600000ns, VDD,
+ 287999.800000ns, VDD,
+ 287999.900000ns, VSS,
+ 288600.300000ns, VSS,
+ 288600.400000ns, VDD,
+ 288840.500000ns, VDD,
+ 288840.600000ns, VSS,
+ 288960.600000ns, VSS,
+ 288960.700000ns, VDD,
+ 290521.900000ns, VDD,
+ 290522.000000ns, VSS,
+ 290762.100000ns, VSS,
+ 290762.200000ns, VDD,
+ 291002.300000ns, VDD,
+ 291002.400000ns, VSS,
+ 291242.500000ns, VSS,
+ 291242.600000ns, VDD,
+ 291963.100000ns, VDD,
+ 291963.200000ns, VSS,
+ 292083.200000ns, VSS,
+ 292083.300000ns, VDD,
+ 292443.500000ns, VDD,
+ 292443.600000ns, VSS,
+ 292563.600000ns, VSS,
+ 292563.700000ns, VDD,
+ 293644.500000ns, VDD,
+ 293644.600000ns, VSS,
+ 294245.000000ns, VSS,
+ 294245.100000ns, VDD,
+ 294605.300000ns, VDD,
+ 294605.400000ns, VSS,
+ 294725.400000ns, VSS,
+ 294725.500000ns, VDD,
+ 294965.600000ns, VDD,
+ 294965.700000ns, VSS,
+ 295325.900000ns, VSS,
+ 295326.000000ns, VDD,
+ 295566.100000ns, VDD,
+ 295566.200000ns, VSS,
+ 295686.200000ns, VSS,
+ 295686.300000ns, VDD,
+ 296286.700000ns, VDD,
+ 296286.800000ns, VSS,
+ 296406.800000ns, VSS,
+ 296406.900000ns, VDD,
+ 296767.100000ns, VDD,
+ 296767.200000ns, VSS,
+ 296887.200000ns, VSS,
+ 296887.300000ns, VDD,
+ 297007.300000ns, VDD,
+ 297007.400000ns, VSS,
+ 297127.400000ns, VSS,
+ 297127.500000ns, VDD,
+ 297487.700000ns, VDD,
+ 297487.800000ns, VSS,
+ 298088.200000ns, VSS,
+ 298088.300000ns, VDD,
+ 298208.300000ns, VDD,
+ 298208.400000ns, VSS,
+ 298328.400000ns, VSS,
+ 298328.500000ns, VDD,
+ 298568.600000ns, VDD,
+ 298568.700000ns, VSS,
+ 299169.100000ns, VSS,
+ 299169.200000ns, VDD,
+ 300129.900000ns, VDD,
+ 300130.000000ns, VSS,
+ 300250.000000ns, VSS,
+ 300250.100000ns, VDD,
+ 300490.200000ns, VDD,
+ 300490.300000ns, VSS,
+ 300610.300000ns, VSS,
+ 300610.400000ns, VDD,
+ 301451.000000ns, VDD,
+ 301451.100000ns, VSS,
+ 301691.200000ns, VSS,
+ 301691.300000ns, VDD,
+ 301931.400000ns, VDD,
+ 301931.500000ns, VSS,
+ 302051.500000ns, VSS,
+ 302051.600000ns, VDD,
+ 302411.800000ns, VDD,
+ 302411.900000ns, VSS,
+ 302531.900000ns, VSS,
+ 302532.000000ns, VDD,
+ 303012.300000ns, VDD,
+ 303012.400000ns, VSS,
+ 303492.700000ns, VSS,
+ 303492.800000ns, VDD,
+ 303612.800000ns, VDD,
+ 303612.900000ns, VSS,
+ 303973.100000ns, VSS,
+ 303973.200000ns, VDD,
+ 304213.300000ns, VDD,
+ 304213.400000ns, VSS,
+ 304333.400000ns, VSS,
+ 304333.500000ns, VDD,
+ 304933.900000ns, VDD,
+ 304934.000000ns, VSS,
+ 305054.000000ns, VSS,
+ 305054.100000ns, VDD,
+ 305894.700000ns, VDD,
+ 305894.800000ns, VSS,
+ 306014.800000ns, VSS,
+ 306014.900000ns, VDD,
+ 306375.100000ns, VDD,
+ 306375.200000ns, VSS,
+ 306495.200000ns, VSS,
+ 306495.300000ns, VDD,
+ 307215.800000ns, VDD,
+ 307215.900000ns, VSS,
+ 307696.200000ns, VSS,
+ 307696.300000ns, VDD,
+ 308777.100000ns, VDD,
+ 308777.200000ns, VSS,
+ 309017.300000ns, VSS,
+ 309017.400000ns, VDD,
+ 309377.600000ns, VDD,
+ 309377.700000ns, VSS,
+ 309617.800000ns, VSS,
+ 309617.900000ns, VDD,
+ 309858.000000ns, VDD,
+ 309858.100000ns, VSS,
+ 310458.500000ns, VSS,
+ 310458.600000ns, VDD,
+ 310818.800000ns, VDD,
+ 310818.900000ns, VSS,
+ 311059.000000ns, VSS,
+ 311059.100000ns, VDD,
+ 311419.300000ns, VDD,
+ 311419.400000ns, VSS,
+ 311659.500000ns, VSS,
+ 311659.600000ns, VDD,
+ 312019.800000ns, VDD,
+ 312019.900000ns, VSS,
+ 312500.200000ns, VSS,
+ 312500.300000ns, VDD,
+ 312620.300000ns, VDD,
+ 312620.400000ns, VSS,
+ 312740.400000ns, VSS,
+ 312740.500000ns, VDD,
+ 312860.500000ns, VDD,
+ 312860.600000ns, VSS,
+ 313100.700000ns, VSS,
+ 313100.800000ns, VDD,
+ 313581.100000ns, VDD,
+ 313581.200000ns, VSS,
+ 314301.700000ns, VSS,
+ 314301.800000ns, VDD,
+ 314541.900000ns, VDD,
+ 314542.000000ns, VSS,
+ 314662.000000ns, VSS,
+ 314662.100000ns, VDD,
+ 315022.300000ns, VDD,
+ 315022.400000ns, VSS,
+ 315142.400000ns, VSS,
+ 315142.500000ns, VDD,
+ 315262.500000ns, VDD,
+ 315262.600000ns, VSS,
+ 315983.100000ns, VSS,
+ 315983.200000ns, VDD,
+ 316223.300000ns, VDD,
+ 316223.400000ns, VSS,
+ 316343.400000ns, VSS,
+ 316343.500000ns, VDD,
+ 316583.600000ns, VDD,
+ 316583.700000ns, VSS,
+ 318024.800000ns, VSS,
+ 318024.900000ns, VDD,
+ 318265.000000ns, VDD,
+ 318265.100000ns, VSS,
+ 318625.300000ns, VSS,
+ 318625.400000ns, VDD,
+ 319105.700000ns, VDD,
+ 319105.800000ns, VSS,
+ 319946.400000ns, VSS,
+ 319946.500000ns, VDD,
+ 320066.500000ns, VDD,
+ 320066.600000ns, VSS,
+ 320306.700000ns, VSS,
+ 320306.800000ns, VDD,
+ 320667.000000ns, VDD,
+ 320667.100000ns, VSS,
+ 321147.400000ns, VSS,
+ 321147.500000ns, VDD,
+ 321267.500000ns, VDD,
+ 321267.600000ns, VSS,
+ 321627.800000ns, VSS,
+ 321627.900000ns, VDD,
+ 321988.100000ns, VDD,
+ 321988.200000ns, VSS,
+ 322108.200000ns, VSS,
+ 322108.300000ns, VDD,
+ 322348.400000ns, VDD,
+ 322348.500000ns, VSS,
+ 322468.500000ns, VSS,
+ 322468.600000ns, VDD,
+ 323309.200000ns, VDD,
+ 323309.300000ns, VSS,
+ 323429.300000ns, VSS,
+ 323429.400000ns, VDD,
+ 323909.700000ns, VDD,
+ 323909.800000ns, VSS,
+ 325230.800000ns, VSS,
+ 325230.900000ns, VDD,
+ 325591.100000ns, VDD,
+ 325591.200000ns, VSS,
+ 325831.300000ns, VSS,
+ 325831.400000ns, VDD,
+ 325951.400000ns, VDD,
+ 325951.500000ns, VSS,
+ 326551.900000ns, VSS,
+ 326552.000000ns, VDD,
+ 326792.100000ns, VDD,
+ 326792.200000ns, VSS,
+ 327152.400000ns, VSS,
+ 327152.500000ns, VDD,
+ 327272.500000ns, VDD,
+ 327272.600000ns, VSS,
+ 327752.900000ns, VSS,
+ 327753.000000ns, VDD,
+ 328233.300000ns, VDD,
+ 328233.400000ns, VSS,
+ 328713.700000ns, VSS,
+ 328713.800000ns, VDD,
+ 329434.300000ns, VDD,
+ 329434.400000ns, VSS,
+ 329794.600000ns, VSS,
+ 329794.700000ns, VDD,
+ 331235.800000ns, VDD,
+ 331235.900000ns, VSS,
+ 331596.100000ns, VSS,
+ 331596.200000ns, VDD,
+ 331836.300000ns, VDD,
+ 331836.400000ns, VSS,
+ 332316.700000ns, VSS,
+ 332316.800000ns, VDD,
+ 332917.200000ns, VDD,
+ 332917.300000ns, VSS,
+ 333277.500000ns, VSS,
+ 333277.600000ns, VDD,
+ 333397.600000ns, VDD,
+ 333397.700000ns, VSS,
+ 333517.700000ns, VSS,
+ 333517.800000ns, VDD,
+ 334598.600000ns, VDD,
+ 334598.700000ns, VSS,
+ 334718.700000ns, VSS,
+ 334718.800000ns, VDD,
+ 335079.000000ns, VDD,
+ 335079.100000ns, VSS,
+ 335199.100000ns, VSS,
+ 335199.200000ns, VDD,
+ 335679.500000ns, VDD,
+ 335679.600000ns, VSS,
+ 335919.700000ns, VSS,
+ 335919.800000ns, VDD,
+ 336640.300000ns, VDD,
+ 336640.400000ns, VSS,
+ 337000.600000ns, VSS,
+ 337000.700000ns, VDD,
+ 337721.200000ns, VDD,
+ 337721.300000ns, VSS,
+ 338201.600000ns, VSS,
+ 338201.700000ns, VDD,
+ 338922.200000ns, VDD,
+ 338922.300000ns, VSS,
+ 339042.300000ns, VSS,
+ 339042.400000ns, VDD,
+ 339522.700000ns, VDD,
+ 339522.800000ns, VSS,
+ 339762.900000ns, VSS,
+ 339763.000000ns, VDD,
+ 340123.200000ns, VDD,
+ 340123.300000ns, VSS,
+ 340483.500000ns, VSS,
+ 340483.600000ns, VDD,
+ 340723.700000ns, VDD,
+ 340723.800000ns, VSS,
+ 340843.800000ns, VSS,
+ 340843.900000ns, VDD,
+ 341564.400000ns, VDD,
+ 341564.500000ns, VSS,
+ 342285.000000ns, VSS,
+ 342285.100000ns, VDD,
+ 343005.600000ns, VDD,
+ 343005.700000ns, VSS,
+ 343245.800000ns, VSS,
+ 343245.900000ns, VDD,
+ 343486.000000ns, VDD,
+ 343486.100000ns, VSS,
+ 343606.100000ns, VSS,
+ 343606.200000ns, VDD,
+ 343726.200000ns, VDD,
+ 343726.300000ns, VSS,
+ 343846.300000ns, VSS,
+ 343846.400000ns, VDD,
+ 344086.500000ns, VDD,
+ 344086.600000ns, VSS,
+ 344687.000000ns, VSS,
+ 344687.100000ns, VDD,
+ 345047.300000ns, VDD,
+ 345047.400000ns, VSS,
+ 345407.600000ns, VSS,
+ 345407.700000ns, VDD,
+ 346128.200000ns, VDD,
+ 346128.300000ns, VSS,
+ 346368.400000ns, VSS,
+ 346368.500000ns, VDD,
+ 346608.600000ns, VDD,
+ 346608.700000ns, VSS,
+ 347089.000000ns, VSS,
+ 347089.100000ns, VDD,
+ 347569.400000ns, VDD,
+ 347569.500000ns, VSS,
+ 347929.700000ns, VSS,
+ 347929.800000ns, VDD,
+ 348169.900000ns, VDD,
+ 348170.000000ns, VSS,
+ 348290.000000ns, VSS,
+ 348290.100000ns, VDD,
+ 348530.200000ns, VDD,
+ 348530.300000ns, VSS,
+ 349130.700000ns, VSS,
+ 349130.800000ns, VDD,
+ 349611.100000ns, VDD,
+ 349611.200000ns, VSS,
+ 349851.300000ns, VSS,
+ 349851.400000ns, VDD,
+ 350211.600000ns, VDD,
+ 350211.700000ns, VSS,
+ 350331.700000ns, VSS,
+ 350331.800000ns, VDD,
+ 350692.000000ns, VDD,
+ 350692.100000ns, VSS,
+ 351172.400000ns, VSS,
+ 351172.500000ns, VDD,
+ 351532.700000ns, VDD,
+ 351532.800000ns, VSS,
+ 352013.100000ns, VSS,
+ 352013.200000ns, VDD,
+ 352253.300000ns, VDD,
+ 352253.400000ns, VSS,
+ 352373.400000ns, VSS,
+ 352373.500000ns, VDD,
+ 352853.800000ns, VDD,
+ 352853.900000ns, VSS,
+ 353214.100000ns, VSS,
+ 353214.200000ns, VDD,
+ 353934.700000ns, VDD,
+ 353934.800000ns, VSS,
+ 354054.800000ns, VSS,
+ 354054.900000ns, VDD,
+ 354415.100000ns, VDD,
+ 354415.200000ns, VSS,
+ 354895.500000ns, VSS,
+ 354895.600000ns, VDD,
+ 355255.800000ns, VDD,
+ 355255.900000ns, VSS,
+ 355856.300000ns, VSS,
+ 355856.400000ns, VDD,
+ 356937.200000ns, VDD,
+ 356937.300000ns, VSS,
+ 357057.300000ns, VSS,
+ 357057.400000ns, VDD,
+ 358618.600000ns, VDD,
+ 358618.700000ns, VSS,
+ 358738.700000ns, VSS,
+ 358738.800000ns, VDD,
+ 358858.800000ns, VDD,
+ 358858.900000ns, VSS,
+ 359579.400000ns, VSS,
+ 359579.500000ns, VDD,
+ 359819.600000ns, VDD,
+ 359819.700000ns, VSS,
+ 359939.700000ns, VSS,
+ 359939.800000ns, VDD,
+ 360780.400000ns, VDD,
+ 360780.500000ns, VSS,
+ 361020.600000ns, VSS,
+ 361020.700000ns, VDD,
+ 361861.300000ns, VDD,
+ 361861.400000ns, VSS,
+ 362341.700000ns, VSS,
+ 362341.800000ns, VDD,
+ 362581.900000ns, VDD,
+ 362582.000000ns, VSS,
+ 362702.000000ns, VSS,
+ 362702.100000ns, VDD,
+ 362822.100000ns, VDD,
+ 362822.200000ns, VSS,
+ 363062.300000ns, VSS,
+ 363062.400000ns, VDD,
+ 363422.600000ns, VDD,
+ 363422.700000ns, VSS,
+ 363662.800000ns, VSS,
+ 363662.900000ns, VDD,
+ 363782.900000ns, VDD,
+ 363783.000000ns, VSS,
+ 363903.000000ns, VSS,
+ 363903.100000ns, VDD,
+ 364503.500000ns, VDD,
+ 364503.600000ns, VSS,
+ 364743.700000ns, VSS,
+ 364743.800000ns, VDD,
+ 365944.700000ns, VDD,
+ 365944.800000ns, VSS,
+ 366064.800000ns, VSS,
+ 366064.900000ns, VDD,
+ 366425.100000ns, VDD,
+ 366425.200000ns, VSS,
+ 366545.200000ns, VSS,
+ 366545.300000ns, VDD,
+ 366785.400000ns, VDD,
+ 366785.500000ns, VSS,
+ 367506.000000ns, VSS,
+ 367506.100000ns, VDD,
+ 367626.100000ns, VDD,
+ 367626.200000ns, VSS,
+ 368586.900000ns, VSS,
+ 368587.000000ns, VDD,
+ 368947.200000ns, VDD,
+ 368947.300000ns, VSS,
+ 369067.300000ns, VSS,
+ 369067.400000ns, VDD,
+ 369667.800000ns, VDD,
+ 369667.900000ns, VSS,
+ 369908.000000ns, VSS,
+ 369908.100000ns, VDD,
+ 370268.300000ns, VDD,
+ 370268.400000ns, VSS,
+ 370508.500000ns, VSS,
+ 370508.600000ns, VDD,
+ 370868.800000ns, VDD,
+ 370868.900000ns, VSS,
+ 370988.900000ns, VSS,
+ 370989.000000ns, VDD,
+ 371229.100000ns, VDD,
+ 371229.200000ns, VSS,
+ 371949.700000ns, VSS,
+ 371949.800000ns, VDD,
+ 372189.900000ns, VDD,
+ 372190.000000ns, VSS,
+ 372550.200000ns, VSS,
+ 372550.300000ns, VDD,
+ 373150.700000ns, VDD,
+ 373150.800000ns, VSS,
+ 373511.000000ns, VSS,
+ 373511.100000ns, VDD,
+ 374111.500000ns, VDD,
+ 374111.600000ns, VSS,
+ 374351.700000ns, VSS,
+ 374351.800000ns, VDD,
+ 374952.200000ns, VDD,
+ 374952.300000ns, VSS,
+ 375432.600000ns, VSS,
+ 375432.700000ns, VDD,
+ 375792.900000ns, VDD,
+ 375793.000000ns, VSS,
+ 376033.100000ns, VSS,
+ 376033.200000ns, VDD,
+ 376993.900000ns, VDD,
+ 376994.000000ns, VSS,
+ 377234.100000ns, VSS,
+ 377234.200000ns, VDD,
+ 377594.400000ns, VDD,
+ 377594.500000ns, VSS,
+ 377834.600000ns, VSS,
+ 377834.700000ns, VDD,
+ 377954.700000ns, VDD,
+ 377954.800000ns, VSS,
+ 378435.100000ns, VSS,
+ 378435.200000ns, VDD,
+ 379155.700000ns, VDD,
+ 379155.800000ns, VSS,
+ 379636.100000ns, VSS,
+ 379636.200000ns, VDD,
+ 379996.400000ns, VDD,
+ 379996.500000ns, VSS,
+ 380356.700000ns, VSS,
+ 380356.800000ns, VDD,
+ 380717.000000ns, VDD,
+ 380717.100000ns, VSS,
+ 380957.200000ns, VSS,
+ 380957.300000ns, VDD,
+ 382278.300000ns, VDD,
+ 382278.400000ns, VSS,
+ 382398.400000ns, VSS,
+ 382398.500000ns, VDD,
+ 384320.000000ns, VDD,
+ 384320.100000ns, VSS,
+ 384560.200000ns, VSS,
+ 384560.300000ns, VDD,
+ 384680.300000ns, VDD,
+ 384680.400000ns, VSS,
+ 385160.700000ns, VSS,
+ 385160.800000ns, VDD,
+ 385280.800000ns, VDD,
+ 385280.900000ns, VSS,
+ 385881.300000ns, VSS,
+ 385881.400000ns, VDD,
+ 387082.300000ns, VDD,
+ 387082.400000ns, VSS,
+ 387562.700000ns, VSS,
+ 387562.800000ns, VDD,
+ 388283.300000ns, VDD,
+ 388283.400000ns, VSS,
+ 388523.500000ns, VSS,
+ 388523.600000ns, VDD,
+ 388883.800000ns, VDD,
+ 388883.900000ns, VSS,
+ 389364.200000ns, VSS,
+ 389364.300000ns, VDD,
+ 389604.400000ns, VDD,
+ 389604.500000ns, VSS,
+ 389964.700000ns, VSS,
+ 389964.800000ns, VDD,
+ 390325.000000ns, VDD,
+ 390325.100000ns, VSS,
+ 390445.100000ns, VSS,
+ 390445.200000ns, VDD,
+ 391045.600000ns, VDD,
+ 391045.700000ns, VSS,
+ 391646.100000ns, VSS,
+ 391646.200000ns, VDD,
+ 392006.400000ns, VDD,
+ 392006.500000ns, VSS,
+ 392246.600000ns, VSS,
+ 392246.700000ns, VDD,
+ 392847.100000ns, VDD,
+ 392847.200000ns, VSS,
+ 392967.200000ns, VSS,
+ 392967.300000ns, VDD,
+ 393207.400000ns, VDD,
+ 393207.500000ns, VSS,
+ 393327.500000ns, VSS,
+ 393327.600000ns, VDD,
+ 393447.600000ns, VDD,
+ 393447.700000ns, VSS,
+ 393567.700000ns, VSS,
+ 393567.800000ns, VDD,
+ 393687.800000ns, VDD,
+ 393687.900000ns, VSS,
+ 394048.100000ns, VSS,
+ 394048.200000ns, VDD,
+ 394408.400000ns, VDD,
+ 394408.500000ns, VSS,
+ 394528.500000ns, VSS,
+ 394528.600000ns, VDD,
+ 395729.500000ns, VDD,
+ 395729.600000ns, VSS,
+ 395969.700000ns, VSS,
+ 395969.800000ns, VDD,
+ 397050.600000ns, VDD,
+ 397050.700000ns, VSS,
+ 397290.800000ns, VSS,
+ 397290.900000ns, VDD,
+ 397771.200000ns, VDD,
+ 397771.300000ns, VSS,
+ 398131.500000ns, VSS,
+ 398131.600000ns, VDD,
+ 398251.600000ns, VDD,
+ 398251.700000ns, VSS,
+ 398491.800000ns, VSS,
+ 398491.900000ns, VDD,
+ 399933.000000ns, VDD,
+ 399933.100000ns, VSS,
+ 400293.300000ns, VSS,
+ 400293.400000ns, VDD,
+ 400773.700000ns, VDD,
+ 400773.800000ns, VSS,
+ 400893.800000ns, VSS,
+ 400893.900000ns, VDD,
+ 401013.900000ns, VDD,
+ 401014.000000ns, VSS,
+ 401254.100000ns, VSS,
+ 401254.200000ns, VDD,
+ 401494.300000ns, VDD,
+ 401494.400000ns, VSS,
+ 401734.500000ns, VSS,
+ 401734.600000ns, VDD,
+ 401854.600000ns, VDD,
+ 401854.700000ns, VSS,
+ 402094.800000ns, VSS,
+ 402094.900000ns, VDD,
+ 402455.100000ns, VDD,
+ 402455.200000ns, VSS,
+ 402575.200000ns, VSS,
+ 402575.300000ns, VDD,
+ 403295.800000ns, VDD,
+ 403295.900000ns, VSS,
+ 403415.900000ns, VSS,
+ 403416.000000ns, VDD,
+ 403776.200000ns, VDD,
+ 403776.300000ns, VSS,
+ 404136.500000ns, VSS,
+ 404136.600000ns, VDD,
+ 404496.800000ns, VDD,
+ 404496.900000ns, VSS,
+ 404737.000000ns, VSS,
+ 404737.100000ns, VDD,
+ 405577.700000ns, VDD,
+ 405577.800000ns, VSS,
+ 405697.800000ns, VSS,
+ 405697.900000ns, VDD,
+ 406418.400000ns, VDD,
+ 406418.500000ns, VSS,
+ 407139.000000ns, VSS,
+ 407139.100000ns, VDD,
+ 407739.500000ns, VDD,
+ 407739.600000ns, VSS,
+ 407979.700000ns, VSS,
+ 407979.800000ns, VDD,
+ 408219.900000ns, VDD,
+ 408220.000000ns, VSS,
+ 408460.100000ns, VSS,
+ 408460.200000ns, VDD,
+ 408820.400000ns, VDD,
+ 408820.500000ns, VSS,
+ 409060.600000ns, VSS,
+ 409060.700000ns, VDD,
+ 409420.900000ns, VDD,
+ 409421.000000ns, VSS,
+ 409541.000000ns, VSS,
+ 409541.100000ns, VDD,
+ 409781.200000ns, VDD,
+ 409781.300000ns, VSS,
+ 409901.300000ns, VSS,
+ 409901.400000ns, VDD,
+ 410141.500000ns, VDD,
+ 410141.600000ns, VSS,
+ 410381.700000ns, VSS,
+ 410381.800000ns, VDD,
+ 410501.800000ns, VDD,
+ 410501.900000ns, VSS,
+ 410982.200000ns, VSS,
+ 410982.300000ns, VDD,
+ 411342.500000ns, VDD,
+ 411342.600000ns, VSS,
+ 411943.000000ns, VSS,
+ 411943.100000ns, VDD,
+ 413384.200000ns, VDD,
+ 413384.300000ns, VSS,
+ 413744.500000ns, VSS,
+ 413744.600000ns, VDD,
+ 414104.800000ns, VDD,
+ 414104.900000ns, VSS,
+ 414705.300000ns, VSS,
+ 414705.400000ns, VDD,
+ 414825.400000ns, VDD,
+ 414825.500000ns, VSS,
+ 415185.700000ns, VSS,
+ 415185.800000ns, VDD,
+ 415425.900000ns, VDD,
+ 415426.000000ns, VSS,
+ 415546.000000ns, VSS,
+ 415546.100000ns, VDD,
+ 415786.200000ns, VDD,
+ 415786.300000ns, VSS,
+ 415906.300000ns, VSS,
+ 415906.400000ns, VDD,
+ 416867.100000ns, VDD,
+ 416867.200000ns, VSS,
+ 416987.200000ns, VSS,
+ 416987.300000ns, VDD,
+ 417227.400000ns, VDD,
+ 417227.500000ns, VSS,
+ 417587.700000ns, VSS,
+ 417587.800000ns, VDD,
+ 417707.800000ns, VDD,
+ 417707.900000ns, VSS,
+ 417948.000000ns, VSS,
+ 417948.100000ns, VDD,
+ 418668.600000ns, VDD,
+ 418668.700000ns, VSS,
+ 418788.700000ns, VSS,
+ 418788.800000ns, VDD,
+ 419869.600000ns, VDD,
+ 419869.700000ns, VSS,
+ 419989.700000ns, VSS,
+ 419989.800000ns, VDD,
+ 420590.200000ns, VDD,
+ 420590.300000ns, VSS,
+ 421310.800000ns, VSS,
+ 421310.900000ns, VDD,
+ 421551.000000ns, VDD,
+ 421551.100000ns, VSS,
+ 421911.300000ns, VSS,
+ 421911.400000ns, VDD,
+ 422271.600000ns, VDD,
+ 422271.700000ns, VSS,
+ 422391.700000ns, VSS,
+ 422391.800000ns, VDD,
+ 422752.000000ns, VDD,
+ 422752.100000ns, VSS,
+ 422992.200000ns, VSS,
+ 422992.300000ns, VDD,
+ 423712.800000ns, VDD,
+ 423712.900000ns, VSS,
+ 423832.900000ns, VSS,
+ 423833.000000ns, VDD,
+ 424313.300000ns, VDD,
+ 424313.400000ns, VSS,
+ 424553.500000ns, VSS,
+ 424553.600000ns, VDD,
+ 424793.700000ns, VDD,
+ 424793.800000ns, VSS,
+ 425033.900000ns, VSS,
+ 425034.000000ns, VDD,
+ 425394.200000ns, VDD,
+ 425394.300000ns, VSS,
+ 425994.700000ns, VSS,
+ 425994.800000ns, VDD,
+ 426114.800000ns, VDD,
+ 426114.900000ns, VSS,
+ 426355.000000ns, VSS,
+ 426355.100000ns, VDD,
+ 426715.300000ns, VDD,
+ 426715.400000ns, VSS,
+ 427556.000000ns, VSS,
+ 427556.100000ns, VDD,
+ 428156.500000ns, VDD,
+ 428156.600000ns, VSS,
+ 428396.700000ns, VSS,
+ 428396.800000ns, VDD,
+ 429117.300000ns, VDD,
+ 429117.400000ns, VSS,
+ 429237.400000ns, VSS,
+ 429237.500000ns, VDD,
+ 430198.200000ns, VDD,
+ 430198.300000ns, VSS,
+ 430798.700000ns, VSS,
+ 430798.800000ns, VDD,
+ 431038.900000ns, VDD,
+ 431039.000000ns, VSS,
+ 431399.200000ns, VSS,
+ 431399.300000ns, VDD,
+ 431999.700000ns, VDD,
+ 431999.800000ns, VSS,
+ 432119.800000ns, VSS,
+ 432119.900000ns, VDD,
+ 432239.900000ns, VDD,
+ 432240.000000ns, VSS,
+ 432480.100000ns, VSS,
+ 432480.200000ns, VDD,
+ 432840.400000ns, VDD,
+ 432840.500000ns, VSS,
+ 432960.500000ns, VSS,
+ 432960.600000ns, VDD,
+ 433921.300000ns, VDD,
+ 433921.400000ns, VSS,
+ 434281.600000ns, VSS,
+ 434281.700000ns, VDD,
+ 435362.500000ns, VDD,
+ 435362.600000ns, VSS,
+ 435963.000000ns, VSS,
+ 435963.100000ns, VDD,
+ 436443.400000ns, VDD,
+ 436443.500000ns, VSS,
+ 436563.500000ns, VSS,
+ 436563.600000ns, VDD,
+ 436683.600000ns, VDD,
+ 436683.700000ns, VSS,
+ 436923.800000ns, VSS,
+ 436923.900000ns, VDD,
+ 437043.900000ns, VDD,
+ 437044.000000ns, VSS,
+ 437764.500000ns, VSS,
+ 437764.600000ns, VDD,
+ 438244.900000ns, VDD,
+ 438245.000000ns, VSS,
+ 439085.600000ns, VSS,
+ 439085.700000ns, VDD,
+ 439806.200000ns, VDD,
+ 439806.300000ns, VSS,
+ 440046.400000ns, VSS,
+ 440046.500000ns, VDD,
+ 440646.900000ns, VDD,
+ 440647.000000ns, VSS,
+ 440767.000000ns, VSS,
+ 440767.100000ns, VDD,
+ 441727.800000ns, VDD,
+ 441727.900000ns, VSS,
+ 442208.200000ns, VSS,
+ 442208.300000ns, VDD,
+ 442568.500000ns, VDD,
+ 442568.600000ns, VSS,
+ 442688.600000ns, VSS,
+ 442688.700000ns, VDD,
+ 443048.900000ns, VDD,
+ 443049.000000ns, VSS,
+ 443169.000000ns, VSS,
+ 443169.100000ns, VDD,
+ 443289.100000ns, VDD,
+ 443289.200000ns, VSS,
+ 443529.300000ns, VSS,
+ 443529.400000ns, VDD,
+ 443769.500000ns, VDD,
+ 443769.600000ns, VSS,
+ 444129.800000ns, VSS,
+ 444129.900000ns, VDD,
+ 444370.000000ns, VDD,
+ 444370.100000ns, VSS,
+ 444490.100000ns, VSS,
+ 444490.200000ns, VDD,
+ 445210.700000ns, VDD,
+ 445210.800000ns, VSS,
+ 445330.800000ns, VSS,
+ 445330.900000ns, VDD,
+ 445811.200000ns, VDD,
+ 445811.300000ns, VSS,
+ 446051.400000ns, VSS,
+ 446051.500000ns, VDD,
+ 446892.100000ns, VDD,
+ 446892.200000ns, VSS,
+ 447012.200000ns, VSS,
+ 447012.300000ns, VDD,
+ 447492.600000ns, VDD,
+ 447492.700000ns, VSS,
+ 447612.700000ns, VSS,
+ 447612.800000ns, VDD,
+ 447852.900000ns, VDD,
+ 447853.000000ns, VSS,
+ 447973.000000ns, VSS,
+ 447973.100000ns, VDD,
+ 448333.300000ns, VDD,
+ 448333.400000ns, VSS,
+ 449534.300000ns, VSS,
+ 449534.400000ns, VDD,
+ 449894.600000ns, VDD,
+ 449894.700000ns, VSS,
+ 450254.900000ns, VSS,
+ 450255.000000ns, VDD,
+ 450495.100000ns, VDD,
+ 450495.200000ns, VSS,
+ 450615.200000ns, VSS,
+ 450615.300000ns, VDD,
+ 450735.300000ns, VDD,
+ 450735.400000ns, VSS,
+ 451095.600000ns, VSS,
+ 451095.700000ns, VDD,
+ 451455.900000ns, VDD,
+ 451456.000000ns, VSS,
+ 451576.000000ns, VSS,
+ 451576.100000ns, VDD,
+ 451816.200000ns, VDD,
+ 451816.300000ns, VSS,
+ 452296.600000ns, VSS,
+ 452296.700000ns, VDD,
+ 452536.800000ns, VDD,
+ 452536.900000ns, VSS,
+ 452656.900000ns, VSS,
+ 452657.000000ns, VDD,
+ 452777.000000ns, VDD,
+ 452777.100000ns, VSS,
+ 453137.300000ns, VSS,
+ 453137.400000ns, VDD,
+ 453497.600000ns, VDD,
+ 453497.700000ns, VSS,
+ 453737.800000ns, VSS,
+ 453737.900000ns, VDD,
+ 453978.000000ns, VDD,
+ 453978.100000ns, VSS,
+ 454218.200000ns, VSS,
+ 454218.300000ns, VDD,
+ 454578.500000ns, VDD,
+ 454578.600000ns, VSS,
+ 454698.600000ns, VSS,
+ 454698.700000ns, VDD,
+ 455058.900000ns, VDD,
+ 455059.000000ns, VSS,
+ 455299.100000ns, VSS,
+ 455299.200000ns, VDD,
+ 456259.900000ns, VDD,
+ 456260.000000ns, VSS,
+ 456620.200000ns, VSS,
+ 456620.300000ns, VDD,
+ 457100.600000ns, VDD,
+ 457100.700000ns, VSS,
+ 457220.700000ns, VSS,
+ 457220.800000ns, VDD,
+ 457821.200000ns, VDD,
+ 457821.300000ns, VSS,
+ 458181.500000ns, VSS,
+ 458181.600000ns, VDD,
+ 458782.000000ns, VDD,
+ 458782.100000ns, VSS,
+ 458902.100000ns, VSS,
+ 458902.200000ns, VDD,
+ 459622.700000ns, VDD,
+ 459622.800000ns, VSS,
+ 460103.100000ns, VSS,
+ 460103.200000ns, VDD,
+ 460343.300000ns, VDD,
+ 460343.400000ns, VSS,
+ 460823.700000ns, VSS,
+ 460823.800000ns, VDD,
+ 461424.200000ns, VDD,
+ 461424.300000ns, VSS,
+ 461544.300000ns, VSS,
+ 461544.400000ns, VDD,
+ 462024.700000ns, VDD,
+ 462024.800000ns, VSS,
+ 462385.000000ns, VSS,
+ 462385.100000ns, VDD,
+ 462505.100000ns, VDD,
+ 462505.200000ns, VSS,
+ 462625.200000ns, VSS,
+ 462625.300000ns, VDD,
+ 463826.200000ns, VDD,
+ 463826.300000ns, VSS,
+ 464066.400000ns, VSS,
+ 464066.500000ns, VDD,
+ 464186.500000ns, VDD,
+ 464186.600000ns, VSS,
+ 464546.800000ns, VSS,
+ 464546.900000ns, VDD,
+ 464787.000000ns, VDD,
+ 464787.100000ns, VSS,
+ 464907.100000ns, VSS,
+ 464907.200000ns, VDD,
+ 465747.800000ns, VDD,
+ 465747.900000ns, VSS,
+ 466108.100000ns, VSS,
+ 466108.200000ns, VDD,
+ 466828.700000ns, VDD,
+ 466828.800000ns, VSS,
+ 466948.800000ns, VSS,
+ 466948.900000ns, VDD,
+ 467309.100000ns, VDD,
+ 467309.200000ns, VSS,
+ 467429.200000ns, VSS,
+ 467429.300000ns, VDD,
+ 467669.400000ns, VDD,
+ 467669.500000ns, VSS,
+ 468029.700000ns, VSS,
+ 468029.800000ns, VDD,
+ 468390.000000ns, VDD,
+ 468390.100000ns, VSS,
+ 469230.700000ns, VSS,
+ 469230.800000ns, VDD,
+ 469470.900000ns, VDD,
+ 469471.000000ns, VSS,
+ 469591.000000ns, VSS,
+ 469591.100000ns, VDD,
+ 470671.900000ns, VDD,
+ 470672.000000ns, VSS,
+ 470792.000000ns, VSS,
+ 470792.100000ns, VDD,
+ 471032.200000ns, VDD,
+ 471032.300000ns, VSS,
+ 471752.800000ns, VSS,
+ 471752.900000ns, VDD,
+ 472113.100000ns, VDD,
+ 472113.200000ns, VSS,
+ 472233.200000ns, VSS,
+ 472233.300000ns, VDD,
+ 472353.300000ns, VDD,
+ 472353.400000ns, VSS,
+ 472713.600000ns, VSS,
+ 472713.700000ns, VDD,
+ 473073.900000ns, VDD,
+ 473074.000000ns, VSS,
+ 473194.000000ns, VSS,
+ 473194.100000ns, VDD,
+ 473674.400000ns, VDD,
+ 473674.500000ns, VSS,
+ 474154.800000ns, VSS,
+ 474154.900000ns, VDD,
+ 475235.700000ns, VDD,
+ 475235.800000ns, VSS,
+ 475836.200000ns, VSS,
+ 475836.300000ns, VDD,
+ 476196.500000ns, VDD,
+ 476196.600000ns, VSS,
+ 476436.700000ns, VSS,
+ 476436.800000ns, VDD,
+ 476797.000000ns, VDD,
+ 476797.100000ns, VSS,
+ 477277.400000ns, VSS,
+ 477277.500000ns, VDD,
+ 477637.700000ns, VDD,
+ 477637.800000ns, VSS,
+ 477998.000000ns, VSS,
+ 477998.100000ns, VDD,
+ 478358.300000ns, VDD,
+ 478358.400000ns, VSS,
+ 478958.800000ns, VSS,
+ 478958.900000ns, VDD,
+ 479199.000000ns, VDD,
+ 479199.100000ns, VSS,
+ 479799.500000ns, VSS,
+ 479799.600000ns, VDD,
+ 480880.400000ns, VDD,
+ 480880.500000ns, VSS,
+ 481000.500000ns, VSS,
+ 481000.600000ns, VDD,
+ 482081.400000ns, VDD,
+ 482081.500000ns, VSS,
+ 482922.100000ns, VSS,
+ 482922.200000ns, VDD,
+ 483162.300000ns, VDD,
+ 483162.400000ns, VSS,
+ 483402.500000ns, VSS,
+ 483402.600000ns, VDD,
+ 483642.700000ns, VDD,
+ 483642.800000ns, VSS,
+ 483762.800000ns, VSS,
+ 483762.900000ns, VDD,
+ 484603.500000ns, VDD,
+ 484603.600000ns, VSS,
+ 486284.900000ns, VSS,
+ 486285.000000ns, VDD,
+ 486405.000000ns, VDD,
+ 486405.100000ns, VSS,
+ 486765.300000ns, VSS,
+ 486765.400000ns, VDD,
+ 487365.800000ns, VDD,
+ 487365.900000ns, VSS,
+ 487726.100000ns, VSS,
+ 487726.200000ns, VDD,
+ 487846.200000ns, VDD,
+ 487846.300000ns, VSS,
+ 488326.600000ns, VSS,
+ 488326.700000ns, VDD,
+ 488566.800000ns, VDD,
+ 488566.900000ns, VSS,
+ 488686.900000ns, VSS,
+ 488687.000000ns, VDD,
+ 488807.000000ns, VDD,
+ 488807.100000ns, VSS,
+ 489047.200000ns, VSS,
+ 489047.300000ns, VDD,
+ 490248.200000ns, VDD,
+ 490248.300000ns, VSS,
+ 490488.400000ns, VSS,
+ 490488.500000ns, VDD,
+ 490608.500000ns, VDD,
+ 490608.600000ns, VSS,
+ 490728.600000ns, VSS,
+ 490728.700000ns, VDD,
+ 491449.200000ns, VDD,
+ 491449.300000ns, VSS,
+ 491689.400000ns, VSS,
+ 491689.500000ns, VDD,
+ 492169.800000ns, VDD,
+ 492169.900000ns, VSS,
+ 492289.900000ns, VSS,
+ 492290.000000ns, VDD,
+ 492530.100000ns, VDD,
+ 492530.200000ns, VSS,
+ 493010.500000ns, VSS,
+ 493010.600000ns, VDD,
+ 493370.800000ns, VDD,
+ 493370.900000ns, VSS,
+ 493611.000000ns, VSS,
+ 493611.100000ns, VDD,
+ 494211.500000ns, VDD,
+ 494211.600000ns, VSS,
+ 494451.700000ns, VSS,
+ 494451.800000ns, VDD,
+ 494812.000000ns, VDD,
+ 494812.100000ns, VSS,
+ 495532.600000ns, VSS,
+ 495532.700000ns, VDD,
+ 496493.400000ns, VDD,
+ 496493.500000ns, VSS,
+ 496733.600000ns, VSS,
+ 496733.700000ns, VDD,
+ 496853.700000ns, VDD,
+ 496853.800000ns, VSS,
+ 497934.600000ns, VSS,
+ 497934.700000ns, VDD,
+ 498294.900000ns, VDD,
+ 498295.000000ns, VSS,
+ 498415.000000ns, VSS,
+ 498415.100000ns, VDD,
+ 498655.200000ns, VDD,
+ 498655.300000ns, VSS,
+ 498895.400000ns, VSS,
+ 498895.500000ns, VDD,
+ 499255.700000ns, VDD,
+ 499255.800000ns, VSS,
+ 499495.900000ns, VSS,
+ 499496.000000ns, VDD,
+ 499616.000000ns, VDD,
+ 499616.100000ns, VSS,
+ 499736.100000ns, VSS,
+ 499736.200000ns, VDD,
+ 499976.300000ns, VDD,
+ 499976.400000ns, VSS,
+ 500096.400000ns, VSS,
+ 500096.500000ns, VDD,
+ 500456.700000ns, VDD,
+ 500456.800000ns, VSS,
+ 500817.000000ns, VSS,
+ 500817.100000ns, VDD,
+ 501657.700000ns, VDD,
+ 501657.800000ns, VSS,
+ 501777.800000ns, VSS,
+ 501777.900000ns, VDD,
+ 501897.900000ns, VDD,
+ 501898.000000ns, VSS,
+ 502018.000000ns, VSS,
+ 502018.100000ns, VDD,
+ 502498.400000ns, VDD,
+ 502498.500000ns, VSS,
+ 502978.800000ns, VSS,
+ 502978.900000ns, VDD,
+ 503339.100000ns, VDD,
+ 503339.200000ns, VSS,
+ 503819.500000ns, VSS,
+ 503819.600000ns, VDD,
+ 503939.600000ns, VDD,
+ 503939.700000ns, VSS,
+ 504420.000000ns, VSS,
+ 504420.100000ns, VDD,
+ 504660.200000ns, VDD,
+ 504660.300000ns, VSS,
+ 505020.500000ns, VSS,
+ 505020.600000ns, VDD,
+ 505140.600000ns, VDD,
+ 505140.700000ns, VSS,
+ 505500.900000ns, VSS,
+ 505501.000000ns, VDD,
+ 506221.500000ns, VDD,
+ 506221.600000ns, VSS,
+ 506461.700000ns, VSS,
+ 506461.800000ns, VDD,
+ 506581.800000ns, VDD,
+ 506581.900000ns, VSS,
+ 506701.900000ns, VSS,
+ 506702.000000ns, VDD,
+ 507062.200000ns, VDD,
+ 507062.300000ns, VSS,
+ 507782.800000ns, VSS,
+ 507782.900000ns, VDD,
+ 507902.900000ns, VDD,
+ 507903.000000ns, VSS,
+ 508383.300000ns, VSS,
+ 508383.400000ns, VDD,
+ 508503.400000ns, VDD,
+ 508503.500000ns, VSS,
+ 508863.700000ns, VSS,
+ 508863.800000ns, VDD,
+ 509224.000000ns, VDD,
+ 509224.100000ns, VSS,
+ 509344.100000ns, VSS,
+ 509344.200000ns, VDD,
+ 509704.400000ns, VDD,
+ 509704.500000ns, VSS,
+ 509824.500000ns, VSS,
+ 509824.600000ns, VDD,
+ 510545.100000ns, VDD,
+ 510545.200000ns, VSS,
+ 511145.600000ns, VSS,
+ 511145.700000ns, VDD,
+ 511385.800000ns, VDD,
+ 511385.900000ns, VSS,
+ 511626.000000ns, VSS,
+ 511626.100000ns, VDD,
+ 511986.300000ns, VDD,
+ 511986.400000ns, VSS,
+ 512106.400000ns, VSS,
+ 512106.500000ns, VDD,
+ 512706.900000ns, VDD,
+ 512707.000000ns, VSS,
+ 512827.000000ns, VSS,
+ 512827.100000ns, VDD,
+ 512947.100000ns, VDD,
+ 512947.200000ns, VSS,
+ 513187.300000ns, VSS,
+ 513187.400000ns, VDD,
+ 513307.400000ns, VDD,
+ 513307.500000ns, VSS,
+ 513427.500000ns, VSS,
+ 513427.600000ns, VDD,
+ 513547.600000ns, VDD,
+ 513547.700000ns, VSS,
+ 513907.900000ns, VSS,
+ 513908.000000ns, VDD,
+ 514268.200000ns, VDD,
+ 514268.300000ns, VSS,
+ 514628.500000ns, VSS,
+ 514628.600000ns, VDD,
+ 515229.000000ns, VDD,
+ 515229.100000ns, VSS,
+ 515349.100000ns, VSS,
+ 515349.200000ns, VDD,
+ 515589.300000ns, VDD,
+ 515589.400000ns, VSS,
+ 515709.400000ns, VSS,
+ 515709.500000ns, VDD,
+ 515829.500000ns, VDD,
+ 515829.600000ns, VSS,
+ 515949.600000ns, VSS,
+ 515949.700000ns, VDD,
+ 517270.700000ns, VDD,
+ 517270.800000ns, VSS,
+ 517751.100000ns, VSS,
+ 517751.200000ns, VDD,
+ 517871.200000ns, VDD,
+ 517871.300000ns, VSS,
+ 517991.300000ns, VSS,
+ 517991.400000ns, VDD,
+ 518351.600000ns, VDD,
+ 518351.700000ns, VSS,
+ 518711.900000ns, VSS,
+ 518712.000000ns, VDD,
+ 518832.000000ns, VDD,
+ 518832.100000ns, VSS,
+ 519072.200000ns, VSS,
+ 519072.300000ns, VDD,
+ 520273.200000ns, VDD,
+ 520273.300000ns, VSS,
+ 520633.500000ns, VSS,
+ 520633.600000ns, VDD,
+ 521113.900000ns, VDD,
+ 521114.000000ns, VSS,
+ 521234.000000ns, VSS,
+ 521234.100000ns, VDD,
+ 521594.300000ns, VDD,
+ 521594.400000ns, VSS,
+ 521954.600000ns, VSS,
+ 521954.700000ns, VDD,
+ 522675.200000ns, VDD,
+ 522675.300000ns, VSS,
+ 522795.300000ns, VSS,
+ 522795.400000ns, VDD,
+ 523155.600000ns, VDD,
+ 523155.700000ns, VSS,
+ 523636.000000ns, VSS,
+ 523636.100000ns, VDD,
+ 523996.300000ns, VDD,
+ 523996.400000ns, VSS,
+ 524236.500000ns, VSS,
+ 524236.600000ns, VDD,
+ 525437.500000ns, VDD,
+ 525437.600000ns, VSS,
+ 525677.700000ns, VSS,
+ 525677.800000ns, VDD,
+ 526038.000000ns, VDD,
+ 526038.100000ns, VSS,
+ 526278.200000ns, VSS,
+ 526278.300000ns, VDD,
+ 526758.600000ns, VDD,
+ 526758.700000ns, VSS,
+ 527239.000000ns, VSS,
+ 527239.100000ns, VDD,
+ 528319.900000ns, VDD,
+ 528320.000000ns, VSS,
+ 529160.600000ns, VSS,
+ 529160.700000ns, VDD,
+ 529400.800000ns, VDD,
+ 529400.900000ns, VSS,
+ 529761.100000ns, VSS,
+ 529761.200000ns, VDD,
+ 530481.700000ns, VDD,
+ 530481.800000ns, VSS,
+ 531442.500000ns, VSS,
+ 531442.600000ns, VDD,
+ 531802.800000ns, VDD,
+ 531802.900000ns, VSS,
+ 532043.000000ns, VSS,
+ 532043.100000ns, VDD,
+ 532403.300000ns, VDD,
+ 532403.400000ns, VSS,
+ 532643.500000ns, VSS,
+ 532643.600000ns, VDD,
+ 532883.700000ns, VDD,
+ 532883.800000ns, VSS,
+ 533003.800000ns, VSS,
+ 533003.900000ns, VDD,
+ 533123.900000ns, VDD,
+ 533124.000000ns, VSS,
+ 533244.000000ns, VSS,
+ 533244.100000ns, VDD,
+ 533364.100000ns, VDD,
+ 533364.200000ns, VSS,
+ 533604.300000ns, VSS,
+ 533604.400000ns, VDD,
+ 534084.700000ns, VDD,
+ 534084.800000ns, VSS,
+ 534445.000000ns, VSS,
+ 534445.100000ns, VDD,
+ 534565.100000ns, VDD,
+ 534565.200000ns, VSS,
+ 535285.700000ns, VSS,
+ 535285.800000ns, VDD,
+ 536967.100000ns, VDD,
+ 536967.200000ns, VSS,
+ 538048.000000ns, VSS,
+ 538048.100000ns, VDD,
+ 538528.400000ns, VDD,
+ 538528.500000ns, VSS,
+ 538648.500000ns, VSS,
+ 538648.600000ns, VDD,
+ 540810.300000ns, VDD,
+ 540810.400000ns, VSS,
+ 541170.600000ns, VSS,
+ 541170.700000ns, VDD,
+ 541290.700000ns, VDD,
+ 541290.800000ns, VSS,
+ 541410.800000ns, VSS,
+ 541410.900000ns, VDD,
+ 541891.200000ns, VDD,
+ 541891.300000ns, VSS,
+ 542251.500000ns, VSS,
+ 542251.600000ns, VDD,
+ 542731.900000ns, VDD,
+ 542732.000000ns, VSS,
+ 542852.000000ns, VSS,
+ 542852.100000ns, VDD,
+ 543212.300000ns, VDD,
+ 543212.400000ns, VSS,
+ 543332.400000ns, VSS,
+ 543332.500000ns, VDD,
+ 543692.700000ns, VDD,
+ 543692.800000ns, VSS,
+ 544053.000000ns, VSS,
+ 544053.100000ns, VDD,
+ 544173.100000ns, VDD,
+ 544173.200000ns, VSS,
+ 544293.200000ns, VSS,
+ 544293.300000ns, VDD,
+ 545734.400000ns, VDD,
+ 545734.500000ns, VSS,
+ 545854.500000ns, VSS,
+ 545854.600000ns, VDD,
+ 545974.600000ns, VDD,
+ 545974.700000ns, VSS,
+ 546334.900000ns, VSS,
+ 546335.000000ns, VDD,
+ 546455.000000ns, VDD,
+ 546455.100000ns, VSS,
+ 546575.100000ns, VSS,
+ 546575.200000ns, VDD,
+ 546935.400000ns, VDD,
+ 546935.500000ns, VSS,
+ 547175.600000ns, VSS,
+ 547175.700000ns, VDD,
+ 548376.600000ns, VDD,
+ 548376.700000ns, VSS,
+ 548857.000000ns, VSS,
+ 548857.100000ns, VDD,
+ 549337.400000ns, VDD,
+ 549337.500000ns, VSS,
+ 549817.800000ns, VSS,
+ 549817.900000ns, VDD,
+ 550538.400000ns, VDD,
+ 550538.500000ns, VSS,
+ 550778.600000ns, VSS,
+ 550778.700000ns, VDD,
+ 551619.300000ns, VDD,
+ 551619.400000ns, VSS,
+ 551859.500000ns, VSS,
+ 551859.600000ns, VDD,
+ 552099.700000ns, VDD,
+ 552099.800000ns, VSS,
+ 552339.900000ns, VSS,
+ 552340.000000ns, VDD,
+ 552580.100000ns, VDD,
+ 552580.200000ns, VSS,
+ 552700.200000ns, VSS,
+ 552700.300000ns, VDD,
+ 553060.500000ns, VDD,
+ 553060.600000ns, VSS,
+ 553180.600000ns, VSS,
+ 553180.700000ns, VDD,
+ 553300.700000ns, VDD,
+ 553300.800000ns, VSS,
+ 553420.800000ns, VSS,
+ 553420.900000ns, VDD,
+ 553540.900000ns, VDD,
+ 553541.000000ns, VSS,
+ 553661.000000ns, VSS,
+ 553661.100000ns, VDD,
+ 554501.700000ns, VDD,
+ 554501.800000ns, VSS,
+ 554862.000000ns, VSS,
+ 554862.100000ns, VDD,
+ 555102.200000ns, VDD,
+ 555102.300000ns, VSS,
+ 556423.300000ns, VSS,
+ 556423.400000ns, VDD,
+ 556903.700000ns, VDD,
+ 556903.800000ns, VSS,
+ 558465.000000ns, VSS,
+ 558465.100000ns, VDD,
+ 558825.300000ns, VDD,
+ 558825.400000ns, VSS,
+ 559425.800000ns, VSS,
+ 559425.900000ns, VDD,
+ 559666.000000ns, VDD,
+ 559666.100000ns, VSS,
+ 559906.200000ns, VSS,
+ 559906.300000ns, VDD,
+ 560026.300000ns, VDD,
+ 560026.400000ns, VSS,
+ 560146.400000ns, VSS,
+ 560146.500000ns, VDD,
+ 562188.100000ns, VDD,
+ 562188.200000ns, VSS,
+ 562308.200000ns, VSS,
+ 562308.300000ns, VDD,
+ 562428.300000ns, VDD,
+ 562428.400000ns, VSS,
+ 562788.600000ns, VSS,
+ 562788.700000ns, VDD,
+ 563028.800000ns, VDD,
+ 563028.900000ns, VSS,
+ 563148.900000ns, VSS,
+ 563149.000000ns, VDD,
+ 563629.300000ns, VDD,
+ 563629.400000ns, VSS,
+ 564349.900000ns, VSS,
+ 564350.000000ns, VDD,
+ 564950.400000ns, VDD,
+ 564950.500000ns, VSS,
+ 565310.700000ns, VSS,
+ 565310.800000ns, VDD,
+ 565911.200000ns, VDD,
+ 565911.300000ns, VSS,
+ 566031.300000ns, VSS,
+ 566031.400000ns, VDD,
+ 566511.700000ns, VDD,
+ 566511.800000ns, VSS,
+ 566751.900000ns, VSS,
+ 566752.000000ns, VDD,
+ 567472.500000ns, VDD,
+ 567472.600000ns, VSS,
+ 567832.800000ns, VSS,
+ 567832.900000ns, VDD,
+ 568193.100000ns, VDD,
+ 568193.200000ns, VSS,
+ 568313.200000ns, VSS,
+ 568313.300000ns, VDD,
+ 568673.500000ns, VDD,
+ 568673.600000ns, VSS,
+ 568793.600000ns, VSS,
+ 568793.700000ns, VDD,
+ 569274.000000ns, VDD,
+ 569274.100000ns, VSS,
+ 569514.200000ns, VSS,
+ 569514.300000ns, VDD,
+ 569634.300000ns, VDD,
+ 569634.400000ns, VSS,
+ 569874.500000ns, VSS,
+ 569874.600000ns, VDD,
+ 569994.600000ns, VDD,
+ 569994.700000ns, VSS,
+ 570114.700000ns, VSS,
+ 570114.800000ns, VDD,
+ 570234.800000ns, VDD,
+ 570234.900000ns, VSS,
+ 570595.100000ns, VSS,
+ 570595.200000ns, VDD,
+ 570715.200000ns, VDD,
+ 570715.300000ns, VSS,
+ 571315.700000ns, VSS,
+ 571315.800000ns, VDD,
+ 572036.300000ns, VDD,
+ 572036.400000ns, VSS,
+ 572636.800000ns, VSS,
+ 572636.900000ns, VDD,
+ 573357.400000ns, VDD,
+ 573357.500000ns, VSS,
+ 574078.000000ns, VSS,
+ 574078.100000ns, VDD,
+ 574318.200000ns, VDD,
+ 574318.300000ns, VSS,
+ 574798.600000ns, VSS,
+ 574798.700000ns, VDD,
+ 575759.400000ns, VDD,
+ 575759.500000ns, VSS,
+ 575999.600000ns, VSS,
+ 575999.700000ns, VDD,
+ 576720.200000ns, VDD,
+ 576720.300000ns, VSS,
+ 576840.300000ns, VSS,
+ 576840.400000ns, VDD,
+ 577200.600000ns, VDD,
+ 577200.700000ns, VSS,
+ 577320.700000ns, VSS,
+ 577320.800000ns, VDD,
+ 577681.000000ns, VDD,
+ 577681.100000ns, VSS,
+ 578041.300000ns, VSS,
+ 578041.400000ns, VDD,
+ 578281.500000ns, VDD,
+ 578281.600000ns, VSS,
+ 578641.800000ns, VSS,
+ 578641.900000ns, VDD,
+ 579122.200000ns, VDD,
+ 579122.300000ns, VSS,
+ 579242.300000ns, VSS,
+ 579242.400000ns, VDD,
+ 579362.400000ns, VDD,
+ 579362.500000ns, VSS,
+ 579602.600000ns, VSS,
+ 579602.700000ns, VDD,
+ 580923.700000ns, VDD,
+ 580923.800000ns, VSS,
+ 581644.300000ns, VSS,
+ 581644.400000ns, VDD,
+ 581764.400000ns, VDD,
+ 581764.500000ns, VSS,
+ 581884.500000ns, VSS,
+ 581884.600000ns, VDD,
+ 582244.800000ns, VDD,
+ 582244.900000ns, VSS,
+ 582364.900000ns, VSS,
+ 582365.000000ns, VDD,
+ 582725.200000ns, VDD,
+ 582725.300000ns, VSS,
+ 582965.400000ns, VSS,
+ 582965.500000ns, VDD,
+ 583085.500000ns, VDD,
+ 583085.600000ns, VSS,
+ 583445.800000ns, VSS,
+ 583445.900000ns, VDD,
+ 583926.200000ns, VDD,
+ 583926.300000ns, VSS,
+ 584046.300000ns, VSS,
+ 584046.400000ns, VDD,
+ 585247.300000ns, VDD,
+ 585247.400000ns, VSS,
+ 585607.600000ns, VSS,
+ 585607.700000ns, VDD,
+ 585847.800000ns, VDD,
+ 585847.900000ns, VSS,
+ 586448.300000ns, VSS,
+ 586448.400000ns, VDD,
+ 587168.900000ns, VDD,
+ 587169.000000ns, VSS,
+ 587769.400000ns, VSS,
+ 587769.500000ns, VDD,
+ 588009.600000ns, VDD,
+ 588009.700000ns, VSS,
+ 588129.700000ns, VSS,
+ 588129.800000ns, VDD,
+ 588369.900000ns, VDD,
+ 588370.000000ns, VSS,
+ 588850.300000ns, VSS,
+ 588850.400000ns, VDD,
+ 588970.400000ns, VDD,
+ 588970.500000ns, VSS,
+ 589330.700000ns, VSS,
+ 589330.800000ns, VDD,
+ 589811.100000ns, VDD,
+ 589811.200000ns, VSS,
+ 590051.300000ns, VSS,
+ 590051.400000ns, VDD,
+ 590771.900000ns, VDD,
+ 590772.000000ns, VSS,
+ 591492.500000ns, VSS,
+ 591492.600000ns, VDD,
+ 591612.600000ns, VDD,
+ 591612.700000ns, VSS,
+ 591852.800000ns, VSS,
+ 591852.900000ns, VDD,
+ 591972.900000ns, VDD,
+ 591973.000000ns, VSS,
+ 592093.000000ns, VSS,
+ 592093.100000ns, VDD,
+ 592333.200000ns, VDD,
+ 592333.300000ns, VSS,
+ 592573.400000ns, VSS,
+ 592573.500000ns, VDD,
+ 593053.800000ns, VDD,
+ 593053.900000ns, VSS,
+ 593173.900000ns, VSS,
+ 593174.000000ns, VDD,
+ 594374.900000ns, VDD,
+ 594375.000000ns, VSS,
+ 594495.000000ns, VSS,
+ 594495.100000ns, VDD,
+ 595215.600000ns, VDD,
+ 595215.700000ns, VSS,
+ 595696.000000ns, VSS,
+ 595696.100000ns, VDD,
+ 596176.400000ns, VDD,
+ 596176.500000ns, VSS,
+ 596296.500000ns, VSS,
+ 596296.600000ns, VDD,
+ 596416.600000ns, VDD,
+ 596416.700000ns, VSS,
+ 596776.900000ns, VSS,
+ 596777.000000ns, VDD,
+ 597137.200000ns, VDD,
+ 597137.300000ns, VSS,
+ 597257.300000ns, VSS,
+ 597257.400000ns, VDD,
+ 597497.500000ns, VDD,
+ 597497.600000ns, VSS,
+ 597617.600000ns, VSS,
+ 597617.700000ns, VDD,
+ 597977.900000ns, VDD,
+ 597978.000000ns, VSS,
+ 598218.100000ns, VSS,
+ 598218.200000ns, VDD,
+ 598698.500000ns, VDD,
+ 598698.600000ns, VSS,
+ 598938.700000ns, VSS,
+ 598938.800000ns, VDD,
+ 599178.900000ns, VDD,
+ 599179.000000ns, VSS,
+ 599299.000000ns, VSS,
+ 599299.100000ns, VDD,
+ 599539.200000ns, VDD,
+ 599539.300000ns, VSS,
+ 599659.300000ns, VSS,
+ 599659.400000ns, VDD,
+ 600259.800000ns, VDD,
+ 600259.900000ns, VSS,
+ 600860.300000ns, VSS,
+ 600860.400000ns, VDD,
+ 600980.400000ns, VDD,
+ 600980.500000ns, VSS,
+ 601100.500000ns, VSS,
+ 601100.600000ns, VDD,
+ 601220.600000ns, VDD,
+ 601220.700000ns, VSS,
+ 602421.600000ns, VSS,
+ 602421.700000ns, VDD,
+ 602661.800000ns, VDD,
+ 602661.900000ns, VSS,
+ 603262.300000ns, VSS,
+ 603262.400000ns, VDD,
+ 604103.000000ns, VDD,
+ 604103.100000ns, VSS,
+ 604223.100000ns, VSS,
+ 604223.200000ns, VDD,
+ 604583.400000ns, VDD,
+ 604583.500000ns, VSS,
+ 604943.700000ns, VSS,
+ 604943.800000ns, VDD,
+ 605304.000000ns, VDD,
+ 605304.100000ns, VSS,
+ 605784.400000ns, VSS,
+ 605784.500000ns, VDD,
+ 606144.700000ns, VDD,
+ 606144.800000ns, VSS,
+ 606264.800000ns, VSS,
+ 606264.900000ns, VDD,
+ 606865.300000ns, VDD,
+ 606865.400000ns, VSS,
+ 606985.400000ns, VSS,
+ 606985.500000ns, VDD,
+ 607105.500000ns, VDD,
+ 607105.600000ns, VSS,
+ 607585.900000ns, VSS,
+ 607586.000000ns, VDD,
+ 607706.000000ns, VDD,
+ 607706.100000ns, VSS,
+ 608306.500000ns, VSS,
+ 608306.600000ns, VDD,
+ 608666.800000ns, VDD,
+ 608666.900000ns, VSS,
+ 609027.100000ns, VSS,
+ 609027.200000ns, VDD,
+ 609147.200000ns, VDD,
+ 609147.300000ns, VSS,
+ 609267.300000ns, VSS,
+ 609267.400000ns, VDD,
+ 609387.400000ns, VDD,
+ 609387.500000ns, VSS,
+ 609507.500000ns, VSS,
+ 609507.600000ns, VDD,
+ 610348.200000ns, VDD,
+ 610348.300000ns, VSS,
+ 610708.500000ns, VSS,
+ 610708.600000ns, VDD,
+ 611309.000000ns, VDD,
+ 611309.100000ns, VSS,
+ 611429.100000ns, VSS,
+ 611429.200000ns, VDD,
+ 611549.200000ns, VDD,
+ 611549.300000ns, VSS,
+ 611789.400000ns, VSS,
+ 611789.500000ns, VDD,
+ 612389.900000ns, VDD,
+ 612390.000000ns, VSS,
+ 612990.400000ns, VSS,
+ 612990.500000ns, VDD,
+ 613590.900000ns, VDD,
+ 613591.000000ns, VSS,
+ 613711.000000ns, VSS,
+ 613711.100000ns, VDD,
+ 613831.100000ns, VDD,
+ 613831.200000ns, VSS,
+ 614311.500000ns, VSS,
+ 614311.600000ns, VDD,
+ 614671.800000ns, VDD,
+ 614671.900000ns, VSS,
+ 614912.000000ns, VSS,
+ 614912.100000ns, VDD,
+ 615512.500000ns, VDD,
+ 615512.600000ns, VSS,
+ 615632.600000ns, VSS,
+ 615632.700000ns, VDD,
+ 615992.900000ns, VDD,
+ 615993.000000ns, VSS,
+ 616473.300000ns, VSS,
+ 616473.400000ns, VDD,
+ 617073.800000ns, VDD,
+ 617073.900000ns, VSS,
+ 617193.900000ns, VSS,
+ 617194.000000ns, VDD,
+ 617554.200000ns, VDD,
+ 617554.300000ns, VSS,
+ 617914.500000ns, VSS,
+ 617914.600000ns, VDD,
+ 618274.800000ns, VDD,
+ 618274.900000ns, VSS,
+ 618394.900000ns, VSS,
+ 618395.000000ns, VDD,
+ 618635.100000ns, VDD,
+ 618635.200000ns, VSS,
+ 618755.200000ns, VSS,
+ 618755.300000ns, VDD,
+ 618875.300000ns, VDD,
+ 618875.400000ns, VSS,
+ 619235.600000ns, VSS,
+ 619235.700000ns, VDD,
+ 620917.000000ns, VDD,
+ 620917.100000ns, VSS,
+ 621037.100000ns, VSS,
+ 621037.200000ns, VDD,
+ 621157.200000ns, VDD,
+ 621157.300000ns, VSS,
+ 621397.400000ns, VSS,
+ 621397.500000ns, VDD,
+ 621637.600000ns, VDD,
+ 621637.700000ns, VSS,
+ 621997.900000ns, VSS,
+ 621998.000000ns, VDD,
+ 622118.000000ns, VDD,
+ 622118.100000ns, VSS,
+ 622238.100000ns, VSS,
+ 622238.200000ns, VDD,
+ 622598.400000ns, VDD,
+ 622598.500000ns, VSS,
+ 622718.500000ns, VSS,
+ 622718.600000ns, VDD,
+ 622838.600000ns, VDD,
+ 622838.700000ns, VSS,
+ 623319.000000ns, VSS,
+ 623319.100000ns, VDD,
+ 623679.300000ns, VDD,
+ 623679.400000ns, VSS,
+ 623799.400000ns, VSS,
+ 623799.500000ns, VDD,
+ 624520.000000ns, VDD,
+ 624520.100000ns, VSS,
+ 624880.300000ns, VSS,
+ 624880.400000ns, VDD,
+ 625000.400000ns, VDD,
+ 625000.500000ns, VSS,
+ 625480.800000ns, VSS,
+ 625480.900000ns, VDD,
+ 625600.900000ns, VDD,
+ 625601.000000ns, VSS,
+ 625961.200000ns, VSS,
+ 625961.300000ns, VDD,
+ 626081.300000ns, VDD,
+ 626081.400000ns, VSS,
+ 626561.700000ns, VSS,
+ 626561.800000ns, VDD,
+ 626922.000000ns, VDD,
+ 626922.100000ns, VSS,
+ 627282.300000ns, VSS,
+ 627282.400000ns, VDD,
+ 627402.400000ns, VDD,
+ 627402.500000ns, VSS,
+ 627522.500000ns, VSS,
+ 627522.600000ns, VDD,
+ 627762.700000ns, VDD,
+ 627762.800000ns, VSS,
+ 628002.900000ns, VSS,
+ 628003.000000ns, VDD,
+ 628243.100000ns, VDD,
+ 628243.200000ns, VSS,
+ 628363.200000ns, VSS,
+ 628363.300000ns, VDD,
+ 629684.300000ns, VDD,
+ 629684.400000ns, VSS,
+ 630765.200000ns, VSS,
+ 630765.300000ns, VDD,
+ 630885.300000ns, VDD,
+ 630885.400000ns, VSS,
+ 631125.500000ns, VSS,
+ 631125.600000ns, VDD,
+ 631966.200000ns, VDD,
+ 631966.300000ns, VSS,
+ 632566.700000ns, VSS,
+ 632566.800000ns, VDD,
+ 632806.900000ns, VDD,
+ 632807.000000ns, VSS,
+ 632927.000000ns, VSS,
+ 632927.100000ns, VDD,
+ 633887.800000ns, VDD,
+ 633887.900000ns, VSS,
+ 634128.000000ns, VSS,
+ 634128.100000ns, VDD,
+ 634248.100000ns, VDD,
+ 634248.200000ns, VSS,
+ 634488.300000ns, VSS,
+ 634488.400000ns, VDD,
+ 634848.600000ns, VDD,
+ 634848.700000ns, VSS,
+ 634968.700000ns, VSS,
+ 634968.800000ns, VDD,
+ 635329.000000ns, VDD,
+ 635329.100000ns, VSS,
+ 635449.100000ns, VSS,
+ 635449.200000ns, VDD,
+ 635809.400000ns, VDD,
+ 635809.500000ns, VSS,
+ 636169.700000ns, VSS,
+ 636169.800000ns, VDD,
+ 636770.200000ns, VDD,
+ 636770.300000ns, VSS,
+ 637010.400000ns, VSS,
+ 637010.500000ns, VDD,
+ 637370.700000ns, VDD,
+ 637370.800000ns, VSS,
+ 637490.800000ns, VSS,
+ 637490.900000ns, VDD,
+ 637851.100000ns, VDD,
+ 637851.200000ns, VSS,
+ 637971.200000ns, VSS,
+ 637971.300000ns, VDD,
+ 638331.500000ns, VDD,
+ 638331.600000ns, VSS,
+ 638451.600000ns, VSS,
+ 638451.700000ns, VDD,
+ 638571.700000ns, VDD,
+ 638571.800000ns, VSS,
+ 639172.200000ns, VSS,
+ 639172.300000ns, VDD,
+ 640373.200000ns, VDD,
+ 640373.300000ns, VSS,
+ 640733.500000ns, VSS,
+ 640733.600000ns, VDD,
+ 640853.600000ns, VDD,
+ 640853.700000ns, VSS,
+ 640973.700000ns, VSS,
+ 640973.800000ns, VDD,
+ 641213.900000ns, VDD,
+ 641214.000000ns, VSS,
+ 641334.000000ns, VSS,
+ 641334.100000ns, VDD,
+ 641454.100000ns, VDD,
+ 641454.200000ns, VSS,
+ 641694.300000ns, VSS,
+ 641694.400000ns, VDD,
+ 641814.400000ns, VDD,
+ 641814.500000ns, VSS,
+ 642294.800000ns, VSS,
+ 642294.900000ns, VDD,
+ 642775.200000ns, VDD,
+ 642775.300000ns, VSS,
+ 642895.300000ns, VSS,
+ 642895.400000ns, VDD,
+ 643255.600000ns, VDD,
+ 643255.700000ns, VSS,
+ 643495.800000ns, VSS,
+ 643495.900000ns, VDD,
+ 644456.600000ns, VDD,
+ 644456.700000ns, VSS,
+ 644696.800000ns, VSS,
+ 644696.900000ns, VDD,
+ 645297.300000ns, VDD,
+ 645297.400000ns, VSS,
+ 645657.600000ns, VSS,
+ 645657.700000ns, VDD,
+ 645897.800000ns, VDD,
+ 645897.900000ns, VSS,
+ 646138.000000ns, VSS,
+ 646138.100000ns, VDD,
+ 646258.100000ns, VDD,
+ 646258.200000ns, VSS,
+ 646618.400000ns, VSS,
+ 646618.500000ns, VDD,
+ 646978.700000ns, VDD,
+ 646978.800000ns, VSS,
+ 647218.900000ns, VSS,
+ 647219.000000ns, VDD,
+ 648059.600000ns, VDD,
+ 648059.700000ns, VSS,
+ 648299.800000ns, VSS,
+ 648299.900000ns, VDD,
+ 648419.900000ns, VDD,
+ 648420.000000ns, VSS,
+ 648660.100000ns, VSS,
+ 648660.200000ns, VDD,
+ 649260.600000ns, VDD,
+ 649260.700000ns, VSS,
+ 649500.800000ns, VSS,
+ 649500.900000ns, VDD,
+ 650701.800000ns, VDD,
+ 650701.900000ns, VSS,
+ 650821.900000ns, VSS,
+ 650822.000000ns, VDD,
+ 652623.400000ns, VDD,
+ 652623.500000ns, VSS,
+ 653464.100000ns, VSS,
+ 653464.200000ns, VDD,
+ 653944.500000ns, VDD,
+ 653944.600000ns, VSS,
+ 654184.700000ns, VSS,
+ 654184.800000ns, VDD,
+ 655385.700000ns, VDD,
+ 655385.800000ns, VSS,
+ 655505.800000ns, VSS,
+ 655505.900000ns, VDD,
+ 655746.000000ns, VDD,
+ 655746.100000ns, VSS,
+ 655986.200000ns, VSS,
+ 655986.300000ns, VDD,
+ 656106.300000ns, VDD,
+ 656106.400000ns, VSS,
+ 656346.500000ns, VSS,
+ 656346.600000ns, VDD,
+ 656466.600000ns, VDD,
+ 656466.700000ns, VSS,
+ 656586.700000ns, VSS,
+ 656586.800000ns, VDD,
+ 656826.900000ns, VDD,
+ 656827.000000ns, VSS,
+ 656947.000000ns, VSS,
+ 656947.100000ns, VDD,
+ 658988.700000ns, VDD,
+ 658988.800000ns, VSS,
+ 659829.400000ns, VSS,
+ 659829.500000ns, VDD,
+ 660069.600000ns, VDD,
+ 660069.700000ns, VSS,
+ 660189.700000ns, VSS,
+ 660189.800000ns, VDD,
+ 661030.400000ns, VDD,
+ 661030.500000ns, VSS,
+ 661510.800000ns, VSS,
+ 661510.900000ns, VDD,
+ 661630.900000ns, VDD,
+ 661631.000000ns, VSS,
+ 661871.100000ns, VSS,
+ 661871.200000ns, VDD,
+ 662831.900000ns, VDD,
+ 662832.000000ns, VSS,
+ 663072.100000ns, VSS,
+ 663072.200000ns, VDD,
+ 663312.300000ns, VDD,
+ 663312.400000ns, VSS,
+ 663792.700000ns, VSS,
+ 663792.800000ns, VDD,
+ 664273.100000ns, VDD,
+ 664273.200000ns, VSS,
+ 664393.200000ns, VSS,
+ 664393.300000ns, VDD,
+ 664633.400000ns, VDD,
+ 664633.500000ns, VSS,
+ 665113.800000ns, VSS,
+ 665113.900000ns, VDD,
+ 665233.900000ns, VDD,
+ 665234.000000ns, VSS,
+ 665354.000000ns, VSS,
+ 665354.100000ns, VDD,
+ 665594.200000ns, VDD,
+ 665594.300000ns, VSS,
+ 665714.300000ns, VSS,
+ 665714.400000ns, VDD,
+ 666314.800000ns, VDD,
+ 666314.900000ns, VSS,
+ 667275.600000ns, VSS,
+ 667275.700000ns, VDD,
+ 667515.800000ns, VDD,
+ 667515.900000ns, VSS,
+ 668116.300000ns, VSS,
+ 668116.400000ns, VDD,
+ 668716.800000ns, VDD,
+ 668716.900000ns, VSS,
+ 668836.900000ns, VSS,
+ 668837.000000ns, VDD,
+ 669317.300000ns, VDD,
+ 669317.400000ns, VSS,
+ 669557.500000ns, VSS,
+ 669557.600000ns, VDD,
+ 669797.700000ns, VDD,
+ 669797.800000ns, VSS,
+ 670158.000000ns, VSS,
+ 670158.100000ns, VDD,
+ 670518.300000ns, VDD,
+ 670518.400000ns, VSS,
+ 670638.400000ns, VSS,
+ 670638.500000ns, VDD,
+ 670998.700000ns, VDD,
+ 670998.800000ns, VSS,
+ 671238.900000ns, VSS,
+ 671239.000000ns, VDD,
+ 671959.500000ns, VDD,
+ 671959.600000ns, VSS,
+ 672079.600000ns, VSS,
+ 672079.700000ns, VDD,
+ 672319.800000ns, VDD,
+ 672319.900000ns, VSS,
+ 672439.900000ns, VSS,
+ 672440.000000ns, VDD,
+ 673280.600000ns, VDD,
+ 673280.700000ns, VSS,
+ 673400.700000ns, VSS,
+ 673400.800000ns, VDD,
+ 674241.400000ns, VDD,
+ 674241.500000ns, VSS,
+ 674601.700000ns, VSS,
+ 674601.800000ns, VDD,
+ 675082.100000ns, VDD,
+ 675082.200000ns, VSS,
+ 675202.200000ns, VSS,
+ 675202.300000ns, VDD,
+ 675322.300000ns, VDD,
+ 675322.400000ns, VSS,
+ 675682.600000ns, VSS,
+ 675682.700000ns, VDD,
+ 676163.000000ns, VDD,
+ 676163.100000ns, VSS,
+ 676403.200000ns, VSS,
+ 676403.300000ns, VDD,
+ 676643.400000ns, VDD,
+ 676643.500000ns, VSS,
+ 677003.700000ns, VSS,
+ 677003.800000ns, VDD,
+ 677364.000000ns, VDD,
+ 677364.100000ns, VSS,
+ 677604.200000ns, VSS,
+ 677604.300000ns, VDD,
+ 679886.100000ns, VDD,
+ 679886.200000ns, VSS,
+ 680246.400000ns, VSS,
+ 680246.500000ns, VDD,
+ 680366.500000ns, VDD,
+ 680366.600000ns, VSS,
+ 680726.800000ns, VSS,
+ 680726.900000ns, VDD,
+ 681087.100000ns, VDD,
+ 681087.200000ns, VSS,
+ 681327.300000ns, VSS,
+ 681327.400000ns, VDD,
+ 681807.700000ns, VDD,
+ 681807.800000ns, VSS,
+ 681927.800000ns, VSS,
+ 681927.900000ns, VDD,
+ 683128.800000ns, VDD,
+ 683128.900000ns, VSS,
+ 684089.600000ns, VSS,
+ 684089.700000ns, VDD,
+ 685650.900000ns, VDD,
+ 685651.000000ns, VSS,
+ 685891.100000ns, VSS,
+ 685891.200000ns, VDD,
+ 686131.300000ns, VDD,
+ 686131.400000ns, VSS,
+ 686251.400000ns, VSS,
+ 686251.500000ns, VDD,
+ 686972.000000ns, VDD,
+ 686972.100000ns, VSS,
+ 687692.600000ns, VSS,
+ 687692.700000ns, VDD,
+ 687812.700000ns, VDD,
+ 687812.800000ns, VSS,
+ 687932.800000ns, VSS,
+ 687932.900000ns, VDD,
+ 688413.200000ns, VDD,
+ 688413.300000ns, VSS,
+ 688653.400000ns, VSS,
+ 688653.500000ns, VDD,
+ 688893.600000ns, VDD,
+ 688893.700000ns, VSS,
+ 689253.900000ns, VSS,
+ 689254.000000ns, VDD,
+ 690334.800000ns, VDD,
+ 690334.900000ns, VSS,
+ 690575.000000ns, VSS,
+ 690575.100000ns, VDD,
+ 691295.600000ns, VDD,
+ 691295.700000ns, VSS,
+ 691415.700000ns, VSS,
+ 691415.800000ns, VDD,
+ 692256.400000ns, VDD,
+ 692256.500000ns, VSS,
+ 692736.800000ns, VSS,
+ 692736.900000ns, VDD,
+ 693097.100000ns, VDD,
+ 693097.200000ns, VSS,
+ 693577.500000ns, VSS,
+ 693577.600000ns, VDD,
+ 693937.800000ns, VDD,
+ 693937.900000ns, VSS,
+ 694418.200000ns, VSS,
+ 694418.300000ns, VDD,
+ 694898.600000ns, VDD,
+ 694898.700000ns, VSS,
+ 695138.800000ns, VSS,
+ 695138.900000ns, VDD,
+ 695859.400000ns, VDD,
+ 695859.500000ns, VSS,
+ 696339.800000ns, VSS,
+ 696339.900000ns, VDD,
+ 696700.100000ns, VDD,
+ 696700.200000ns, VSS,
+ 696820.200000ns, VSS,
+ 696820.300000ns, VDD,
+ 697180.500000ns, VDD,
+ 697180.600000ns, VSS,
+ 698381.500000ns, VSS,
+ 698381.600000ns, VDD,
+ 698621.700000ns, VDD,
+ 698621.800000ns, VSS,
+ 698861.900000ns, VSS,
+ 698862.000000ns, VDD,
+ 698982.000000ns, VDD,
+ 698982.100000ns, VSS,
+ 699102.100000ns, VSS,
+ 699102.200000ns, VDD,
+ 699222.200000ns, VDD,
+ 699222.300000ns, VSS,
+ 699462.400000ns, VSS,
+ 699462.500000ns, VDD,
+ 700783.500000ns, VDD,
+ 700783.600000ns, VSS,
+ 700903.600000ns, VSS,
+ 700903.700000ns, VDD,
+ 701143.800000ns, VDD,
+ 701143.900000ns, VSS,
+ 701384.000000ns, VSS,
+ 701384.100000ns, VDD,
+ 701624.200000ns, VDD,
+ 701624.300000ns, VSS,
+ 701744.300000ns, VSS,
+ 701744.400000ns, VDD,
+ 702104.600000ns, VDD,
+ 702104.700000ns, VSS,
+ 702224.700000ns, VSS,
+ 702224.800000ns, VDD,
+ 702344.800000ns, VDD,
+ 702344.900000ns, VSS,
+ 702825.200000ns, VSS,
+ 702825.300000ns, VDD,
+ 702945.300000ns, VDD,
+ 702945.400000ns, VSS,
+ 703665.900000ns, VSS,
+ 703666.000000ns, VDD,
+ 704026.200000ns, VDD,
+ 704026.300000ns, VSS,
+ 704626.700000ns, VSS,
+ 704626.800000ns, VDD,
+ 704866.900000ns, VDD,
+ 704867.000000ns, VSS,
+ 704987.000000ns, VSS,
+ 704987.100000ns, VDD,
+ 705107.100000ns, VDD,
+ 705107.200000ns, VSS,
+ 705227.200000ns, VSS,
+ 705227.300000ns, VDD,
+ 705467.400000ns, VDD,
+ 705467.500000ns, VSS,
+ 705707.600000ns, VSS,
+ 705707.700000ns, VDD,
+ 706188.000000ns, VDD,
+ 706188.100000ns, VSS,
+ 706308.100000ns, VSS,
+ 706308.200000ns, VDD,
+ 706428.200000ns, VDD,
+ 706428.300000ns, VSS,
+ 706548.300000ns, VSS,
+ 706548.400000ns, VDD,
+ 706788.500000ns, VDD,
+ 706788.600000ns, VSS,
+ 707148.800000ns, VSS,
+ 707148.900000ns, VDD,
+ 708349.800000ns, VDD,
+ 708349.900000ns, VSS,
+ 708590.000000ns, VSS,
+ 708590.100000ns, VDD,
+ 708950.300000ns, VDD,
+ 708950.400000ns, VSS,
+ 709070.400000ns, VSS,
+ 709070.500000ns, VDD,
+ 710031.200000ns, VDD,
+ 710031.300000ns, VSS,
+ 710391.500000ns, VSS,
+ 710391.600000ns, VDD,
+ 710751.800000ns, VDD,
+ 710751.900000ns, VSS,
+ 711232.200000ns, VSS,
+ 711232.300000ns, VDD,
+ 711832.700000ns, VDD,
+ 711832.800000ns, VSS,
+ 712072.900000ns, VSS,
+ 712073.000000ns, VDD,
+ 713033.700000ns, VDD,
+ 713033.800000ns, VSS,
+ 714114.600000ns, VSS,
+ 714114.700000ns, VDD,
+ 714474.900000ns, VDD,
+ 714475.000000ns, VSS,
+ 714715.100000ns, VSS,
+ 714715.200000ns, VDD,
+ 715075.400000ns, VDD,
+ 715075.500000ns, VSS,
+ 715195.500000ns, VSS,
+ 715195.600000ns, VDD,
+ 715315.600000ns, VDD,
+ 715315.700000ns, VSS,
+ 715435.700000ns, VSS,
+ 715435.800000ns, VDD,
+ 715916.100000ns, VDD,
+ 715916.200000ns, VSS,
+ 716396.500000ns, VSS,
+ 716396.600000ns, VDD,
+ 716636.700000ns, VDD,
+ 716636.800000ns, VSS,
+ 717237.200000ns, VSS,
+ 717237.300000ns, VDD,
+ 717717.600000ns, VDD,
+ 717717.700000ns, VSS,
+ 718438.200000ns, VSS,
+ 718438.300000ns, VDD,
+ 718918.600000ns, VDD,
+ 718918.700000ns, VSS,
+ 719278.900000ns, VSS,
+ 719279.000000ns, VDD,
+ 719519.100000ns, VDD,
+ 719519.200000ns, VSS,
+ 719639.200000ns, VSS,
+ 719639.300000ns, VDD,
+ 719759.300000ns, VDD,
+ 719759.400000ns, VSS,
+ 720359.800000ns, VSS,
+ 720359.900000ns, VDD,
+ 720479.900000ns, VDD,
+ 720480.000000ns, VSS,
+ 720840.200000ns, VSS,
+ 720840.300000ns, VDD,
+ 722041.200000ns, VDD,
+ 722041.300000ns, VSS,
+ 722281.400000ns, VSS,
+ 722281.500000ns, VDD,
+ 722521.600000ns, VDD,
+ 722521.700000ns, VSS,
+ 722761.800000ns, VSS,
+ 722761.900000ns, VDD,
+ 722881.900000ns, VDD,
+ 722882.000000ns, VSS,
+ 723002.000000ns, VSS,
+ 723002.100000ns, VDD,
+ 723362.300000ns, VDD,
+ 723362.400000ns, VSS,
+ 723722.600000ns, VSS,
+ 723722.700000ns, VDD,
+ 724923.600000ns, VDD,
+ 724923.700000ns, VSS,
+ 725043.700000ns, VSS,
+ 725043.800000ns, VDD,
+ 726004.500000ns, VDD,
+ 726004.600000ns, VSS,
+ 726484.900000ns, VSS,
+ 726485.000000ns, VDD,
+ 726605.000000ns, VDD,
+ 726605.100000ns, VSS,
+ 726965.300000ns, VSS,
+ 726965.400000ns, VDD,
+ 727565.800000ns, VDD,
+ 727565.900000ns, VSS,
+ 727685.900000ns, VSS,
+ 727686.000000ns, VDD,
+ 727806.000000ns, VDD,
+ 727806.100000ns, VSS,
+ 728166.300000ns, VSS,
+ 728166.400000ns, VDD,
+ 729727.600000ns, VDD,
+ 729727.700000ns, VSS,
+ 729967.800000ns, VSS,
+ 729967.900000ns, VDD,
+ 730208.000000ns, VDD,
+ 730208.100000ns, VSS,
+ 730808.500000ns, VSS,
+ 730808.600000ns, VDD,
+ 731168.800000ns, VDD,
+ 731168.900000ns, VSS,
+ 732009.500000ns, VSS,
+ 732009.600000ns, VDD,
+ 732249.700000ns, VDD,
+ 732249.800000ns, VSS,
+ 732369.800000ns, VSS,
+ 732369.900000ns, VDD,
+ 732489.900000ns, VDD,
+ 732490.000000ns, VSS,
+ 732610.000000ns, VSS,
+ 732610.100000ns, VDD,
+ 732970.300000ns, VDD,
+ 732970.400000ns, VSS,
+ 733330.600000ns, VSS,
+ 733330.700000ns, VDD,
+ 733450.700000ns, VDD,
+ 733450.800000ns, VSS,
+ 733690.900000ns, VSS,
+ 733691.000000ns, VDD,
+ 734051.200000ns, VDD,
+ 734051.300000ns, VSS,
+ 734411.500000ns, VSS,
+ 734411.600000ns, VDD,
+ 734651.700000ns, VDD,
+ 734651.800000ns, VSS,
+ 734771.800000ns, VSS,
+ 734771.900000ns, VDD,
+ 735012.000000ns, VDD,
+ 735012.100000ns, VSS,
+ 735612.500000ns, VSS,
+ 735612.600000ns, VDD,
+ 737894.400000ns, VDD,
+ 737894.500000ns, VSS,
+ 738254.700000ns, VSS,
+ 738254.800000ns, VDD,
+ 739816.000000ns, VDD,
+ 739816.100000ns, VSS,
+ 740416.500000ns, VSS,
+ 740416.600000ns, VDD,
+ 740776.800000ns, VDD,
+ 740776.900000ns, VSS,
+ 741017.000000ns, VSS,
+ 741017.100000ns, VDD,
+ 741497.400000ns, VDD,
+ 741497.500000ns, VSS,
+ 741857.700000ns, VSS,
+ 741857.800000ns, VDD,
+ 742218.000000ns, VDD,
+ 742218.100000ns, VSS,
+ 742458.200000ns, VSS,
+ 742458.300000ns, VDD,
+ 743058.700000ns, VDD,
+ 743058.800000ns, VSS,
+ 743779.300000ns, VSS,
+ 743779.400000ns, VDD,
+ 744259.700000ns, VDD,
+ 744259.800000ns, VSS,
+ 744379.800000ns, VSS,
+ 744379.900000ns, VDD,
+ 744499.900000ns, VDD,
+ 744500.000000ns, VSS,
+ 744980.300000ns, VSS,
+ 744980.400000ns, VDD,
+ 746301.400000ns, VDD,
+ 746301.500000ns, VSS,
+ 746421.500000ns, VSS,
+ 746421.600000ns, VDD,
+ 746541.600000ns, VDD,
+ 746541.700000ns, VSS,
+ 746781.800000ns, VSS,
+ 746781.900000ns, VDD,
+ 746901.900000ns, VDD,
+ 746902.000000ns, VSS,
+ 747262.200000ns, VSS,
+ 747262.300000ns, VDD,
+ 748583.300000ns, VDD,
+ 748583.400000ns, VSS,
+ 748943.600000ns, VSS,
+ 748943.700000ns, VDD,
+ 749063.700000ns, VDD,
+ 749063.800000ns, VSS,
+ 749303.900000ns, VSS,
+ 749304.000000ns, VDD,
+ 749424.000000ns, VDD,
+ 749424.100000ns, VSS,
+ 749784.300000ns, VSS,
+ 749784.400000ns, VDD,
+ 750024.500000ns, VDD,
+ 750024.600000ns, VSS,
+ 750144.600000ns, VSS,
+ 750144.700000ns, VDD,
+ 750625.000000ns, VDD,
+ 750625.100000ns, VSS,
+ 751705.900000ns, VSS,
+ 751706.000000ns, VDD,
+ 751946.100000ns, VDD,
+ 751946.200000ns, VSS,
+ 752066.200000ns, VSS,
+ 752066.300000ns, VDD,
+ 752426.500000ns, VDD,
+ 752426.600000ns, VSS,
+ 753027.000000ns, VSS,
+ 753027.100000ns, VDD,
+ 753507.400000ns, VDD,
+ 753507.500000ns, VSS,
+ 753747.600000ns, VSS,
+ 753747.700000ns, VDD,
+ 753867.700000ns, VDD,
+ 753867.800000ns, VSS,
+ 753987.800000ns, VSS,
+ 753987.900000ns, VDD,
+ 754107.900000ns, VDD,
+ 754108.000000ns, VSS,
+ 754468.200000ns, VSS,
+ 754468.300000ns, VDD,
+ 754828.500000ns, VDD,
+ 754828.600000ns, VSS,
+ 755549.100000ns, VSS,
+ 755549.200000ns, VDD,
+ 755789.300000ns, VDD,
+ 755789.400000ns, VSS,
+ 755909.400000ns, VSS,
+ 755909.500000ns, VDD,
+ 756029.500000ns, VDD,
+ 756029.600000ns, VSS,
+ 756750.100000ns, VSS,
+ 756750.200000ns, VDD,
+ 756870.200000ns, VDD,
+ 756870.300000ns, VSS,
+ 756990.300000ns, VSS,
+ 756990.400000ns, VDD,
+ 757230.500000ns, VDD,
+ 757230.600000ns, VSS,
+ 757951.100000ns, VSS,
+ 757951.200000ns, VDD,
+ 758191.300000ns, VDD,
+ 758191.400000ns, VSS,
+ 758431.500000ns, VSS,
+ 758431.600000ns, VDD,
+ 759152.100000ns, VDD,
+ 759152.200000ns, VSS,
+ 759392.300000ns, VSS,
+ 759392.400000ns, VDD,
+ 759512.400000ns, VDD,
+ 759512.500000ns, VSS,
+ 759872.700000ns, VSS,
+ 759872.800000ns, VDD,
+ 760473.200000ns, VDD,
+ 760473.300000ns, VSS,
+ 761073.700000ns, VSS,
+ 761073.800000ns, VDD,
+ 761434.000000ns, VDD,
+ 761434.100000ns, VSS,
+ 761914.400000ns, VSS,
+ 761914.500000ns, VDD,
+ 762394.800000ns, VDD,
+ 762394.900000ns, VSS,
+ 762995.300000ns, VSS,
+ 762995.400000ns, VDD,
+ 763355.600000ns, VDD,
+ 763355.700000ns, VSS,
+ 763595.800000ns, VSS,
+ 763595.900000ns, VDD,
+ 764436.500000ns, VDD,
+ 764436.600000ns, VSS,
+ 764796.800000ns, VSS,
+ 764796.900000ns, VDD,
+ 765037.000000ns, VDD,
+ 765037.100000ns, VSS,
+ 765637.500000ns, VSS,
+ 765637.600000ns, VDD,
+ 765757.600000ns, VDD,
+ 765757.700000ns, VSS,
+ 765877.700000ns, VSS,
+ 765877.800000ns, VDD,
+ 766718.400000ns, VDD,
+ 766718.500000ns, VSS,
+ 766838.500000ns, VSS,
+ 766838.600000ns, VDD,
+ 767318.900000ns, VDD,
+ 767319.000000ns, VSS,
+ 767679.200000ns, VSS,
+ 767679.300000ns, VDD,
+ 768279.700000ns, VDD,
+ 768279.800000ns, VSS,
+ 768399.800000ns, VSS,
+ 768399.900000ns, VDD,
+ 768760.100000ns, VDD,
+ 768760.200000ns, VSS,
+ 769120.400000ns, VSS,
+ 769120.500000ns, VDD,
+ 769961.100000ns, VDD,
+ 769961.200000ns, VSS,
+ 770081.200000ns, VSS,
+ 770081.300000ns, VDD,
+ 770441.500000ns, VDD,
+ 770441.600000ns, VSS,
+ 770921.900000ns, VSS,
+ 770922.000000ns, VDD,
+ 771282.200000ns, VDD,
+ 771282.300000ns, VSS,
+ 771402.300000ns, VSS,
+ 771402.400000ns, VDD,
+ 771642.500000ns, VDD,
+ 771642.600000ns, VSS,
+ 771762.600000ns, VSS,
+ 771762.700000ns, VDD,
+ 772122.900000ns, VDD,
+ 772123.000000ns, VSS,
+ 772723.400000ns, VSS,
+ 772723.500000ns, VDD,
+ 773684.200000ns, VDD,
+ 773684.300000ns, VSS,
+ 773804.300000ns, VSS,
+ 773804.400000ns, VDD,
+ 774164.600000ns, VDD,
+ 774164.700000ns, VSS,
+ 774404.800000ns, VSS,
+ 774404.900000ns, VDD,
+ 775245.500000ns, VDD,
+ 775245.600000ns, VSS,
+ 775365.600000ns, VSS,
+ 775365.700000ns, VDD,
+ 775605.800000ns, VDD,
+ 775605.900000ns, VSS,
+ 776086.200000ns, VSS,
+ 776086.300000ns, VDD,
+ 776446.500000ns, VDD,
+ 776446.600000ns, VSS,
+ 776566.600000ns, VSS,
+ 776566.700000ns, VDD,
+ 777167.100000ns, VDD,
+ 777167.200000ns, VSS,
+ 777527.400000ns, VSS,
+ 777527.500000ns, VDD,
+ 777647.500000ns, VDD,
+ 777647.600000ns, VSS,
+ 777887.700000ns, VSS,
+ 777887.800000ns, VDD,
+ 778127.900000ns, VDD,
+ 778128.000000ns, VSS,
+ 779328.900000ns, VSS,
+ 779329.000000ns, VDD,
+ 781971.100000ns, VDD,
+ 781971.200000ns, VSS,
+ 782211.300000ns, VSS,
+ 782211.400000ns, VDD,
+ 782571.600000ns, VDD,
+ 782571.700000ns, VSS,
+ 782691.700000ns, VSS,
+ 782691.800000ns, VDD,
+ 783292.200000ns, VDD,
+ 783292.300000ns, VSS,
+ 783532.400000ns, VSS,
+ 783532.500000ns, VDD,
+ 785093.700000ns, VDD,
+ 785093.800000ns, VSS,
+ 785333.900000ns, VSS,
+ 785334.000000ns, VDD,
+ 786534.900000ns, VDD,
+ 786535.000000ns, VSS,
+ 786655.000000ns, VSS,
+ 786655.100000ns, VDD,
+ 786775.100000ns, VDD,
+ 786775.200000ns, VSS,
+ 787015.300000ns, VSS,
+ 787015.400000ns, VDD,
+ 787135.400000ns, VDD,
+ 787135.500000ns, VSS,
+ 787255.500000ns, VSS,
+ 787255.600000ns, VDD,
+ 788216.300000ns, VDD,
+ 788216.400000ns, VSS,
+ 788456.500000ns, VSS,
+ 788456.600000ns, VDD,
+ 788576.600000ns, VDD,
+ 788576.700000ns, VSS,
+ 788936.900000ns, VSS,
+ 788937.000000ns, VDD,
+ 789057.000000ns, VDD,
+ 789057.100000ns, VSS,
+ 789657.500000ns, VSS,
+ 789657.600000ns, VDD,
+ 790017.800000ns, VDD,
+ 790017.900000ns, VSS,
+ 790258.000000ns, VSS,
+ 790258.100000ns, VDD,
+ 790618.300000ns, VDD,
+ 790618.400000ns, VSS,
+ 790978.600000ns, VSS,
+ 790978.700000ns, VDD,
+ 791819.300000ns, VDD,
+ 791819.400000ns, VSS,
+ 792059.500000ns, VSS,
+ 792059.600000ns, VDD,
+ 792419.800000ns, VDD,
+ 792419.900000ns, VSS,
+ 792780.100000ns, VSS,
+ 792780.200000ns, VDD,
+ 792900.200000ns, VDD,
+ 792900.300000ns, VSS,
+ 793020.300000ns, VSS,
+ 793020.400000ns, VDD,
+ 793140.400000ns, VDD,
+ 793140.500000ns, VSS,
+ 793260.500000ns, VSS,
+ 793260.600000ns, VDD,
+ 793380.600000ns, VDD,
+ 793380.700000ns, VSS,
+ 793861.000000ns, VSS,
+ 793861.100000ns, VDD,
+ 795182.100000ns, VDD,
+ 795182.200000ns, VSS,
+ 795422.300000ns, VSS,
+ 795422.400000ns, VDD,
+ 795782.600000ns, VDD,
+ 795782.700000ns, VSS,
+ 796142.900000ns, VSS,
+ 796143.000000ns, VDD,
+ 796503.200000ns, VDD,
+ 796503.300000ns, VSS,
+ 796623.300000ns, VSS,
+ 796623.400000ns, VDD,
+ 796743.400000ns, VDD,
+ 796743.500000ns, VSS,
+ 796863.500000ns, VSS,
+ 796863.600000ns, VDD,
+ 797584.100000ns, VDD,
+ 797584.200000ns, VSS,
+ 797824.300000ns, VSS,
+ 797824.400000ns, VDD,
+ 798304.700000ns, VDD,
+ 798304.800000ns, VSS,
+ 798544.900000ns, VSS,
+ 798545.000000ns, VDD,
+ 798665.000000ns, VDD,
+ 798665.100000ns, VSS,
+ 799145.400000ns, VSS,
+ 799145.500000ns, VDD,
+ 799505.700000ns, VDD,
+ 799505.800000ns, VSS,
+ 799866.000000ns, VSS,
+ 799866.100000ns, VDD,
+ 800826.800000ns, VDD,
+ 800826.900000ns, VSS,
+ 801067.000000ns, VSS,
+ 801067.100000ns, VDD,
+ 801187.100000ns, VDD,
+ 801187.200000ns, VSS,
+ 802268.000000ns, VSS,
+ 802268.100000ns, VDD,
+ 803589.100000ns, VDD,
+ 803589.200000ns, VSS,
+ 803709.200000ns, VSS,
+ 803709.300000ns, VDD,
+ 803829.300000ns, VDD,
+ 803829.400000ns, VSS,
+ 804069.500000ns, VSS,
+ 804069.600000ns, VDD,
+ 805030.300000ns, VDD,
+ 805030.400000ns, VSS,
+ 805750.900000ns, VSS,
+ 805751.000000ns, VDD,
+ 806231.300000ns, VDD,
+ 806231.400000ns, VSS,
+ 806351.400000ns, VSS,
+ 806351.500000ns, VDD,
+ 806711.700000ns, VDD,
+ 806711.800000ns, VSS,
+ 806951.900000ns, VSS,
+ 806952.000000ns, VDD,
+ 807672.500000ns, VDD,
+ 807672.600000ns, VSS,
+ 807792.600000ns, VSS,
+ 807792.700000ns, VDD,
+ 807912.700000ns, VDD,
+ 807912.800000ns, VSS,
+ 808393.100000ns, VSS,
+ 808393.200000ns, VDD,
+ 808633.300000ns, VDD,
+ 808633.400000ns, VSS,
+ 809353.900000ns, VSS,
+ 809354.000000ns, VDD,
+ 809594.100000ns, VDD,
+ 809594.200000ns, VSS,
+ 810074.500000ns, VSS,
+ 810074.600000ns, VDD,
+ 810554.900000ns, VDD,
+ 810555.000000ns, VSS,
+ 810915.200000ns, VSS,
+ 810915.300000ns, VDD,
+ 811275.500000ns, VDD,
+ 811275.600000ns, VSS,
+ 811755.900000ns, VSS,
+ 811756.000000ns, VDD,
+ 812116.200000ns, VDD,
+ 812116.300000ns, VSS,
+ 812356.400000ns, VSS,
+ 812356.500000ns, VDD,
+ 812596.600000ns, VDD,
+ 812596.700000ns, VSS,
+ 812836.800000ns, VSS,
+ 812836.900000ns, VDD,
+ 813197.100000ns, VDD,
+ 813197.200000ns, VSS,
+ 813317.200000ns, VSS,
+ 813317.300000ns, VDD,
+ 813677.500000ns, VDD,
+ 813677.600000ns, VSS,
+ 813797.600000ns, VSS,
+ 813797.700000ns, VDD,
+ 814157.900000ns, VDD,
+ 814158.000000ns, VSS,
+ 814278.000000ns, VSS,
+ 814278.100000ns, VDD,
+ 815118.700000ns, VDD,
+ 815118.800000ns, VSS,
+ 815238.800000ns, VSS,
+ 815238.900000ns, VDD,
+ 815358.900000ns, VDD,
+ 815359.000000ns, VSS,
+ 815479.000000ns, VSS,
+ 815479.100000ns, VDD,
+ 815839.300000ns, VDD,
+ 815839.400000ns, VSS,
+ 816559.900000ns, VSS,
+ 816560.000000ns, VDD,
+ 816680.000000ns, VDD,
+ 816680.100000ns, VSS,
+ 817040.300000ns, VSS,
+ 817040.400000ns, VDD,
+ 817881.000000ns, VDD,
+ 817881.100000ns, VSS,
+ 818121.200000ns, VSS,
+ 818121.300000ns, VDD,
+ 818481.500000ns, VDD,
+ 818481.600000ns, VSS,
+ 818601.600000ns, VSS,
+ 818601.700000ns, VDD,
+ 819322.200000ns, VDD,
+ 819322.300000ns, VSS,
+ 819442.300000ns, VSS,
+ 819442.400000ns, VDD,
+ 819922.700000ns, VDD,
+ 819922.800000ns, VSS,
+ 820042.800000ns, VSS,
+ 820042.900000ns, VDD,
+ 820883.500000ns, VDD,
+ 820883.600000ns, VSS,
+ 821363.900000ns, VSS,
+ 821364.000000ns, VDD,
+ 821724.200000ns, VDD,
+ 821724.300000ns, VSS,
+ 822204.600000ns, VSS,
+ 822204.700000ns, VDD,
+ 822444.800000ns, VDD,
+ 822444.900000ns, VSS,
+ 822685.000000ns, VSS,
+ 822685.100000ns, VDD,
+ 823045.300000ns, VDD,
+ 823045.400000ns, VSS,
+ 823525.700000ns, VSS,
+ 823525.800000ns, VDD,
+ 823886.000000ns, VDD,
+ 823886.100000ns, VSS,
+ 824126.200000ns, VSS,
+ 824126.300000ns, VDD,
+ 824246.300000ns, VDD,
+ 824246.400000ns, VSS,
+ 824606.600000ns, VSS,
+ 824606.700000ns, VDD,
+ 824966.900000ns, VDD,
+ 824967.000000ns, VSS,
+ 825087.000000ns, VSS,
+ 825087.100000ns, VDD,
+ 825447.300000ns, VDD,
+ 825447.400000ns, VSS,
+ 825567.400000ns, VSS,
+ 825567.500000ns, VDD,
+ 825687.500000ns, VDD,
+ 825687.600000ns, VSS,
+ 825807.600000ns, VSS,
+ 825807.700000ns, VDD,
+ 826167.900000ns, VDD,
+ 826168.000000ns, VSS,
+ 826528.200000ns, VSS,
+ 826528.300000ns, VDD,
+ 826768.400000ns, VDD,
+ 826768.500000ns, VSS,
+ 827248.800000ns, VSS,
+ 827248.900000ns, VDD,
+ 829410.600000ns, VDD,
+ 829410.700000ns, VSS,
+ 830251.300000ns, VSS,
+ 830251.400000ns, VDD,
+ 831572.400000ns, VDD,
+ 831572.500000ns, VSS,
+ 831812.600000ns, VSS,
+ 831812.700000ns, VDD,
+ 832052.800000ns, VDD,
+ 832052.900000ns, VSS,
+ 832413.100000ns, VSS,
+ 832413.200000ns, VDD,
+ 832653.300000ns, VDD,
+ 832653.400000ns, VSS,
+ 833013.600000ns, VSS,
+ 833013.700000ns, VDD,
+ 834094.500000ns, VDD,
+ 834094.600000ns, VSS,
+ 834214.600000ns, VSS,
+ 834214.700000ns, VDD,
+ 834334.700000ns, VDD,
+ 834334.800000ns, VSS,
+ 834574.900000ns, VSS,
+ 834575.000000ns, VDD,
+ 834815.100000ns, VDD,
+ 834815.200000ns, VSS,
+ 835055.300000ns, VSS,
+ 835055.400000ns, VDD,
+ 835295.500000ns, VDD,
+ 835295.600000ns, VSS,
+ 835655.800000ns, VSS,
+ 835655.900000ns, VDD,
+ 836136.200000ns, VDD,
+ 836136.300000ns, VSS,
+ 836496.500000ns, VSS,
+ 836496.600000ns, VDD,
+ 836736.700000ns, VDD,
+ 836736.800000ns, VSS,
+ 836856.800000ns, VSS,
+ 836856.900000ns, VDD,
+ 836976.900000ns, VDD,
+ 836977.000000ns, VSS,
+ 837217.100000ns, VSS,
+ 837217.200000ns, VDD,
+ 838177.900000ns, VDD,
+ 838178.000000ns, VSS,
+ 838298.000000ns, VSS,
+ 838298.100000ns, VDD,
+ 839138.700000ns, VDD,
+ 839138.800000ns, VSS,
+ 839258.800000ns, VSS,
+ 839258.900000ns, VDD,
+ 839619.100000ns, VDD,
+ 839619.200000ns, VSS,
+ 841180.400000ns, VSS,
+ 841180.500000ns, VDD,
+ 841901.000000ns, VDD,
+ 841901.100000ns, VSS,
+ 842621.600000ns, VSS,
+ 842621.700000ns, VDD,
+ 843822.600000ns, VDD,
+ 843822.700000ns, VSS,
+ 844182.900000ns, VSS,
+ 844183.000000ns, VDD,
+ 844783.400000ns, VDD,
+ 844783.500000ns, VSS,
+ 845143.700000ns, VSS,
+ 845143.800000ns, VDD,
+ 845984.400000ns, VDD,
+ 845984.500000ns, VSS,
+ 846705.000000ns, VSS,
+ 846705.100000ns, VDD,
+ 847065.300000ns, VDD,
+ 847065.400000ns, VSS,
+ 847425.600000ns, VSS,
+ 847425.700000ns, VDD,
+ 847665.800000ns, VDD,
+ 847665.900000ns, VSS,
+ 847785.900000ns, VSS,
+ 847786.000000ns, VDD,
+ 848026.100000ns, VDD,
+ 848026.200000ns, VSS,
+ 848266.300000ns, VSS,
+ 848266.400000ns, VDD,
+ 849467.300000ns, VDD,
+ 849467.400000ns, VSS,
+ 849587.400000ns, VSS,
+ 849587.500000ns, VDD,
+ 850187.900000ns, VDD,
+ 850188.000000ns, VSS,
+ 850668.300000ns, VSS,
+ 850668.400000ns, VDD,
+ 851028.600000ns, VDD,
+ 851028.700000ns, VSS,
+ 851268.800000ns, VSS,
+ 851268.900000ns, VDD,
+ 852830.100000ns, VDD,
+ 852830.200000ns, VSS,
+ 853070.300000ns, VSS,
+ 853070.400000ns, VDD,
+ 853550.700000ns, VDD,
+ 853550.800000ns, VSS,
+ 853911.000000ns, VSS,
+ 853911.100000ns, VDD,
+ 854511.500000ns, VDD,
+ 854511.600000ns, VSS,
+ 854991.900000ns, VSS,
+ 854992.000000ns, VDD,
+ 855352.200000ns, VDD,
+ 855352.300000ns, VSS,
+ 855952.700000ns, VSS,
+ 855952.800000ns, VDD,
+ 856313.000000ns, VDD,
+ 856313.100000ns, VSS,
+ 856913.500000ns, VSS,
+ 856913.600000ns, VDD,
+ 857033.600000ns, VDD,
+ 857033.700000ns, VSS,
+ 857514.000000ns, VSS,
+ 857514.100000ns, VDD,
+ 857994.400000ns, VDD,
+ 857994.500000ns, VSS,
+ 858234.600000ns, VSS,
+ 858234.700000ns, VDD,
+ 859435.600000ns, VDD,
+ 859435.700000ns, VSS,
+ 859555.700000ns, VSS,
+ 859555.800000ns, VDD,
+ 859916.000000ns, VDD,
+ 859916.100000ns, VSS,
+ 860276.300000ns, VSS,
+ 860276.400000ns, VDD,
+ 860636.600000ns, VDD,
+ 860636.700000ns, VSS,
+ 860996.900000ns, VSS,
+ 860997.000000ns, VDD,
+ 861357.200000ns, VDD,
+ 861357.300000ns, VSS,
+ 861597.400000ns, VSS,
+ 861597.500000ns, VDD,
+ 862077.800000ns, VDD,
+ 862077.900000ns, VSS,
+ 862197.900000ns, VSS,
+ 862198.000000ns, VDD,
+ 862438.100000ns, VDD,
+ 862438.200000ns, VSS,
+ 862678.300000ns, VSS,
+ 862678.400000ns, VDD,
+ 862798.400000ns, VDD,
+ 862798.500000ns, VSS,
+ 863158.700000ns, VSS,
+ 863158.800000ns, VDD,
+ 863519.000000ns, VDD,
+ 863519.100000ns, VSS,
+ 863879.300000ns, VSS,
+ 863879.400000ns, VDD,
+ 864599.900000ns, VDD,
+ 864600.000000ns, VSS,
+ 864720.000000ns, VSS,
+ 864720.100000ns, VDD,
+ 864840.100000ns, VDD,
+ 864840.200000ns, VSS,
+ 864960.200000ns, VSS,
+ 864960.300000ns, VDD,
+ 865320.500000ns, VDD,
+ 865320.600000ns, VSS,
+ 865680.800000ns, VSS,
+ 865680.900000ns, VDD,
+ 866041.100000ns, VDD,
+ 866041.200000ns, VSS,
+ 866401.400000ns, VSS,
+ 866401.500000ns, VDD,
+ 866761.700000ns, VDD,
+ 866761.800000ns, VSS,
+ 867242.100000ns, VSS,
+ 867242.200000ns, VDD,
+ 867362.200000ns, VDD,
+ 867362.300000ns, VSS,
+ 867842.600000ns, VSS,
+ 867842.700000ns, VDD,
+ 867962.700000ns, VDD,
+ 867962.800000ns, VSS,
+ 868202.900000ns, VSS,
+ 868203.000000ns, VDD,
+ 869403.900000ns, VDD,
+ 869404.000000ns, VSS,
+ 869764.200000ns, VSS,
+ 869764.300000ns, VDD,
+ 870604.900000ns, VDD,
+ 870605.000000ns, VSS,
+ 870965.200000ns, VSS,
+ 870965.300000ns, VDD,
+ 872166.200000ns, VDD,
+ 872166.300000ns, VSS,
+ 872886.800000ns, VSS,
+ 872886.900000ns, VDD,
+ 873127.000000ns, VDD,
+ 873127.100000ns, VSS,
+ 873607.400000ns, VSS,
+ 873607.500000ns, VDD,
+ 874328.000000ns, VDD,
+ 874328.100000ns, VSS,
+ 875529.000000ns, VSS,
+ 875529.100000ns, VDD,
+ 876249.600000ns, VDD,
+ 876249.700000ns, VSS,
+ 876369.700000ns, VSS,
+ 876369.800000ns, VDD,
+ 876850.100000ns, VDD,
+ 876850.200000ns, VSS,
+ 876970.200000ns, VSS,
+ 876970.300000ns, VDD,
+ 877090.300000ns, VDD,
+ 877090.400000ns, VSS,
+ 877450.600000ns, VSS,
+ 877450.700000ns, VDD,
+ 877931.000000ns, VDD,
+ 877931.100000ns, VSS,
+ 878171.200000ns, VSS,
+ 878171.300000ns, VDD,
+ 878651.600000ns, VDD,
+ 878651.700000ns, VSS,
+ 878891.800000ns, VSS,
+ 878891.900000ns, VDD,
+ 879372.200000ns, VDD,
+ 879372.300000ns, VSS,
+ 879972.700000ns, VSS,
+ 879972.800000ns, VDD,
+ 880333.000000ns, VDD,
+ 880333.100000ns, VSS,
+ 880453.100000ns, VSS,
+ 880453.200000ns, VDD,
+ 880573.200000ns, VDD,
+ 880573.300000ns, VSS,
+ 880813.400000ns, VSS,
+ 880813.500000ns, VDD,
+ 881173.700000ns, VDD,
+ 881173.800000ns, VSS,
+ 881293.800000ns, VSS,
+ 881293.900000ns, VDD,
+ 881534.000000ns, VDD,
+ 881534.100000ns, VSS,
+ 881654.100000ns, VSS,
+ 881654.200000ns, VDD,
+ 881894.300000ns, VDD,
+ 881894.400000ns, VSS,
+ 882014.400000ns, VSS,
+ 882014.500000ns, VDD,
+ 882374.700000ns, VDD,
+ 882374.800000ns, VSS,
+ 882614.900000ns, VSS,
+ 882615.000000ns, VDD,
+ 882735.000000ns, VDD,
+ 882735.100000ns, VSS,
+ 882855.100000ns, VSS,
+ 882855.200000ns, VDD,
+ 883215.400000ns, VDD,
+ 883215.500000ns, VSS,
+ 883575.700000ns, VSS,
+ 883575.800000ns, VDD,
+ 884296.300000ns, VDD,
+ 884296.400000ns, VSS,
+ 884776.700000ns, VSS,
+ 884776.800000ns, VDD,
+ 885737.500000ns, VDD,
+ 885737.600000ns, VSS,
+ 885857.600000ns, VSS,
+ 885857.700000ns, VDD,
+ 886217.900000ns, VDD,
+ 886218.000000ns, VSS,
+ 886338.000000ns, VSS,
+ 886338.100000ns, VDD,
+ 886458.100000ns, VDD,
+ 886458.200000ns, VSS,
+ 886578.200000ns, VSS,
+ 886578.300000ns, VDD,
+ 887058.600000ns, VDD,
+ 887058.700000ns, VSS,
+ 887298.800000ns, VSS,
+ 887298.900000ns, VDD,
+ 888019.400000ns, VDD,
+ 888019.500000ns, VSS,
+ 888259.600000ns, VSS,
+ 888259.700000ns, VDD,
+ 888619.900000ns, VDD,
+ 888620.000000ns, VSS,
+ 888980.200000ns, VSS,
+ 888980.300000ns, VDD,
+ 889220.400000ns, VDD,
+ 889220.500000ns, VSS,
+ 889580.700000ns, VSS,
+ 889580.800000ns, VDD,
+ 890061.100000ns, VDD,
+ 890061.200000ns, VSS,
+ 890421.400000ns, VSS,
+ 890421.500000ns, VDD,
+ 890661.600000ns, VDD,
+ 890661.700000ns, VSS,
+ 891021.900000ns, VSS,
+ 891022.000000ns, VDD,
+ 891382.200000ns, VDD,
+ 891382.300000ns, VSS,
+ 891862.600000ns, VSS,
+ 891862.700000ns, VDD,
+ 892343.000000ns, VDD,
+ 892343.100000ns, VSS,
+ 892583.200000ns, VSS,
+ 892583.300000ns, VDD,
+ 892823.400000ns, VDD,
+ 892823.500000ns, VSS,
+ 893423.900000ns, VSS,
+ 893424.000000ns, VDD,
+ 893544.000000ns, VDD,
+ 893544.100000ns, VSS,
+ 894024.400000ns, VSS,
+ 894024.500000ns, VDD,
+ 894384.700000ns, VDD,
+ 894384.800000ns, VSS,
+ 894745.000000ns, VSS,
+ 894745.100000ns, VDD,
+ 894865.100000ns, VDD,
+ 894865.200000ns, VSS,
+ 894985.200000ns, VSS,
+ 894985.300000ns, VDD,
+ 895225.400000ns, VDD,
+ 895225.500000ns, VSS,
+ 895345.500000ns, VSS,
+ 895345.600000ns, VDD,
+ 895465.600000ns, VDD,
+ 895465.700000ns, VSS,
+ 895585.700000ns, VSS,
+ 895585.800000ns, VDD,
+ 896306.300000ns, VDD,
+ 896306.400000ns, VSS,
+ 896426.400000ns, VSS,
+ 896426.500000ns, VDD,
+ 897507.300000ns, VDD,
+ 897507.400000ns, VSS,
+ 897867.600000ns, VSS,
+ 897867.700000ns, VDD,
+ 898828.400000ns, VDD,
+ 898828.500000ns, VSS,
+ 899068.600000ns, VSS,
+ 899068.700000ns, VDD,
+ 899428.900000ns, VDD,
+ 899429.000000ns, VSS,
+ 899909.300000ns, VSS,
+ 899909.400000ns, VDD,
+ 900269.600000ns, VDD,
+ 900269.700000ns, VSS,
+ 900750.000000ns, VSS,
+ 900750.100000ns, VDD,
+ 901110.300000ns, VDD,
+ 901110.400000ns, VSS,
+ 901590.700000ns, VSS,
+ 901590.800000ns, VDD,
+ 901951.000000ns, VDD,
+ 901951.100000ns, VSS,
+ 902791.700000ns, VSS,
+ 902791.800000ns, VDD,
+ 902911.800000ns, VDD,
+ 902911.900000ns, VSS,
+ 903031.900000ns, VSS,
+ 903032.000000ns, VDD,
+ 903392.200000ns, VDD,
+ 903392.300000ns, VSS,
+ 903512.300000ns, VSS,
+ 903512.400000ns, VDD,
+ 903752.500000ns, VDD,
+ 903752.600000ns, VSS,
+ 903872.600000ns, VSS,
+ 903872.700000ns, VDD,
+ 903992.700000ns, VDD,
+ 903992.800000ns, VSS,
+ 904232.900000ns, VSS,
+ 904233.000000ns, VDD,
+ 904713.300000ns, VDD,
+ 904713.400000ns, VSS,
+ 905193.700000ns, VSS,
+ 905193.800000ns, VDD,
+ 905554.000000ns, VDD,
+ 905554.100000ns, VSS,
+ 905794.200000ns, VSS,
+ 905794.300000ns, VDD,
+ 906154.500000ns, VDD,
+ 906154.600000ns, VSS,
+ 906514.800000ns, VSS,
+ 906514.900000ns, VDD,
+ 906634.900000ns, VDD,
+ 906635.000000ns, VSS,
+ 906875.100000ns, VSS,
+ 906875.200000ns, VDD,
+ 909757.500000ns, VDD,
+ 909757.600000ns, VSS,
+ 909877.600000ns, VSS,
+ 909877.700000ns, VDD,
+ 910237.900000ns, VDD,
+ 910238.000000ns, VSS,
+ 910478.100000ns, VSS,
+ 910478.200000ns, VDD,
+ 911679.100000ns, VDD,
+ 911679.200000ns, VSS,
+ 912039.400000ns, VSS,
+ 912039.500000ns, VDD,
+ 912399.700000ns, VDD,
+ 912399.800000ns, VSS,
+ 912519.800000ns, VSS,
+ 912519.900000ns, VDD,
+ 913720.800000ns, VDD,
+ 913720.900000ns, VSS,
+ 914081.100000ns, VSS,
+ 914081.200000ns, VDD,
+ 915162.000000ns, VDD,
+ 915162.100000ns, VSS,
+ 915282.100000ns, VSS,
+ 915282.200000ns, VDD,
+ 915642.400000ns, VDD,
+ 915642.500000ns, VSS,
+ 915882.600000ns, VSS,
+ 915882.700000ns, VDD,
+ 916002.700000ns, VDD,
+ 916002.800000ns, VSS,
+ 916483.100000ns, VSS,
+ 916483.200000ns, VDD,
+ 916843.400000ns, VDD,
+ 916843.500000ns, VSS,
+ 917323.800000ns, VSS,
+ 917323.900000ns, VDD,
+ 919125.300000ns, VDD,
+ 919125.400000ns, VSS,
+ 919605.700000ns, VSS,
+ 919605.800000ns, VDD,
+ 919966.000000ns, VDD,
+ 919966.100000ns, VSS,
+ 920206.200000ns, VSS,
+ 920206.300000ns, VDD,
+ 920566.500000ns, VDD,
+ 920566.600000ns, VSS,
+ 920926.800000ns, VSS,
+ 920926.900000ns, VDD,
+ 922488.100000ns, VDD,
+ 922488.200000ns, VSS,
+ 922848.400000ns, VSS,
+ 922848.500000ns, VDD,
+ 923208.700000ns, VDD,
+ 923208.800000ns, VSS,
+ 923448.900000ns, VSS,
+ 923449.000000ns, VDD,
+ 923569.000000ns, VDD,
+ 923569.100000ns, VSS,
+ 923689.100000ns, VSS,
+ 923689.200000ns, VDD,
+ 923809.200000ns, VDD,
+ 923809.300000ns, VSS,
+ 924409.700000ns, VSS,
+ 924409.800000ns, VDD,
+ 924890.100000ns, VDD,
+ 924890.200000ns, VSS,
+ 925130.300000ns, VSS,
+ 925130.400000ns, VDD,
+ 925250.400000ns, VDD,
+ 925250.500000ns, VSS,
+ 925610.700000ns, VSS,
+ 925610.800000ns, VDD,
+ 925971.000000ns, VDD,
+ 925971.100000ns, VSS,
+ 926331.300000ns, VSS,
+ 926331.400000ns, VDD,
+ 927772.500000ns, VDD,
+ 927772.600000ns, VSS,
+ 928493.100000ns, VSS,
+ 928493.200000ns, VDD,
+ 929453.900000ns, VDD,
+ 929454.000000ns, VSS,
+ 929934.300000ns, VSS,
+ 929934.400000ns, VDD,
+ 930174.500000ns, VDD,
+ 930174.600000ns, VSS,
+ 930534.800000ns, VSS,
+ 930534.900000ns, VDD,
+ 930654.900000ns, VDD,
+ 930655.000000ns, VSS,
+ 930895.100000ns, VSS,
+ 930895.200000ns, VDD,
+ 931135.300000ns, VDD,
+ 931135.400000ns, VSS,
+ 931495.600000ns, VSS,
+ 931495.700000ns, VDD,
+ 931855.900000ns, VDD,
+ 931856.000000ns, VSS,
+ 932216.200000ns, VSS,
+ 932216.300000ns, VDD,
+ 932576.500000ns, VDD,
+ 932576.600000ns, VSS,
+ 932816.700000ns, VSS,
+ 932816.800000ns, VDD,
+ 933056.900000ns, VDD,
+ 933057.000000ns, VSS,
+ 933177.000000ns, VSS,
+ 933177.100000ns, VDD,
+ 933297.100000ns, VDD,
+ 933297.200000ns, VSS,
+ 933657.400000ns, VSS,
+ 933657.500000ns, VDD,
+ 934017.700000ns, VDD,
+ 934017.800000ns, VSS,
+ 934257.900000ns, VSS,
+ 934258.000000ns, VDD,
+ 934498.100000ns, VDD,
+ 934498.200000ns, VSS,
+ 934858.400000ns, VSS,
+ 934858.500000ns, VDD,
+ 935218.700000ns, VDD,
+ 935218.800000ns, VSS,
+ 935458.900000ns, VSS,
+ 935459.000000ns, VDD,
+ 935819.200000ns, VDD,
+ 935819.300000ns, VSS,
+ 936179.500000ns, VSS,
+ 936179.600000ns, VDD,
+ 936900.100000ns, VDD,
+ 936900.200000ns, VSS,
+ 937380.500000ns, VSS,
+ 937380.600000ns, VDD,
+ 938221.200000ns, VDD,
+ 938221.300000ns, VSS,
+ 938701.600000ns, VSS,
+ 938701.700000ns, VDD,
+ 938821.700000ns, VDD,
+ 938821.800000ns, VSS,
+ 939182.000000ns, VSS,
+ 939182.100000ns, VDD,
+ 939302.100000ns, VDD,
+ 939302.200000ns, VSS,
+ 939422.200000ns, VSS,
+ 939422.300000ns, VDD,
+ 939782.500000ns, VDD,
+ 939782.600000ns, VSS,
+ 940383.000000ns, VSS,
+ 940383.100000ns, VDD,
+ 940743.300000ns, VDD,
+ 940743.400000ns, VSS,
+ 941103.600000ns, VSS,
+ 941103.700000ns, VDD,
+ 941463.900000ns, VDD,
+ 941464.000000ns, VSS,
+ 942184.500000ns, VSS,
+ 942184.600000ns, VDD,
+ 942424.700000ns, VDD,
+ 942424.800000ns, VSS,
+ 942785.000000ns, VSS,
+ 942785.100000ns, VDD,
+ 943385.500000ns, VDD,
+ 943385.600000ns, VSS,
+ 943865.900000ns, VSS,
+ 943866.000000ns, VDD,
+ 943986.000000ns, VDD,
+ 943986.100000ns, VSS,
+ 944106.100000ns, VSS,
+ 944106.200000ns, VDD,
+ 944466.400000ns, VDD,
+ 944466.500000ns, VSS,
+ 944586.500000ns, VSS,
+ 944586.600000ns, VDD,
+ 945307.100000ns, VDD,
+ 945307.200000ns, VSS,
+ 945667.400000ns, VSS,
+ 945667.500000ns, VDD,
+ 946027.700000ns, VDD,
+ 946027.800000ns, VSS,
+ 946388.000000ns, VSS,
+ 946388.100000ns, VDD,
+ 946508.100000ns, VDD,
+ 946508.200000ns, VSS,
+ 946628.200000ns, VSS,
+ 946628.300000ns, VDD,
+ 946868.400000ns, VDD,
+ 946868.500000ns, VSS,
+ 946988.500000ns, VSS,
+ 946988.600000ns, VDD,
+ 947348.800000ns, VDD,
+ 947348.900000ns, VSS,
+ 947468.900000ns, VSS,
+ 947469.000000ns, VDD,
+ 948309.600000ns, VDD,
+ 948309.700000ns, VSS,
+ 948429.700000ns, VSS,
+ 948429.800000ns, VDD,
+ 949030.200000ns, VDD,
+ 949030.300000ns, VSS,
+ 949270.400000ns, VSS,
+ 949270.500000ns, VDD,
+ 949390.500000ns, VDD,
+ 949390.600000ns, VSS,
+ 949510.600000ns, VSS,
+ 949510.700000ns, VDD,
+ 949870.900000ns, VDD,
+ 949871.000000ns, VSS,
+ 950111.100000ns, VSS,
+ 950111.200000ns, VDD,
+ 950231.200000ns, VDD,
+ 950231.300000ns, VSS,
+ 950351.300000ns, VSS,
+ 950351.400000ns, VDD,
+ 950951.800000ns, VDD,
+ 950951.900000ns, VSS,
+ 951192.000000ns, VSS,
+ 951192.100000ns, VDD,
+ 951432.200000ns, VDD,
+ 951432.300000ns, VSS,
+ 951672.400000ns, VSS,
+ 951672.500000ns, VDD,
+ 951912.600000ns, VDD,
+ 951912.700000ns, VSS,
+ 952272.900000ns, VSS,
+ 952273.000000ns, VDD,
+ 952513.100000ns, VDD,
+ 952513.200000ns, VSS,
+ 952873.400000ns, VSS,
+ 952873.500000ns, VDD,
+ 953594.000000ns, VDD,
+ 953594.100000ns, VSS,
+ 953714.100000ns, VSS,
+ 953714.200000ns, VDD,
+ 953834.200000ns, VDD,
+ 953834.300000ns, VSS,
+ 954314.600000ns, VSS,
+ 954314.700000ns, VDD,
+ 955275.400000ns, VDD,
+ 955275.500000ns, VSS,
+ 955395.500000ns, VSS,
+ 955395.600000ns, VDD,
+ 955515.600000ns, VDD,
+ 955515.700000ns, VSS,
+ 955755.800000ns, VSS,
+ 955755.900000ns, VDD,
+ 955875.900000ns, VDD,
+ 955876.000000ns, VSS,
+ 955996.000000ns, VSS,
+ 955996.100000ns, VDD,
+ 956356.300000ns, VDD,
+ 956356.400000ns, VSS,
+ 956596.500000ns, VSS,
+ 956596.600000ns, VDD,
+ 957076.900000ns, VDD,
+ 957077.000000ns, VSS,
+ 957437.200000ns, VSS,
+ 957437.300000ns, VDD,
+ 957557.300000ns, VDD,
+ 957557.400000ns, VSS,
+ 957797.500000ns, VSS,
+ 957797.600000ns, VDD,
+ 957917.600000ns, VDD,
+ 957917.700000ns, VSS,
+ 958758.300000ns, VSS,
+ 958758.400000ns, VDD,
+ 958998.500000ns, VDD,
+ 958998.600000ns, VSS,
+ 959118.600000ns, VSS,
+ 959118.700000ns, VDD,
+ 959238.700000ns, VDD,
+ 959238.800000ns, VSS,
+ 959358.800000ns, VSS,
+ 959358.900000ns, VDD,
+ 960439.700000ns, VDD,
+ 960439.800000ns, VSS,
+ 961040.200000ns, VSS,
+ 961040.300000ns, VDD,
+ 962961.800000ns, VDD,
+ 962961.900000ns, VSS,
+ 963322.100000ns, VSS,
+ 963322.200000ns, VDD,
+ 963562.300000ns, VDD,
+ 963562.400000ns, VSS,
+ 963682.400000ns, VSS,
+ 963682.500000ns, VDD,
+ 964042.700000ns, VDD,
+ 964042.800000ns, VSS,
+ 964162.800000ns, VSS,
+ 964162.900000ns, VDD,
+ 964282.900000ns, VDD,
+ 964283.000000ns, VSS,
+ 964403.000000ns, VSS,
+ 964403.100000ns, VDD,
+ 965604.000000ns, VDD,
+ 965604.100000ns, VSS,
+ 965724.100000ns, VSS,
+ 965724.200000ns, VDD,
+ 965964.300000ns, VDD,
+ 965964.400000ns, VSS,
+ 966084.400000ns, VSS,
+ 966084.500000ns, VDD,
+ 966204.500000ns, VDD,
+ 966204.600000ns, VSS,
+ 966324.600000ns, VSS,
+ 966324.700000ns, VDD,
+ 967045.200000ns, VDD,
+ 967045.300000ns, VSS,
+ 967165.300000ns, VSS,
+ 967165.400000ns, VDD,
+ 967885.900000ns, VDD,
+ 967886.000000ns, VSS,
+ 968006.000000ns, VSS,
+ 968006.100000ns, VDD,
+ 968366.300000ns, VDD,
+ 968366.400000ns, VSS,
+ 968606.500000ns, VSS,
+ 968606.600000ns, VDD,
+ 968846.700000ns, VDD,
+ 968846.800000ns, VSS,
+ 969447.200000ns, VSS,
+ 969447.300000ns, VDD,
+ 969567.300000ns, VDD,
+ 969567.400000ns, VSS,
+ 969807.500000ns, VSS,
+ 969807.600000ns, VDD,
+ 969927.600000ns, VDD,
+ 969927.700000ns, VSS,
+ 970047.700000ns, VSS,
+ 970047.800000ns, VDD,
+ 970287.900000ns, VDD,
+ 970288.000000ns, VSS,
+ 970408.000000ns, VSS,
+ 970408.100000ns, VDD,
+ 970528.100000ns, VDD,
+ 970528.200000ns, VSS,
+ 971729.100000ns, VSS,
+ 971729.200000ns, VDD,
+ 972089.400000ns, VDD,
+ 972089.500000ns, VSS,
+ 972329.600000ns, VSS,
+ 972329.700000ns, VDD,
+ 972810.000000ns, VDD,
+ 972810.100000ns, VSS,
+ 972930.100000ns, VSS,
+ 972930.200000ns, VDD,
+ 973170.300000ns, VDD,
+ 973170.400000ns, VSS,
+ 973410.500000ns, VSS,
+ 973410.600000ns, VDD,
+ 973530.600000ns, VDD,
+ 973530.700000ns, VSS,
+ 973650.700000ns, VSS,
+ 973650.800000ns, VDD,
+ 973890.900000ns, VDD,
+ 973891.000000ns, VSS,
+ 974011.000000ns, VSS,
+ 974011.100000ns, VDD,
+ 974371.300000ns, VDD,
+ 974371.400000ns, VSS,
+ 974491.400000ns, VSS,
+ 974491.500000ns, VDD,
+ 974611.500000ns, VDD,
+ 974611.600000ns, VSS,
+ 974731.600000ns, VSS,
+ 974731.700000ns, VDD,
+ 975091.900000ns, VDD,
+ 975092.000000ns, VSS,
+ 975452.200000ns, VSS,
+ 975452.300000ns, VDD,
+ 975692.400000ns, VDD,
+ 975692.500000ns, VSS,
+ 975932.600000ns, VSS,
+ 975932.700000ns, VDD,
+ 976172.800000ns, VDD,
+ 976172.900000ns, VSS,
+ 976533.100000ns, VSS,
+ 976533.200000ns, VDD,
+ 976773.300000ns, VDD,
+ 976773.400000ns, VSS,
+ 976893.400000ns, VSS,
+ 976893.500000ns, VDD,
+ 978094.400000ns, VDD,
+ 978094.500000ns, VSS,
+ 978334.600000ns, VSS,
+ 978334.700000ns, VDD,
+ 978574.800000ns, VDD,
+ 978574.900000ns, VSS,
+ 978815.000000ns, VSS,
+ 978815.100000ns, VDD,
+ 979175.300000ns, VDD,
+ 979175.400000ns, VSS,
+ 979295.400000ns, VSS,
+ 979295.500000ns, VDD,
+ 979535.600000ns, VDD,
+ 979535.700000ns, VSS,
+ 979655.700000ns, VSS,
+ 979655.800000ns, VDD,
+ 979775.800000ns, VDD,
+ 979775.900000ns, VSS,
+ 980136.100000ns, VSS,
+ 980136.200000ns, VDD,
+ 980616.500000ns, VDD,
+ 980616.600000ns, VSS,
+ 980736.600000ns, VSS,
+ 980736.700000ns, VDD,
+ 980976.800000ns, VDD,
+ 980976.900000ns, VSS,
+ 981096.900000ns, VSS,
+ 981097.000000ns, VDD,
+ 981217.000000ns, VDD,
+ 981217.100000ns, VSS,
+ 981577.300000ns, VSS,
+ 981577.400000ns, VDD,
+ 982177.800000ns, VDD,
+ 982177.900000ns, VSS,
+ 982297.900000ns, VSS,
+ 982298.000000ns, VDD,
+ 982538.100000ns, VDD,
+ 982538.200000ns, VSS,
+ 982658.200000ns, VSS,
+ 982658.300000ns, VDD,
+ 982898.400000ns, VDD,
+ 982898.500000ns, VSS,
+ 983498.900000ns, VSS,
+ 983499.000000ns, VDD,
+ 983859.200000ns, VDD,
+ 983859.300000ns, VSS,
+ 984219.500000ns, VSS,
+ 984219.600000ns, VDD,
+ 984459.700000ns, VDD,
+ 984459.800000ns, VSS,
+ 984579.800000ns, VSS,
+ 984579.900000ns, VDD,
+ 984699.900000ns, VDD,
+ 984700.000000ns, VSS,
+ 985180.300000ns, VSS,
+ 985180.400000ns, VDD,
+ 985540.600000ns, VDD,
+ 985540.700000ns, VSS,
+ 985780.800000ns, VSS,
+ 985780.900000ns, VDD,
+ 986141.100000ns, VDD,
+ 986141.200000ns, VSS,
+ 986741.600000ns, VSS,
+ 986741.700000ns, VDD,
+ 987101.900000ns, VDD,
+ 987102.000000ns, VSS,
+ 987702.400000ns, VSS,
+ 987702.500000ns, VDD,
+ 988062.700000ns, VDD,
+ 988062.800000ns, VSS,
+ 988182.800000ns, VSS,
+ 988182.900000ns, VDD,
+ 988302.900000ns, VDD,
+ 988303.000000ns, VSS,
+ 988783.300000ns, VSS,
+ 988783.400000ns, VDD,
+ 989383.800000ns, VDD,
+ 989383.900000ns, VSS,
+ 989503.900000ns, VSS,
+ 989504.000000ns, VDD,
+ 991065.200000ns, VDD,
+ 991065.300000ns, VSS,
+ 991425.500000ns, VSS,
+ 991425.600000ns, VDD,
+ 991665.700000ns, VDD,
+ 991665.800000ns, VSS,
+ 991905.900000ns, VSS,
+ 991906.000000ns, VDD,
+ 992026.000000ns, VDD,
+ 992026.100000ns, VSS,
+ 992386.300000ns, VSS,
+ 992386.400000ns, VDD,
+ 992626.500000ns, VDD,
+ 992626.600000ns, VSS,
+ 992746.600000ns, VSS,
+ 992746.700000ns, VDD,
+ 992986.800000ns, VDD,
+ 992986.900000ns, VSS,
+ 993707.400000ns, VSS,
+ 993707.500000ns, VDD,
+ 993947.600000ns, VDD,
+ 993947.700000ns, VSS,
+ 994307.900000ns, VSS,
+ 994308.000000ns, VDD,
+ 995148.600000ns, VDD,
+ 995148.700000ns, VSS,
+ 995268.700000ns, VSS,
+ 995268.800000ns, VDD,
+ 996349.600000ns, VDD,
+ 996349.700000ns, VSS,
+ 996469.700000ns, VSS,
+ 996469.800000ns, VDD,
+ 996589.800000ns, VDD,
+ 996589.900000ns, VSS,
+ 997070.200000ns, VSS,
+ 997070.300000ns, VDD,
+ 998751.600000ns, VDD,
+ 998751.700000ns, VSS,
+ 998871.700000ns, VSS,
+ 998871.800000ns, VDD,
+ 999232.000000ns, VDD,
+ 999232.100000ns, VSS,
+ 999352.100000ns, VSS,
+ 999352.200000ns, VDD,
+ 999592.300000ns, VDD,
+ 999592.400000ns, VSS,
+ 999832.500000ns, VSS,
+ 999832.600000ns, VDD,
+ 999952.600000ns, VDD,
+ 999952.700000ns, VSS,
+ 1000312.900000ns, VSS,
+ 1000313.000000ns, VDD,
+ 1000553.100000ns, VDD,
+ 1000553.200000ns, VSS,
+ 1000673.200000ns, VSS,
+ 1000673.300000ns, VDD,
+ 1001513.900000ns, VDD,
+ 1001514.000000ns, VSS,
+ 1001634.000000ns, VSS,
+ 1001634.100000ns, VDD,
+ 1001874.200000ns, VDD,
+ 1001874.300000ns, VSS,
+ 1002114.400000ns, VSS,
+ 1002114.500000ns, VDD,
+ 1002474.700000ns, VDD,
+ 1002474.800000ns, VSS,
+ 1002835.000000ns, VSS,
+ 1002835.100000ns, VDD,
+ 1002955.100000ns, VDD,
+ 1002955.200000ns, VSS,
+ 1003075.200000ns, VSS,
+ 1003075.300000ns, VDD,
+ 1003315.400000ns, VDD,
+ 1003315.500000ns, VSS,
+ 1003435.500000ns, VSS,
+ 1003435.600000ns, VDD,
+ 1003675.700000ns, VDD,
+ 1003675.800000ns, VSS,
+ 1003795.800000ns, VSS,
+ 1003795.900000ns, VDD,
+ 1003915.900000ns, VDD,
+ 1003916.000000ns, VSS,
+ 1004276.200000ns, VSS,
+ 1004276.300000ns, VDD,
+ 1004996.800000ns, VDD,
+ 1004996.900000ns, VSS,
+ 1005237.000000ns, VSS,
+ 1005237.100000ns, VDD,
+ 1006317.900000ns, VDD,
+ 1006318.000000ns, VSS,
+ 1006678.200000ns, VSS,
+ 1006678.300000ns, VDD,
+ 1007759.100000ns, VDD,
+ 1007759.200000ns, VSS,
+ 1008239.500000ns, VSS,
+ 1008239.600000ns, VDD,
+ 1008719.900000ns, VDD,
+ 1008720.000000ns, VSS,
+ 1009920.900000ns, VSS,
+ 1009921.000000ns, VDD,
+ 1010041.000000ns, VDD,
+ 1010041.100000ns, VSS,
+ 1010281.200000ns, VSS,
+ 1010281.300000ns, VDD,
+ 1011001.800000ns, VDD,
+ 1011001.900000ns, VSS,
+ 1011121.900000ns, VSS,
+ 1011122.000000ns, VDD,
+ 1011602.300000ns, VDD,
+ 1011602.400000ns, VSS,
+ 1011962.600000ns, VSS,
+ 1011962.700000ns, VDD,
+ 1012322.900000ns, VDD,
+ 1012323.000000ns, VSS,
+ 1012563.100000ns, VSS,
+ 1012563.200000ns, VDD,
+ 1012803.300000ns, VDD,
+ 1012803.400000ns, VSS,
+ 1013283.700000ns, VSS,
+ 1013283.800000ns, VDD,
+ 1013644.000000ns, VDD,
+ 1013644.100000ns, VSS,
+ 1014004.300000ns, VSS,
+ 1014004.400000ns, VDD,
+ 1014364.600000ns, VDD,
+ 1014364.700000ns, VSS,
+ 1014724.900000ns, VSS,
+ 1014725.000000ns, VDD,
+ 1015685.700000ns, VDD,
+ 1015685.800000ns, VSS,
+ 1015925.900000ns, VSS,
+ 1015926.000000ns, VDD,
+ 1016166.100000ns, VDD,
+ 1016166.200000ns, VSS,
+ 1016406.300000ns, VSS,
+ 1016406.400000ns, VDD,
+ 1016526.400000ns, VDD,
+ 1016526.500000ns, VSS,
+ 1016766.600000ns, VSS,
+ 1016766.700000ns, VDD,
+ 1017006.800000ns, VDD,
+ 1017006.900000ns, VSS,
+ 1017126.900000ns, VSS,
+ 1017127.000000ns, VDD,
+ 1017847.500000ns, VDD,
+ 1017847.600000ns, VSS,
+ 1017967.600000ns, VSS,
+ 1017967.700000ns, VDD,
+ 1018087.700000ns, VDD,
+ 1018087.800000ns, VSS,
+ 1018448.000000ns, VSS,
+ 1018448.100000ns, VDD,
+ 1018688.200000ns, VDD,
+ 1018688.300000ns, VSS,
+ 1018808.300000ns, VSS,
+ 1018808.400000ns, VDD,
+ 1019168.600000ns, VDD,
+ 1019168.700000ns, VSS,
+ 1019288.700000ns, VSS,
+ 1019288.800000ns, VDD,
+ 1020609.800000ns, VDD,
+ 1020609.900000ns, VSS,
+ 1020729.900000ns, VSS,
+ 1020730.000000ns, VDD,
+ 1020850.000000ns, VDD,
+ 1020850.100000ns, VSS,
+ 1020970.100000ns, VSS,
+ 1020970.200000ns, VDD,
+ 1021690.700000ns, VDD,
+ 1021690.800000ns, VSS,
+ 1021930.900000ns, VSS,
+ 1021931.000000ns, VDD,
+ 1022171.100000ns, VDD,
+ 1022171.200000ns, VSS,
+ 1023131.900000ns, VSS,
+ 1023132.000000ns, VDD,
+ 1024453.000000ns, VDD,
+ 1024453.100000ns, VSS,
+ 1024573.100000ns, VSS,
+ 1024573.200000ns, VDD,
+ 1025173.600000ns, VDD,
+ 1025173.700000ns, VSS,
+ 1025413.800000ns, VSS,
+ 1025413.900000ns, VDD,
+ 1025894.200000ns, VDD,
+ 1025894.300000ns, VSS,
+ 1026374.600000ns, VSS,
+ 1026374.700000ns, VDD,
+ 1026734.900000ns, VDD,
+ 1026735.000000ns, VSS,
+ 1027455.500000ns, VSS,
+ 1027455.600000ns, VDD,
+ 1027695.700000ns, VDD,
+ 1027695.800000ns, VSS,
+ 1027815.800000ns, VSS,
+ 1027815.900000ns, VDD,
+ 1028176.100000ns, VDD,
+ 1028176.200000ns, VSS,
+ 1028416.300000ns, VSS,
+ 1028416.400000ns, VDD,
+ 1029617.300000ns, VDD,
+ 1029617.400000ns, VSS,
+ 1030217.800000ns, VSS,
+ 1030217.900000ns, VDD,
+ 1031418.800000ns, VDD,
+ 1031418.900000ns, VSS,
+ 1031538.900000ns, VSS,
+ 1031539.000000ns, VDD,
+ 1031659.000000ns, VDD,
+ 1031659.100000ns, VSS,
+ 1031779.100000ns, VSS,
+ 1031779.200000ns, VDD,
+ 1032019.300000ns, VDD,
+ 1032019.400000ns, VSS,
+ 1032860.000000ns, VSS,
+ 1032860.100000ns, VDD,
+ 1033220.300000ns, VDD,
+ 1033220.400000ns, VSS,
+ 1033580.600000ns, VSS,
+ 1033580.700000ns, VDD,
+ 1035502.200000ns, VDD,
+ 1035502.300000ns, VSS,
+ 1035862.500000ns, VSS,
+ 1035862.600000ns, VDD,
+ 1036102.700000ns, VDD,
+ 1036102.800000ns, VSS,
+ 1036463.000000ns, VSS,
+ 1036463.100000ns, VDD,
+ 1036943.400000ns, VDD,
+ 1036943.500000ns, VSS,
+ 1037063.500000ns, VSS,
+ 1037063.600000ns, VDD,
+ 1037543.900000ns, VDD,
+ 1037544.000000ns, VSS,
+ 1037784.100000ns, VSS,
+ 1037784.200000ns, VDD,
+ 1038985.100000ns, VDD,
+ 1038985.200000ns, VSS,
+ 1039585.600000ns, VSS,
+ 1039585.700000ns, VDD,
+ 1039945.900000ns, VDD,
+ 1039946.000000ns, VSS,
+ 1040066.000000ns, VSS,
+ 1040066.100000ns, VDD,
+ 1041146.900000ns, VDD,
+ 1041147.000000ns, VSS,
+ 1041507.200000ns, VSS,
+ 1041507.300000ns, VDD,
+ 1041867.500000ns, VDD,
+ 1041867.600000ns, VSS,
+ 1042468.000000ns, VSS,
+ 1042468.100000ns, VDD,
+ 1042828.300000ns, VDD,
+ 1042828.400000ns, VSS,
+ 1043068.500000ns, VSS,
+ 1043068.600000ns, VDD,
+ 1043669.000000ns, VDD,
+ 1043669.100000ns, VSS,
+ 1043789.100000ns, VSS,
+ 1043789.200000ns, VDD,
+ 1043909.200000ns, VDD,
+ 1043909.300000ns, VSS,
+ 1044149.400000ns, VSS,
+ 1044149.500000ns, VDD,
+ 1044749.900000ns, VDD,
+ 1044750.000000ns, VSS,
+ 1045110.200000ns, VSS,
+ 1045110.300000ns, VDD,
+ 1045230.300000ns, VDD,
+ 1045230.400000ns, VSS,
+ 1045350.400000ns, VSS,
+ 1045350.500000ns, VDD,
+ 1045950.900000ns, VDD,
+ 1045951.000000ns, VSS,
+ 1046071.000000ns, VSS,
+ 1046071.100000ns, VDD,
+ 1046191.100000ns, VDD,
+ 1046191.200000ns, VSS,
+ 1046311.200000ns, VSS,
+ 1046311.300000ns, VDD,
+ 1046431.300000ns, VDD,
+ 1046431.400000ns, VSS,
+ 1046551.400000ns, VSS,
+ 1046551.500000ns, VDD,
+ 1046911.700000ns, VDD,
+ 1046911.800000ns, VSS,
+ 1047272.000000ns, VSS,
+ 1047272.100000ns, VDD,
+ 1047992.600000ns, VDD,
+ 1047992.700000ns, VSS,
+ 1048593.100000ns, VSS,
+ 1048593.200000ns, VDD,
+ 1048833.300000ns, VDD,
+ 1048833.400000ns, VSS,
+ 1049193.600000ns, VSS,
+ 1049193.700000ns, VDD,
+ 1049313.700000ns, VDD,
+ 1049313.800000ns, VSS,
+ 1049433.800000ns, VSS,
+ 1049433.900000ns, VDD,
+ 1050514.700000ns, VDD,
+ 1050514.800000ns, VSS,
+ 1050995.100000ns, VSS,
+ 1050995.200000ns, VDD,
+ 1051475.500000ns, VDD,
+ 1051475.600000ns, VSS,
+ 1051595.600000ns, VSS,
+ 1051595.700000ns, VDD,
+ 1051955.900000ns, VDD,
+ 1051956.000000ns, VSS,
+ 1052076.000000ns, VSS,
+ 1052076.100000ns, VDD,
+ 1052436.300000ns, VDD,
+ 1052436.400000ns, VSS,
+ 1052916.700000ns, VSS,
+ 1052916.800000ns, VDD,
+ 1053036.800000ns, VDD,
+ 1053036.900000ns, VSS,
+ 1053517.200000ns, VSS,
+ 1053517.300000ns, VDD,
+ 1053877.500000ns, VDD,
+ 1053877.600000ns, VSS,
+ 1054117.700000ns, VSS,
+ 1054117.800000ns, VDD,
+ 1054357.900000ns, VDD,
+ 1054358.000000ns, VSS,
+ 1054718.200000ns, VSS,
+ 1054718.300000ns, VDD,
+ 1055679.000000ns, VDD,
+ 1055679.100000ns, VSS,
+ 1056039.300000ns, VSS,
+ 1056039.400000ns, VDD,
+ 1056399.600000ns, VDD,
+ 1056399.700000ns, VSS,
+ 1057120.200000ns, VSS,
+ 1057120.300000ns, VDD,
+ 1057240.300000ns, VDD,
+ 1057240.400000ns, VSS,
+ 1057360.400000ns, VSS,
+ 1057360.500000ns, VDD,
+ 1057600.600000ns, VDD,
+ 1057600.700000ns, VSS,
+ 1057840.800000ns, VSS,
+ 1057840.900000ns, VDD,
+ 1058081.000000ns, VDD,
+ 1058081.100000ns, VSS,
+ 1058201.100000ns, VSS,
+ 1058201.200000ns, VDD,
+ 1058321.200000ns, VDD,
+ 1058321.300000ns, VSS,
+ 1058561.400000ns, VSS,
+ 1058561.500000ns, VDD,
+ 1058801.600000ns, VDD,
+ 1058801.700000ns, VSS,
+ 1059041.800000ns, VSS,
+ 1059041.900000ns, VDD,
+ 1059282.000000ns, VDD,
+ 1059282.100000ns, VSS,
+ 1059402.100000ns, VSS,
+ 1059402.200000ns, VDD,
+ 1059762.400000ns, VDD,
+ 1059762.500000ns, VSS,
+ 1060002.600000ns, VSS,
+ 1060002.700000ns, VDD,
+ 1060122.700000ns, VDD,
+ 1060122.800000ns, VSS,
+ 1060963.400000ns, VSS,
+ 1060963.500000ns, VDD,
+ 1061684.000000ns, VDD,
+ 1061684.100000ns, VSS,
+ 1061924.200000ns, VSS,
+ 1061924.300000ns, VDD,
+ 1062164.400000ns, VDD,
+ 1062164.500000ns, VSS,
+ 1063125.200000ns, VSS,
+ 1063125.300000ns, VDD,
+ 1063725.700000ns, VDD,
+ 1063725.800000ns, VSS,
+ 1064206.100000ns, VSS,
+ 1064206.200000ns, VDD,
+ 1065287.000000ns, VDD,
+ 1065287.100000ns, VSS,
+ 1065647.300000ns, VSS,
+ 1065647.400000ns, VDD,
+ 1066007.600000ns, VDD,
+ 1066007.700000ns, VSS,
+ 1066367.900000ns, VSS,
+ 1066368.000000ns, VDD,
+ 1066728.200000ns, VDD,
+ 1066728.300000ns, VSS,
+ 1066968.400000ns, VSS,
+ 1066968.500000ns, VDD,
+ 1067088.500000ns, VDD,
+ 1067088.600000ns, VSS,
+ 1067328.700000ns, VSS,
+ 1067328.800000ns, VDD,
+ 1067689.000000ns, VDD,
+ 1067689.100000ns, VSS,
+ 1068409.600000ns, VSS,
+ 1068409.700000ns, VDD,
+ 1070211.100000ns, VDD,
+ 1070211.200000ns, VSS,
+ 1070331.200000ns, VSS,
+ 1070331.300000ns, VDD,
+ 1070811.600000ns, VDD,
+ 1070811.700000ns, VSS,
+ 1071171.900000ns, VSS,
+ 1071172.000000ns, VDD,
+ 1072252.800000ns, VDD,
+ 1072252.900000ns, VSS,
+ 1073213.600000ns, VSS,
+ 1073213.700000ns, VDD,
+ 1073573.900000ns, VDD,
+ 1073574.000000ns, VSS,
+ 1073934.200000ns, VSS,
+ 1073934.300000ns, VDD,
+ 1074054.300000ns, VDD,
+ 1074054.400000ns, VSS,
+ 1074414.600000ns, VSS,
+ 1074414.700000ns, VDD,
+ 1074895.000000ns, VDD,
+ 1074895.100000ns, VSS,
+ 1075135.200000ns, VSS,
+ 1075135.300000ns, VDD,
+ 1075495.500000ns, VDD,
+ 1075495.600000ns, VSS,
+ 1075975.900000ns, VSS,
+ 1075976.000000ns, VDD,
+ 1077056.800000ns, VDD,
+ 1077056.900000ns, VSS,
+ 1077897.500000ns, VSS,
+ 1077897.600000ns, VDD,
+ 1078618.100000ns, VDD,
+ 1078618.200000ns, VSS,
+ 1078858.300000ns, VSS,
+ 1078858.400000ns, VDD,
+ 1079338.700000ns, VDD,
+ 1079338.800000ns, VSS,
+ 1079458.800000ns, VSS,
+ 1079458.900000ns, VDD,
+ 1080179.400000ns, VDD,
+ 1080179.500000ns, VSS,
+ 1080299.500000ns, VSS,
+ 1080299.600000ns, VDD,
+ 1080419.600000ns, VDD,
+ 1080419.700000ns, VSS,
+ 1080779.900000ns, VSS,
+ 1080780.000000ns, VDD,
+ 1082341.200000ns, VDD,
+ 1082341.300000ns, VSS,
+ 1082461.300000ns, VSS,
+ 1082461.400000ns, VDD,
+ 1082941.700000ns, VDD,
+ 1082941.800000ns, VSS,
+ 1083662.300000ns, VSS,
+ 1083662.400000ns, VDD,
+ 1083902.500000ns, VDD,
+ 1083902.600000ns, VSS,
+ 1084022.600000ns, VSS,
+ 1084022.700000ns, VDD,
+ 1084142.700000ns, VDD,
+ 1084142.800000ns, VSS,
+ 1084262.800000ns, VSS,
+ 1084262.900000ns, VDD,
+ 1084863.300000ns, VDD,
+ 1084863.400000ns, VSS,
+ 1084983.400000ns, VSS,
+ 1084983.500000ns, VDD,
+ 1085343.700000ns, VDD,
+ 1085343.800000ns, VSS,
+ 1085704.000000ns, VSS,
+ 1085704.100000ns, VDD,
+ 1086064.300000ns, VDD,
+ 1086064.400000ns, VSS,
+ 1086424.600000ns, VSS,
+ 1086424.700000ns, VDD,
+ 1086664.800000ns, VDD,
+ 1086664.900000ns, VSS,
+ 1086784.900000ns, VSS,
+ 1086785.000000ns, VDD,
+ 1087145.200000ns, VDD,
+ 1087145.300000ns, VSS,
+ 1087265.300000ns, VSS,
+ 1087265.400000ns, VDD,
+ 1087385.400000ns, VDD,
+ 1087385.500000ns, VSS,
+ 1088106.000000ns, VSS,
+ 1088106.100000ns, VDD,
+ 1088706.500000ns, VDD,
+ 1088706.600000ns, VSS,
+ 1088946.700000ns, VSS,
+ 1088946.800000ns, VDD,
+ 1089307.000000ns, VDD,
+ 1089307.100000ns, VSS,
+ 1089547.200000ns, VSS,
+ 1089547.300000ns, VDD,
+ 1089787.400000ns, VDD,
+ 1089787.500000ns, VSS,
+ 1089907.500000ns, VSS,
+ 1089907.600000ns, VDD,
+ 1090628.100000ns, VDD,
+ 1090628.200000ns, VSS,
+ 1091228.600000ns, VSS,
+ 1091228.700000ns, VDD,
+ 1091588.900000ns, VDD,
+ 1091589.000000ns, VSS,
+ 1091709.000000ns, VSS,
+ 1091709.100000ns, VDD,
+ 1092069.300000ns, VDD,
+ 1092069.400000ns, VSS,
+ 1092429.600000ns, VSS,
+ 1092429.700000ns, VDD,
+ 1092789.900000ns, VDD,
+ 1092790.000000ns, VSS,
+ 1093150.200000ns, VSS,
+ 1093150.300000ns, VDD,
+ 1094711.500000ns, VDD,
+ 1094711.600000ns, VSS,
+ 1094831.600000ns, VSS,
+ 1094831.700000ns, VDD,
+ 1095191.900000ns, VDD,
+ 1095192.000000ns, VSS,
+ 1095552.200000ns, VSS,
+ 1095552.300000ns, VDD,
+ 1095792.400000ns, VDD,
+ 1095792.500000ns, VSS,
+ 1096753.200000ns, VSS,
+ 1096753.300000ns, VDD,
+ 1097113.500000ns, VDD,
+ 1097113.600000ns, VSS,
+ 1097593.900000ns, VSS,
+ 1097594.000000ns, VDD,
+ 1097834.100000ns, VDD,
+ 1097834.200000ns, VSS,
+ 1098794.900000ns, VSS,
+ 1098795.000000ns, VDD,
+ 1099155.200000ns, VDD,
+ 1099155.300000ns, VSS,
+ 1099635.600000ns, VSS,
+ 1099635.700000ns, VDD,
+ 1099995.900000ns, VDD,
+ 1099996.000000ns, VSS,
+ 1100836.600000ns, VSS,
+ 1100836.700000ns, VDD,
+ 1101196.900000ns, VDD,
+ 1101197.000000ns, VSS,
+ 1101437.100000ns, VSS,
+ 1101437.200000ns, VDD,
+ 1101557.200000ns, VDD,
+ 1101557.300000ns, VSS,
+ 1101677.300000ns, VSS,
+ 1101677.400000ns, VDD,
+ 1103358.700000ns, VDD,
+ 1103358.800000ns, VSS,
+ 1104439.600000ns, VSS,
+ 1104439.700000ns, VDD,
+ 1105160.200000ns, VDD,
+ 1105160.300000ns, VSS,
+ 1105280.300000ns, VSS,
+ 1105280.400000ns, VDD,
+ 1106361.200000ns, VDD,
+ 1106361.300000ns, VSS,
+ 1106721.500000ns, VSS,
+ 1106721.600000ns, VDD,
+ 1107562.200000ns, VDD,
+ 1107562.300000ns, VSS,
+ 1108042.600000ns, VSS,
+ 1108042.700000ns, VDD,
+ 1108162.700000ns, VDD,
+ 1108162.800000ns, VSS,
+ 1108282.800000ns, VSS,
+ 1108282.900000ns, VDD,
+ 1108523.000000ns, VDD,
+ 1108523.100000ns, VSS,
+ 1108643.100000ns, VSS,
+ 1108643.200000ns, VDD,
+ 1108883.300000ns, VDD,
+ 1108883.400000ns, VSS,
+ 1109123.500000ns, VSS,
+ 1109123.600000ns, VDD,
+ 1110084.300000ns, VDD,
+ 1110084.400000ns, VSS,
+ 1110324.500000ns, VSS,
+ 1110324.600000ns, VDD,
+ 1111045.100000ns, VDD,
+ 1111045.200000ns, VSS,
+ 1111525.500000ns, VSS,
+ 1111525.600000ns, VDD,
+ 1111765.700000ns, VDD,
+ 1111765.800000ns, VSS,
+ 1111885.800000ns, VSS,
+ 1111885.900000ns, VDD,
+ 1112005.900000ns, VDD,
+ 1112006.000000ns, VSS,
+ 1112126.000000ns, VSS,
+ 1112126.100000ns, VDD,
+ 1113086.800000ns, VDD,
+ 1113086.900000ns, VSS,
+ 1113327.000000ns, VSS,
+ 1113327.100000ns, VDD,
+ 1114167.700000ns, VDD,
+ 1114167.800000ns, VSS,
+ 1114287.800000ns, VSS,
+ 1114287.900000ns, VDD,
+ 1114648.100000ns, VDD,
+ 1114648.200000ns, VSS,
+ 1115488.800000ns, VSS,
+ 1115488.900000ns, VDD,
+ 1115729.000000ns, VDD,
+ 1115729.100000ns, VSS,
+ 1115849.100000ns, VSS,
+ 1115849.200000ns, VDD,
+ 1116930.000000ns, VDD,
+ 1116930.100000ns, VSS,
+ 1117170.200000ns, VSS,
+ 1117170.300000ns, VDD,
+ 1117410.400000ns, VDD,
+ 1117410.500000ns, VSS,
+ 1117530.500000ns, VSS,
+ 1117530.600000ns, VDD,
+ 1117890.800000ns, VDD,
+ 1117890.900000ns, VSS,
+ 1118131.000000ns, VSS,
+ 1118131.100000ns, VDD,
+ 1119091.800000ns, VDD,
+ 1119091.900000ns, VSS,
+ 1119572.200000ns, VSS,
+ 1119572.300000ns, VDD,
+ 1119932.500000ns, VDD,
+ 1119932.600000ns, VSS,
+ 1120052.600000ns, VSS,
+ 1120052.700000ns, VDD,
+ 1120292.800000ns, VDD,
+ 1120292.900000ns, VSS,
+ 1120412.900000ns, VSS,
+ 1120413.000000ns, VDD,
+ 1120533.000000ns, VDD,
+ 1120533.100000ns, VSS,
+ 1120653.100000ns, VSS,
+ 1120653.200000ns, VDD,
+ 1121253.600000ns, VDD,
+ 1121253.700000ns, VSS,
+ 1121373.700000ns, VSS,
+ 1121373.800000ns, VDD,
+ 1121854.100000ns, VDD,
+ 1121854.200000ns, VSS,
+ 1122214.400000ns, VSS,
+ 1122214.500000ns, VDD,
+ 1122574.700000ns, VDD,
+ 1122574.800000ns, VSS,
+ 1122694.800000ns, VSS,
+ 1122694.900000ns, VDD,
+ 1122935.000000ns, VDD,
+ 1122935.100000ns, VSS,
+ 1123295.300000ns, VSS,
+ 1123295.400000ns, VDD,
+ 1124015.900000ns, VDD,
+ 1124016.000000ns, VSS,
+ 1124496.300000ns, VSS,
+ 1124496.400000ns, VDD,
+ 1125817.400000ns, VDD,
+ 1125817.500000ns, VSS,
+ 1126057.600000ns, VSS,
+ 1126057.700000ns, VDD,
+ 1126297.800000ns, VDD,
+ 1126297.900000ns, VSS,
+ 1126538.000000ns, VSS,
+ 1126538.100000ns, VDD,
+ 1127138.500000ns, VDD,
+ 1127138.600000ns, VSS,
+ 1127498.800000ns, VSS,
+ 1127498.900000ns, VDD,
+ 1128459.600000ns, VDD,
+ 1128459.700000ns, VSS,
+ 1128699.800000ns, VSS,
+ 1128699.900000ns, VDD,
+ 1129540.500000ns, VDD,
+ 1129540.600000ns, VSS,
+ 1129900.800000ns, VSS,
+ 1129900.900000ns, VDD,
+ 1130141.000000ns, VDD,
+ 1130141.100000ns, VSS,
+ 1130981.700000ns, VSS,
+ 1130981.800000ns, VDD,
+ 1131221.900000ns, VDD,
+ 1131222.000000ns, VSS,
+ 1131582.200000ns, VSS,
+ 1131582.300000ns, VDD,
+ 1131942.500000ns, VDD,
+ 1131942.600000ns, VSS,
+ 1132302.800000ns, VSS,
+ 1132302.900000ns, VDD,
+ 1132422.900000ns, VDD,
+ 1132423.000000ns, VSS,
+ 1132543.000000ns, VSS,
+ 1132543.100000ns, VDD,
+ 1132783.200000ns, VDD,
+ 1132783.300000ns, VSS,
+ 1132903.300000ns, VSS,
+ 1132903.400000ns, VDD,
+ 1133023.400000ns, VDD,
+ 1133023.500000ns, VSS,
+ 1133744.000000ns, VSS,
+ 1133744.100000ns, VDD,
+ 1133984.200000ns, VDD,
+ 1133984.300000ns, VSS,
+ 1134224.400000ns, VSS,
+ 1134224.500000ns, VDD,
+ 1134344.500000ns, VDD,
+ 1134344.600000ns, VSS,
+ 1134464.600000ns, VSS,
+ 1134464.700000ns, VDD,
+ 1134704.800000ns, VDD,
+ 1134704.900000ns, VSS,
+ 1134945.000000ns, VSS,
+ 1134945.100000ns, VDD,
+ 1135305.300000ns, VDD,
+ 1135305.400000ns, VSS,
+ 1135425.400000ns, VSS,
+ 1135425.500000ns, VDD,
+ 1136025.900000ns, VDD,
+ 1136026.000000ns, VSS,
+ 1136266.100000ns, VSS,
+ 1136266.200000ns, VDD,
+ 1136386.200000ns, VDD,
+ 1136386.300000ns, VSS,
+ 1136506.300000ns, VSS,
+ 1136506.400000ns, VDD,
+ 1136986.700000ns, VDD,
+ 1136986.800000ns, VSS,
+ 1137827.400000ns, VSS,
+ 1137827.500000ns, VDD,
+ 1137947.500000ns, VDD,
+ 1137947.600000ns, VSS,
+ 1138548.000000ns, VSS,
+ 1138548.100000ns, VDD,
+ 1138668.100000ns, VDD,
+ 1138668.200000ns, VSS,
+ 1139028.400000ns, VSS,
+ 1139028.500000ns, VDD,
+ 1139989.200000ns, VDD,
+ 1139989.300000ns, VSS,
+ 1140469.600000ns, VSS,
+ 1140469.700000ns, VDD,
+ 1140950.000000ns, VDD,
+ 1140950.100000ns, VSS,
+ 1141070.100000ns, VSS,
+ 1141070.200000ns, VDD,
+ 1141190.200000ns, VDD,
+ 1141190.300000ns, VSS,
+ 1141310.300000ns, VSS,
+ 1141310.400000ns, VDD,
+ 1141550.500000ns, VDD,
+ 1141550.600000ns, VSS,
+ 1141790.700000ns, VSS,
+ 1141790.800000ns, VDD,
+ 1142391.200000ns, VDD,
+ 1142391.300000ns, VSS,
+ 1143352.000000ns, VSS,
+ 1143352.100000ns, VDD,
+ 1143592.200000ns, VDD,
+ 1143592.300000ns, VSS,
+ 1144072.600000ns, VSS,
+ 1144072.700000ns, VDD,
+ 1144432.900000ns, VDD,
+ 1144433.000000ns, VSS,
+ 1144553.000000ns, VSS,
+ 1144553.100000ns, VDD,
+ 1145153.500000ns, VDD,
+ 1145153.600000ns, VSS,
+ 1145633.900000ns, VSS,
+ 1145634.000000ns, VDD,
+ 1145994.200000ns, VDD,
+ 1145994.300000ns, VSS,
+ 1146234.400000ns, VSS,
+ 1146234.500000ns, VDD,
+ 1146714.800000ns, VDD,
+ 1146714.900000ns, VSS,
+ 1147075.100000ns, VSS,
+ 1147075.200000ns, VDD,
+ 1147315.300000ns, VDD,
+ 1147315.400000ns, VSS,
+ 1147555.500000ns, VSS,
+ 1147555.600000ns, VDD,
+ 1148156.000000ns, VDD,
+ 1148156.100000ns, VSS,
+ 1148636.400000ns, VSS,
+ 1148636.500000ns, VDD,
+ 1149837.400000ns, VDD,
+ 1149837.500000ns, VSS,
+ 1150437.900000ns, VSS,
+ 1150438.000000ns, VDD,
+ 1151038.400000ns, VDD,
+ 1151038.500000ns, VSS,
+ 1151158.500000ns, VSS,
+ 1151158.600000ns, VDD,
+ 1151518.800000ns, VDD,
+ 1151518.900000ns, VSS,
+ 1151638.900000ns, VSS,
+ 1151639.000000ns, VDD,
+ 1151759.000000ns, VDD,
+ 1151759.100000ns, VSS,
+ 1151879.100000ns, VSS,
+ 1151879.200000ns, VDD,
+ 1152599.700000ns, VDD,
+ 1152599.800000ns, VSS,
+ 1152719.800000ns, VSS,
+ 1152719.900000ns, VDD,
+ 1152839.900000ns, VDD,
+ 1152840.000000ns, VSS,
+ 1153080.100000ns, VSS,
+ 1153080.200000ns, VDD,
+ 1153560.500000ns, VDD,
+ 1153560.600000ns, VSS,
+ 1153680.600000ns, VSS,
+ 1153680.700000ns, VDD,
+ 1154521.300000ns, VDD,
+ 1154521.400000ns, VSS,
+ 1154761.500000ns, VSS,
+ 1154761.600000ns, VDD,
+ 1155482.100000ns, VDD,
+ 1155482.200000ns, VSS,
+ 1155602.200000ns, VSS,
+ 1155602.300000ns, VDD,
+ 1155842.400000ns, VDD,
+ 1155842.500000ns, VSS,
+ 1155962.500000ns, VSS,
+ 1155962.600000ns, VDD,
+ 1157043.400000ns, VDD,
+ 1157043.500000ns, VSS,
+ 1157283.600000ns, VSS,
+ 1157283.700000ns, VDD,
+ 1157764.000000ns, VDD,
+ 1157764.100000ns, VSS,
+ 1158004.200000ns, VSS,
+ 1158004.300000ns, VDD,
+ 1158124.300000ns, VDD,
+ 1158124.400000ns, VSS,
+ 1158844.900000ns, VSS,
+ 1158845.000000ns, VDD,
+ 1159085.100000ns, VDD,
+ 1159085.200000ns, VSS,
+ 1159445.400000ns, VSS,
+ 1159445.500000ns, VDD,
+ 1159685.600000ns, VDD,
+ 1159685.700000ns, VSS,
+ 1159805.700000ns, VSS,
+ 1159805.800000ns, VDD,
+ 1160166.000000ns, VDD,
+ 1160166.100000ns, VSS,
+ 1160286.100000ns, VSS,
+ 1160286.200000ns, VDD,
+ 1160526.300000ns, VDD,
+ 1160526.400000ns, VSS,
+ 1160766.500000ns, VSS,
+ 1160766.600000ns, VDD,
+ 1160886.600000ns, VDD,
+ 1160886.700000ns, VSS,
+ 1161006.700000ns, VSS,
+ 1161006.800000ns, VDD,
+ 1161487.100000ns, VDD,
+ 1161487.200000ns, VSS,
+ 1161607.200000ns, VSS,
+ 1161607.300000ns, VDD,
+ 1161727.300000ns, VDD,
+ 1161727.400000ns, VSS,
+ 1161847.400000ns, VSS,
+ 1161847.500000ns, VDD,
+ 1162087.600000ns, VDD,
+ 1162087.700000ns, VSS,
+ 1162207.700000ns, VSS,
+ 1162207.800000ns, VDD,
+ 1162327.800000ns, VDD,
+ 1162327.900000ns, VSS,
+ 1162928.300000ns, VSS,
+ 1162928.400000ns, VDD,
+ 1163288.600000ns, VDD,
+ 1163288.700000ns, VSS,
+ 1163408.700000ns, VSS,
+ 1163408.800000ns, VDD,
+ 1164009.200000ns, VDD,
+ 1164009.300000ns, VSS,
+ 1164129.300000ns, VSS,
+ 1164129.400000ns, VDD,
+ 1164249.400000ns, VDD,
+ 1164249.500000ns, VSS,
+ 1164729.800000ns, VSS,
+ 1164729.900000ns, VDD,
+ 1165090.100000ns, VDD,
+ 1165090.200000ns, VSS,
+ 1165690.600000ns, VSS,
+ 1165690.700000ns, VDD,
+ 1165930.800000ns, VDD,
+ 1165930.900000ns, VSS,
+ 1166291.100000ns, VSS,
+ 1166291.200000ns, VDD,
+ 1166771.500000ns, VDD,
+ 1166771.600000ns, VSS,
+ 1167852.400000ns, VSS,
+ 1167852.500000ns, VDD,
+ 1168332.800000ns, VDD,
+ 1168332.900000ns, VSS,
+ 1168452.900000ns, VSS,
+ 1168453.000000ns, VDD,
+ 1168813.200000ns, VDD,
+ 1168813.300000ns, VSS,
+ 1169173.500000ns, VSS,
+ 1169173.600000ns, VDD,
+ 1170134.300000ns, VDD,
+ 1170134.400000ns, VSS,
+ 1170374.500000ns, VSS,
+ 1170374.600000ns, VDD,
+ 1171095.100000ns, VDD,
+ 1171095.200000ns, VSS,
+ 1171215.200000ns, VSS,
+ 1171215.300000ns, VDD,
+ 1171935.800000ns, VDD,
+ 1171935.900000ns, VSS,
+ 1172055.900000ns, VSS,
+ 1172056.000000ns, VDD,
+ 1173136.800000ns, VDD,
+ 1173136.900000ns, VSS,
+ 1173256.900000ns, VSS,
+ 1173257.000000ns, VDD,
+ 1173377.000000ns, VDD,
+ 1173377.100000ns, VSS,
+ 1173617.200000ns, VSS,
+ 1173617.300000ns, VDD,
+ 1173977.500000ns, VDD,
+ 1173977.600000ns, VSS,
+ 1174818.200000ns, VSS,
+ 1174818.300000ns, VDD,
+ 1176379.500000ns, VDD,
+ 1176379.600000ns, VSS,
+ 1176739.800000ns, VSS,
+ 1176739.900000ns, VDD,
+ 1176980.000000ns, VDD,
+ 1176980.100000ns, VSS,
+ 1177340.300000ns, VSS,
+ 1177340.400000ns, VDD,
+ 1177700.600000ns, VDD,
+ 1177700.700000ns, VSS,
+ 1178181.000000ns, VSS,
+ 1178181.100000ns, VDD,
+ 1178301.100000ns, VDD,
+ 1178301.200000ns, VSS,
+ 1178421.200000ns, VSS,
+ 1178421.300000ns, VDD,
+ 1178901.600000ns, VDD,
+ 1178901.700000ns, VSS,
+ 1179261.900000ns, VSS,
+ 1179262.000000ns, VDD,
+ 1179502.100000ns, VDD,
+ 1179502.200000ns, VSS,
+ 1180462.900000ns, VSS,
+ 1180463.000000ns, VDD,
+ 1180703.100000ns, VDD,
+ 1180703.200000ns, VSS,
+ 1180943.300000ns, VSS,
+ 1180943.400000ns, VDD,
+ 1181303.600000ns, VDD,
+ 1181303.700000ns, VSS,
+ 1181663.900000ns, VSS,
+ 1181664.000000ns, VDD,
+ 1182144.300000ns, VDD,
+ 1182144.400000ns, VSS,
+ 1182264.400000ns, VSS,
+ 1182264.500000ns, VDD,
+ 1182384.500000ns, VDD,
+ 1182384.600000ns, VSS,
+ 1182624.700000ns, VSS,
+ 1182624.800000ns, VDD,
+ 1183825.700000ns, VDD,
+ 1183825.800000ns, VSS,
+ 1183945.800000ns, VSS,
+ 1183945.900000ns, VDD,
+ 1184065.900000ns, VDD,
+ 1184066.000000ns, VSS,
+ 1184546.300000ns, VSS,
+ 1184546.400000ns, VDD,
+ 1185026.700000ns, VDD,
+ 1185026.800000ns, VSS,
+ 1185146.800000ns, VSS,
+ 1185146.900000ns, VDD,
+ 1185387.000000ns, VDD,
+ 1185387.100000ns, VSS,
+ 1185507.100000ns, VSS,
+ 1185507.200000ns, VDD,
+ 1185627.200000ns, VDD,
+ 1185627.300000ns, VSS,
+ 1185747.300000ns, VSS,
+ 1185747.400000ns, VDD,
+ 1187548.800000ns, VDD,
+ 1187548.900000ns, VSS,
+ 1187668.900000ns, VSS,
+ 1187669.000000ns, VDD,
+ 1188149.300000ns, VDD,
+ 1188149.400000ns, VSS,
+ 1188269.400000ns, VSS,
+ 1188269.500000ns, VDD,
+ 1188389.500000ns, VDD,
+ 1188389.600000ns, VSS,
+ 1188629.700000ns, VSS,
+ 1188629.800000ns, VDD,
+ 1188990.000000ns, VDD,
+ 1188990.100000ns, VSS,
+ 1189110.100000ns, VSS,
+ 1189110.200000ns, VDD,
+ 1189350.300000ns, VDD,
+ 1189350.400000ns, VSS,
+ 1189710.600000ns, VSS,
+ 1189710.700000ns, VDD,
+ 1190551.300000ns, VDD,
+ 1190551.400000ns, VSS,
+ 1190791.500000ns, VSS,
+ 1190791.600000ns, VDD,
+ 1191632.200000ns, VDD,
+ 1191632.300000ns, VSS,
+ 1191992.500000ns, VSS,
+ 1191992.600000ns, VDD,
+ 1192352.800000ns, VDD,
+ 1192352.900000ns, VSS,
+ 1193073.400000ns, VSS,
+ 1193073.500000ns, VDD,
+ 1193914.100000ns, VDD,
+ 1193914.200000ns, VSS,
+ 1194154.300000ns, VSS,
+ 1194154.400000ns, VDD,
+ 1194874.900000ns, VDD,
+ 1194875.000000ns, VSS,
+ 1194995.000000ns, VSS,
+ 1194995.100000ns, VDD,
+ 1195235.200000ns, VDD,
+ 1195235.300000ns, VSS,
+ 1195475.400000ns, VSS,
+ 1195475.500000ns, VDD,
+ 1195835.700000ns, VDD,
+ 1195835.800000ns, VSS,
+ 1196075.900000ns, VSS,
+ 1196076.000000ns, VDD,
+ 1196196.000000ns, VDD,
+ 1196196.100000ns, VSS,
+ 1197036.700000ns, VSS,
+ 1197036.800000ns, VDD,
+ 1197397.000000ns, VDD,
+ 1197397.100000ns, VSS,
+ 1197877.400000ns, VSS,
+ 1197877.500000ns, VDD,
+ 1198477.900000ns, VDD,
+ 1198478.000000ns, VSS,
+ 1198718.100000ns, VSS,
+ 1198718.200000ns, VDD,
+ 1199078.400000ns, VDD,
+ 1199078.500000ns, VSS,
+ 1199799.000000ns, VSS,
+ 1199799.100000ns, VDD,
+ 1200519.600000ns, VDD,
+ 1200519.700000ns, VSS,
+ 1200879.900000ns, VSS,
+ 1200880.000000ns, VDD,
+ 1201120.100000ns, VDD,
+ 1201120.200000ns, VSS,
+ 1201840.700000ns, VSS,
+ 1201840.800000ns, VDD,
+ 1202921.600000ns, VDD,
+ 1202921.700000ns, VSS,
+ 1203281.900000ns, VSS,
+ 1203282.000000ns, VDD,
+ 1203402.000000ns, VDD,
+ 1203402.100000ns, VSS,
+ 1203522.100000ns, VSS,
+ 1203522.200000ns, VDD,
+ 1204002.500000ns, VDD,
+ 1204002.600000ns, VSS,
+ 1204242.700000ns, VSS,
+ 1204242.800000ns, VDD,
+ 1204603.000000ns, VDD,
+ 1204603.100000ns, VSS,
+ 1205203.500000ns, VSS,
+ 1205203.600000ns, VDD,
+ 1205563.800000ns, VDD,
+ 1205563.900000ns, VSS,
+ 1206044.200000ns, VSS,
+ 1206044.300000ns, VDD,
+ 1206404.500000ns, VDD,
+ 1206404.600000ns, VSS,
+ 1207125.100000ns, VSS,
+ 1207125.200000ns, VDD,
+ 1207365.300000ns, VDD,
+ 1207365.400000ns, VSS,
+ 1207725.600000ns, VSS,
+ 1207725.700000ns, VDD,
+ 1208085.900000ns, VDD,
+ 1208086.000000ns, VSS,
+ 1208446.200000ns, VSS,
+ 1208446.300000ns, VDD,
+ 1208806.500000ns, VDD,
+ 1208806.600000ns, VSS,
+ 1209166.800000ns, VSS,
+ 1209166.900000ns, VDD,
+ 1209887.400000ns, VDD,
+ 1209887.500000ns, VSS,
+ 1210127.600000ns, VSS,
+ 1210127.700000ns, VDD,
+ 1210608.000000ns, VDD,
+ 1210608.100000ns, VSS,
+ 1210848.200000ns, VSS,
+ 1210848.300000ns, VDD,
+ 1211448.700000ns, VDD,
+ 1211448.800000ns, VSS,
+ 1211568.800000ns, VSS,
+ 1211568.900000ns, VDD,
+ 1212289.400000ns, VDD,
+ 1212289.500000ns, VSS,
+ 1212529.600000ns, VSS,
+ 1212529.700000ns, VDD,
+ 1213130.100000ns, VDD,
+ 1213130.200000ns, VSS,
+ 1213490.400000ns, VSS,
+ 1213490.500000ns, VDD,
+ 1213850.700000ns, VDD,
+ 1213850.800000ns, VSS,
+ 1214451.200000ns, VSS,
+ 1214451.300000ns, VDD,
+ 1214811.500000ns, VDD,
+ 1214811.600000ns, VSS,
+ 1214931.600000ns, VSS,
+ 1214931.700000ns, VDD,
+ 1215291.900000ns, VDD,
+ 1215292.000000ns, VSS,
+ 1216132.600000ns, VSS,
+ 1216132.700000ns, VDD,
+ 1216252.700000ns, VDD,
+ 1216252.800000ns, VSS,
+ 1216372.800000ns, VSS,
+ 1216372.900000ns, VDD,
+ 1218654.700000ns, VDD,
+ 1218654.800000ns, VSS,
+ 1218894.900000ns, VSS,
+ 1218895.000000ns, VDD,
+ 1219615.500000ns, VDD,
+ 1219615.600000ns, VSS,
+ 1219855.700000ns, VSS,
+ 1219855.800000ns, VDD,
+ 1220336.100000ns, VDD,
+ 1220336.200000ns, VSS,
+ 1220576.300000ns, VSS,
+ 1220576.400000ns, VDD,
+ 1220696.400000ns, VDD,
+ 1220696.500000ns, VSS,
+ 1220936.600000ns, VSS,
+ 1220936.700000ns, VDD,
+ 1221296.900000ns, VDD,
+ 1221297.000000ns, VSS,
+ 1221417.000000ns, VSS,
+ 1221417.100000ns, VDD,
+ 1221537.100000ns, VDD,
+ 1221537.200000ns, VSS,
+ 1221657.200000ns, VSS,
+ 1221657.300000ns, VDD,
+ 1222017.500000ns, VDD,
+ 1222017.600000ns, VSS,
+ 1222137.600000ns, VSS,
+ 1222137.700000ns, VDD,
+ 1223698.900000ns, VDD,
+ 1223699.000000ns, VSS,
+ 1223819.000000ns, VSS,
+ 1223819.100000ns, VDD,
+ 1224299.400000ns, VDD,
+ 1224299.500000ns, VSS,
+ 1224899.900000ns, VSS,
+ 1224900.000000ns, VDD,
+ 1225020.000000ns, VDD,
+ 1225020.100000ns, VSS,
+ 1225260.200000ns, VSS,
+ 1225260.300000ns, VDD,
+ 1225620.500000ns, VDD,
+ 1225620.600000ns, VSS,
+ 1225860.700000ns, VSS,
+ 1225860.800000ns, VDD,
+ 1226221.000000ns, VDD,
+ 1226221.100000ns, VSS,
+ 1226341.100000ns, VSS,
+ 1226341.200000ns, VDD,
+ 1226581.300000ns, VDD,
+ 1226581.400000ns, VSS,
+ 1226941.600000ns, VSS,
+ 1226941.700000ns, VDD,
+ 1227061.700000ns, VDD,
+ 1227061.800000ns, VSS,
+ 1227181.800000ns, VSS,
+ 1227181.900000ns, VDD,
+ 1227301.900000ns, VDD,
+ 1227302.000000ns, VSS,
+ 1227662.200000ns, VSS,
+ 1227662.300000ns, VDD,
+ 1227782.300000ns, VDD,
+ 1227782.400000ns, VSS,
+ 1227902.400000ns, VSS,
+ 1227902.500000ns, VDD,
+ 1229103.400000ns, VDD,
+ 1229103.500000ns, VSS,
+ 1229223.500000ns, VSS,
+ 1229223.600000ns, VDD,
+ 1229583.800000ns, VDD,
+ 1229583.900000ns, VSS,
+ 1229944.100000ns, VSS,
+ 1229944.200000ns, VDD,
+ 1230784.800000ns, VDD,
+ 1230784.900000ns, VSS,
+ 1231145.100000ns, VSS,
+ 1231145.200000ns, VDD,
+ 1231265.200000ns, VDD,
+ 1231265.300000ns, VSS,
+ 1231505.400000ns, VSS,
+ 1231505.500000ns, VDD,
+ 1231865.700000ns, VDD,
+ 1231865.800000ns, VSS,
+ 1231985.800000ns, VSS,
+ 1231985.900000ns, VDD,
+ 1232706.400000ns, VDD,
+ 1232706.500000ns, VSS,
+ 1233066.700000ns, VSS,
+ 1233066.800000ns, VDD,
+ 1233306.900000ns, VDD,
+ 1233307.000000ns, VSS,
+ 1233787.300000ns, VSS,
+ 1233787.400000ns, VDD,
+ 1234147.600000ns, VDD,
+ 1234147.700000ns, VSS,
+ 1234387.800000ns, VSS,
+ 1234387.900000ns, VDD,
+ 1234507.900000ns, VDD,
+ 1234508.000000ns, VSS,
+ 1234628.000000ns, VSS,
+ 1234628.100000ns, VDD,
+ 1234988.300000ns, VDD,
+ 1234988.400000ns, VSS,
+ 1235108.400000ns, VSS,
+ 1235108.500000ns, VDD,
+ 1235228.500000ns, VDD,
+ 1235228.600000ns, VSS,
+ 1235348.600000ns, VSS,
+ 1235348.700000ns, VDD,
+ 1235708.900000ns, VDD,
+ 1235709.000000ns, VSS,
+ 1236309.400000ns, VSS,
+ 1236309.500000ns, VDD,
+ 1236549.600000ns, VDD,
+ 1236549.700000ns, VSS,
+ 1236909.900000ns, VSS,
+ 1236910.000000ns, VDD,
+ 1237510.400000ns, VDD,
+ 1237510.500000ns, VSS,
+ 1237630.500000ns, VSS,
+ 1237630.600000ns, VDD,
+ 1237750.600000ns, VDD,
+ 1237750.700000ns, VSS,
+ 1237990.800000ns, VSS,
+ 1237990.900000ns, VDD,
+ 1239311.900000ns, VDD,
+ 1239312.000000ns, VSS,
+ 1239432.000000ns, VSS,
+ 1239432.100000ns, VDD,
+ 1239912.400000ns, VDD,
+ 1239912.500000ns, VSS,
+ 1240152.600000ns, VSS,
+ 1240152.700000ns, VDD,
+ 1241233.500000ns, VDD,
+ 1241233.600000ns, VSS,
+ 1241713.900000ns, VSS,
+ 1241714.000000ns, VDD,
+ 1241954.100000ns, VDD,
+ 1241954.200000ns, VSS,
+ 1242554.600000ns, VSS,
+ 1242554.700000ns, VDD,
+ 1242674.700000ns, VDD,
+ 1242674.800000ns, VSS,
+ 1243155.100000ns, VSS,
+ 1243155.200000ns, VDD,
+ 1243515.400000ns, VDD,
+ 1243515.500000ns, VSS,
+ 1243875.700000ns, VSS,
+ 1243875.800000ns, VDD,
+ 1243995.800000ns, VDD,
+ 1243995.900000ns, VSS,
+ 1244476.200000ns, VSS,
+ 1244476.300000ns, VDD,
+ 1244836.500000ns, VDD,
+ 1244836.600000ns, VSS,
+ 1245076.700000ns, VSS,
+ 1245076.800000ns, VDD,
+ 1245917.400000ns, VDD,
+ 1245917.500000ns, VSS,
+ 1246397.800000ns, VSS,
+ 1246397.900000ns, VDD,
+ 1247118.400000ns, VDD,
+ 1247118.500000ns, VSS,
+ 1247478.700000ns, VSS,
+ 1247478.800000ns, VDD,
+ 1247839.000000ns, VDD,
+ 1247839.100000ns, VSS,
+ 1248199.300000ns, VSS,
+ 1248199.400000ns, VDD,
+ 1248799.800000ns, VDD,
+ 1248799.900000ns, VSS,
+ 1248919.900000ns, VSS,
+ 1248920.000000ns, VDD,
+ 1249040.000000ns, VDD,
+ 1249040.100000ns, VSS,
+ 1249160.100000ns, VSS,
+ 1249160.200000ns, VDD,
+ 1249520.400000ns, VDD,
+ 1249520.500000ns, VSS,
+ 1250000.800000ns, VSS,
+ 1250000.900000ns, VDD,
+ 1250481.200000ns, VDD,
+ 1250481.300000ns, VSS,
+ 1250721.400000ns, VSS,
+ 1250721.500000ns, VDD,
+ 1251081.700000ns, VDD,
+ 1251081.800000ns, VSS,
+ 1251442.000000ns, VSS,
+ 1251442.100000ns, VDD,
+ 1251562.100000ns, VDD,
+ 1251562.200000ns, VSS,
+ 1252042.500000ns, VSS,
+ 1252042.600000ns, VDD,
+ 1252162.600000ns, VDD,
+ 1252162.700000ns, VSS,
+ 1252402.800000ns, VSS,
+ 1252402.900000ns, VDD,
+ 1253003.300000ns, VDD,
+ 1253003.400000ns, VSS,
+ 1253123.400000ns, VSS,
+ 1253123.500000ns, VDD,
+ 1253483.700000ns, VDD,
+ 1253483.800000ns, VSS,
+ 1253723.900000ns, VSS,
+ 1253724.000000ns, VDD,
+ 1255405.300000ns, VDD,
+ 1255405.400000ns, VSS,
+ 1255525.400000ns, VSS,
+ 1255525.500000ns, VDD,
+ 1256246.000000ns, VDD,
+ 1256246.100000ns, VSS,
+ 1256486.200000ns, VSS,
+ 1256486.300000ns, VDD,
+ 1256846.500000ns, VDD,
+ 1256846.600000ns, VSS,
+ 1257206.800000ns, VSS,
+ 1257206.900000ns, VDD,
+ 1257807.300000ns, VDD,
+ 1257807.400000ns, VSS,
+ 1258047.500000ns, VSS,
+ 1258047.600000ns, VDD,
+ 1258768.100000ns, VDD,
+ 1258768.200000ns, VSS,
+ 1259008.300000ns, VSS,
+ 1259008.400000ns, VDD,
+ 1259368.600000ns, VDD,
+ 1259368.700000ns, VSS,
+ 1259728.900000ns, VSS,
+ 1259729.000000ns, VDD,
+ 1259969.100000ns, VDD,
+ 1259969.200000ns, VSS,
+ 1260449.500000ns, VSS,
+ 1260449.600000ns, VDD,
+ 1261170.100000ns, VDD,
+ 1261170.200000ns, VSS,
+ 1261530.400000ns, VSS,
+ 1261530.500000ns, VDD,
+ 1262010.800000ns, VDD,
+ 1262010.900000ns, VSS,
+ 1262731.400000ns, VSS,
+ 1262731.500000ns, VDD,
+ 1263091.700000ns, VDD,
+ 1263091.800000ns, VSS,
+ 1263331.900000ns, VSS,
+ 1263332.000000ns, VDD,
+ 1263812.300000ns, VDD,
+ 1263812.400000ns, VSS,
+ 1263932.400000ns, VSS,
+ 1263932.500000ns, VDD,
+ 1264292.700000ns, VDD,
+ 1264292.800000ns, VSS,
+ 1265373.600000ns, VSS,
+ 1265373.700000ns, VDD,
+ 1265613.800000ns, VDD,
+ 1265613.900000ns, VSS,
+ 1265733.900000ns, VSS,
+ 1265734.000000ns, VDD,
+ 1265854.000000ns, VDD,
+ 1265854.100000ns, VSS,
+ 1266094.200000ns, VSS,
+ 1266094.300000ns, VDD,
+ 1266334.400000ns, VDD,
+ 1266334.500000ns, VSS,
+ 1266454.500000ns, VSS,
+ 1266454.600000ns, VDD,
+ 1268256.000000ns, VDD,
+ 1268256.100000ns, VSS,
+ 1268736.400000ns, VSS,
+ 1268736.500000ns, VDD,
+ 1269457.000000ns, VDD,
+ 1269457.100000ns, VSS,
+ 1269697.200000ns, VSS,
+ 1269697.300000ns, VDD,
+ 1269937.400000ns, VDD,
+ 1269937.500000ns, VSS,
+ 1270057.500000ns, VSS,
+ 1270057.600000ns, VDD,
+ 1270177.600000ns, VDD,
+ 1270177.700000ns, VSS,
+ 1270297.700000ns, VSS,
+ 1270297.800000ns, VDD,
+ 1270537.900000ns, VDD,
+ 1270538.000000ns, VSS,
+ 1270898.200000ns, VSS,
+ 1270898.300000ns, VDD,
+ 1271738.900000ns, VDD,
+ 1271739.000000ns, VSS,
+ 1272579.600000ns, VSS,
+ 1272579.700000ns, VDD,
+ 1272939.900000ns, VDD,
+ 1272940.000000ns, VSS,
+ 1273060.000000ns, VSS,
+ 1273060.100000ns, VDD,
+ 1273180.100000ns, VDD,
+ 1273180.200000ns, VSS,
+ 1273300.200000ns, VSS,
+ 1273300.300000ns, VDD,
+ 1273540.400000ns, VDD,
+ 1273540.500000ns, VSS,
+ 1274020.800000ns, VSS,
+ 1274020.900000ns, VDD,
+ 1274501.200000ns, VDD,
+ 1274501.300000ns, VSS,
+ 1274861.500000ns, VSS,
+ 1274861.600000ns, VDD,
+ 1274981.600000ns, VDD,
+ 1274981.700000ns, VSS,
+ 1275822.300000ns, VSS,
+ 1275822.400000ns, VDD,
+ 1276182.600000ns, VDD,
+ 1276182.700000ns, VSS,
+ 1277503.700000ns, VSS,
+ 1277503.800000ns, VDD,
+ 1277864.000000ns, VDD,
+ 1277864.100000ns, VSS,
+ 1278344.400000ns, VSS,
+ 1278344.500000ns, VDD,
+ 1278464.500000ns, VDD,
+ 1278464.600000ns, VSS,
+ 1278584.600000ns, VSS,
+ 1278584.700000ns, VDD,
+ 1278824.800000ns, VDD,
+ 1278824.900000ns, VSS,
+ 1279425.300000ns, VSS,
+ 1279425.400000ns, VDD,
+ 1279545.400000ns, VDD,
+ 1279545.500000ns, VSS,
+ 1279905.700000ns, VSS,
+ 1279905.800000ns, VDD,
+ 1280506.200000ns, VDD,
+ 1280506.300000ns, VSS,
+ 1280626.300000ns, VSS,
+ 1280626.400000ns, VDD,
+ 1281226.800000ns, VDD,
+ 1281226.900000ns, VSS,
+ 1281587.100000ns, VSS,
+ 1281587.200000ns, VDD,
+ 1281827.300000ns, VDD,
+ 1281827.400000ns, VSS,
+ 1282307.700000ns, VSS,
+ 1282307.800000ns, VDD,
+ 1283508.700000ns, VDD,
+ 1283508.800000ns, VSS,
+ 1283628.800000ns, VSS,
+ 1283628.900000ns, VDD,
+ 1286150.900000ns, VDD,
+ 1286151.000000ns, VSS,
+ 1286991.600000ns, VSS,
+ 1286991.700000ns, VDD,
+ 1287832.300000ns, VDD,
+ 1287832.400000ns, VSS,
+ 1287952.400000ns, VSS,
+ 1287952.500000ns, VDD,
+ 1289633.800000ns, VDD,
+ 1289633.900000ns, VSS,
+ 1289753.900000ns, VSS,
+ 1289754.000000ns, VDD,
+ 1289874.000000ns, VDD,
+ 1289874.100000ns, VSS,
+ 1290474.500000ns, VSS,
+ 1290474.600000ns, VDD,
+ 1290834.800000ns, VDD,
+ 1290834.900000ns, VSS,
+ 1291195.100000ns, VSS,
+ 1291195.200000ns, VDD,
+ 1291675.500000ns, VDD,
+ 1291675.600000ns, VSS,
+ 1291915.700000ns, VSS,
+ 1291915.800000ns, VDD,
+ 1292876.500000ns, VDD,
+ 1292876.600000ns, VSS,
+ 1292996.600000ns, VSS,
+ 1292996.700000ns, VDD,
+ 1293717.200000ns, VDD,
+ 1293717.300000ns, VSS,
+ 1293837.300000ns, VSS,
+ 1293837.400000ns, VDD,
+ 1294197.600000ns, VDD,
+ 1294197.700000ns, VSS,
+ 1294317.700000ns, VSS,
+ 1294317.800000ns, VDD,
+ 1294798.100000ns, VDD,
+ 1294798.200000ns, VSS,
+ 1294918.200000ns, VSS,
+ 1294918.300000ns, VDD,
+ 1295038.300000ns, VDD,
+ 1295038.400000ns, VSS,
+ 1295398.600000ns, VSS,
+ 1295398.700000ns, VDD,
+ 1295999.100000ns, VDD,
+ 1295999.200000ns, VSS,
+ 1296359.400000ns, VSS,
+ 1296359.500000ns, VDD,
+ 1296599.600000ns, VDD,
+ 1296599.700000ns, VSS,
+ 1296839.800000ns, VSS,
+ 1296839.900000ns, VDD,
+ 1298160.900000ns, VDD,
+ 1298161.000000ns, VSS,
+ 1298761.400000ns, VSS,
+ 1298761.500000ns, VDD,
+ 1299602.100000ns, VDD,
+ 1299602.200000ns, VSS,
+ 1299842.300000ns, VSS,
+ 1299842.400000ns, VDD,
+ 1300082.500000ns, VDD,
+ 1300082.600000ns, VSS,
+ 1300202.600000ns, VSS,
+ 1300202.700000ns, VDD,
+ 1300683.000000ns, VDD,
+ 1300683.100000ns, VSS,
+ 1301163.400000ns, VSS,
+ 1301163.500000ns, VDD,
+ 1301523.700000ns, VDD,
+ 1301523.800000ns, VSS,
+ 1301643.800000ns, VSS,
+ 1301643.900000ns, VDD,
+ 1301763.900000ns, VDD,
+ 1301764.000000ns, VSS,
+ 1301884.000000ns, VSS,
+ 1301884.100000ns, VDD,
+ 1302004.100000ns, VDD,
+ 1302004.200000ns, VSS,
+ 1302484.500000ns, VSS,
+ 1302484.600000ns, VDD,
+ 1302604.600000ns, VDD,
+ 1302604.700000ns, VSS,
+ 1302724.700000ns, VSS,
+ 1302724.800000ns, VDD,
+ 1303205.100000ns, VDD,
+ 1303205.200000ns, VSS,
+ 1304165.900000ns, VSS,
+ 1304166.000000ns, VDD,
+ 1304886.500000ns, VDD,
+ 1304886.600000ns, VSS,
+ 1305126.700000ns, VSS,
+ 1305126.800000ns, VDD,
+ 1305246.800000ns, VDD,
+ 1305246.900000ns, VSS,
+ 1305366.900000ns, VSS,
+ 1305367.000000ns, VDD,
+ 1305487.000000ns, VDD,
+ 1305487.100000ns, VSS,
+ 1305967.400000ns, VSS,
+ 1305967.500000ns, VDD,
+ 1306087.500000ns, VDD,
+ 1306087.600000ns, VSS,
+ 1306327.700000ns, VSS,
+ 1306327.800000ns, VDD,
+ 1306808.100000ns, VDD,
+ 1306808.200000ns, VSS,
+ 1307288.500000ns, VSS,
+ 1307288.600000ns, VDD,
+ 1308609.600000ns, VDD,
+ 1308609.700000ns, VSS,
+ 1308969.900000ns, VSS,
+ 1308970.000000ns, VDD,
+ 1309210.100000ns, VDD,
+ 1309210.200000ns, VSS,
+ 1309570.400000ns, VSS,
+ 1309570.500000ns, VDD,
+ 1310050.800000ns, VDD,
+ 1310050.900000ns, VSS,
+ 1310291.000000ns, VSS,
+ 1310291.100000ns, VDD,
+ 1310531.200000ns, VDD,
+ 1310531.300000ns, VSS,
+ 1310651.300000ns, VSS,
+ 1310651.400000ns, VDD,
+ 1310771.400000ns, VDD,
+ 1310771.500000ns, VSS,
+ 1311251.800000ns, VSS,
+ 1311251.900000ns, VDD,
+ 1311371.900000ns, VDD,
+ 1311372.000000ns, VSS,
+ 1311492.000000ns, VSS,
+ 1311492.100000ns, VDD,
+ 1311732.200000ns, VDD,
+ 1311732.300000ns, VSS,
+ 1311972.400000ns, VSS,
+ 1311972.500000ns, VDD,
+ 1312693.000000ns, VDD,
+ 1312693.100000ns, VSS,
+ 1312933.200000ns, VSS,
+ 1312933.300000ns, VDD,
+ 1313293.500000ns, VDD,
+ 1313293.600000ns, VSS,
+ 1313413.600000ns, VSS,
+ 1313413.700000ns, VDD,
+ 1313533.700000ns, VDD,
+ 1313533.800000ns, VSS,
+ 1313773.900000ns, VSS,
+ 1313774.000000ns, VDD,
+ 1314974.900000ns, VDD,
+ 1314975.000000ns, VSS,
+ 1315575.400000ns, VSS,
+ 1315575.500000ns, VDD,
+ 1315935.700000ns, VDD,
+ 1315935.800000ns, VSS,
+ 1316296.000000ns, VSS,
+ 1316296.100000ns, VDD,
+ 1316536.200000ns, VDD,
+ 1316536.300000ns, VSS,
+ 1316656.300000ns, VSS,
+ 1316656.400000ns, VDD,
+ 1316896.500000ns, VDD,
+ 1316896.600000ns, VSS,
+ 1317617.100000ns, VSS,
+ 1317617.200000ns, VDD,
+ 1317857.300000ns, VDD,
+ 1317857.400000ns, VSS,
+ 1318097.500000ns, VSS,
+ 1318097.600000ns, VDD,
+ 1318818.100000ns, VDD,
+ 1318818.200000ns, VSS,
+ 1319658.800000ns, VSS,
+ 1319658.900000ns, VDD,
+ 1319778.900000ns, VDD,
+ 1319779.000000ns, VSS,
+ 1319899.000000ns, VSS,
+ 1319899.100000ns, VDD,
+ 1320019.100000ns, VDD,
+ 1320019.200000ns, VSS,
+ 1320499.500000ns, VSS,
+ 1320499.600000ns, VDD,
+ 1321340.200000ns, VDD,
+ 1321340.300000ns, VSS,
+ 1322180.900000ns, VSS,
+ 1322181.000000ns, VDD,
+ 1322301.000000ns, VDD,
+ 1322301.100000ns, VSS,
+ 1322421.100000ns, VSS,
+ 1322421.200000ns, VDD,
+ 1322661.300000ns, VDD,
+ 1322661.400000ns, VSS,
+ 1322781.400000ns, VSS,
+ 1322781.500000ns, VDD,
+ 1323502.000000ns, VDD,
+ 1323502.100000ns, VSS,
+ 1323742.200000ns, VSS,
+ 1323742.300000ns, VDD,
+ 1324222.600000ns, VDD,
+ 1324222.700000ns, VSS,
+ 1324342.700000ns, VSS,
+ 1324342.800000ns, VDD,
+ 1324462.800000ns, VDD,
+ 1324462.900000ns, VSS,
+ 1324582.900000ns, VSS,
+ 1324583.000000ns, VDD,
+ 1324823.100000ns, VDD,
+ 1324823.200000ns, VSS,
+ 1324943.200000ns, VSS,
+ 1324943.300000ns, VDD,
+ 1325303.500000ns, VDD,
+ 1325303.600000ns, VSS,
+ 1325783.900000ns, VSS,
+ 1325784.000000ns, VDD,
+ 1326264.300000ns, VDD,
+ 1326264.400000ns, VSS,
+ 1326384.400000ns, VSS,
+ 1326384.500000ns, VDD,
+ 1326624.600000ns, VDD,
+ 1326624.700000ns, VSS,
+ 1327465.300000ns, VSS,
+ 1327465.400000ns, VDD,
+ 1328065.800000ns, VDD,
+ 1328065.900000ns, VSS,
+ 1328306.000000ns, VSS,
+ 1328306.100000ns, VDD,
+ 1329146.700000ns, VDD,
+ 1329146.800000ns, VSS,
+ 1329266.800000ns, VSS,
+ 1329266.900000ns, VDD,
+ 1329386.900000ns, VDD,
+ 1329387.000000ns, VSS,
+ 1329507.000000ns, VSS,
+ 1329507.100000ns, VDD,
+ 1329627.100000ns, VDD,
+ 1329627.200000ns, VSS,
+ 1330347.700000ns, VSS,
+ 1330347.800000ns, VDD,
+ 1330708.000000ns, VDD,
+ 1330708.100000ns, VSS,
+ 1331068.300000ns, VSS,
+ 1331068.400000ns, VDD,
+ 1332269.300000ns, VDD,
+ 1332269.400000ns, VSS,
+ 1332749.700000ns, VSS,
+ 1332749.800000ns, VDD,
+ 1333110.000000ns, VDD,
+ 1333110.100000ns, VSS,
+ 1333470.300000ns, VSS,
+ 1333470.400000ns, VDD,
+ 1333590.400000ns, VDD,
+ 1333590.500000ns, VSS,
+ 1333830.600000ns, VSS,
+ 1333830.700000ns, VDD,
+ 1335151.700000ns, VDD,
+ 1335151.800000ns, VSS,
+ 1335391.900000ns, VSS,
+ 1335392.000000ns, VDD,
+ 1335992.400000ns, VDD,
+ 1335992.500000ns, VSS,
+ 1336592.900000ns, VSS,
+ 1336593.000000ns, VDD,
+ 1336953.200000ns, VDD,
+ 1336953.300000ns, VSS,
+ 1337073.300000ns, VSS,
+ 1337073.400000ns, VDD,
+ 1337313.500000ns, VDD,
+ 1337313.600000ns, VSS,
+ 1337433.600000ns, VSS,
+ 1337433.700000ns, VDD,
+ 1337914.000000ns, VDD,
+ 1337914.100000ns, VSS,
+ 1338274.300000ns, VSS,
+ 1338274.400000ns, VDD,
+ 1338514.500000ns, VDD,
+ 1338514.600000ns, VSS,
+ 1338874.800000ns, VSS,
+ 1338874.900000ns, VDD,
+ 1339115.000000ns, VDD,
+ 1339115.100000ns, VSS,
+ 1339715.500000ns, VSS,
+ 1339715.600000ns, VDD,
+ 1340075.800000ns, VDD,
+ 1340075.900000ns, VSS,
+ 1341036.600000ns, VSS,
+ 1341036.700000ns, VDD,
+ 1341396.900000ns, VDD,
+ 1341397.000000ns, VSS,
+ 1341757.200000ns, VSS,
+ 1341757.300000ns, VDD,
+ 1342718.000000ns, VDD,
+ 1342718.100000ns, VSS,
+ 1343078.300000ns, VSS,
+ 1343078.400000ns, VDD,
+ 1343318.500000ns, VDD,
+ 1343318.600000ns, VSS,
+ 1343438.600000ns, VSS,
+ 1343438.700000ns, VDD,
+ 1345360.200000ns, VDD,
+ 1345360.300000ns, VSS,
+ 1346321.000000ns, VSS,
+ 1346321.100000ns, VDD,
+ 1346681.300000ns, VDD,
+ 1346681.400000ns, VSS,
+ 1346801.400000ns, VSS,
+ 1346801.500000ns, VDD,
+ 1346921.500000ns, VDD,
+ 1346921.600000ns, VSS,
+ 1347041.600000ns, VSS,
+ 1347041.700000ns, VDD,
+ 1347281.800000ns, VDD,
+ 1347281.900000ns, VSS,
+ 1347762.200000ns, VSS,
+ 1347762.300000ns, VDD,
+ 1347882.300000ns, VDD,
+ 1347882.400000ns, VSS,
+ 1348843.100000ns, VSS,
+ 1348843.200000ns, VDD,
+ 1349683.800000ns, VDD,
+ 1349683.900000ns, VSS,
+ 1350284.300000ns, VSS,
+ 1350284.400000ns, VDD,
+ 1350644.600000ns, VDD,
+ 1350644.700000ns, VSS,
+ 1350764.700000ns, VSS,
+ 1350764.800000ns, VDD,
+ 1351605.400000ns, VDD,
+ 1351605.500000ns, VSS,
+ 1351845.600000ns, VSS,
+ 1351845.700000ns, VDD,
+ 1352926.500000ns, VDD,
+ 1352926.600000ns, VSS,
+ 1353046.600000ns, VSS,
+ 1353046.700000ns, VDD,
+ 1353166.700000ns, VDD,
+ 1353166.800000ns, VSS,
+ 1353527.000000ns, VSS,
+ 1353527.100000ns, VDD,
+ 1354007.400000ns, VDD,
+ 1354007.500000ns, VSS,
+ 1354367.700000ns, VSS,
+ 1354367.800000ns, VDD,
+ 1355208.400000ns, VDD,
+ 1355208.500000ns, VSS,
+ 1355328.500000ns, VSS,
+ 1355328.600000ns, VDD,
+ 1355568.700000ns, VDD,
+ 1355568.800000ns, VSS,
+ 1355688.800000ns, VSS,
+ 1355688.900000ns, VDD,
+ 1355808.900000ns, VDD,
+ 1355809.000000ns, VSS,
+ 1355929.000000ns, VSS,
+ 1355929.100000ns, VDD,
+ 1356169.200000ns, VDD,
+ 1356169.300000ns, VSS,
+ 1356649.600000ns, VSS,
+ 1356649.700000ns, VDD,
+ 1357009.900000ns, VDD,
+ 1357010.000000ns, VSS,
+ 1357130.000000ns, VSS,
+ 1357130.100000ns, VDD,
+ 1357250.100000ns, VDD,
+ 1357250.200000ns, VSS,
+ 1357970.700000ns, VSS,
+ 1357970.800000ns, VDD,
+ 1358090.800000ns, VDD,
+ 1358090.900000ns, VSS,
+ 1358691.300000ns, VSS,
+ 1358691.400000ns, VDD,
+ 1359051.600000ns, VDD,
+ 1359051.700000ns, VSS,
+ 1359171.700000ns, VSS,
+ 1359171.800000ns, VDD,
+ 1360252.600000ns, VDD,
+ 1360252.700000ns, VSS,
+ 1360372.700000ns, VSS,
+ 1360372.800000ns, VDD,
+ 1360733.000000ns, VDD,
+ 1360733.100000ns, VSS,
+ 1360973.200000ns, VSS,
+ 1360973.300000ns, VDD,
+ 1362414.400000ns, VDD,
+ 1362414.500000ns, VSS,
+ 1362534.500000ns, VSS,
+ 1362534.600000ns, VDD,
+ 1362774.700000ns, VDD,
+ 1362774.800000ns, VSS,
+ 1362894.800000ns, VSS,
+ 1362894.900000ns, VDD,
+ 1363014.900000ns, VDD,
+ 1363015.000000ns, VSS,
+ 1363255.100000ns, VSS,
+ 1363255.200000ns, VDD,
+ 1363975.700000ns, VDD,
+ 1363975.800000ns, VSS,
+ 1364095.800000ns, VSS,
+ 1364095.900000ns, VDD,
+ 1364215.900000ns, VDD,
+ 1364216.000000ns, VSS,
+ 1364576.200000ns, VSS,
+ 1364576.300000ns, VDD,
+ 1364696.300000ns, VDD,
+ 1364696.400000ns, VSS,
+ 1365176.700000ns, VSS,
+ 1365176.800000ns, VDD,
+ 1365416.900000ns, VDD,
+ 1365417.000000ns, VSS,
+ 1365537.000000ns, VSS,
+ 1365537.100000ns, VDD,
+ 1365657.100000ns, VDD,
+ 1365657.200000ns, VSS,
+ 1366377.700000ns, VSS,
+ 1366377.800000ns, VDD,
+ 1366738.000000ns, VDD,
+ 1366738.100000ns, VSS,
+ 1366858.100000ns, VSS,
+ 1366858.200000ns, VDD,
+ 1367338.500000ns, VDD,
+ 1367338.600000ns, VSS,
+ 1367698.800000ns, VSS,
+ 1367698.900000ns, VDD,
+ 1368059.100000ns, VDD,
+ 1368059.200000ns, VSS,
+ 1368779.700000ns, VSS,
+ 1368779.800000ns, VDD,
+ 1369140.000000ns, VDD,
+ 1369140.100000ns, VSS,
+ 1369260.100000ns, VSS,
+ 1369260.200000ns, VDD,
+ 1369620.400000ns, VDD,
+ 1369620.500000ns, VSS,
+ 1369860.600000ns, VSS,
+ 1369860.700000ns, VDD,
+ 1370341.000000ns, VDD,
+ 1370341.100000ns, VSS,
+ 1370581.200000ns, VSS,
+ 1370581.300000ns, VDD,
+ 1371181.700000ns, VDD,
+ 1371181.800000ns, VSS,
+ 1371662.100000ns, VSS,
+ 1371662.200000ns, VDD,
+ 1372142.500000ns, VDD,
+ 1372142.600000ns, VSS,
+ 1372382.700000ns, VSS,
+ 1372382.800000ns, VDD,
+ 1372983.200000ns, VDD,
+ 1372983.300000ns, VSS,
+ 1373223.400000ns, VSS,
+ 1373223.500000ns, VDD,
+ 1373583.700000ns, VDD,
+ 1373583.800000ns, VSS,
+ 1373944.000000ns, VSS,
+ 1373944.100000ns, VDD,
+ 1374664.600000ns, VDD,
+ 1374664.700000ns, VSS,
+ 1374904.800000ns, VSS,
+ 1374904.900000ns, VDD,
+ 1375145.000000ns, VDD,
+ 1375145.100000ns, VSS,
+ 1375625.400000ns, VSS,
+ 1375625.500000ns, VDD,
+ 1376706.300000ns, VDD,
+ 1376706.400000ns, VSS,
+ 1376826.400000ns, VSS,
+ 1376826.500000ns, VDD,
+ 1377186.700000ns, VDD,
+ 1377186.800000ns, VSS,
+ 1377306.800000ns, VSS,
+ 1377306.900000ns, VDD,
+ 1378868.100000ns, VDD,
+ 1378868.200000ns, VSS,
+ 1378988.200000ns, VSS,
+ 1378988.300000ns, VDD,
+ 1379348.500000ns, VDD,
+ 1379348.600000ns, VSS,
+ 1379708.800000ns, VSS,
+ 1379708.900000ns, VDD,
+ 1380429.400000ns, VDD,
+ 1380429.500000ns, VSS,
+ 1380669.600000ns, VSS,
+ 1380669.700000ns, VDD,
+ 1382591.200000ns, VDD,
+ 1382591.300000ns, VSS,
+ 1382711.300000ns, VSS,
+ 1382711.400000ns, VDD,
+ 1383431.900000ns, VDD,
+ 1383432.000000ns, VSS,
+ 1383792.200000ns, VSS,
+ 1383792.300000ns, VDD,
+ 1384152.500000ns, VDD,
+ 1384152.600000ns, VSS,
+ 1384512.800000ns, VSS,
+ 1384512.900000ns, VDD,
+ 1385113.300000ns, VDD,
+ 1385113.400000ns, VSS,
+ 1385233.400000ns, VSS,
+ 1385233.500000ns, VDD,
+ 1385713.800000ns, VDD,
+ 1385713.900000ns, VSS,
+ 1385954.000000ns, VSS,
+ 1385954.100000ns, VDD,
+ 1386074.100000ns, VDD,
+ 1386074.200000ns, VSS,
+ 1386194.200000ns, VSS,
+ 1386194.300000ns, VDD,
+ 1386554.500000ns, VDD,
+ 1386554.600000ns, VSS,
+ 1386674.600000ns, VSS,
+ 1386674.700000ns, VDD,
+ 1387275.100000ns, VDD,
+ 1387275.200000ns, VSS,
+ 1387395.200000ns, VSS,
+ 1387395.300000ns, VDD,
+ 1387515.300000ns, VDD,
+ 1387515.400000ns, VSS,
+ 1388115.800000ns, VSS,
+ 1388115.900000ns, VDD,
+ 1388476.100000ns, VDD,
+ 1388476.200000ns, VSS,
+ 1388596.200000ns, VSS,
+ 1388596.300000ns, VDD,
+ 1388836.400000ns, VDD,
+ 1388836.500000ns, VSS,
+ 1389436.900000ns, VSS,
+ 1389437.000000ns, VDD,
+ 1390037.400000ns, VDD,
+ 1390037.500000ns, VSS,
+ 1390157.500000ns, VSS,
+ 1390157.600000ns, VDD,
+ 1390397.700000ns, VDD,
+ 1390397.800000ns, VSS,
+ 1390517.800000ns, VSS,
+ 1390517.900000ns, VDD,
+ 1390637.900000ns, VDD,
+ 1390638.000000ns, VSS,
+ 1390998.200000ns, VSS,
+ 1390998.300000ns, VDD,
+ 1391118.300000ns, VDD,
+ 1391118.400000ns, VSS,
+ 1391238.400000ns, VSS,
+ 1391238.500000ns, VDD,
+ 1392199.200000ns, VDD,
+ 1392199.300000ns, VSS,
+ 1392319.300000ns, VSS,
+ 1392319.400000ns, VDD,
+ 1392679.600000ns, VDD,
+ 1392679.700000ns, VSS,
+ 1392799.700000ns, VSS,
+ 1392799.800000ns, VDD,
+ 1392919.800000ns, VDD,
+ 1392919.900000ns, VSS,
+ 1393400.200000ns, VSS,
+ 1393400.300000ns, VDD,
+ 1393760.500000ns, VDD,
+ 1393760.600000ns, VSS,
+ 1394000.700000ns, VSS,
+ 1394000.800000ns, VDD,
+ 1394240.900000ns, VDD,
+ 1394241.000000ns, VSS,
+ 1394601.200000ns, VSS,
+ 1394601.300000ns, VDD,
+ 1395201.700000ns, VDD,
+ 1395201.800000ns, VSS,
+ 1395321.800000ns, VSS,
+ 1395321.900000ns, VDD,
+ 1395441.900000ns, VDD,
+ 1395442.000000ns, VSS,
+ 1395682.100000ns, VSS,
+ 1395682.200000ns, VDD,
+ 1395922.300000ns, VDD,
+ 1395922.400000ns, VSS,
+ 1396042.400000ns, VSS,
+ 1396042.500000ns, VDD,
+ 1397363.500000ns, VDD,
+ 1397363.600000ns, VSS,
+ 1397483.600000ns, VSS,
+ 1397483.700000ns, VDD,
+ 1397603.700000ns, VDD,
+ 1397603.800000ns, VSS,
+ 1397964.000000ns, VSS,
+ 1397964.100000ns, VDD,
+ 1398324.300000ns, VDD,
+ 1398324.400000ns, VSS,
+ 1398444.400000ns, VSS,
+ 1398444.500000ns, VDD,
+ 1398684.600000ns, VDD,
+ 1398684.700000ns, VSS,
+ 1398804.700000ns, VSS,
+ 1398804.800000ns, VDD,
+ 1399165.000000ns, VDD,
+ 1399165.100000ns, VSS,
+ 1399525.300000ns, VSS,
+ 1399525.400000ns, VDD,
+ 1399645.400000ns, VDD,
+ 1399645.500000ns, VSS,
+ 1399765.500000ns, VSS,
+ 1399765.600000ns, VDD,
+ 1400125.800000ns, VDD,
+ 1400125.900000ns, VSS,
+ 1400245.900000ns, VSS,
+ 1400246.000000ns, VDD,
+ 1400606.200000ns, VDD,
+ 1400606.300000ns, VSS,
+ 1401086.600000ns, VSS,
+ 1401086.700000ns, VDD,
+ 1401326.800000ns, VDD,
+ 1401326.900000ns, VSS,
+ 1401807.200000ns, VSS,
+ 1401807.300000ns, VDD,
+ 1402167.500000ns, VDD,
+ 1402167.600000ns, VSS,
+ 1402287.600000ns, VSS,
+ 1402287.700000ns, VDD,
+ 1402888.100000ns, VDD,
+ 1402888.200000ns, VSS,
+ 1403008.200000ns, VSS,
+ 1403008.300000ns, VDD,
+ 1403128.300000ns, VDD,
+ 1403128.400000ns, VSS,
+ 1403248.400000ns, VSS,
+ 1403248.500000ns, VDD,
+ 1403488.600000ns, VDD,
+ 1403488.700000ns, VSS,
+ 1403848.900000ns, VSS,
+ 1403849.000000ns, VDD,
+ 1405530.300000ns, VDD,
+ 1405530.400000ns, VSS,
+ 1406010.700000ns, VSS,
+ 1406010.800000ns, VDD,
+ 1406731.300000ns, VDD,
+ 1406731.400000ns, VSS,
+ 1406851.400000ns, VSS,
+ 1406851.500000ns, VDD,
+ 1407451.900000ns, VDD,
+ 1407452.000000ns, VSS,
+ 1407692.100000ns, VSS,
+ 1407692.200000ns, VDD,
+ 1408292.600000ns, VDD,
+ 1408292.700000ns, VSS,
+ 1408532.800000ns, VSS,
+ 1408532.900000ns, VDD,
+ 1409853.900000ns, VDD,
+ 1409854.000000ns, VSS,
+ 1409974.000000ns, VSS,
+ 1409974.100000ns, VDD,
+ 1410094.100000ns, VDD,
+ 1410094.200000ns, VSS,
+ 1410214.200000ns, VSS,
+ 1410214.300000ns, VDD,
+ 1410454.400000ns, VDD,
+ 1410454.500000ns, VSS,
+ 1410814.700000ns, VSS,
+ 1410814.800000ns, VDD,
+ 1412736.300000ns, VDD,
+ 1412736.400000ns, VSS,
+ 1412856.400000ns, VSS,
+ 1412856.500000ns, VDD,
+ 1413096.600000ns, VDD,
+ 1413096.700000ns, VSS,
+ 1413216.700000ns, VSS,
+ 1413216.800000ns, VDD,
+ 1413336.800000ns, VDD,
+ 1413336.900000ns, VSS,
+ 1413817.200000ns, VSS,
+ 1413817.300000ns, VDD,
+ 1413937.300000ns, VDD,
+ 1413937.400000ns, VSS,
+ 1414297.600000ns, VSS,
+ 1414297.700000ns, VDD,
+ 1414537.800000ns, VDD,
+ 1414537.900000ns, VSS,
+ 1414778.000000ns, VSS,
+ 1414778.100000ns, VDD,
+ 1415618.700000ns, VDD,
+ 1415618.800000ns, VSS,
+ 1415738.800000ns, VSS,
+ 1415738.900000ns, VDD,
+ 1415979.000000ns, VDD,
+ 1415979.100000ns, VSS,
+ 1416099.100000ns, VSS,
+ 1416099.200000ns, VDD,
+ 1416219.200000ns, VDD,
+ 1416219.300000ns, VSS,
+ 1416579.500000ns, VSS,
+ 1416579.600000ns, VDD,
+ 1417420.200000ns, VDD,
+ 1417420.300000ns, VSS,
+ 1417540.300000ns, VSS,
+ 1417540.400000ns, VDD,
+ 1417660.400000ns, VDD,
+ 1417660.500000ns, VSS,
+ 1417780.500000ns, VSS,
+ 1417780.600000ns, VDD,
+ 1418140.800000ns, VDD,
+ 1418140.900000ns, VSS,
+ 1418260.900000ns, VSS,
+ 1418261.000000ns, VDD,
+ 1418981.500000ns, VDD,
+ 1418981.600000ns, VSS,
+ 1419702.100000ns, VSS,
+ 1419702.200000ns, VDD,
+ 1421503.600000ns, VDD,
+ 1421503.700000ns, VSS,
+ 1421623.700000ns, VSS,
+ 1421623.800000ns, VDD,
+ 1421984.000000ns, VDD,
+ 1421984.100000ns, VSS,
+ 1422104.100000ns, VSS,
+ 1422104.200000ns, VDD,
+ 1422464.400000ns, VDD,
+ 1422464.500000ns, VSS,
+ 1422824.700000ns, VSS,
+ 1422824.800000ns, VDD,
+ 1423064.900000ns, VDD,
+ 1423065.000000ns, VSS,
+ 1423305.100000ns, VSS,
+ 1423305.200000ns, VDD,
+ 1423425.200000ns, VDD,
+ 1423425.300000ns, VSS,
+ 1423545.300000ns, VSS,
+ 1423545.400000ns, VDD,
+ 1423905.600000ns, VDD,
+ 1423905.700000ns, VSS,
+ 1424866.400000ns, VSS,
+ 1424866.500000ns, VDD,
+ 1425106.600000ns, VDD,
+ 1425106.700000ns, VSS,
+ 1425346.800000ns, VSS,
+ 1425346.900000ns, VDD,
+ 1425466.900000ns, VDD,
+ 1425467.000000ns, VSS,
+ 1425587.000000ns, VSS,
+ 1425587.100000ns, VDD,
+ 1425827.200000ns, VDD,
+ 1425827.300000ns, VSS,
+ 1425947.300000ns, VSS,
+ 1425947.400000ns, VDD,
+ 1426307.600000ns, VDD,
+ 1426307.700000ns, VSS,
+ 1426427.700000ns, VSS,
+ 1426427.800000ns, VDD,
+ 1426667.900000ns, VDD,
+ 1426668.000000ns, VSS,
+ 1426908.100000ns, VSS,
+ 1426908.200000ns, VDD,
+ 1427268.400000ns, VDD,
+ 1427268.500000ns, VSS,
+ 1427388.500000ns, VSS,
+ 1427388.600000ns, VDD,
+ 1427508.600000ns, VDD,
+ 1427508.700000ns, VSS,
+ 1427628.700000ns, VSS,
+ 1427628.800000ns, VDD,
+ 1428469.400000ns, VDD,
+ 1428469.500000ns, VSS,
+ 1428829.700000ns, VSS,
+ 1428829.800000ns, VDD,
+ 1429190.000000ns, VDD,
+ 1429190.100000ns, VSS,
+ 1429430.200000ns, VSS,
+ 1429430.300000ns, VDD,
+ 1429790.500000ns, VDD,
+ 1429790.600000ns, VSS,
+ 1430150.800000ns, VSS,
+ 1430150.900000ns, VDD,
+ 1430631.200000ns, VDD,
+ 1430631.300000ns, VSS,
+ 1430751.300000ns, VSS,
+ 1430751.400000ns, VDD,
+ 1431111.600000ns, VDD,
+ 1431111.700000ns, VSS,
+ 1431471.900000ns, VSS,
+ 1431472.000000ns, VDD,
+ 1431952.300000ns, VDD,
+ 1431952.400000ns, VSS,
+ 1432072.400000ns, VSS,
+ 1432072.500000ns, VDD,
+ 1432432.700000ns, VDD,
+ 1432432.800000ns, VSS,
+ 1433033.200000ns, VSS,
+ 1433033.300000ns, VDD,
+ 1433633.700000ns, VDD,
+ 1433633.800000ns, VSS,
+ 1433873.900000ns, VSS,
+ 1433874.000000ns, VDD,
+ 1433994.000000ns, VDD,
+ 1433994.100000ns, VSS,
+ 1434234.200000ns, VSS,
+ 1434234.300000ns, VDD,
+ 1435074.900000ns, VDD,
+ 1435075.000000ns, VSS,
+ 1435435.200000ns, VSS,
+ 1435435.300000ns, VDD,
+ 1435675.400000ns, VDD,
+ 1435675.500000ns, VSS,
+ 1435795.500000ns, VSS,
+ 1435795.600000ns, VDD,
+ 1436155.800000ns, VDD,
+ 1436155.900000ns, VSS,
+ 1436516.100000ns, VSS,
+ 1436516.200000ns, VDD,
+ 1436756.300000ns, VDD,
+ 1436756.400000ns, VSS,
+ 1436996.500000ns, VSS,
+ 1436996.600000ns, VDD,
+ 1438197.500000ns, VDD,
+ 1438197.600000ns, VSS,
+ 1438317.600000ns, VSS,
+ 1438317.700000ns, VDD,
+ 1438557.800000ns, VDD,
+ 1438557.900000ns, VSS,
+ 1438677.900000ns, VSS,
+ 1438678.000000ns, VDD,
+ 1438798.000000ns, VDD,
+ 1438798.100000ns, VSS,
+ 1439518.600000ns, VSS,
+ 1439518.700000ns, VDD,
+ 1439638.700000ns, VDD,
+ 1439638.800000ns, VSS,
+ 1440599.500000ns, VSS,
+ 1440599.600000ns, VDD,
+ 1441320.100000ns, VDD,
+ 1441320.200000ns, VSS,
+ 1441680.400000ns, VSS,
+ 1441680.500000ns, VDD,
+ 1441920.600000ns, VDD,
+ 1441920.700000ns, VSS,
+ 1442280.900000ns, VSS,
+ 1442281.000000ns, VDD,
+ 1442881.400000ns, VDD,
+ 1442881.500000ns, VSS,
+ 1443121.600000ns, VSS,
+ 1443121.700000ns, VDD,
+ 1443602.000000ns, VDD,
+ 1443602.100000ns, VSS,
+ 1443722.100000ns, VSS,
+ 1443722.200000ns, VDD,
+ 1443842.200000ns, VDD,
+ 1443842.300000ns, VSS,
+ 1444322.600000ns, VSS,
+ 1444322.700000ns, VDD,
+ 1444442.700000ns, VDD,
+ 1444442.800000ns, VSS,
+ 1444562.800000ns, VSS,
+ 1444562.900000ns, VDD,
+ 1444682.900000ns, VDD,
+ 1444683.000000ns, VSS,
+ 1445403.500000ns, VSS,
+ 1445403.600000ns, VDD,
+ 1446124.100000ns, VDD,
+ 1446124.200000ns, VSS,
+ 1446244.200000ns, VSS,
+ 1446244.300000ns, VDD,
+ 1446724.600000ns, VDD,
+ 1446724.700000ns, VSS,
+ 1447205.000000ns, VSS,
+ 1447205.100000ns, VDD,
+ 1448165.800000ns, VDD,
+ 1448165.900000ns, VSS,
+ 1448406.000000ns, VSS,
+ 1448406.100000ns, VDD,
+ 1448526.100000ns, VDD,
+ 1448526.200000ns, VSS,
+ 1449607.000000ns, VSS,
+ 1449607.100000ns, VDD,
+ 1450687.900000ns, VDD,
+ 1450688.000000ns, VSS,
+ 1451048.200000ns, VSS,
+ 1451048.300000ns, VDD,
+ 1451288.400000ns, VDD,
+ 1451288.500000ns, VSS,
+ 1451408.500000ns, VSS,
+ 1451408.600000ns, VDD,
+ 1451888.900000ns, VDD,
+ 1451889.000000ns, VSS,
+ 1452129.100000ns, VSS,
+ 1452129.200000ns, VDD,
+ 1452609.500000ns, VDD,
+ 1452609.600000ns, VSS,
+ 1452729.600000ns, VSS,
+ 1452729.700000ns, VDD,
+ 1453089.900000ns, VDD,
+ 1453090.000000ns, VSS,
+ 1453450.200000ns, VSS,
+ 1453450.300000ns, VDD,
+ 1453690.400000ns, VDD,
+ 1453690.500000ns, VSS,
+ 1454050.700000ns, VSS,
+ 1454050.800000ns, VDD,
+ 1454411.000000ns, VDD,
+ 1454411.100000ns, VSS,
+ 1454651.200000ns, VSS,
+ 1454651.300000ns, VDD,
+ 1454771.300000ns, VDD,
+ 1454771.400000ns, VSS,
+ 1454891.400000ns, VSS,
+ 1454891.500000ns, VDD,
+ 1455251.700000ns, VDD,
+ 1455251.800000ns, VSS,
+ 1455612.000000ns, VSS,
+ 1455612.100000ns, VDD,
+ 1455852.200000ns, VDD,
+ 1455852.300000ns, VSS,
+ 1456092.400000ns, VSS,
+ 1456092.500000ns, VDD,
+ 1456212.500000ns, VDD,
+ 1456212.600000ns, VSS,
+ 1456452.700000ns, VSS,
+ 1456452.800000ns, VDD,
+ 1456933.100000ns, VDD,
+ 1456933.200000ns, VSS,
+ 1457533.600000ns, VSS,
+ 1457533.700000ns, VDD,
+ 1457653.700000ns, VDD,
+ 1457653.800000ns, VSS,
+ 1457893.900000ns, VSS,
+ 1457894.000000ns, VDD,
+ 1458614.500000ns, VDD,
+ 1458614.600000ns, VSS,
+ 1458974.800000ns, VSS,
+ 1458974.900000ns, VDD,
+ 1459094.900000ns, VDD,
+ 1459095.000000ns, VSS,
+ 1459455.200000ns, VSS,
+ 1459455.300000ns, VDD,
+ 1459575.300000ns, VDD,
+ 1459575.400000ns, VSS,
+ 1459695.400000ns, VSS,
+ 1459695.500000ns, VDD,
+ 1459935.600000ns, VDD,
+ 1459935.700000ns, VSS,
+ 1460536.100000ns, VSS,
+ 1460536.200000ns, VDD,
+ 1460896.400000ns, VDD,
+ 1460896.500000ns, VSS,
+ 1461136.600000ns, VSS,
+ 1461136.700000ns, VDD,
+ 1461496.900000ns, VDD,
+ 1461497.000000ns, VSS,
+ 1462217.500000ns, VSS,
+ 1462217.600000ns, VDD,
+ 1462577.800000ns, VDD,
+ 1462577.900000ns, VSS,
+ 1462818.000000ns, VSS,
+ 1462818.100000ns, VDD,
+ 1463898.900000ns, VDD,
+ 1463899.000000ns, VSS,
+ 1464139.100000ns, VSS,
+ 1464139.200000ns, VDD,
+ 1464379.300000ns, VDD,
+ 1464379.400000ns, VSS,
+ 1464499.400000ns, VSS,
+ 1464499.500000ns, VDD,
+ 1464739.600000ns, VDD,
+ 1464739.700000ns, VSS,
+ 1464859.700000ns, VSS,
+ 1464859.800000ns, VDD,
+ 1464979.800000ns, VDD,
+ 1464979.900000ns, VSS,
+ 1465460.200000ns, VSS,
+ 1465460.300000ns, VDD,
+ 1465700.400000ns, VDD,
+ 1465700.500000ns, VSS,
+ 1465820.500000ns, VSS,
+ 1465820.600000ns, VDD,
+ 1466421.000000ns, VDD,
+ 1466421.100000ns, VSS,
+ 1466661.200000ns, VSS,
+ 1466661.300000ns, VDD,
+ 1467501.900000ns, VDD,
+ 1467502.000000ns, VSS,
+ 1467622.000000ns, VSS,
+ 1467622.100000ns, VDD,
+ 1467742.100000ns, VDD,
+ 1467742.200000ns, VSS,
+ 1468102.400000ns, VSS,
+ 1468102.500000ns, VDD,
+ 1468342.600000ns, VDD,
+ 1468342.700000ns, VSS,
+ 1468823.000000ns, VSS,
+ 1468823.100000ns, VDD,
+ 1468943.100000ns, VDD,
+ 1468943.200000ns, VSS,
+ 1469543.600000ns, VSS,
+ 1469543.700000ns, VDD,
+ 1470024.000000ns, VDD,
+ 1470024.100000ns, VSS,
+ 1470384.300000ns, VSS,
+ 1470384.400000ns, VDD,
+ 1470744.600000ns, VDD,
+ 1470744.700000ns, VSS,
+ 1470864.700000ns, VSS,
+ 1470864.800000ns, VDD,
+ 1472065.700000ns, VDD,
+ 1472065.800000ns, VSS,
+ 1472185.800000ns, VSS,
+ 1472185.900000ns, VDD,
+ 1472305.900000ns, VDD,
+ 1472306.000000ns, VSS,
+ 1472666.200000ns, VSS,
+ 1472666.300000ns, VDD,
+ 1472906.400000ns, VDD,
+ 1472906.500000ns, VSS,
+ 1473026.500000ns, VSS,
+ 1473026.600000ns, VDD,
+ 1473146.600000ns, VDD,
+ 1473146.700000ns, VSS,
+ 1473266.700000ns, VSS,
+ 1473266.800000ns, VDD,
+ 1473747.100000ns, VDD,
+ 1473747.200000ns, VSS,
+ 1473867.200000ns, VSS,
+ 1473867.300000ns, VDD,
+ 1474227.500000ns, VDD,
+ 1474227.600000ns, VSS,
+ 1474347.600000ns, VSS,
+ 1474347.700000ns, VDD,
+ 1474707.900000ns, VDD,
+ 1474708.000000ns, VSS,
+ 1475068.200000ns, VSS,
+ 1475068.300000ns, VDD,
+ 1475548.600000ns, VDD,
+ 1475548.700000ns, VSS,
+ 1475788.800000ns, VSS,
+ 1475788.900000ns, VDD,
+ 1477590.300000ns, VDD,
+ 1477590.400000ns, VSS,
+ 1477710.400000ns, VSS,
+ 1477710.500000ns, VDD,
+ 1477830.500000ns, VDD,
+ 1477830.600000ns, VSS,
+ 1477950.600000ns, VSS,
+ 1477950.700000ns, VDD,
+ 1478310.900000ns, VDD,
+ 1478311.000000ns, VSS,
+ 1478431.000000ns, VSS,
+ 1478431.100000ns, VDD,
+ 1479151.600000ns, VDD,
+ 1479151.700000ns, VSS,
+ 1479391.800000ns, VSS,
+ 1479391.900000ns, VDD,
+ 1480232.500000ns, VDD,
+ 1480232.600000ns, VSS,
+ 1480472.700000ns, VSS,
+ 1480472.800000ns, VDD,
+ 1480953.100000ns, VDD,
+ 1480953.200000ns, VSS,
+ 1481553.600000ns, VSS,
+ 1481553.700000ns, VDD,
+ 1481913.900000ns, VDD,
+ 1481914.000000ns, VSS,
+ 1482154.100000ns, VSS,
+ 1482154.200000ns, VDD,
+ 1482994.800000ns, VDD,
+ 1482994.900000ns, VSS,
+ 1483355.100000ns, VSS,
+ 1483355.200000ns, VDD,
+ 1483715.400000ns, VDD,
+ 1483715.500000ns, VSS,
+ 1484436.000000ns, VSS,
+ 1484436.100000ns, VDD,
+ 1485637.000000ns, VDD,
+ 1485637.100000ns, VSS,
+ 1486237.500000ns, VSS,
+ 1486237.600000ns, VDD,
+ 1486717.900000ns, VDD,
+ 1486718.000000ns, VSS,
+ 1486838.000000ns, VSS,
+ 1486838.100000ns, VDD,
+ 1487198.300000ns, VDD,
+ 1487198.400000ns, VSS,
+ 1487318.400000ns, VSS,
+ 1487318.500000ns, VDD,
+ 1487678.700000ns, VDD,
+ 1487678.800000ns, VSS,
+ 1488039.000000ns, VSS,
+ 1488039.100000ns, VDD,
+ 1488639.500000ns, VDD,
+ 1488639.600000ns, VSS,
+ 1488999.800000ns, VSS,
+ 1488999.900000ns, VDD,
+ 1490200.800000ns, VDD,
+ 1490200.900000ns, VSS,
+ 1490561.100000ns, VSS,
+ 1490561.200000ns, VDD,
+ 1491041.500000ns, VDD,
+ 1491041.600000ns, VSS,
+ 1491401.800000ns, VSS,
+ 1491401.900000ns, VDD,
+ 1492122.400000ns, VDD,
+ 1492122.500000ns, VSS,
+ 1492482.700000ns, VSS,
+ 1492482.800000ns, VDD,
+ 1493323.400000ns, VDD,
+ 1493323.500000ns, VSS,
+ 1493443.500000ns, VSS,
+ 1493443.600000ns, VDD,
+ 1494524.400000ns, VDD,
+ 1494524.500000ns, VSS,
+ 1494764.600000ns, VSS,
+ 1494764.700000ns, VDD,
+ 1494884.700000ns, VDD,
+ 1494884.800000ns, VSS,
+ 1495004.800000ns, VSS,
+ 1495004.900000ns, VDD,
+ 1495124.900000ns, VDD,
+ 1495125.000000ns, VSS,
+ 1495245.000000ns, VSS,
+ 1495245.100000ns, VDD,
+ 1495365.100000ns, VDD,
+ 1495365.200000ns, VSS,
+ 1495605.300000ns, VSS,
+ 1495605.400000ns, VDD,
+ 1495965.600000ns, VDD,
+ 1495965.700000ns, VSS,
+ 1496205.800000ns, VSS,
+ 1496205.900000ns, VDD,
+ 1496566.100000ns, VDD,
+ 1496566.200000ns, VSS,
+ 1497166.600000ns, VSS,
+ 1497166.700000ns, VDD,
+ 1497526.900000ns, VDD,
+ 1497527.000000ns, VSS,
+ 1497647.000000ns, VSS,
+ 1497647.100000ns, VDD,
+ 1498367.600000ns, VDD,
+ 1498367.700000ns, VSS,
+ 1498607.800000ns, VSS,
+ 1498607.900000ns, VDD,
+ 1498968.100000ns, VDD,
+ 1498968.200000ns, VSS,
+ 1499328.400000ns, VSS,
+ 1499328.500000ns, VDD,
+ 1499808.800000ns, VDD,
+ 1499808.900000ns, VSS,
+ 1500049.000000ns, VSS,
+ 1500049.100000ns, VDD,
+ 1500409.300000ns, VDD,
+ 1500409.400000ns, VSS,
+ 1501009.800000ns, VSS,
+ 1501009.900000ns, VDD,
+ 1501129.900000ns, VDD,
+ 1501130.000000ns, VSS,
+ 1501490.200000ns, VSS,
+ 1501490.300000ns, VDD,
+ 1503171.600000ns, VDD,
+ 1503171.700000ns, VSS,
+ 1503291.700000ns, VSS,
+ 1503291.800000ns, VDD,
+ 1504012.300000ns, VDD,
+ 1504012.400000ns, VSS,
+ 1504132.400000ns, VSS,
+ 1504132.500000ns, VDD,
+ 1504252.500000ns, VDD,
+ 1504252.600000ns, VSS,
+ 1504732.900000ns, VSS,
+ 1504733.000000ns, VDD,
+ 1505333.400000ns, VDD,
+ 1505333.500000ns, VSS,
+ 1505813.800000ns, VSS,
+ 1505813.900000ns, VDD,
+ 1506294.200000ns, VDD,
+ 1506294.300000ns, VSS,
+ 1506414.300000ns, VSS,
+ 1506414.400000ns, VDD,
+ 1506774.600000ns, VDD,
+ 1506774.700000ns, VSS,
+ 1506894.700000ns, VSS,
+ 1506894.800000ns, VDD,
+ 1507014.800000ns, VDD,
+ 1507014.900000ns, VSS,
+ 1507375.100000ns, VSS,
+ 1507375.200000ns, VDD,
+ 1507735.400000ns, VDD,
+ 1507735.500000ns, VSS,
+ 1507855.500000ns, VSS,
+ 1507855.600000ns, VDD,
+ 1507975.600000ns, VDD,
+ 1507975.700000ns, VSS,
+ 1508335.900000ns, VSS,
+ 1508336.000000ns, VDD,
+ 1508816.300000ns, VDD,
+ 1508816.400000ns, VSS,
+ 1508936.400000ns, VSS,
+ 1508936.500000ns, VDD,
+ 1509176.600000ns, VDD,
+ 1509176.700000ns, VSS,
+ 1509296.700000ns, VSS,
+ 1509296.800000ns, VDD,
+ 1510017.300000ns, VDD,
+ 1510017.400000ns, VSS,
+ 1510377.600000ns, VSS,
+ 1510377.700000ns, VDD,
+ 1510858.000000ns, VDD,
+ 1510858.100000ns, VSS,
+ 1510978.100000ns, VSS,
+ 1510978.200000ns, VDD,
+ 1511098.200000ns, VDD,
+ 1511098.300000ns, VSS,
+ 1511458.500000ns, VSS,
+ 1511458.600000ns, VDD,
+ 1512779.600000ns, VDD,
+ 1512779.700000ns, VSS,
+ 1512899.700000ns, VSS,
+ 1512899.800000ns, VDD,
+ 1513260.000000ns, VDD,
+ 1513260.100000ns, VSS,
+ 1513620.300000ns, VSS,
+ 1513620.400000ns, VDD,
+ 1513860.500000ns, VDD,
+ 1513860.600000ns, VSS,
+ 1514100.700000ns, VSS,
+ 1514100.800000ns, VDD,
+ 1514821.300000ns, VDD,
+ 1514821.400000ns, VSS,
+ 1515301.700000ns, VSS,
+ 1515301.800000ns, VDD,
+ 1515541.900000ns, VDD,
+ 1515542.000000ns, VSS,
+ 1515782.100000ns, VSS,
+ 1515782.200000ns, VDD,
+ 1516142.400000ns, VDD,
+ 1516142.500000ns, VSS,
+ 1516742.900000ns, VSS,
+ 1516743.000000ns, VDD,
+ 1517103.200000ns, VDD,
+ 1517103.300000ns, VSS,
+ 1517223.300000ns, VSS,
+ 1517223.400000ns, VDD,
+ 1517343.400000ns, VDD,
+ 1517343.500000ns, VSS,
+ 1517703.700000ns, VSS,
+ 1517703.800000ns, VDD,
+ 1518184.100000ns, VDD,
+ 1518184.200000ns, VSS,
+ 1518304.200000ns, VSS,
+ 1518304.300000ns, VDD,
+ 1518424.300000ns, VDD,
+ 1518424.400000ns, VSS,
+ 1518664.500000ns, VSS,
+ 1518664.600000ns, VDD,
+ 1519505.200000ns, VDD,
+ 1519505.300000ns, VSS,
+ 1519745.400000ns, VSS,
+ 1519745.500000ns, VDD,
+ 1519985.600000ns, VDD,
+ 1519985.700000ns, VSS,
+ 1520225.800000ns, VSS,
+ 1520225.900000ns, VDD,
+ 1520826.300000ns, VDD,
+ 1520826.400000ns, VSS,
+ 1521066.500000ns, VSS,
+ 1521066.600000ns, VDD,
+ 1521426.800000ns, VDD,
+ 1521426.900000ns, VSS,
+ 1521787.100000ns, VSS,
+ 1521787.200000ns, VDD,
+ 1522267.500000ns, VDD,
+ 1522267.600000ns, VSS,
+ 1522507.700000ns, VSS,
+ 1522507.800000ns, VDD,
+ 1522627.800000ns, VDD,
+ 1522627.900000ns, VSS,
+ 1522747.900000ns, VSS,
+ 1522748.000000ns, VDD,
+ 1522868.000000ns, VDD,
+ 1522868.100000ns, VSS,
+ 1522988.100000ns, VSS,
+ 1522988.200000ns, VDD,
+ 1523588.600000ns, VDD,
+ 1523588.700000ns, VSS,
+ 1523708.700000ns, VSS,
+ 1523708.800000ns, VDD,
+ 1524549.400000ns, VDD,
+ 1524549.500000ns, VSS,
+ 1525029.800000ns, VSS,
+ 1525029.900000ns, VDD,
+ 1525270.000000ns, VDD,
+ 1525270.100000ns, VSS,
+ 1525990.600000ns, VSS,
+ 1525990.700000ns, VDD,
+ 1526350.900000ns, VDD,
+ 1526351.000000ns, VSS,
+ 1527431.800000ns, VSS,
+ 1527431.900000ns, VDD,
+ 1528032.300000ns, VDD,
+ 1528032.400000ns, VSS,
+ 1528632.800000ns, VSS,
+ 1528632.900000ns, VDD,
+ 1528873.000000ns, VDD,
+ 1528873.100000ns, VSS,
+ 1528993.100000ns, VSS,
+ 1528993.200000ns, VDD,
+ 1529833.800000ns, VDD,
+ 1529833.900000ns, VSS,
+ 1530074.000000ns, VSS,
+ 1530074.100000ns, VDD,
+ 1530314.200000ns, VDD,
+ 1530314.300000ns, VSS,
+ 1530674.500000ns, VSS,
+ 1530674.600000ns, VDD,
+ 1531034.800000ns, VDD,
+ 1531034.900000ns, VSS,
+ 1531755.400000ns, VSS,
+ 1531755.500000ns, VDD,
+ 1532716.200000ns, VDD,
+ 1532716.300000ns, VSS,
+ 1532956.400000ns, VSS,
+ 1532956.500000ns, VDD,
+ 1533076.500000ns, VDD,
+ 1533076.600000ns, VSS,
+ 1533196.600000ns, VSS,
+ 1533196.700000ns, VDD,
+ 1533677.000000ns, VDD,
+ 1533677.100000ns, VSS,
+ 1533797.100000ns, VSS,
+ 1533797.200000ns, VDD,
+ 1534277.500000ns, VDD,
+ 1534277.600000ns, VSS,
+ 1534517.700000ns, VSS,
+ 1534517.800000ns, VDD,
+ 1534637.800000ns, VDD,
+ 1534637.900000ns, VSS,
+ 1534998.100000ns, VSS,
+ 1534998.200000ns, VDD,
+ 1535118.200000ns, VDD,
+ 1535118.300000ns, VSS,
+ 1535358.400000ns, VSS,
+ 1535358.500000ns, VDD,
+ 1535958.900000ns, VDD,
+ 1535959.000000ns, VSS,
+ 1536079.000000ns, VSS,
+ 1536079.100000ns, VDD,
+ 1536799.600000ns, VDD,
+ 1536799.700000ns, VSS,
+ 1536919.700000ns, VSS,
+ 1536919.800000ns, VDD,
+ 1537039.800000ns, VDD,
+ 1537039.900000ns, VSS,
+ 1537159.900000ns, VSS,
+ 1537160.000000ns, VDD,
+ 1538000.600000ns, VDD,
+ 1538000.700000ns, VSS,
+ 1538481.000000ns, VSS,
+ 1538481.100000ns, VDD,
+ 1538601.100000ns, VDD,
+ 1538601.200000ns, VSS,
+ 1538841.300000ns, VSS,
+ 1538841.400000ns, VDD,
+ 1539321.700000ns, VDD,
+ 1539321.800000ns, VSS,
+ 1539802.100000ns, VSS,
+ 1539802.200000ns, VDD,
+ 1541243.300000ns, VDD,
+ 1541243.400000ns, VSS,
+ 1541963.900000ns, VSS,
+ 1541964.000000ns, VDD,
+ 1542324.200000ns, VDD,
+ 1542324.300000ns, VSS,
+ 1542444.300000ns, VSS,
+ 1542444.400000ns, VDD,
+ 1542804.600000ns, VDD,
+ 1542804.700000ns, VSS,
+ 1542924.700000ns, VSS,
+ 1542924.800000ns, VDD,
+ 1543405.100000ns, VDD,
+ 1543405.200000ns, VSS,
+ 1543885.500000ns, VSS,
+ 1543885.600000ns, VDD,
+ 1544245.800000ns, VDD,
+ 1544245.900000ns, VSS,
+ 1545086.500000ns, VSS,
+ 1545086.600000ns, VDD,
+ 1545326.700000ns, VDD,
+ 1545326.800000ns, VSS,
+ 1545807.100000ns, VSS,
+ 1545807.200000ns, VDD,
+ 1547008.100000ns, VDD,
+ 1547008.200000ns, VSS,
+ 1547368.400000ns, VSS,
+ 1547368.500000ns, VDD,
+ 1547728.700000ns, VDD,
+ 1547728.800000ns, VSS,
+ 1547968.900000ns, VSS,
+ 1547969.000000ns, VDD,
+ 1548089.000000ns, VDD,
+ 1548089.100000ns, VSS,
+ 1548929.700000ns, VSS,
+ 1548929.800000ns, VDD,
+ 1549049.800000ns, VDD,
+ 1549049.900000ns, VSS,
+ 1549169.900000ns, VSS,
+ 1549170.000000ns, VDD,
+ 1550130.700000ns, VDD,
+ 1550130.800000ns, VSS
+)}


RCDN in_CDN 0 1.0
BCDN in_CDN 0 V={table(time,
+ 0.100000ns, VSS,
+ 840.700000ns, VSS,
+ 840.800000ns, VDD,
+ 960.800000ns, VDD,
+ 960.900000ns, VSS,
+ 1921.600000ns, VSS,
+ 1921.700000ns, VDD,
+ 2402.000000ns, VDD,
+ 2402.100000ns, VSS,
+ 2642.200000ns, VSS,
+ 2642.300000ns, VDD,
+ 2762.300000ns, VDD,
+ 2762.400000ns, VSS,
+ 3002.500000ns, VSS,
+ 3002.600000ns, VDD,
+ 3362.800000ns, VDD,
+ 3362.900000ns, VSS,
+ 3843.200000ns, VSS,
+ 3843.300000ns, VDD,
+ 4083.400000ns, VDD,
+ 4083.500000ns, VSS,
+ 4323.600000ns, VSS,
+ 4323.700000ns, VDD,
+ 4443.700000ns, VDD,
+ 4443.800000ns, VSS,
+ 4563.800000ns, VSS,
+ 4563.900000ns, VDD,
+ 4804.000000ns, VDD,
+ 4804.100000ns, VSS,
+ 5044.200000ns, VSS,
+ 5044.300000ns, VDD,
+ 5644.700000ns, VDD,
+ 5644.800000ns, VSS,
+ 5884.900000ns, VSS,
+ 5885.000000ns, VDD,
+ 6005.000000ns, VDD,
+ 6005.100000ns, VSS,
+ 6365.300000ns, VSS,
+ 6365.400000ns, VDD,
+ 6845.700000ns, VDD,
+ 6845.800000ns, VSS,
+ 7326.100000ns, VSS,
+ 7326.200000ns, VDD,
+ 7446.200000ns, VDD,
+ 7446.300000ns, VSS,
+ 8286.900000ns, VSS,
+ 8287.000000ns, VDD,
+ 8527.100000ns, VDD,
+ 8527.200000ns, VSS,
+ 8647.200000ns, VSS,
+ 8647.300000ns, VDD,
+ 9127.600000ns, VDD,
+ 9127.700000ns, VSS,
+ 9367.800000ns, VSS,
+ 9367.900000ns, VDD,
+ 9608.000000ns, VDD,
+ 9608.100000ns, VSS,
+ 9968.300000ns, VSS,
+ 9968.400000ns, VDD,
+ 10088.400000ns, VDD,
+ 10088.500000ns, VSS,
+ 10568.800000ns, VSS,
+ 10568.900000ns, VDD,
+ 10929.100000ns, VDD,
+ 10929.200000ns, VSS,
+ 11169.300000ns, VSS,
+ 11169.400000ns, VDD,
+ 11769.800000ns, VDD,
+ 11769.900000ns, VSS,
+ 12490.400000ns, VSS,
+ 12490.500000ns, VDD,
+ 12850.700000ns, VDD,
+ 12850.800000ns, VSS,
+ 13691.400000ns, VSS,
+ 13691.500000ns, VDD,
+ 15492.900000ns, VDD,
+ 15493.000000ns, VSS,
+ 15613.000000ns, VSS,
+ 15613.100000ns, VDD,
+ 16453.700000ns, VDD,
+ 16453.800000ns, VSS,
+ 16573.800000ns, VSS,
+ 16573.900000ns, VDD,
+ 17534.600000ns, VDD,
+ 17534.700000ns, VSS,
+ 17654.700000ns, VSS,
+ 17654.800000ns, VDD,
+ 18855.700000ns, VDD,
+ 18855.800000ns, VSS,
+ 20056.700000ns, VSS,
+ 20056.800000ns, VDD,
+ 20176.800000ns, VDD,
+ 20176.900000ns, VSS,
+ 20417.000000ns, VSS,
+ 20417.100000ns, VDD,
+ 20657.200000ns, VDD,
+ 20657.300000ns, VSS,
+ 21137.600000ns, VSS,
+ 21137.700000ns, VDD,
+ 21497.900000ns, VDD,
+ 21498.000000ns, VSS,
+ 22218.500000ns, VSS,
+ 22218.600000ns, VDD,
+ 22819.000000ns, VDD,
+ 22819.100000ns, VSS,
+ 23419.500000ns, VSS,
+ 23419.600000ns, VDD,
+ 23779.800000ns, VDD,
+ 23779.900000ns, VSS,
+ 24020.000000ns, VSS,
+ 24020.100000ns, VDD,
+ 24380.300000ns, VDD,
+ 24380.400000ns, VSS,
+ 25341.100000ns, VSS,
+ 25341.200000ns, VDD,
+ 25701.400000ns, VDD,
+ 25701.500000ns, VSS,
+ 25941.600000ns, VSS,
+ 25941.700000ns, VDD,
+ 26422.000000ns, VDD,
+ 26422.100000ns, VSS,
+ 27502.900000ns, VSS,
+ 27503.000000ns, VDD,
+ 27743.100000ns, VDD,
+ 27743.200000ns, VSS,
+ 27863.200000ns, VSS,
+ 27863.300000ns, VDD,
+ 27983.300000ns, VDD,
+ 27983.400000ns, VSS,
+ 28583.800000ns, VSS,
+ 28583.900000ns, VDD,
+ 29304.400000ns, VDD,
+ 29304.500000ns, VSS,
+ 29664.700000ns, VSS,
+ 29664.800000ns, VDD,
+ 29904.900000ns, VDD,
+ 29905.000000ns, VSS,
+ 30145.100000ns, VSS,
+ 30145.200000ns, VDD,
+ 30625.500000ns, VDD,
+ 30625.600000ns, VSS,
+ 31105.900000ns, VSS,
+ 31106.000000ns, VDD,
+ 31466.200000ns, VDD,
+ 31466.300000ns, VSS,
+ 31586.300000ns, VSS,
+ 31586.400000ns, VDD,
+ 31826.500000ns, VDD,
+ 31826.600000ns, VSS,
+ 31946.600000ns, VSS,
+ 31946.700000ns, VDD,
+ 32186.800000ns, VDD,
+ 32186.900000ns, VSS,
+ 32547.100000ns, VSS,
+ 32547.200000ns, VDD,
+ 32667.200000ns, VDD,
+ 32667.300000ns, VSS,
+ 33748.100000ns, VSS,
+ 33748.200000ns, VDD,
+ 34468.700000ns, VDD,
+ 34468.800000ns, VSS,
+ 35069.200000ns, VSS,
+ 35069.300000ns, VDD,
+ 35789.800000ns, VDD,
+ 35789.900000ns, VSS,
+ 35909.900000ns, VSS,
+ 35910.000000ns, VDD,
+ 36030.000000ns, VDD,
+ 36030.100000ns, VSS,
+ 36390.300000ns, VSS,
+ 36390.400000ns, VDD,
+ 38311.900000ns, VDD,
+ 38312.000000ns, VSS,
+ 39032.500000ns, VSS,
+ 39032.600000ns, VDD,
+ 39272.700000ns, VDD,
+ 39272.800000ns, VSS,
+ 40353.600000ns, VSS,
+ 40353.700000ns, VDD,
+ 40473.700000ns, VDD,
+ 40473.800000ns, VSS,
+ 40593.800000ns, VSS,
+ 40593.900000ns, VDD,
+ 41074.200000ns, VDD,
+ 41074.300000ns, VSS,
+ 41434.500000ns, VSS,
+ 41434.600000ns, VDD,
+ 41554.600000ns, VDD,
+ 41554.700000ns, VSS,
+ 42035.000000ns, VSS,
+ 42035.100000ns, VDD,
+ 42155.100000ns, VDD,
+ 42155.200000ns, VSS,
+ 42395.300000ns, VSS,
+ 42395.400000ns, VDD,
+ 42515.400000ns, VDD,
+ 42515.500000ns, VSS,
+ 43115.900000ns, VSS,
+ 43116.000000ns, VDD,
+ 43476.200000ns, VDD,
+ 43476.300000ns, VSS,
+ 43596.300000ns, VSS,
+ 43596.400000ns, VDD,
+ 44076.700000ns, VDD,
+ 44076.800000ns, VSS,
+ 44557.100000ns, VSS,
+ 44557.200000ns, VDD,
+ 44917.400000ns, VDD,
+ 44917.500000ns, VSS,
+ 45037.500000ns, VSS,
+ 45037.600000ns, VDD,
+ 45277.700000ns, VDD,
+ 45277.800000ns, VSS,
+ 46118.400000ns, VSS,
+ 46118.500000ns, VDD,
+ 46598.800000ns, VDD,
+ 46598.900000ns, VSS,
+ 46959.100000ns, VSS,
+ 46959.200000ns, VDD,
+ 47319.400000ns, VDD,
+ 47319.500000ns, VSS,
+ 47439.500000ns, VSS,
+ 47439.600000ns, VDD,
+ 47919.900000ns, VDD,
+ 47920.000000ns, VSS,
+ 48160.100000ns, VSS,
+ 48160.200000ns, VDD,
+ 48280.200000ns, VDD,
+ 48280.300000ns, VSS,
+ 48400.300000ns, VSS,
+ 48400.400000ns, VDD,
+ 49601.300000ns, VDD,
+ 49601.400000ns, VSS,
+ 49721.400000ns, VSS,
+ 49721.500000ns, VDD,
+ 50442.000000ns, VDD,
+ 50442.100000ns, VSS,
+ 50562.100000ns, VSS,
+ 50562.200000ns, VDD,
+ 51282.700000ns, VDD,
+ 51282.800000ns, VSS,
+ 51883.200000ns, VSS,
+ 51883.300000ns, VDD,
+ 52003.300000ns, VDD,
+ 52003.400000ns, VSS,
+ 52483.700000ns, VSS,
+ 52483.800000ns, VDD,
+ 52723.900000ns, VDD,
+ 52724.000000ns, VSS,
+ 53444.500000ns, VSS,
+ 53444.600000ns, VDD,
+ 54405.300000ns, VDD,
+ 54405.400000ns, VSS,
+ 54765.600000ns, VSS,
+ 54765.700000ns, VDD,
+ 55966.600000ns, VDD,
+ 55966.700000ns, VSS,
+ 56567.100000ns, VSS,
+ 56567.200000ns, VDD,
+ 56687.200000ns, VDD,
+ 56687.300000ns, VSS,
+ 57047.500000ns, VSS,
+ 57047.600000ns, VDD,
+ 57167.600000ns, VDD,
+ 57167.700000ns, VSS,
+ 57527.900000ns, VSS,
+ 57528.000000ns, VDD,
+ 57888.200000ns, VDD,
+ 57888.300000ns, VSS,
+ 58008.300000ns, VSS,
+ 58008.400000ns, VDD,
+ 58248.500000ns, VDD,
+ 58248.600000ns, VSS,
+ 58728.900000ns, VSS,
+ 58729.000000ns, VDD,
+ 59209.300000ns, VDD,
+ 59209.400000ns, VSS,
+ 59689.700000ns, VSS,
+ 59689.800000ns, VDD,
+ 59929.900000ns, VDD,
+ 59930.000000ns, VSS,
+ 60050.000000ns, VSS,
+ 60050.100000ns, VDD,
+ 60170.100000ns, VDD,
+ 60170.200000ns, VSS,
+ 61130.900000ns, VSS,
+ 61131.000000ns, VDD,
+ 61371.100000ns, VDD,
+ 61371.200000ns, VSS,
+ 61851.500000ns, VSS,
+ 61851.600000ns, VDD,
+ 62211.800000ns, VDD,
+ 62211.900000ns, VSS,
+ 62572.100000ns, VSS,
+ 62572.200000ns, VDD,
+ 62812.300000ns, VDD,
+ 62812.400000ns, VSS,
+ 63412.800000ns, VSS,
+ 63412.900000ns, VDD,
+ 63893.200000ns, VDD,
+ 63893.300000ns, VSS,
+ 64493.700000ns, VSS,
+ 64493.800000ns, VDD,
+ 64854.000000ns, VDD,
+ 64854.100000ns, VSS,
+ 65094.200000ns, VSS,
+ 65094.300000ns, VDD,
+ 65574.600000ns, VDD,
+ 65574.700000ns, VSS,
+ 66655.500000ns, VSS,
+ 66655.600000ns, VDD,
+ 66895.700000ns, VDD,
+ 66895.800000ns, VSS,
+ 67135.900000ns, VSS,
+ 67136.000000ns, VDD,
+ 68096.700000ns, VDD,
+ 68096.800000ns, VSS,
+ 68336.900000ns, VSS,
+ 68337.000000ns, VDD,
+ 68457.000000ns, VDD,
+ 68457.100000ns, VSS,
+ 68697.200000ns, VSS,
+ 68697.300000ns, VDD,
+ 68937.400000ns, VDD,
+ 68937.500000ns, VSS,
+ 69417.800000ns, VSS,
+ 69417.900000ns, VDD,
+ 69898.200000ns, VDD,
+ 69898.300000ns, VSS,
+ 70138.400000ns, VSS,
+ 70138.500000ns, VDD,
+ 70618.800000ns, VDD,
+ 70618.900000ns, VSS,
+ 71219.300000ns, VSS,
+ 71219.400000ns, VDD,
+ 71699.700000ns, VDD,
+ 71699.800000ns, VSS,
+ 72180.100000ns, VSS,
+ 72180.200000ns, VDD,
+ 72660.500000ns, VDD,
+ 72660.600000ns, VSS,
+ 73140.900000ns, VSS,
+ 73141.000000ns, VDD,
+ 73381.100000ns, VDD,
+ 73381.200000ns, VSS,
+ 73981.600000ns, VSS,
+ 73981.700000ns, VDD,
+ 74341.900000ns, VDD,
+ 74342.000000ns, VSS,
+ 74462.000000ns, VSS,
+ 74462.100000ns, VDD,
+ 75062.500000ns, VDD,
+ 75062.600000ns, VSS,
+ 75903.200000ns, VSS,
+ 75903.300000ns, VDD,
+ 76143.400000ns, VDD,
+ 76143.500000ns, VSS,
+ 76503.700000ns, VSS,
+ 76503.800000ns, VDD,
+ 76623.800000ns, VDD,
+ 76623.900000ns, VSS,
+ 77104.200000ns, VSS,
+ 77104.300000ns, VDD,
+ 77824.800000ns, VDD,
+ 77824.900000ns, VSS,
+ 78065.000000ns, VSS,
+ 78065.100000ns, VDD,
+ 78185.100000ns, VDD,
+ 78185.200000ns, VSS,
+ 78305.200000ns, VSS,
+ 78305.300000ns, VDD,
+ 79266.000000ns, VDD,
+ 79266.100000ns, VSS,
+ 79746.400000ns, VSS,
+ 79746.500000ns, VDD,
+ 80106.700000ns, VDD,
+ 80106.800000ns, VSS,
+ 80827.300000ns, VSS,
+ 80827.400000ns, VDD,
+ 81427.800000ns, VDD,
+ 81427.900000ns, VSS,
+ 81668.000000ns, VSS,
+ 81668.100000ns, VDD,
+ 81788.100000ns, VDD,
+ 81788.200000ns, VSS,
+ 81908.200000ns, VSS,
+ 81908.300000ns, VDD,
+ 82148.400000ns, VDD,
+ 82148.500000ns, VSS,
+ 82268.500000ns, VSS,
+ 82268.600000ns, VDD,
+ 82388.600000ns, VDD,
+ 82388.700000ns, VSS,
+ 82508.700000ns, VSS,
+ 82508.800000ns, VDD,
+ 82748.900000ns, VDD,
+ 82749.000000ns, VSS,
+ 83469.500000ns, VSS,
+ 83469.600000ns, VDD,
+ 83829.800000ns, VDD,
+ 83829.900000ns, VSS,
+ 84070.000000ns, VSS,
+ 84070.100000ns, VDD,
+ 84310.200000ns, VDD,
+ 84310.300000ns, VSS,
+ 84790.600000ns, VSS,
+ 84790.700000ns, VDD,
+ 85271.000000ns, VDD,
+ 85271.100000ns, VSS,
+ 85511.200000ns, VSS,
+ 85511.300000ns, VDD,
+ 85751.400000ns, VDD,
+ 85751.500000ns, VSS,
+ 86111.700000ns, VSS,
+ 86111.800000ns, VDD,
+ 86351.900000ns, VDD,
+ 86352.000000ns, VSS,
+ 87312.700000ns, VSS,
+ 87312.800000ns, VDD,
+ 87913.200000ns, VDD,
+ 87913.300000ns, VSS,
+ 88033.300000ns, VSS,
+ 88033.400000ns, VDD,
+ 88273.500000ns, VDD,
+ 88273.600000ns, VSS,
+ 88393.600000ns, VSS,
+ 88393.700000ns, VDD,
+ 88874.000000ns, VDD,
+ 88874.100000ns, VSS,
+ 88994.100000ns, VSS,
+ 88994.200000ns, VDD,
+ 89354.400000ns, VDD,
+ 89354.500000ns, VSS,
+ 89474.500000ns, VSS,
+ 89474.600000ns, VDD,
+ 89714.700000ns, VDD,
+ 89714.800000ns, VSS,
+ 91516.200000ns, VSS,
+ 91516.300000ns, VDD,
+ 91876.500000ns, VDD,
+ 91876.600000ns, VSS,
+ 91996.600000ns, VSS,
+ 91996.700000ns, VDD,
+ 92356.900000ns, VDD,
+ 92357.000000ns, VSS,
+ 92957.400000ns, VSS,
+ 92957.500000ns, VDD,
+ 93557.900000ns, VDD,
+ 93558.000000ns, VSS,
+ 93798.100000ns, VSS,
+ 93798.200000ns, VDD,
+ 94278.500000ns, VDD,
+ 94278.600000ns, VSS,
+ 94398.600000ns, VSS,
+ 94398.700000ns, VDD,
+ 95719.700000ns, VDD,
+ 95719.800000ns, VSS,
+ 95959.900000ns, VSS,
+ 95960.000000ns, VDD,
+ 96200.100000ns, VDD,
+ 96200.200000ns, VSS,
+ 96320.200000ns, VSS,
+ 96320.300000ns, VDD,
+ 96680.500000ns, VDD,
+ 96680.600000ns, VSS,
+ 97160.900000ns, VSS,
+ 97161.000000ns, VDD,
+ 98001.600000ns, VDD,
+ 98001.700000ns, VSS,
+ 98121.700000ns, VSS,
+ 98121.800000ns, VDD,
+ 98241.800000ns, VDD,
+ 98241.900000ns, VSS,
+ 99202.600000ns, VSS,
+ 99202.700000ns, VDD,
+ 99683.000000ns, VDD,
+ 99683.100000ns, VSS,
+ 100163.400000ns, VSS,
+ 100163.500000ns, VDD,
+ 100523.700000ns, VDD,
+ 100523.800000ns, VSS,
+ 100643.800000ns, VSS,
+ 100643.900000ns, VDD,
+ 100763.900000ns, VDD,
+ 100764.000000ns, VSS,
+ 101364.400000ns, VSS,
+ 101364.500000ns, VDD,
+ 101844.800000ns, VDD,
+ 101844.900000ns, VSS,
+ 101964.900000ns, VSS,
+ 101965.000000ns, VDD,
+ 102805.600000ns, VDD,
+ 102805.700000ns, VSS,
+ 103045.800000ns, VSS,
+ 103045.900000ns, VDD,
+ 103286.000000ns, VDD,
+ 103286.100000ns, VSS,
+ 103646.300000ns, VSS,
+ 103646.400000ns, VDD,
+ 104006.600000ns, VDD,
+ 104006.700000ns, VSS,
+ 104847.300000ns, VSS,
+ 104847.400000ns, VDD,
+ 105447.800000ns, VDD,
+ 105447.900000ns, VSS,
+ 105688.000000ns, VSS,
+ 105688.100000ns, VDD,
+ 105808.100000ns, VDD,
+ 105808.200000ns, VSS,
+ 107969.900000ns, VSS,
+ 107970.000000ns, VDD,
+ 108090.000000ns, VDD,
+ 108090.100000ns, VSS,
+ 109651.300000ns, VSS,
+ 109651.400000ns, VDD,
+ 110011.600000ns, VDD,
+ 110011.700000ns, VSS,
+ 110251.800000ns, VSS,
+ 110251.900000ns, VDD,
+ 110732.200000ns, VDD,
+ 110732.300000ns, VSS,
+ 110972.400000ns, VSS,
+ 110972.500000ns, VDD,
+ 111092.500000ns, VDD,
+ 111092.600000ns, VSS,
+ 111332.700000ns, VSS,
+ 111332.800000ns, VDD,
+ 111452.800000ns, VDD,
+ 111452.900000ns, VSS,
+ 111572.900000ns, VSS,
+ 111573.000000ns, VDD,
+ 111813.100000ns, VDD,
+ 111813.200000ns, VSS,
+ 112173.400000ns, VSS,
+ 112173.500000ns, VDD,
+ 112894.000000ns, VDD,
+ 112894.100000ns, VSS,
+ 113014.100000ns, VSS,
+ 113014.200000ns, VDD,
+ 113134.200000ns, VDD,
+ 113134.300000ns, VSS,
+ 113974.900000ns, VSS,
+ 113975.000000ns, VDD,
+ 114215.100000ns, VDD,
+ 114215.200000ns, VSS,
+ 115055.800000ns, VSS,
+ 115055.900000ns, VDD,
+ 115536.200000ns, VDD,
+ 115536.300000ns, VSS,
+ 116016.600000ns, VSS,
+ 116016.700000ns, VDD,
+ 116136.700000ns, VDD,
+ 116136.800000ns, VSS,
+ 116256.800000ns, VSS,
+ 116256.900000ns, VDD,
+ 116737.200000ns, VDD,
+ 116737.300000ns, VSS,
+ 117217.600000ns, VSS,
+ 117217.700000ns, VDD,
+ 117818.100000ns, VDD,
+ 117818.200000ns, VSS,
+ 118178.400000ns, VSS,
+ 118178.500000ns, VDD,
+ 118418.600000ns, VDD,
+ 118418.700000ns, VSS,
+ 119619.600000ns, VSS,
+ 119619.700000ns, VDD,
+ 119859.800000ns, VDD,
+ 119859.900000ns, VSS,
+ 119979.900000ns, VSS,
+ 119980.000000ns, VDD,
+ 120100.000000ns, VDD,
+ 120100.100000ns, VSS,
+ 120340.200000ns, VSS,
+ 120340.300000ns, VDD,
+ 120580.400000ns, VDD,
+ 120580.500000ns, VSS,
+ 120940.700000ns, VSS,
+ 120940.800000ns, VDD,
+ 121541.200000ns, VDD,
+ 121541.300000ns, VSS,
+ 122021.600000ns, VSS,
+ 122021.700000ns, VDD,
+ 122381.900000ns, VDD,
+ 122382.000000ns, VSS,
+ 122622.100000ns, VSS,
+ 122622.200000ns, VDD,
+ 122742.200000ns, VDD,
+ 122742.300000ns, VSS,
+ 123342.700000ns, VSS,
+ 123342.800000ns, VDD,
+ 123703.000000ns, VDD,
+ 123703.100000ns, VSS,
+ 124183.400000ns, VSS,
+ 124183.500000ns, VDD,
+ 124663.800000ns, VDD,
+ 124663.900000ns, VSS,
+ 124904.000000ns, VSS,
+ 124904.100000ns, VDD,
+ 125024.100000ns, VDD,
+ 125024.200000ns, VSS,
+ 125144.200000ns, VSS,
+ 125144.300000ns, VDD,
+ 125504.500000ns, VDD,
+ 125504.600000ns, VSS,
+ 126225.100000ns, VSS,
+ 126225.200000ns, VDD,
+ 128026.600000ns, VDD,
+ 128026.700000ns, VSS,
+ 128867.300000ns, VSS,
+ 128867.400000ns, VDD,
+ 129107.500000ns, VDD,
+ 129107.600000ns, VSS,
+ 129347.700000ns, VSS,
+ 129347.800000ns, VDD,
+ 129587.900000ns, VDD,
+ 129588.000000ns, VSS,
+ 129828.100000ns, VSS,
+ 129828.200000ns, VDD,
+ 130188.400000ns, VDD,
+ 130188.500000ns, VSS,
+ 130428.600000ns, VSS,
+ 130428.700000ns, VDD,
+ 130548.700000ns, VDD,
+ 130548.800000ns, VSS,
+ 130668.800000ns, VSS,
+ 130668.900000ns, VDD,
+ 131389.400000ns, VDD,
+ 131389.500000ns, VSS,
+ 131989.900000ns, VSS,
+ 131990.000000ns, VDD,
+ 132710.500000ns, VDD,
+ 132710.600000ns, VSS,
+ 132830.600000ns, VSS,
+ 132830.700000ns, VDD,
+ 133311.000000ns, VDD,
+ 133311.100000ns, VSS,
+ 133671.300000ns, VSS,
+ 133671.400000ns, VDD,
+ 133791.400000ns, VDD,
+ 133791.500000ns, VSS,
+ 134512.000000ns, VSS,
+ 134512.100000ns, VDD,
+ 134992.400000ns, VDD,
+ 134992.500000ns, VSS,
+ 135592.900000ns, VSS,
+ 135593.000000ns, VDD,
+ 135713.000000ns, VDD,
+ 135713.100000ns, VSS,
+ 136073.300000ns, VSS,
+ 136073.400000ns, VDD,
+ 136433.600000ns, VDD,
+ 136433.700000ns, VSS,
+ 137034.100000ns, VSS,
+ 137034.200000ns, VDD,
+ 137274.300000ns, VDD,
+ 137274.400000ns, VSS,
+ 137634.600000ns, VSS,
+ 137634.700000ns, VDD,
+ 137874.800000ns, VDD,
+ 137874.900000ns, VSS,
+ 138355.200000ns, VSS,
+ 138355.300000ns, VDD,
+ 139556.200000ns, VDD,
+ 139556.300000ns, VSS,
+ 139676.300000ns, VSS,
+ 139676.400000ns, VDD,
+ 140156.700000ns, VDD,
+ 140156.800000ns, VSS,
+ 140637.100000ns, VSS,
+ 140637.200000ns, VDD,
+ 141237.600000ns, VDD,
+ 141237.700000ns, VSS,
+ 141357.700000ns, VSS,
+ 141357.800000ns, VDD,
+ 141477.800000ns, VDD,
+ 141477.900000ns, VSS,
+ 141597.900000ns, VSS,
+ 141598.000000ns, VDD,
+ 141838.100000ns, VDD,
+ 141838.200000ns, VSS,
+ 141958.200000ns, VSS,
+ 141958.300000ns, VDD,
+ 142318.500000ns, VDD,
+ 142318.600000ns, VSS,
+ 142558.700000ns, VSS,
+ 142558.800000ns, VDD,
+ 143039.100000ns, VDD,
+ 143039.200000ns, VSS,
+ 143639.600000ns, VSS,
+ 143639.700000ns, VDD,
+ 143879.800000ns, VDD,
+ 143879.900000ns, VSS,
+ 144120.000000ns, VSS,
+ 144120.100000ns, VDD,
+ 144240.100000ns, VDD,
+ 144240.200000ns, VSS,
+ 144720.500000ns, VSS,
+ 144720.600000ns, VDD,
+ 145321.000000ns, VDD,
+ 145321.100000ns, VSS,
+ 145441.100000ns, VSS,
+ 145441.200000ns, VDD,
+ 145801.400000ns, VDD,
+ 145801.500000ns, VSS,
+ 146161.700000ns, VSS,
+ 146161.800000ns, VDD,
+ 147002.400000ns, VDD,
+ 147002.500000ns, VSS,
+ 147122.500000ns, VSS,
+ 147122.600000ns, VDD,
+ 147242.600000ns, VDD,
+ 147242.700000ns, VSS,
+ 148083.300000ns, VSS,
+ 148083.400000ns, VDD,
+ 149404.400000ns, VDD,
+ 149404.500000ns, VSS,
+ 149644.600000ns, VSS,
+ 149644.700000ns, VDD,
+ 150125.000000ns, VDD,
+ 150125.100000ns, VSS,
+ 150485.300000ns, VSS,
+ 150485.400000ns, VDD,
+ 151326.000000ns, VDD,
+ 151326.100000ns, VSS,
+ 151446.100000ns, VSS,
+ 151446.200000ns, VDD,
+ 152286.800000ns, VDD,
+ 152286.900000ns, VSS,
+ 152887.300000ns, VSS,
+ 152887.400000ns, VDD,
+ 153607.900000ns, VDD,
+ 153608.000000ns, VSS,
+ 154208.400000ns, VSS,
+ 154208.500000ns, VDD,
+ 154688.800000ns, VDD,
+ 154688.900000ns, VSS,
+ 154929.000000ns, VSS,
+ 154929.100000ns, VDD,
+ 157811.400000ns, VDD,
+ 157811.500000ns, VSS,
+ 159252.600000ns, VSS,
+ 159252.700000ns, VDD,
+ 159973.200000ns, VDD,
+ 159973.300000ns, VSS,
+ 160213.400000ns, VSS,
+ 160213.500000ns, VDD,
+ 160693.800000ns, VDD,
+ 160693.900000ns, VSS,
+ 161174.200000ns, VSS,
+ 161174.300000ns, VDD,
+ 161414.400000ns, VDD,
+ 161414.500000ns, VSS,
+ 161534.500000ns, VSS,
+ 161534.600000ns, VDD,
+ 162135.000000ns, VDD,
+ 162135.100000ns, VSS,
+ 162375.200000ns, VSS,
+ 162375.300000ns, VDD,
+ 162975.700000ns, VDD,
+ 162975.800000ns, VSS,
+ 163336.000000ns, VSS,
+ 163336.100000ns, VDD,
+ 164537.000000ns, VDD,
+ 164537.100000ns, VSS,
+ 164657.100000ns, VSS,
+ 164657.200000ns, VDD,
+ 165017.400000ns, VDD,
+ 165017.500000ns, VSS,
+ 165497.800000ns, VSS,
+ 165497.900000ns, VDD,
+ 165858.100000ns, VDD,
+ 165858.200000ns, VSS,
+ 166218.400000ns, VSS,
+ 166218.500000ns, VDD,
+ 166338.500000ns, VDD,
+ 166338.600000ns, VSS,
+ 166578.700000ns, VSS,
+ 166578.800000ns, VDD,
+ 168140.000000ns, VDD,
+ 168140.100000ns, VSS,
+ 168500.300000ns, VSS,
+ 168500.400000ns, VDD,
+ 169100.800000ns, VDD,
+ 169100.900000ns, VSS,
+ 169461.100000ns, VSS,
+ 169461.200000ns, VDD,
+ 169821.400000ns, VDD,
+ 169821.500000ns, VSS,
+ 170061.600000ns, VSS,
+ 170061.700000ns, VDD,
+ 170421.900000ns, VDD,
+ 170422.000000ns, VSS,
+ 170662.100000ns, VSS,
+ 170662.200000ns, VDD,
+ 171142.500000ns, VDD,
+ 171142.600000ns, VSS,
+ 171743.000000ns, VSS,
+ 171743.100000ns, VDD,
+ 171863.100000ns, VDD,
+ 171863.200000ns, VSS,
+ 171983.200000ns, VSS,
+ 171983.300000ns, VDD,
+ 172223.400000ns, VDD,
+ 172223.500000ns, VSS,
+ 172703.800000ns, VSS,
+ 172703.900000ns, VDD,
+ 173064.100000ns, VDD,
+ 173064.200000ns, VSS,
+ 173184.200000ns, VSS,
+ 173184.300000ns, VDD,
+ 174024.900000ns, VDD,
+ 174025.000000ns, VSS,
+ 174505.300000ns, VSS,
+ 174505.400000ns, VDD,
+ 174985.700000ns, VDD,
+ 174985.800000ns, VSS,
+ 175346.000000ns, VSS,
+ 175346.100000ns, VDD,
+ 175946.500000ns, VDD,
+ 175946.600000ns, VSS,
+ 176667.100000ns, VSS,
+ 176667.200000ns, VDD,
+ 176907.300000ns, VDD,
+ 176907.400000ns, VSS,
+ 178708.800000ns, VSS,
+ 178708.900000ns, VDD,
+ 178949.000000ns, VDD,
+ 178949.100000ns, VSS,
+ 179069.100000ns, VSS,
+ 179069.200000ns, VDD,
+ 179549.500000ns, VDD,
+ 179549.600000ns, VSS,
+ 179669.600000ns, VSS,
+ 179669.700000ns, VDD,
+ 180270.100000ns, VDD,
+ 180270.200000ns, VSS,
+ 180390.200000ns, VSS,
+ 180390.300000ns, VDD,
+ 180510.300000ns, VDD,
+ 180510.400000ns, VSS,
+ 180750.500000ns, VSS,
+ 180750.600000ns, VDD,
+ 181471.100000ns, VDD,
+ 181471.200000ns, VSS,
+ 181591.200000ns, VSS,
+ 181591.300000ns, VDD,
+ 181831.400000ns, VDD,
+ 181831.500000ns, VSS,
+ 182311.800000ns, VSS,
+ 182311.900000ns, VDD,
+ 183272.600000ns, VDD,
+ 183272.700000ns, VSS,
+ 183753.000000ns, VSS,
+ 183753.100000ns, VDD,
+ 184113.300000ns, VDD,
+ 184113.400000ns, VSS,
+ 184833.900000ns, VSS,
+ 184834.000000ns, VDD,
+ 185194.200000ns, VDD,
+ 185194.300000ns, VSS,
+ 185314.300000ns, VSS,
+ 185314.400000ns, VDD,
+ 185554.500000ns, VDD,
+ 185554.600000ns, VSS,
+ 185794.700000ns, VSS,
+ 185794.800000ns, VDD,
+ 186155.000000ns, VDD,
+ 186155.100000ns, VSS,
+ 186635.400000ns, VSS,
+ 186635.500000ns, VDD,
+ 186875.600000ns, VDD,
+ 186875.700000ns, VSS,
+ 187476.100000ns, VSS,
+ 187476.200000ns, VDD,
+ 187716.300000ns, VDD,
+ 187716.400000ns, VSS,
+ 187836.400000ns, VSS,
+ 187836.500000ns, VDD,
+ 188196.700000ns, VDD,
+ 188196.800000ns, VSS,
+ 188316.800000ns, VSS,
+ 188316.900000ns, VDD,
+ 188436.900000ns, VDD,
+ 188437.000000ns, VSS,
+ 188557.000000ns, VSS,
+ 188557.100000ns, VDD,
+ 189758.000000ns, VDD,
+ 189758.100000ns, VSS,
+ 190238.400000ns, VSS,
+ 190238.500000ns, VDD,
+ 190598.700000ns, VDD,
+ 190598.800000ns, VSS,
+ 191799.700000ns, VSS,
+ 191799.800000ns, VDD,
+ 192039.900000ns, VDD,
+ 192040.000000ns, VSS,
+ 192280.100000ns, VSS,
+ 192280.200000ns, VDD,
+ 192400.200000ns, VDD,
+ 192400.300000ns, VSS,
+ 192760.500000ns, VSS,
+ 192760.600000ns, VDD,
+ 192880.600000ns, VDD,
+ 192880.700000ns, VSS,
+ 193000.700000ns, VSS,
+ 193000.800000ns, VDD,
+ 193361.000000ns, VDD,
+ 193361.100000ns, VSS,
+ 193841.400000ns, VSS,
+ 193841.500000ns, VDD,
+ 193961.500000ns, VDD,
+ 193961.600000ns, VSS,
+ 194441.900000ns, VSS,
+ 194442.000000ns, VDD,
+ 194682.100000ns, VDD,
+ 194682.200000ns, VSS,
+ 194922.300000ns, VSS,
+ 194922.400000ns, VDD,
+ 195763.000000ns, VDD,
+ 195763.100000ns, VSS,
+ 196243.400000ns, VSS,
+ 196243.500000ns, VDD,
+ 196363.500000ns, VDD,
+ 196363.600000ns, VSS,
+ 196843.900000ns, VSS,
+ 196844.000000ns, VDD,
+ 197084.100000ns, VDD,
+ 197084.200000ns, VSS,
+ 197204.200000ns, VSS,
+ 197204.300000ns, VDD,
+ 197564.500000ns, VDD,
+ 197564.600000ns, VSS,
+ 197684.600000ns, VSS,
+ 197684.700000ns, VDD,
+ 197804.700000ns, VDD,
+ 197804.800000ns, VSS,
+ 198165.000000ns, VSS,
+ 198165.100000ns, VDD,
+ 198645.400000ns, VDD,
+ 198645.500000ns, VSS,
+ 198765.500000ns, VSS,
+ 198765.600000ns, VDD,
+ 199005.700000ns, VDD,
+ 199005.800000ns, VSS,
+ 199125.800000ns, VSS,
+ 199125.900000ns, VDD,
+ 199245.900000ns, VDD,
+ 199246.000000ns, VSS,
+ 200086.600000ns, VSS,
+ 200086.700000ns, VDD,
+ 200807.200000ns, VDD,
+ 200807.300000ns, VSS,
+ 200927.300000ns, VSS,
+ 200927.400000ns, VDD,
+ 201768.000000ns, VDD,
+ 201768.100000ns, VSS,
+ 202008.200000ns, VSS,
+ 202008.300000ns, VDD,
+ 202368.500000ns, VDD,
+ 202368.600000ns, VSS,
+ 202608.700000ns, VSS,
+ 202608.800000ns, VDD,
+ 203569.500000ns, VDD,
+ 203569.600000ns, VSS,
+ 203929.800000ns, VSS,
+ 203929.900000ns, VDD,
+ 206211.700000ns, VDD,
+ 206211.800000ns, VSS,
+ 206331.800000ns, VSS,
+ 206331.900000ns, VDD,
+ 206451.900000ns, VDD,
+ 206452.000000ns, VSS,
+ 206932.300000ns, VSS,
+ 206932.400000ns, VDD,
+ 207893.100000ns, VDD,
+ 207893.200000ns, VSS,
+ 208253.400000ns, VSS,
+ 208253.500000ns, VDD,
+ 208493.600000ns, VDD,
+ 208493.700000ns, VSS,
+ 209334.300000ns, VSS,
+ 209334.400000ns, VDD,
+ 209574.500000ns, VDD,
+ 209574.600000ns, VSS,
+ 210295.100000ns, VSS,
+ 210295.200000ns, VDD,
+ 210655.400000ns, VDD,
+ 210655.500000ns, VSS,
+ 210775.500000ns, VSS,
+ 210775.600000ns, VDD,
+ 211135.800000ns, VDD,
+ 211135.900000ns, VSS,
+ 211496.100000ns, VSS,
+ 211496.200000ns, VDD,
+ 211856.400000ns, VDD,
+ 211856.500000ns, VSS,
+ 212096.600000ns, VSS,
+ 212096.700000ns, VDD,
+ 213177.500000ns, VDD,
+ 213177.600000ns, VSS,
+ 213417.700000ns, VSS,
+ 213417.800000ns, VDD,
+ 213537.800000ns, VDD,
+ 213537.900000ns, VSS,
+ 213898.100000ns, VSS,
+ 213898.200000ns, VDD,
+ 214378.500000ns, VDD,
+ 214378.600000ns, VSS,
+ 214618.700000ns, VSS,
+ 214618.800000ns, VDD,
+ 214858.900000ns, VDD,
+ 214859.000000ns, VSS,
+ 215219.200000ns, VSS,
+ 215219.300000ns, VDD,
+ 215939.800000ns, VDD,
+ 215939.900000ns, VSS,
+ 216059.900000ns, VSS,
+ 216060.000000ns, VDD,
+ 217020.700000ns, VDD,
+ 217020.800000ns, VSS,
+ 217381.000000ns, VSS,
+ 217381.100000ns, VDD,
+ 217741.300000ns, VDD,
+ 217741.400000ns, VSS,
+ 217861.400000ns, VSS,
+ 217861.500000ns, VDD,
+ 218341.800000ns, VDD,
+ 218341.900000ns, VSS,
+ 218702.100000ns, VSS,
+ 218702.200000ns, VDD,
+ 219062.400000ns, VDD,
+ 219062.500000ns, VSS,
+ 219182.500000ns, VSS,
+ 219182.600000ns, VDD,
+ 219422.700000ns, VDD,
+ 219422.800000ns, VSS,
+ 219783.000000ns, VSS,
+ 219783.100000ns, VDD,
+ 219903.100000ns, VDD,
+ 219903.200000ns, VSS,
+ 220863.900000ns, VSS,
+ 220864.000000ns, VDD,
+ 221224.200000ns, VDD,
+ 221224.300000ns, VSS,
+ 221464.400000ns, VSS,
+ 221464.500000ns, VDD,
+ 221584.500000ns, VDD,
+ 221584.600000ns, VSS,
+ 221704.600000ns, VSS,
+ 221704.700000ns, VDD,
+ 222305.100000ns, VDD,
+ 222305.200000ns, VSS,
+ 223866.400000ns, VSS,
+ 223866.500000ns, VDD,
+ 224226.700000ns, VDD,
+ 224226.800000ns, VSS,
+ 224346.800000ns, VSS,
+ 224346.900000ns, VDD,
+ 224466.900000ns, VDD,
+ 224467.000000ns, VSS,
+ 224587.000000ns, VSS,
+ 224587.100000ns, VDD,
+ 225908.100000ns, VDD,
+ 225908.200000ns, VSS,
+ 226148.300000ns, VSS,
+ 226148.400000ns, VDD,
+ 226508.600000ns, VDD,
+ 226508.700000ns, VSS,
+ 226628.700000ns, VSS,
+ 226628.800000ns, VDD,
+ 227109.100000ns, VDD,
+ 227109.200000ns, VSS,
+ 227469.400000ns, VSS,
+ 227469.500000ns, VDD,
+ 227949.800000ns, VDD,
+ 227949.900000ns, VSS,
+ 228550.300000ns, VSS,
+ 228550.400000ns, VDD,
+ 229150.800000ns, VDD,
+ 229150.900000ns, VSS,
+ 229631.200000ns, VSS,
+ 229631.300000ns, VDD,
+ 230111.600000ns, VDD,
+ 230111.700000ns, VSS,
+ 230231.700000ns, VSS,
+ 230231.800000ns, VDD,
+ 230592.000000ns, VDD,
+ 230592.100000ns, VSS,
+ 230712.100000ns, VSS,
+ 230712.200000ns, VDD,
+ 231192.500000ns, VDD,
+ 231192.600000ns, VSS,
+ 231432.700000ns, VSS,
+ 231432.800000ns, VDD,
+ 231552.800000ns, VDD,
+ 231552.900000ns, VSS,
+ 232513.600000ns, VSS,
+ 232513.700000ns, VDD,
+ 232633.700000ns, VDD,
+ 232633.800000ns, VSS,
+ 233234.200000ns, VSS,
+ 233234.300000ns, VDD,
+ 233474.400000ns, VDD,
+ 233474.500000ns, VSS,
+ 233594.500000ns, VSS,
+ 233594.600000ns, VDD,
+ 233714.600000ns, VDD,
+ 233714.700000ns, VSS,
+ 234315.100000ns, VSS,
+ 234315.200000ns, VDD,
+ 234435.200000ns, VDD,
+ 234435.300000ns, VSS,
+ 234675.400000ns, VSS,
+ 234675.500000ns, VDD,
+ 234795.500000ns, VDD,
+ 234795.600000ns, VSS,
+ 235275.900000ns, VSS,
+ 235276.000000ns, VDD,
+ 235516.100000ns, VDD,
+ 235516.200000ns, VSS,
+ 236236.700000ns, VSS,
+ 236236.800000ns, VDD,
+ 236476.900000ns, VDD,
+ 236477.000000ns, VSS,
+ 237677.900000ns, VSS,
+ 237678.000000ns, VDD,
+ 238398.500000ns, VDD,
+ 238398.600000ns, VSS,
+ 238518.600000ns, VSS,
+ 238518.700000ns, VDD,
+ 238638.700000ns, VDD,
+ 238638.800000ns, VSS,
+ 239119.100000ns, VSS,
+ 239119.200000ns, VDD,
+ 239239.200000ns, VDD,
+ 239239.300000ns, VSS,
+ 239839.700000ns, VSS,
+ 239839.800000ns, VDD,
+ 240800.500000ns, VDD,
+ 240800.600000ns, VSS,
+ 241761.300000ns, VSS,
+ 241761.400000ns, VDD,
+ 242361.800000ns, VDD,
+ 242361.900000ns, VSS,
+ 242602.000000ns, VSS,
+ 242602.100000ns, VDD,
+ 244043.200000ns, VDD,
+ 244043.300000ns, VSS,
+ 244163.300000ns, VSS,
+ 244163.400000ns, VDD,
+ 244523.600000ns, VDD,
+ 244523.700000ns, VSS,
+ 244643.700000ns, VSS,
+ 244643.800000ns, VDD,
+ 245124.100000ns, VDD,
+ 245124.200000ns, VSS,
+ 245364.300000ns, VSS,
+ 245364.400000ns, VDD,
+ 245484.400000ns, VDD,
+ 245484.500000ns, VSS,
+ 245844.700000ns, VSS,
+ 245844.800000ns, VDD,
+ 246565.300000ns, VDD,
+ 246565.400000ns, VSS,
+ 247165.800000ns, VSS,
+ 247165.900000ns, VDD,
+ 247526.100000ns, VDD,
+ 247526.200000ns, VSS,
+ 247646.200000ns, VSS,
+ 247646.300000ns, VDD,
+ 248126.600000ns, VDD,
+ 248126.700000ns, VSS,
+ 248486.900000ns, VSS,
+ 248487.000000ns, VDD,
+ 249327.600000ns, VDD,
+ 249327.700000ns, VSS,
+ 249687.900000ns, VSS,
+ 249688.000000ns, VDD,
+ 250288.400000ns, VDD,
+ 250288.500000ns, VSS,
+ 250408.500000ns, VSS,
+ 250408.600000ns, VDD,
+ 250648.700000ns, VDD,
+ 250648.800000ns, VSS,
+ 251009.000000ns, VSS,
+ 251009.100000ns, VDD,
+ 253050.700000ns, VDD,
+ 253050.800000ns, VSS,
+ 254131.600000ns, VSS,
+ 254131.700000ns, VDD,
+ 254371.800000ns, VDD,
+ 254371.900000ns, VSS,
+ 254732.100000ns, VSS,
+ 254732.200000ns, VDD,
+ 255692.900000ns, VDD,
+ 255693.000000ns, VSS,
+ 255813.000000ns, VSS,
+ 255813.100000ns, VDD,
+ 255933.100000ns, VDD,
+ 255933.200000ns, VSS,
+ 257014.000000ns, VSS,
+ 257014.100000ns, VDD,
+ 257374.300000ns, VDD,
+ 257374.400000ns, VSS,
+ 257614.500000ns, VSS,
+ 257614.600000ns, VDD,
+ 258094.900000ns, VDD,
+ 258095.000000ns, VSS,
+ 258215.000000ns, VSS,
+ 258215.100000ns, VDD,
+ 258575.300000ns, VDD,
+ 258575.400000ns, VSS,
+ 258815.500000ns, VSS,
+ 258815.600000ns, VDD,
+ 259776.300000ns, VDD,
+ 259776.400000ns, VSS,
+ 260376.800000ns, VSS,
+ 260376.900000ns, VDD,
+ 261217.500000ns, VDD,
+ 261217.600000ns, VSS,
+ 261457.700000ns, VSS,
+ 261457.800000ns, VDD,
+ 261818.000000ns, VDD,
+ 261818.100000ns, VSS,
+ 261938.100000ns, VSS,
+ 261938.200000ns, VDD,
+ 262058.200000ns, VDD,
+ 262058.300000ns, VSS,
+ 263379.300000ns, VSS,
+ 263379.400000ns, VDD,
+ 263859.700000ns, VDD,
+ 263859.800000ns, VSS,
+ 264099.900000ns, VSS,
+ 264100.000000ns, VDD,
+ 264220.000000ns, VDD,
+ 264220.100000ns, VSS,
+ 264340.100000ns, VSS,
+ 264340.200000ns, VDD,
+ 264700.400000ns, VDD,
+ 264700.500000ns, VSS,
+ 265060.700000ns, VSS,
+ 265060.800000ns, VDD,
+ 265541.100000ns, VDD,
+ 265541.200000ns, VSS,
+ 265661.200000ns, VSS,
+ 265661.300000ns, VDD,
+ 266021.500000ns, VDD,
+ 266021.600000ns, VSS,
+ 266141.600000ns, VSS,
+ 266141.700000ns, VDD,
+ 266501.900000ns, VDD,
+ 266502.000000ns, VSS,
+ 266622.000000ns, VSS,
+ 266622.100000ns, VDD,
+ 266982.300000ns, VDD,
+ 266982.400000ns, VSS,
+ 267462.700000ns, VSS,
+ 267462.800000ns, VDD,
+ 268423.500000ns, VDD,
+ 268423.600000ns, VSS,
+ 268663.700000ns, VSS,
+ 268663.800000ns, VDD,
+ 268903.900000ns, VDD,
+ 268904.000000ns, VSS,
+ 269024.000000ns, VSS,
+ 269024.100000ns, VDD,
+ 269384.300000ns, VDD,
+ 269384.400000ns, VSS,
+ 269504.400000ns, VSS,
+ 269504.500000ns, VDD,
+ 270104.900000ns, VDD,
+ 270105.000000ns, VSS,
+ 270585.300000ns, VSS,
+ 270585.400000ns, VDD,
+ 271185.800000ns, VDD,
+ 271185.900000ns, VSS,
+ 271666.200000ns, VSS,
+ 271666.300000ns, VDD,
+ 271906.400000ns, VDD,
+ 271906.500000ns, VSS,
+ 272386.800000ns, VSS,
+ 272386.900000ns, VDD,
+ 272627.000000ns, VDD,
+ 272627.100000ns, VSS,
+ 273347.600000ns, VSS,
+ 273347.700000ns, VDD,
+ 273828.000000ns, VDD,
+ 273828.100000ns, VSS,
+ 274428.500000ns, VSS,
+ 274428.600000ns, VDD,
+ 275629.500000ns, VDD,
+ 275629.600000ns, VSS,
+ 275869.700000ns, VSS,
+ 275869.800000ns, VDD,
+ 276590.300000ns, VDD,
+ 276590.400000ns, VSS,
+ 276710.400000ns, VSS,
+ 276710.500000ns, VDD,
+ 277911.400000ns, VDD,
+ 277911.500000ns, VSS,
+ 278391.800000ns, VSS,
+ 278391.900000ns, VDD,
+ 278632.000000ns, VDD,
+ 278632.100000ns, VSS,
+ 279112.400000ns, VSS,
+ 279112.500000ns, VDD,
+ 279352.600000ns, VDD,
+ 279352.700000ns, VSS,
+ 279472.700000ns, VSS,
+ 279472.800000ns, VDD,
+ 279592.800000ns, VDD,
+ 279592.900000ns, VSS,
+ 279712.900000ns, VSS,
+ 279713.000000ns, VDD,
+ 280313.400000ns, VDD,
+ 280313.500000ns, VSS,
+ 280433.500000ns, VSS,
+ 280433.600000ns, VDD,
+ 281274.200000ns, VDD,
+ 281274.300000ns, VSS,
+ 281514.400000ns, VSS,
+ 281514.500000ns, VDD,
+ 281874.700000ns, VDD,
+ 281874.800000ns, VSS,
+ 282475.200000ns, VSS,
+ 282475.300000ns, VDD,
+ 282715.400000ns, VDD,
+ 282715.500000ns, VSS,
+ 282835.500000ns, VSS,
+ 282835.600000ns, VDD,
+ 283075.700000ns, VDD,
+ 283075.800000ns, VSS,
+ 284036.500000ns, VSS,
+ 284036.600000ns, VDD,
+ 284516.900000ns, VDD,
+ 284517.000000ns, VSS,
+ 284637.000000ns, VSS,
+ 284637.100000ns, VDD,
+ 284997.300000ns, VDD,
+ 284997.400000ns, VSS,
+ 285477.700000ns, VSS,
+ 285477.800000ns, VDD,
+ 285838.000000ns, VDD,
+ 285838.100000ns, VSS,
+ 286558.600000ns, VSS,
+ 286558.700000ns, VDD,
+ 287519.400000ns, VDD,
+ 287519.500000ns, VSS,
+ 288240.000000ns, VSS,
+ 288240.100000ns, VDD,
+ 288480.200000ns, VDD,
+ 288480.300000ns, VSS,
+ 289200.800000ns, VSS,
+ 289200.900000ns, VDD,
+ 290161.600000ns, VDD,
+ 290161.700000ns, VSS,
+ 290401.800000ns, VSS,
+ 290401.900000ns, VDD,
+ 290762.100000ns, VDD,
+ 290762.200000ns, VSS,
+ 291002.300000ns, VSS,
+ 291002.400000ns, VDD,
+ 291122.400000ns, VDD,
+ 291122.500000ns, VSS,
+ 291362.600000ns, VSS,
+ 291362.700000ns, VDD,
+ 291602.800000ns, VDD,
+ 291602.900000ns, VSS,
+ 291843.000000ns, VSS,
+ 291843.100000ns, VDD,
+ 292203.300000ns, VDD,
+ 292203.400000ns, VSS,
+ 292323.400000ns, VSS,
+ 292323.500000ns, VDD,
+ 293644.500000ns, VDD,
+ 293644.600000ns, VSS,
+ 294124.900000ns, VSS,
+ 294125.000000ns, VDD,
+ 294485.200000ns, VDD,
+ 294485.300000ns, VSS,
+ 294845.500000ns, VSS,
+ 294845.600000ns, VDD,
+ 294965.600000ns, VDD,
+ 294965.700000ns, VSS,
+ 295926.400000ns, VSS,
+ 295926.500000ns, VDD,
+ 296526.900000ns, VDD,
+ 296527.000000ns, VSS,
+ 296647.000000ns, VSS,
+ 296647.100000ns, VDD,
+ 297007.300000ns, VDD,
+ 297007.400000ns, VSS,
+ 297487.700000ns, VSS,
+ 297487.800000ns, VDD,
+ 297968.100000ns, VDD,
+ 297968.200000ns, VSS,
+ 298208.300000ns, VSS,
+ 298208.400000ns, VDD,
+ 298448.500000ns, VDD,
+ 298448.600000ns, VSS,
+ 299169.100000ns, VSS,
+ 299169.200000ns, VDD,
+ 299409.300000ns, VDD,
+ 299409.400000ns, VSS,
+ 299529.400000ns, VSS,
+ 299529.500000ns, VDD,
+ 299649.500000ns, VDD,
+ 299649.600000ns, VSS,
+ 299889.700000ns, VSS,
+ 299889.800000ns, VDD,
+ 300250.000000ns, VDD,
+ 300250.100000ns, VSS,
+ 300490.200000ns, VSS,
+ 300490.300000ns, VDD,
+ 300730.400000ns, VDD,
+ 300730.500000ns, VSS,
+ 300850.500000ns, VSS,
+ 300850.600000ns, VDD,
+ 300970.600000ns, VDD,
+ 300970.700000ns, VSS,
+ 301210.800000ns, VSS,
+ 301210.900000ns, VDD,
+ 301571.100000ns, VDD,
+ 301571.200000ns, VSS,
+ 302291.700000ns, VSS,
+ 302291.800000ns, VDD,
+ 302892.200000ns, VDD,
+ 302892.300000ns, VSS,
+ 303612.800000ns, VSS,
+ 303612.900000ns, VDD,
+ 303853.000000ns, VDD,
+ 303853.100000ns, VSS,
+ 304093.200000ns, VSS,
+ 304093.300000ns, VDD,
+ 304573.600000ns, VDD,
+ 304573.700000ns, VSS,
+ 304813.800000ns, VSS,
+ 304813.900000ns, VDD,
+ 305174.100000ns, VDD,
+ 305174.200000ns, VSS,
+ 305294.200000ns, VSS,
+ 305294.300000ns, VDD,
+ 305894.700000ns, VDD,
+ 305894.800000ns, VSS,
+ 306855.500000ns, VSS,
+ 306855.600000ns, VDD,
+ 307215.800000ns, VDD,
+ 307215.900000ns, VSS,
+ 307936.400000ns, VSS,
+ 307936.500000ns, VDD,
+ 308056.500000ns, VDD,
+ 308056.600000ns, VSS,
+ 308657.000000ns, VSS,
+ 308657.100000ns, VDD,
+ 309017.300000ns, VDD,
+ 309017.400000ns, VSS,
+ 309257.500000ns, VSS,
+ 309257.600000ns, VDD,
+ 309497.700000ns, VDD,
+ 309497.800000ns, VSS,
+ 309858.000000ns, VSS,
+ 309858.100000ns, VDD,
+ 310338.400000ns, VDD,
+ 310338.500000ns, VSS,
+ 310818.800000ns, VSS,
+ 310818.900000ns, VDD,
+ 310938.900000ns, VDD,
+ 310939.000000ns, VSS,
+ 311419.300000ns, VSS,
+ 311419.400000ns, VDD,
+ 311539.400000ns, VDD,
+ 311539.500000ns, VSS,
+ 313340.900000ns, VSS,
+ 313341.000000ns, VDD,
+ 313461.000000ns, VDD,
+ 313461.100000ns, VSS,
+ 314181.600000ns, VSS,
+ 314181.700000ns, VDD,
+ 314301.700000ns, VDD,
+ 314301.800000ns, VSS,
+ 314421.800000ns, VSS,
+ 314421.900000ns, VDD,
+ 314782.100000ns, VDD,
+ 314782.200000ns, VSS,
+ 314902.200000ns, VSS,
+ 314902.300000ns, VDD,
+ 315142.400000ns, VDD,
+ 315142.500000ns, VSS,
+ 315742.900000ns, VSS,
+ 315743.000000ns, VDD,
+ 315863.000000ns, VDD,
+ 315863.100000ns, VSS,
+ 316223.300000ns, VSS,
+ 316223.400000ns, VDD,
+ 316463.500000ns, VDD,
+ 316463.600000ns, VSS,
+ 316583.600000ns, VSS,
+ 316583.700000ns, VDD,
+ 316823.800000ns, VDD,
+ 316823.900000ns, VSS,
+ 317064.000000ns, VSS,
+ 317064.100000ns, VDD,
+ 317904.700000ns, VDD,
+ 317904.800000ns, VSS,
+ 318144.900000ns, VSS,
+ 318145.000000ns, VDD,
+ 318505.200000ns, VDD,
+ 318505.300000ns, VSS,
+ 318985.600000ns, VSS,
+ 318985.700000ns, VDD,
+ 319826.300000ns, VDD,
+ 319826.400000ns, VSS,
+ 320186.600000ns, VSS,
+ 320186.700000ns, VDD,
+ 320546.900000ns, VDD,
+ 320547.000000ns, VSS,
+ 321747.900000ns, VSS,
+ 321748.000000ns, VDD,
+ 322108.200000ns, VDD,
+ 322108.300000ns, VSS,
+ 322228.300000ns, VSS,
+ 322228.400000ns, VDD,
+ 322588.600000ns, VDD,
+ 322588.700000ns, VSS,
+ 322828.800000ns, VSS,
+ 322828.900000ns, VDD,
+ 323429.300000ns, VDD,
+ 323429.400000ns, VSS,
+ 324149.900000ns, VSS,
+ 324150.000000ns, VDD,
+ 324270.000000ns, VDD,
+ 324270.100000ns, VSS,
+ 325110.700000ns, VSS,
+ 325110.800000ns, VDD,
+ 325471.000000ns, VDD,
+ 325471.100000ns, VSS,
+ 325591.100000ns, VSS,
+ 325591.200000ns, VDD,
+ 326551.900000ns, VDD,
+ 326552.000000ns, VSS,
+ 326672.000000ns, VSS,
+ 326672.100000ns, VDD,
+ 326912.200000ns, VDD,
+ 326912.300000ns, VSS,
+ 327512.700000ns, VSS,
+ 327512.800000ns, VDD,
+ 327632.800000ns, VDD,
+ 327632.900000ns, VSS,
+ 328113.200000ns, VSS,
+ 328113.300000ns, VDD,
+ 328953.900000ns, VDD,
+ 328954.000000ns, VSS,
+ 329314.200000ns, VSS,
+ 329314.300000ns, VDD,
+ 329554.400000ns, VDD,
+ 329554.500000ns, VSS,
+ 329674.500000ns, VSS,
+ 329674.600000ns, VDD,
+ 330154.900000ns, VDD,
+ 330155.000000ns, VSS,
+ 330635.300000ns, VSS,
+ 330635.400000ns, VDD,
+ 331476.000000ns, VDD,
+ 331476.100000ns, VSS,
+ 331836.300000ns, VSS,
+ 331836.400000ns, VDD,
+ 332076.500000ns, VDD,
+ 332076.600000ns, VSS,
+ 332316.700000ns, VSS,
+ 332316.800000ns, VDD,
+ 333157.400000ns, VDD,
+ 333157.500000ns, VSS,
+ 333517.700000ns, VSS,
+ 333517.800000ns, VDD,
+ 334358.400000ns, VDD,
+ 334358.500000ns, VSS,
+ 334478.500000ns, VSS,
+ 334478.600000ns, VDD,
+ 334718.700000ns, VDD,
+ 334718.800000ns, VSS,
+ 334838.800000ns, VSS,
+ 334838.900000ns, VDD,
+ 335799.600000ns, VDD,
+ 335799.700000ns, VSS,
+ 336520.200000ns, VSS,
+ 336520.300000ns, VDD,
+ 337000.600000ns, VDD,
+ 337000.700000ns, VSS,
+ 337601.100000ns, VSS,
+ 337601.200000ns, VDD,
+ 338081.500000ns, VDD,
+ 338081.600000ns, VSS,
+ 338441.800000ns, VSS,
+ 338441.900000ns, VDD,
+ 339162.400000ns, VDD,
+ 339162.500000ns, VSS,
+ 339402.600000ns, VSS,
+ 339402.700000ns, VDD,
+ 339762.900000ns, VDD,
+ 339763.000000ns, VSS,
+ 340003.100000ns, VSS,
+ 340003.200000ns, VDD,
+ 340843.800000ns, VDD,
+ 340843.900000ns, VSS,
+ 340963.900000ns, VSS,
+ 340964.000000ns, VDD,
+ 341324.200000ns, VDD,
+ 341324.300000ns, VSS,
+ 341444.300000ns, VSS,
+ 341444.400000ns, VDD,
+ 342285.000000ns, VDD,
+ 342285.100000ns, VSS,
+ 342525.200000ns, VSS,
+ 342525.300000ns, VDD,
+ 342885.500000ns, VDD,
+ 342885.600000ns, VSS,
+ 343005.600000ns, VSS,
+ 343005.700000ns, VDD,
+ 343245.800000ns, VDD,
+ 343245.900000ns, VSS,
+ 344566.900000ns, VSS,
+ 344567.000000ns, VDD,
+ 344687.000000ns, VDD,
+ 344687.100000ns, VSS,
+ 344807.100000ns, VSS,
+ 344807.200000ns, VDD,
+ 345167.400000ns, VDD,
+ 345167.500000ns, VSS,
+ 345647.800000ns, VSS,
+ 345647.900000ns, VDD,
+ 346968.900000ns, VDD,
+ 346969.000000ns, VSS,
+ 347209.100000ns, VSS,
+ 347209.200000ns, VDD,
+ 347329.200000ns, VDD,
+ 347329.300000ns, VSS,
+ 347449.300000ns, VSS,
+ 347449.400000ns, VDD,
+ 347929.700000ns, VDD,
+ 347929.800000ns, VSS,
+ 348650.300000ns, VSS,
+ 348650.400000ns, VDD,
+ 349370.900000ns, VDD,
+ 349371.000000ns, VSS,
+ 349971.400000ns, VSS,
+ 349971.500000ns, VDD,
+ 350331.700000ns, VDD,
+ 350331.800000ns, VSS,
+ 350451.800000ns, VSS,
+ 350451.900000ns, VDD,
+ 350812.100000ns, VDD,
+ 350812.200000ns, VSS,
+ 352133.200000ns, VSS,
+ 352133.300000ns, VDD,
+ 352613.600000ns, VDD,
+ 352613.700000ns, VSS,
+ 352733.700000ns, VSS,
+ 352733.800000ns, VDD,
+ 353094.000000ns, VDD,
+ 353094.100000ns, VSS,
+ 353334.200000ns, VSS,
+ 353334.300000ns, VDD,
+ 353934.700000ns, VDD,
+ 353934.800000ns, VSS,
+ 354174.900000ns, VSS,
+ 354175.000000ns, VDD,
+ 354295.000000ns, VDD,
+ 354295.100000ns, VSS,
+ 354535.200000ns, VSS,
+ 354535.300000ns, VDD,
+ 354655.300000ns, VDD,
+ 354655.400000ns, VSS,
+ 355736.200000ns, VSS,
+ 355736.300000ns, VDD,
+ 356096.500000ns, VDD,
+ 356096.600000ns, VSS,
+ 356216.600000ns, VSS,
+ 356216.700000ns, VDD,
+ 356697.000000ns, VDD,
+ 356697.100000ns, VSS,
+ 356817.100000ns, VSS,
+ 356817.200000ns, VDD,
+ 358378.400000ns, VDD,
+ 358378.500000ns, VSS,
+ 358498.500000ns, VSS,
+ 358498.600000ns, VDD,
+ 358978.900000ns, VDD,
+ 358979.000000ns, VSS,
+ 359099.000000ns, VSS,
+ 359099.100000ns, VDD,
+ 359459.300000ns, VDD,
+ 359459.400000ns, VSS,
+ 360059.800000ns, VSS,
+ 360059.900000ns, VDD,
+ 360179.900000ns, VDD,
+ 360180.000000ns, VSS,
+ 360540.200000ns, VSS,
+ 360540.300000ns, VDD,
+ 360660.300000ns, VDD,
+ 360660.400000ns, VSS,
+ 360780.400000ns, VSS,
+ 360780.500000ns, VDD,
+ 361020.600000ns, VDD,
+ 361020.700000ns, VSS,
+ 361140.700000ns, VSS,
+ 361140.800000ns, VDD,
+ 361501.000000ns, VDD,
+ 361501.100000ns, VSS,
+ 361621.100000ns, VSS,
+ 361621.200000ns, VDD,
+ 362221.600000ns, VDD,
+ 362221.700000ns, VSS,
+ 362461.800000ns, VSS,
+ 362461.900000ns, VDD,
+ 362581.900000ns, VDD,
+ 362582.000000ns, VSS,
+ 362822.100000ns, VSS,
+ 362822.200000ns, VDD,
+ 362942.200000ns, VDD,
+ 362942.300000ns, VSS,
+ 364383.400000ns, VSS,
+ 364383.500000ns, VDD,
+ 365824.600000ns, VDD,
+ 365824.700000ns, VSS,
+ 366305.000000ns, VSS,
+ 366305.100000ns, VDD,
+ 366665.300000ns, VDD,
+ 366665.400000ns, VSS,
+ 367145.700000ns, VSS,
+ 367145.800000ns, VDD,
+ 367385.900000ns, VDD,
+ 367386.000000ns, VSS,
+ 367746.200000ns, VSS,
+ 367746.300000ns, VDD,
+ 368226.600000ns, VDD,
+ 368226.700000ns, VSS,
+ 369307.500000ns, VSS,
+ 369307.600000ns, VDD,
+ 369787.900000ns, VDD,
+ 369788.000000ns, VSS,
+ 370028.100000ns, VSS,
+ 370028.200000ns, VDD,
+ 370388.400000ns, VDD,
+ 370388.500000ns, VSS,
+ 370628.600000ns, VSS,
+ 370628.700000ns, VDD,
+ 370988.900000ns, VDD,
+ 370989.000000ns, VSS,
+ 371109.000000ns, VSS,
+ 371109.100000ns, VDD,
+ 371829.600000ns, VDD,
+ 371829.700000ns, VSS,
+ 372189.900000ns, VSS,
+ 372190.000000ns, VDD,
+ 372430.100000ns, VDD,
+ 372430.200000ns, VSS,
+ 373030.600000ns, VSS,
+ 373030.700000ns, VDD,
+ 373390.900000ns, VDD,
+ 373391.000000ns, VSS,
+ 373991.400000ns, VSS,
+ 373991.500000ns, VDD,
+ 374231.600000ns, VDD,
+ 374231.700000ns, VSS,
+ 374351.700000ns, VSS,
+ 374351.800000ns, VDD,
+ 374952.200000ns, VDD,
+ 374952.300000ns, VSS,
+ 375192.400000ns, VSS,
+ 375192.500000ns, VDD,
+ 375552.700000ns, VDD,
+ 375552.800000ns, VSS,
+ 375672.800000ns, VSS,
+ 375672.900000ns, VDD,
+ 375913.000000ns, VDD,
+ 375913.100000ns, VSS,
+ 376033.100000ns, VSS,
+ 376033.200000ns, VDD,
+ 376633.600000ns, VDD,
+ 376633.700000ns, VSS,
+ 377234.100000ns, VSS,
+ 377234.200000ns, VDD,
+ 377474.300000ns, VDD,
+ 377474.400000ns, VSS,
+ 378915.500000ns, VSS,
+ 378915.600000ns, VDD,
+ 379516.000000ns, VDD,
+ 379516.100000ns, VSS,
+ 379996.400000ns, VSS,
+ 379996.500000ns, VDD,
+ 380236.600000ns, VDD,
+ 380236.700000ns, VSS,
+ 380476.800000ns, VSS,
+ 380476.900000ns, VDD,
+ 380596.900000ns, VDD,
+ 380597.000000ns, VSS,
+ 380717.000000ns, VSS,
+ 380717.100000ns, VDD,
+ 380837.100000ns, VDD,
+ 380837.200000ns, VSS,
+ 381077.300000ns, VSS,
+ 381077.400000ns, VDD,
+ 384320.000000ns, VDD,
+ 384320.100000ns, VSS,
+ 385641.100000ns, VSS,
+ 385641.200000ns, VDD,
+ 385761.200000ns, VDD,
+ 385761.300000ns, VSS,
+ 386241.600000ns, VSS,
+ 386241.700000ns, VDD,
+ 387082.300000ns, VDD,
+ 387082.400000ns, VSS,
+ 387562.700000ns, VSS,
+ 387562.800000ns, VDD,
+ 387802.900000ns, VDD,
+ 387803.000000ns, VSS,
+ 387923.000000ns, VSS,
+ 387923.100000ns, VDD,
+ 388043.100000ns, VDD,
+ 388043.200000ns, VSS,
+ 388283.300000ns, VSS,
+ 388283.400000ns, VDD,
+ 388403.400000ns, VDD,
+ 388403.500000ns, VSS,
+ 388643.600000ns, VSS,
+ 388643.700000ns, VDD,
+ 388763.700000ns, VDD,
+ 388763.800000ns, VSS,
+ 388883.800000ns, VSS,
+ 388883.900000ns, VDD,
+ 389364.200000ns, VDD,
+ 389364.300000ns, VSS,
+ 389484.300000ns, VSS,
+ 389484.400000ns, VDD,
+ 389844.600000ns, VDD,
+ 389844.700000ns, VSS,
+ 390325.000000ns, VSS,
+ 390325.100000ns, VDD,
+ 390685.300000ns, VDD,
+ 390685.400000ns, VSS,
+ 390925.500000ns, VSS,
+ 390925.600000ns, VDD,
+ 391526.000000ns, VDD,
+ 391526.100000ns, VSS,
+ 392606.900000ns, VSS,
+ 392607.000000ns, VDD,
+ 392967.200000ns, VDD,
+ 392967.300000ns, VSS,
+ 393087.300000ns, VSS,
+ 393087.400000ns, VDD,
+ 393327.500000ns, VDD,
+ 393327.600000ns, VSS,
+ 393807.900000ns, VSS,
+ 393808.000000ns, VDD,
+ 393928.000000ns, VDD,
+ 393928.100000ns, VSS,
+ 394168.200000ns, VSS,
+ 394168.300000ns, VDD,
+ 394288.300000ns, VDD,
+ 394288.400000ns, VSS,
+ 394408.400000ns, VSS,
+ 394408.500000ns, VDD,
+ 394648.600000ns, VDD,
+ 394648.700000ns, VSS,
+ 394768.700000ns, VSS,
+ 394768.800000ns, VDD,
+ 396089.800000ns, VDD,
+ 396089.900000ns, VSS,
+ 396209.900000ns, VSS,
+ 396210.000000ns, VDD,
+ 396810.400000ns, VDD,
+ 396810.500000ns, VSS,
+ 396930.500000ns, VSS,
+ 396930.600000ns, VDD,
+ 397531.000000ns, VDD,
+ 397531.100000ns, VSS,
+ 397651.100000ns, VSS,
+ 397651.200000ns, VDD,
+ 398011.400000ns, VDD,
+ 398011.500000ns, VSS,
+ 398371.700000ns, VSS,
+ 398371.800000ns, VDD,
+ 398732.000000ns, VDD,
+ 398732.100000ns, VSS,
+ 398852.100000ns, VSS,
+ 398852.200000ns, VDD,
+ 399572.700000ns, VDD,
+ 399572.800000ns, VSS,
+ 399692.800000ns, VSS,
+ 399692.900000ns, VDD,
+ 400053.100000ns, VDD,
+ 400053.200000ns, VSS,
+ 400173.200000ns, VSS,
+ 400173.300000ns, VDD,
+ 400413.400000ns, VDD,
+ 400413.500000ns, VSS,
+ 400653.600000ns, VSS,
+ 400653.700000ns, VDD,
+ 401134.000000ns, VDD,
+ 401134.100000ns, VSS,
+ 401494.300000ns, VSS,
+ 401494.400000ns, VDD,
+ 401614.400000ns, VDD,
+ 401614.500000ns, VSS,
+ 401854.600000ns, VSS,
+ 401854.700000ns, VDD,
+ 401974.700000ns, VDD,
+ 401974.800000ns, VSS,
+ 402455.100000ns, VSS,
+ 402455.200000ns, VDD,
+ 402815.400000ns, VDD,
+ 402815.500000ns, VSS,
+ 403055.600000ns, VSS,
+ 403055.700000ns, VDD,
+ 403656.100000ns, VDD,
+ 403656.200000ns, VSS,
+ 403896.300000ns, VSS,
+ 403896.400000ns, VDD,
+ 404376.700000ns, VDD,
+ 404376.800000ns, VSS,
+ 404496.800000ns, VSS,
+ 404496.900000ns, VDD,
+ 404616.900000ns, VDD,
+ 404617.000000ns, VSS,
+ 404857.100000ns, VSS,
+ 404857.200000ns, VDD,
+ 405817.900000ns, VDD,
+ 405818.000000ns, VSS,
+ 405938.000000ns, VSS,
+ 405938.100000ns, VDD,
+ 406058.100000ns, VDD,
+ 406058.200000ns, VSS,
+ 406658.600000ns, VSS,
+ 406658.700000ns, VDD,
+ 406778.700000ns, VDD,
+ 406778.800000ns, VSS,
+ 406898.800000ns, VSS,
+ 406898.900000ns, VDD,
+ 407018.900000ns, VDD,
+ 407019.000000ns, VSS,
+ 407259.100000ns, VSS,
+ 407259.200000ns, VDD,
+ 408099.800000ns, VDD,
+ 408099.900000ns, VSS,
+ 408219.900000ns, VSS,
+ 408220.000000ns, VDD,
+ 408460.100000ns, VDD,
+ 408460.200000ns, VSS,
+ 408700.300000ns, VSS,
+ 408700.400000ns, VDD,
+ 409060.600000ns, VDD,
+ 409060.700000ns, VSS,
+ 409180.700000ns, VSS,
+ 409180.800000ns, VDD,
+ 409541.000000ns, VDD,
+ 409541.100000ns, VSS,
+ 409661.100000ns, VSS,
+ 409661.200000ns, VDD,
+ 410021.400000ns, VDD,
+ 410021.500000ns, VSS,
+ 410862.100000ns, VSS,
+ 410862.200000ns, VDD,
+ 411102.300000ns, VDD,
+ 411102.400000ns, VSS,
+ 411222.400000ns, VSS,
+ 411222.500000ns, VDD,
+ 411342.500000ns, VDD,
+ 411342.600000ns, VSS,
+ 411822.900000ns, VSS,
+ 411823.000000ns, VDD,
+ 412183.200000ns, VDD,
+ 412183.300000ns, VSS,
+ 412423.400000ns, VSS,
+ 412423.500000ns, VDD,
+ 413023.900000ns, VDD,
+ 413024.000000ns, VSS,
+ 413264.100000ns, VSS,
+ 413264.200000ns, VDD,
+ 413504.300000ns, VDD,
+ 413504.400000ns, VSS,
+ 413624.400000ns, VSS,
+ 413624.500000ns, VDD,
+ 413744.500000ns, VDD,
+ 413744.600000ns, VSS,
+ 413864.600000ns, VSS,
+ 413864.700000ns, VDD,
+ 414224.900000ns, VDD,
+ 414225.000000ns, VSS,
+ 414945.500000ns, VSS,
+ 414945.600000ns, VDD,
+ 415065.600000ns, VDD,
+ 415065.700000ns, VSS,
+ 415305.800000ns, VSS,
+ 415305.900000ns, VDD,
+ 415666.100000ns, VDD,
+ 415666.200000ns, VSS,
+ 415906.300000ns, VSS,
+ 415906.400000ns, VDD,
+ 417107.300000ns, VDD,
+ 417107.400000ns, VSS,
+ 417227.400000ns, VSS,
+ 417227.500000ns, VDD,
+ 417467.600000ns, VDD,
+ 417467.700000ns, VSS,
+ 417707.800000ns, VSS,
+ 417707.900000ns, VDD,
+ 417827.900000ns, VDD,
+ 417828.000000ns, VSS,
+ 418068.100000ns, VSS,
+ 418068.200000ns, VDD,
+ 418188.200000ns, VDD,
+ 418188.300000ns, VSS,
+ 418428.400000ns, VSS,
+ 418428.500000ns, VDD,
+ 418788.700000ns, VDD,
+ 418788.800000ns, VSS,
+ 418908.800000ns, VSS,
+ 418908.900000ns, VDD,
+ 419269.100000ns, VDD,
+ 419269.200000ns, VSS,
+ 419389.200000ns, VSS,
+ 419389.300000ns, VDD,
+ 419509.300000ns, VDD,
+ 419509.400000ns, VSS,
+ 419629.400000ns, VSS,
+ 419629.500000ns, VDD,
+ 419989.700000ns, VDD,
+ 419989.800000ns, VSS,
+ 420350.000000ns, VSS,
+ 420350.100000ns, VDD,
+ 421190.700000ns, VDD,
+ 421190.800000ns, VSS,
+ 421430.900000ns, VSS,
+ 421431.000000ns, VDD,
+ 421791.200000ns, VDD,
+ 421791.300000ns, VSS,
+ 422271.600000ns, VSS,
+ 422271.700000ns, VDD,
+ 422511.800000ns, VDD,
+ 422511.900000ns, VSS,
+ 422631.900000ns, VSS,
+ 422632.000000ns, VDD,
+ 423592.700000ns, VDD,
+ 423592.800000ns, VSS,
+ 424313.300000ns, VSS,
+ 424313.400000ns, VDD,
+ 424553.500000ns, VDD,
+ 424553.600000ns, VSS,
+ 424673.600000ns, VSS,
+ 424673.700000ns, VDD,
+ 424913.800000ns, VDD,
+ 424913.900000ns, VSS,
+ 425274.100000ns, VSS,
+ 425274.200000ns, VDD,
+ 425754.500000ns, VDD,
+ 425754.600000ns, VSS,
+ 426234.900000ns, VSS,
+ 426235.000000ns, VDD,
+ 426355.000000ns, VDD,
+ 426355.100000ns, VSS,
+ 426715.300000ns, VSS,
+ 426715.400000ns, VDD,
+ 427075.600000ns, VDD,
+ 427075.700000ns, VSS,
+ 427315.800000ns, VSS,
+ 427315.900000ns, VDD,
+ 427796.200000ns, VDD,
+ 427796.300000ns, VSS,
+ 428036.400000ns, VSS,
+ 428036.500000ns, VDD,
+ 428396.700000ns, VDD,
+ 428396.800000ns, VSS,
+ 428516.800000ns, VSS,
+ 428516.900000ns, VDD,
+ 429357.500000ns, VDD,
+ 429357.600000ns, VSS,
+ 429477.600000ns, VSS,
+ 429477.700000ns, VDD,
+ 429597.700000ns, VDD,
+ 429597.800000ns, VSS,
+ 429717.800000ns, VSS,
+ 429717.900000ns, VDD,
+ 430078.100000ns, VDD,
+ 430078.200000ns, VSS,
+ 430438.400000ns, VSS,
+ 430438.500000ns, VDD,
+ 430678.600000ns, VDD,
+ 430678.700000ns, VSS,
+ 431038.900000ns, VSS,
+ 431039.000000ns, VDD,
+ 431279.100000ns, VDD,
+ 431279.200000ns, VSS,
+ 431879.600000ns, VSS,
+ 431879.700000ns, VDD,
+ 432720.300000ns, VDD,
+ 432720.400000ns, VSS,
+ 432840.400000ns, VSS,
+ 432840.500000ns, VDD,
+ 433200.700000ns, VDD,
+ 433200.800000ns, VSS,
+ 433681.100000ns, VSS,
+ 433681.200000ns, VDD,
+ 434161.500000ns, VDD,
+ 434161.600000ns, VSS,
+ 434641.900000ns, VSS,
+ 434642.000000ns, VDD,
+ 434882.100000ns, VDD,
+ 434882.200000ns, VSS,
+ 435242.400000ns, VSS,
+ 435242.500000ns, VDD,
+ 435842.900000ns, VDD,
+ 435843.000000ns, VSS,
+ 436683.600000ns, VSS,
+ 436683.700000ns, VDD,
+ 436923.800000ns, VDD,
+ 436923.900000ns, VSS,
+ 437644.400000ns, VSS,
+ 437644.500000ns, VDD,
+ 437884.600000ns, VDD,
+ 437884.700000ns, VSS,
+ 438004.700000ns, VSS,
+ 438004.800000ns, VDD,
+ 438124.800000ns, VDD,
+ 438124.900000ns, VSS,
+ 439566.000000ns, VSS,
+ 439566.100000ns, VDD,
+ 440166.500000ns, VDD,
+ 440166.600000ns, VSS,
+ 440286.600000ns, VSS,
+ 440286.700000ns, VDD,
+ 440406.700000ns, VDD,
+ 440406.800000ns, VSS,
+ 440526.800000ns, VSS,
+ 440526.900000ns, VDD,
+ 440887.100000ns, VDD,
+ 440887.200000ns, VSS,
+ 441727.800000ns, VSS,
+ 441727.900000ns, VDD,
+ 441968.000000ns, VDD,
+ 441968.100000ns, VSS,
+ 442088.100000ns, VSS,
+ 442088.200000ns, VDD,
+ 442448.400000ns, VDD,
+ 442448.500000ns, VSS,
+ 442928.800000ns, VSS,
+ 442928.900000ns, VDD,
+ 443409.200000ns, VDD,
+ 443409.300000ns, VSS,
+ 444610.200000ns, VSS,
+ 444610.300000ns, VDD,
+ 444970.500000ns, VDD,
+ 444970.600000ns, VSS,
+ 445090.600000ns, VSS,
+ 445090.700000ns, VDD,
+ 445450.900000ns, VDD,
+ 445451.000000ns, VSS,
+ 445571.000000ns, VSS,
+ 445571.100000ns, VDD,
+ 445931.300000ns, VDD,
+ 445931.400000ns, VSS,
+ 446171.500000ns, VSS,
+ 446171.600000ns, VDD,
+ 446291.600000ns, VDD,
+ 446291.700000ns, VSS,
+ 446411.700000ns, VSS,
+ 446411.800000ns, VDD,
+ 447132.300000ns, VDD,
+ 447132.400000ns, VSS,
+ 447252.400000ns, VSS,
+ 447252.500000ns, VDD,
+ 447372.500000ns, VDD,
+ 447372.600000ns, VSS,
+ 447732.800000ns, VSS,
+ 447732.900000ns, VDD,
+ 447852.900000ns, VDD,
+ 447853.000000ns, VSS,
+ 449414.200000ns, VSS,
+ 449414.300000ns, VDD,
+ 450615.200000ns, VDD,
+ 450615.300000ns, VSS,
+ 451095.600000ns, VSS,
+ 451095.700000ns, VDD,
+ 451576.000000ns, VDD,
+ 451576.100000ns, VSS,
+ 451696.100000ns, VSS,
+ 451696.200000ns, VDD,
+ 451936.300000ns, VDD,
+ 451936.400000ns, VSS,
+ 452176.500000ns, VSS,
+ 452176.600000ns, VDD,
+ 452296.600000ns, VDD,
+ 452296.700000ns, VSS,
+ 452416.700000ns, VSS,
+ 452416.800000ns, VDD,
+ 453137.300000ns, VDD,
+ 453137.400000ns, VSS,
+ 453617.700000ns, VSS,
+ 453617.800000ns, VDD,
+ 453737.800000ns, VDD,
+ 453737.900000ns, VSS,
+ 453978.000000ns, VSS,
+ 453978.100000ns, VDD,
+ 454098.100000ns, VDD,
+ 454098.200000ns, VSS,
+ 454578.500000ns, VSS,
+ 454578.600000ns, VDD,
+ 454938.800000ns, VDD,
+ 454938.900000ns, VSS,
+ 455058.900000ns, VSS,
+ 455059.000000ns, VDD,
+ 455179.000000ns, VDD,
+ 455179.100000ns, VSS,
+ 456259.900000ns, VSS,
+ 456260.000000ns, VDD,
+ 456500.100000ns, VDD,
+ 456500.200000ns, VSS,
+ 456860.400000ns, VSS,
+ 456860.500000ns, VDD,
+ 457941.300000ns, VDD,
+ 457941.400000ns, VSS,
+ 459022.200000ns, VSS,
+ 459022.300000ns, VDD,
+ 459382.500000ns, VDD,
+ 459382.600000ns, VSS,
+ 459502.600000ns, VSS,
+ 459502.700000ns, VDD,
+ 460103.100000ns, VDD,
+ 460103.200000ns, VSS,
+ 460463.400000ns, VSS,
+ 460463.500000ns, VDD,
+ 460703.600000ns, VDD,
+ 460703.700000ns, VSS,
+ 461304.100000ns, VSS,
+ 461304.200000ns, VDD,
+ 461664.400000ns, VDD,
+ 461664.500000ns, VSS,
+ 461904.600000ns, VSS,
+ 461904.700000ns, VDD,
+ 462264.900000ns, VDD,
+ 462265.000000ns, VSS,
+ 462625.200000ns, VSS,
+ 462625.300000ns, VDD,
+ 462865.400000ns, VDD,
+ 462865.500000ns, VSS,
+ 462985.500000ns, VSS,
+ 462985.600000ns, VDD,
+ 463586.000000ns, VDD,
+ 463586.100000ns, VSS,
+ 463706.100000ns, VSS,
+ 463706.200000ns, VDD,
+ 464066.400000ns, VDD,
+ 464066.500000ns, VSS,
+ 464666.900000ns, VSS,
+ 464667.000000ns, VDD,
+ 464907.100000ns, VDD,
+ 464907.200000ns, VSS,
+ 465027.200000ns, VSS,
+ 465027.300000ns, VDD,
+ 465627.700000ns, VDD,
+ 465627.800000ns, VSS,
+ 465988.000000ns, VSS,
+ 465988.100000ns, VDD,
+ 466348.300000ns, VDD,
+ 466348.400000ns, VSS,
+ 466468.400000ns, VSS,
+ 466468.500000ns, VDD,
+ 466948.800000ns, VDD,
+ 466948.900000ns, VSS,
+ 467068.900000ns, VSS,
+ 467069.000000ns, VDD,
+ 467429.200000ns, VDD,
+ 467429.300000ns, VSS,
+ 467549.300000ns, VSS,
+ 467549.400000ns, VDD,
+ 468029.700000ns, VDD,
+ 468029.800000ns, VSS,
+ 468149.800000ns, VSS,
+ 468149.900000ns, VDD,
+ 469230.700000ns, VDD,
+ 469230.800000ns, VSS,
+ 469350.800000ns, VSS,
+ 469350.900000ns, VDD,
+ 470912.100000ns, VDD,
+ 470912.200000ns, VSS,
+ 471392.500000ns, VSS,
+ 471392.600000ns, VDD,
+ 471872.900000ns, VDD,
+ 471873.000000ns, VSS,
+ 471993.000000ns, VSS,
+ 471993.100000ns, VDD,
+ 472113.100000ns, VDD,
+ 472113.200000ns, VSS,
+ 472473.400000ns, VSS,
+ 472473.500000ns, VDD,
+ 472713.600000ns, VDD,
+ 472713.700000ns, VSS,
+ 472833.700000ns, VSS,
+ 472833.800000ns, VDD,
+ 473194.000000ns, VDD,
+ 473194.100000ns, VSS,
+ 473674.400000ns, VSS,
+ 473674.500000ns, VDD,
+ 473914.600000ns, VDD,
+ 473914.700000ns, VSS,
+ 474034.700000ns, VSS,
+ 474034.800000ns, VDD,
+ 474154.800000ns, VDD,
+ 474154.900000ns, VSS,
+ 474274.900000ns, VSS,
+ 474275.000000ns, VDD,
+ 475235.700000ns, VDD,
+ 475235.800000ns, VSS,
+ 475716.100000ns, VSS,
+ 475716.200000ns, VDD,
+ 475956.300000ns, VDD,
+ 475956.400000ns, VSS,
+ 476316.600000ns, VSS,
+ 476316.700000ns, VDD,
+ 476556.800000ns, VDD,
+ 476556.900000ns, VSS,
+ 476676.900000ns, VSS,
+ 476677.000000ns, VDD,
+ 476797.000000ns, VDD,
+ 476797.100000ns, VSS,
+ 477277.400000ns, VSS,
+ 477277.500000ns, VDD,
+ 477517.600000ns, VDD,
+ 477517.700000ns, VSS,
+ 477757.800000ns, VSS,
+ 477757.900000ns, VDD,
+ 477877.900000ns, VDD,
+ 477878.000000ns, VSS,
+ 478838.700000ns, VSS,
+ 478838.800000ns, VDD,
+ 478958.800000ns, VDD,
+ 478958.900000ns, VSS,
+ 479078.900000ns, VSS,
+ 479079.000000ns, VDD,
+ 479679.400000ns, VDD,
+ 479679.500000ns, VSS,
+ 480279.900000ns, VSS,
+ 480280.000000ns, VDD,
+ 480760.300000ns, VDD,
+ 480760.400000ns, VSS,
+ 481000.500000ns, VSS,
+ 481000.600000ns, VDD,
+ 481841.200000ns, VDD,
+ 481841.300000ns, VSS,
+ 482561.800000ns, VSS,
+ 482561.900000ns, VDD,
+ 482802.000000ns, VDD,
+ 482802.100000ns, VSS,
+ 483522.600000ns, VSS,
+ 483522.700000ns, VDD,
+ 483762.800000ns, VDD,
+ 483762.900000ns, VSS,
+ 484003.000000ns, VSS,
+ 484003.100000ns, VDD,
+ 484363.300000ns, VDD,
+ 484363.400000ns, VSS,
+ 484483.400000ns, VSS,
+ 484483.500000ns, VDD,
+ 486284.900000ns, VDD,
+ 486285.000000ns, VSS,
+ 489047.200000ns, VSS,
+ 489047.300000ns, VDD,
+ 489407.500000ns, VDD,
+ 489407.600000ns, VSS,
+ 489527.600000ns, VSS,
+ 489527.700000ns, VDD,
+ 490128.100000ns, VDD,
+ 490128.200000ns, VSS,
+ 490728.600000ns, VSS,
+ 490728.700000ns, VDD,
+ 491569.300000ns, VDD,
+ 491569.400000ns, VSS,
+ 491929.600000ns, VSS,
+ 491929.700000ns, VDD,
+ 492289.900000ns, VDD,
+ 492290.000000ns, VSS,
+ 492410.000000ns, VSS,
+ 492410.100000ns, VDD,
+ 493250.700000ns, VDD,
+ 493250.800000ns, VSS,
+ 493490.900000ns, VSS,
+ 493491.000000ns, VDD,
+ 493611.000000ns, VDD,
+ 493611.100000ns, VSS,
+ 494091.400000ns, VSS,
+ 494091.500000ns, VDD,
+ 494691.900000ns, VDD,
+ 494692.000000ns, VSS,
+ 494812.000000ns, VSS,
+ 494812.100000ns, VDD,
+ 496013.000000ns, VDD,
+ 496013.100000ns, VSS,
+ 496373.300000ns, VSS,
+ 496373.400000ns, VDD,
+ 496733.600000ns, VDD,
+ 496733.700000ns, VSS,
+ 497214.000000ns, VSS,
+ 497214.100000ns, VDD,
+ 497814.500000ns, VDD,
+ 497814.600000ns, VSS,
+ 498054.700000ns, VSS,
+ 498054.800000ns, VDD,
+ 498174.800000ns, VDD,
+ 498174.900000ns, VSS,
+ 499255.700000ns, VSS,
+ 499255.800000ns, VDD,
+ 499375.800000ns, VDD,
+ 499375.900000ns, VSS,
+ 499856.200000ns, VSS,
+ 499856.300000ns, VDD,
+ 500096.400000ns, VDD,
+ 500096.500000ns, VSS,
+ 500336.600000ns, VSS,
+ 500336.700000ns, VDD,
+ 500817.000000ns, VDD,
+ 500817.100000ns, VSS,
+ 501057.200000ns, VSS,
+ 501057.300000ns, VDD,
+ 501417.500000ns, VDD,
+ 501417.600000ns, VSS,
+ 501537.600000ns, VSS,
+ 501537.700000ns, VDD,
+ 502258.200000ns, VDD,
+ 502258.300000ns, VSS,
+ 502378.300000ns, VSS,
+ 502378.400000ns, VDD,
+ 502978.800000ns, VDD,
+ 502978.900000ns, VSS,
+ 503219.000000ns, VSS,
+ 503219.100000ns, VDD,
+ 503819.500000ns, VDD,
+ 503819.600000ns, VSS,
+ 504179.800000ns, VSS,
+ 504179.900000ns, VDD,
+ 504299.900000ns, VDD,
+ 504300.000000ns, VSS,
+ 504540.100000ns, VSS,
+ 504540.200000ns, VDD,
+ 504900.400000ns, VDD,
+ 504900.500000ns, VSS,
+ 505260.700000ns, VSS,
+ 505260.800000ns, VDD,
+ 505380.800000ns, VDD,
+ 505380.900000ns, VSS,
+ 506221.500000ns, VSS,
+ 506221.600000ns, VDD,
+ 506822.000000ns, VDD,
+ 506822.100000ns, VSS,
+ 506942.100000ns, VSS,
+ 506942.200000ns, VDD,
+ 507302.400000ns, VDD,
+ 507302.500000ns, VSS,
+ 508743.600000ns, VSS,
+ 508743.700000ns, VDD,
+ 508983.800000ns, VDD,
+ 508983.900000ns, VSS,
+ 509103.900000ns, VSS,
+ 509104.000000ns, VDD,
+ 509584.300000ns, VDD,
+ 509584.400000ns, VSS,
+ 509704.400000ns, VSS,
+ 509704.500000ns, VDD,
+ 510064.700000ns, VDD,
+ 510064.800000ns, VSS,
+ 510425.000000ns, VSS,
+ 510425.100000ns, VDD,
+ 511025.500000ns, VDD,
+ 511025.600000ns, VSS,
+ 511265.700000ns, VSS,
+ 511265.800000ns, VDD,
+ 511505.900000ns, VDD,
+ 511506.000000ns, VSS,
+ 511986.300000ns, VSS,
+ 511986.400000ns, VDD,
+ 512706.900000ns, VDD,
+ 512707.000000ns, VSS,
+ 512947.100000ns, VSS,
+ 512947.200000ns, VDD,
+ 513187.300000ns, VDD,
+ 513187.400000ns, VSS,
+ 513547.600000ns, VSS,
+ 513547.700000ns, VDD,
+ 514148.100000ns, VDD,
+ 514148.200000ns, VSS,
+ 514388.300000ns, VSS,
+ 514388.400000ns, VDD,
+ 514508.400000ns, VDD,
+ 514508.500000ns, VSS,
+ 514868.700000ns, VSS,
+ 514868.800000ns, VDD,
+ 515349.100000ns, VDD,
+ 515349.200000ns, VSS,
+ 515469.200000ns, VSS,
+ 515469.300000ns, VDD,
+ 516189.800000ns, VDD,
+ 516189.900000ns, VSS,
+ 516309.900000ns, VSS,
+ 516310.000000ns, VDD,
+ 517751.100000ns, VDD,
+ 517751.200000ns, VSS,
+ 518231.500000ns, VSS,
+ 518231.600000ns, VDD,
+ 518711.900000ns, VDD,
+ 518712.000000ns, VSS,
+ 518952.100000ns, VSS,
+ 518952.200000ns, VDD,
+ 519312.400000ns, VDD,
+ 519312.500000ns, VSS,
+ 520273.200000ns, VSS,
+ 520273.300000ns, VDD,
+ 520513.400000ns, VDD,
+ 520513.500000ns, VSS,
+ 520873.700000ns, VSS,
+ 520873.800000ns, VDD,
+ 521474.200000ns, VDD,
+ 521474.300000ns, VSS,
+ 521714.400000ns, VSS,
+ 521714.500000ns, VDD,
+ 521834.500000ns, VDD,
+ 521834.600000ns, VSS,
+ 521954.600000ns, VSS,
+ 521954.700000ns, VDD,
+ 522915.400000ns, VDD,
+ 522915.500000ns, VSS,
+ 523035.500000ns, VSS,
+ 523035.600000ns, VDD,
+ 523756.100000ns, VDD,
+ 523756.200000ns, VSS,
+ 523876.200000ns, VSS,
+ 523876.300000ns, VDD,
+ 524116.400000ns, VDD,
+ 524116.500000ns, VSS,
+ 524356.600000ns, VSS,
+ 524356.700000ns, VDD,
+ 524837.000000ns, VDD,
+ 524837.100000ns, VSS,
+ 524957.100000ns, VSS,
+ 524957.200000ns, VDD,
+ 525077.200000ns, VDD,
+ 525077.300000ns, VSS,
+ 525557.600000ns, VSS,
+ 525557.700000ns, VDD,
+ 525677.700000ns, VDD,
+ 525677.800000ns, VSS,
+ 525797.800000ns, VSS,
+ 525797.900000ns, VDD,
+ 526398.300000ns, VDD,
+ 526398.400000ns, VSS,
+ 526518.400000ns, VSS,
+ 526518.500000ns, VDD,
+ 526638.500000ns, VDD,
+ 526638.600000ns, VSS,
+ 526998.800000ns, VSS,
+ 526998.900000ns, VDD,
+ 527118.900000ns, VDD,
+ 527119.000000ns, VSS,
+ 527719.400000ns, VSS,
+ 527719.500000ns, VDD,
+ 528560.100000ns, VDD,
+ 528560.200000ns, VSS,
+ 528800.300000ns, VSS,
+ 528800.400000ns, VDD,
+ 529040.500000ns, VDD,
+ 529040.600000ns, VSS,
+ 529400.800000ns, VSS,
+ 529400.900000ns, VDD,
+ 529641.000000ns, VDD,
+ 529641.100000ns, VSS,
+ 529881.200000ns, VSS,
+ 529881.300000ns, VDD,
+ 530001.300000ns, VDD,
+ 530001.400000ns, VSS,
+ 530361.600000ns, VSS,
+ 530361.700000ns, VDD,
+ 530842.000000ns, VDD,
+ 530842.100000ns, VSS,
+ 530962.100000ns, VSS,
+ 530962.200000ns, VDD,
+ 531322.400000ns, VDD,
+ 531322.500000ns, VSS,
+ 531802.800000ns, VSS,
+ 531802.900000ns, VDD,
+ 532283.200000ns, VDD,
+ 532283.300000ns, VSS,
+ 532523.400000ns, VSS,
+ 532523.500000ns, VDD,
+ 533123.900000ns, VDD,
+ 533124.000000ns, VSS,
+ 533844.500000ns, VSS,
+ 533844.600000ns, VDD,
+ 533964.600000ns, VDD,
+ 533964.700000ns, VSS,
+ 534084.700000ns, VSS,
+ 534084.800000ns, VDD,
+ 534445.000000ns, VDD,
+ 534445.100000ns, VSS,
+ 534685.200000ns, VSS,
+ 534685.300000ns, VDD,
+ 534805.300000ns, VDD,
+ 534805.400000ns, VSS,
+ 534925.400000ns, VSS,
+ 534925.500000ns, VDD,
+ 536126.400000ns, VDD,
+ 536126.500000ns, VSS,
+ 536486.700000ns, VSS,
+ 536486.800000ns, VDD,
+ 536726.900000ns, VDD,
+ 536727.000000ns, VSS,
+ 536847.000000ns, VSS,
+ 536847.100000ns, VDD,
+ 537447.500000ns, VDD,
+ 537447.600000ns, VSS,
+ 537927.900000ns, VSS,
+ 537928.000000ns, VDD,
+ 538168.100000ns, VDD,
+ 538168.200000ns, VSS,
+ 538648.500000ns, VSS,
+ 538648.600000ns, VDD,
+ 539609.300000ns, VDD,
+ 539609.400000ns, VSS,
+ 539969.600000ns, VSS,
+ 539969.700000ns, VDD,
+ 540690.200000ns, VDD,
+ 540690.300000ns, VSS,
+ 540930.400000ns, VSS,
+ 540930.500000ns, VDD,
+ 541050.500000ns, VDD,
+ 541050.600000ns, VSS,
+ 541530.900000ns, VSS,
+ 541531.000000ns, VDD,
+ 542131.400000ns, VDD,
+ 542131.500000ns, VSS,
+ 543212.300000ns, VSS,
+ 543212.400000ns, VDD,
+ 543452.500000ns, VDD,
+ 543452.600000ns, VSS,
+ 543572.600000ns, VSS,
+ 543572.700000ns, VDD,
+ 543932.900000ns, VDD,
+ 543933.000000ns, VSS,
+ 544293.200000ns, VSS,
+ 544293.300000ns, VDD,
+ 545133.900000ns, VDD,
+ 545134.000000ns, VSS,
+ 545494.200000ns, VSS,
+ 545494.300000ns, VDD,
+ 545854.500000ns, VDD,
+ 545854.600000ns, VSS,
+ 546815.300000ns, VSS,
+ 546815.400000ns, VDD,
+ 547055.500000ns, VDD,
+ 547055.600000ns, VSS,
+ 547295.700000ns, VSS,
+ 547295.800000ns, VDD,
+ 547415.800000ns, VDD,
+ 547415.900000ns, VSS,
+ 547535.900000ns, VSS,
+ 547536.000000ns, VDD,
+ 548376.600000ns, VDD,
+ 548376.700000ns, VSS,
+ 548736.900000ns, VSS,
+ 548737.000000ns, VDD,
+ 548977.100000ns, VDD,
+ 548977.200000ns, VSS,
+ 549097.200000ns, VSS,
+ 549097.300000ns, VDD,
+ 549217.300000ns, VDD,
+ 549217.400000ns, VSS,
+ 549577.600000ns, VSS,
+ 549577.700000ns, VDD,
+ 549697.700000ns, VDD,
+ 549697.800000ns, VSS,
+ 549817.800000ns, VSS,
+ 549817.900000ns, VDD,
+ 550058.000000ns, VDD,
+ 550058.100000ns, VSS,
+ 550178.100000ns, VSS,
+ 550178.200000ns, VDD,
+ 550298.200000ns, VDD,
+ 550298.300000ns, VSS,
+ 551018.800000ns, VSS,
+ 551018.900000ns, VDD,
+ 551739.400000ns, VDD,
+ 551739.500000ns, VSS,
+ 551979.600000ns, VSS,
+ 551979.700000ns, VDD,
+ 552339.900000ns, VDD,
+ 552340.000000ns, VSS,
+ 552460.000000ns, VSS,
+ 552460.100000ns, VDD,
+ 552820.300000ns, VDD,
+ 552820.400000ns, VSS,
+ 552940.400000ns, VSS,
+ 552940.500000ns, VDD,
+ 553420.800000ns, VDD,
+ 553420.900000ns, VSS,
+ 553781.100000ns, VSS,
+ 553781.200000ns, VDD,
+ 554381.600000ns, VDD,
+ 554381.700000ns, VSS,
+ 554982.100000ns, VSS,
+ 554982.200000ns, VDD,
+ 555222.300000ns, VDD,
+ 555222.400000ns, VSS,
+ 555342.400000ns, VSS,
+ 555342.500000ns, VDD,
+ 555462.500000ns, VDD,
+ 555462.600000ns, VSS,
+ 557143.900000ns, VSS,
+ 557144.000000ns, VDD,
+ 558104.700000ns, VDD,
+ 558104.800000ns, VSS,
+ 558344.900000ns, VSS,
+ 558345.000000ns, VDD,
+ 558705.200000ns, VDD,
+ 558705.300000ns, VSS,
+ 558825.300000ns, VSS,
+ 558825.400000ns, VDD,
+ 559305.700000ns, VDD,
+ 559305.800000ns, VSS,
+ 559666.000000ns, VSS,
+ 559666.100000ns, VDD,
+ 559786.100000ns, VDD,
+ 559786.200000ns, VSS,
+ 560987.100000ns, VSS,
+ 560987.200000ns, VDD,
+ 562188.100000ns, VDD,
+ 562188.200000ns, VSS,
+ 562548.400000ns, VSS,
+ 562548.500000ns, VDD,
+ 562668.500000ns, VDD,
+ 562668.600000ns, VSS,
+ 563269.000000ns, VSS,
+ 563269.100000ns, VDD,
+ 563389.100000ns, VDD,
+ 563389.200000ns, VSS,
+ 563509.200000ns, VSS,
+ 563509.300000ns, VDD,
+ 563749.400000ns, VDD,
+ 563749.500000ns, VSS,
+ 563869.500000ns, VSS,
+ 563869.600000ns, VDD,
+ 564229.800000ns, VDD,
+ 564229.900000ns, VSS,
+ 564830.300000ns, VSS,
+ 564830.400000ns, VDD,
+ 565310.700000ns, VDD,
+ 565310.800000ns, VSS,
+ 565550.900000ns, VSS,
+ 565551.000000ns, VDD,
+ 566271.500000ns, VDD,
+ 566271.600000ns, VSS,
+ 566391.600000ns, VSS,
+ 566391.700000ns, VDD,
+ 566511.700000ns, VDD,
+ 566511.800000ns, VSS,
+ 566872.000000ns, VSS,
+ 566872.100000ns, VDD,
+ 567352.400000ns, VDD,
+ 567352.500000ns, VSS,
+ 567472.500000ns, VSS,
+ 567472.600000ns, VDD,
+ 567712.700000ns, VDD,
+ 567712.800000ns, VSS,
+ 568553.400000ns, VSS,
+ 568553.500000ns, VDD,
+ 569754.400000ns, VDD,
+ 569754.500000ns, VSS,
+ 571195.600000ns, VSS,
+ 571195.700000ns, VDD,
+ 571555.900000ns, VDD,
+ 571556.000000ns, VSS,
+ 571916.200000ns, VSS,
+ 571916.300000ns, VDD,
+ 572516.700000ns, VDD,
+ 572516.800000ns, VSS,
+ 572877.000000ns, VSS,
+ 572877.100000ns, VDD,
+ 573357.400000ns, VDD,
+ 573357.500000ns, VSS,
+ 574198.100000ns, VSS,
+ 574198.200000ns, VDD,
+ 575038.800000ns, VDD,
+ 575038.900000ns, VSS,
+ 575759.400000ns, VSS,
+ 575759.500000ns, VDD,
+ 575879.500000ns, VDD,
+ 575879.600000ns, VSS,
+ 576119.700000ns, VSS,
+ 576119.800000ns, VDD,
+ 576239.800000ns, VDD,
+ 576239.900000ns, VSS,
+ 577440.800000ns, VSS,
+ 577440.900000ns, VDD,
+ 577560.900000ns, VDD,
+ 577561.000000ns, VSS,
+ 577681.000000ns, VSS,
+ 577681.100000ns, VDD,
+ 577921.200000ns, VDD,
+ 577921.300000ns, VSS,
+ 578281.500000ns, VSS,
+ 578281.600000ns, VDD,
+ 578521.700000ns, VDD,
+ 578521.800000ns, VSS,
+ 579002.100000ns, VSS,
+ 579002.200000ns, VDD,
+ 579482.500000ns, VDD,
+ 579482.600000ns, VSS,
+ 579962.900000ns, VSS,
+ 579963.000000ns, VDD,
+ 580803.600000ns, VDD,
+ 580803.700000ns, VSS,
+ 581284.000000ns, VSS,
+ 581284.100000ns, VDD,
+ 581524.200000ns, VDD,
+ 581524.300000ns, VSS,
+ 582004.600000ns, VSS,
+ 582004.700000ns, VDD,
+ 582364.900000ns, VDD,
+ 582365.000000ns, VSS,
+ 582605.100000ns, VSS,
+ 582605.200000ns, VDD,
+ 582845.300000ns, VDD,
+ 582845.400000ns, VSS,
+ 583085.500000ns, VSS,
+ 583085.600000ns, VDD,
+ 583325.700000ns, VDD,
+ 583325.800000ns, VSS,
+ 583445.800000ns, VSS,
+ 583445.900000ns, VDD,
+ 584166.400000ns, VDD,
+ 584166.500000ns, VSS,
+ 584286.500000ns, VSS,
+ 584286.600000ns, VDD,
+ 585247.300000ns, VDD,
+ 585247.400000ns, VSS,
+ 585487.500000ns, VSS,
+ 585487.600000ns, VDD,
+ 585727.700000ns, VDD,
+ 585727.800000ns, VSS,
+ 586208.100000ns, VSS,
+ 586208.200000ns, VDD,
+ 586328.200000ns, VDD,
+ 586328.300000ns, VSS,
+ 587048.800000ns, VSS,
+ 587048.900000ns, VDD,
+ 587289.000000ns, VDD,
+ 587289.100000ns, VSS,
+ 587529.200000ns, VSS,
+ 587529.300000ns, VDD,
+ 588249.800000ns, VDD,
+ 588249.900000ns, VSS,
+ 588490.000000ns, VSS,
+ 588490.100000ns, VDD,
+ 588730.200000ns, VDD,
+ 588730.300000ns, VSS,
+ 589090.500000ns, VSS,
+ 589090.600000ns, VDD,
+ 589210.600000ns, VDD,
+ 589210.700000ns, VSS,
+ 590411.600000ns, VSS,
+ 590411.700000ns, VDD,
+ 590771.900000ns, VDD,
+ 590772.000000ns, VSS,
+ 591252.300000ns, VSS,
+ 591252.400000ns, VDD,
+ 591372.400000ns, VDD,
+ 591372.500000ns, VSS,
+ 591612.600000ns, VSS,
+ 591612.700000ns, VDD,
+ 592093.000000ns, VDD,
+ 592093.100000ns, VSS,
+ 592453.300000ns, VSS,
+ 592453.400000ns, VDD,
+ 592693.500000ns, VDD,
+ 592693.600000ns, VSS,
+ 592813.600000ns, VSS,
+ 592813.700000ns, VDD,
+ 592933.700000ns, VDD,
+ 592933.800000ns, VSS,
+ 593053.800000ns, VSS,
+ 593053.900000ns, VDD,
+ 593414.100000ns, VDD,
+ 593414.200000ns, VSS,
+ 593534.200000ns, VSS,
+ 593534.300000ns, VDD,
+ 593774.400000ns, VDD,
+ 593774.500000ns, VSS,
+ 593894.500000ns, VSS,
+ 593894.600000ns, VDD,
+ 594735.200000ns, VDD,
+ 594735.300000ns, VSS,
+ 594975.400000ns, VSS,
+ 594975.500000ns, VDD,
+ 595696.000000ns, VDD,
+ 595696.100000ns, VSS,
+ 596056.300000ns, VSS,
+ 596056.400000ns, VDD,
+ 596776.900000ns, VDD,
+ 596777.000000ns, VSS,
+ 596897.000000ns, VSS,
+ 596897.100000ns, VDD,
+ 597257.300000ns, VDD,
+ 597257.400000ns, VSS,
+ 597377.400000ns, VSS,
+ 597377.500000ns, VDD,
+ 597737.700000ns, VDD,
+ 597737.800000ns, VSS,
+ 597857.800000ns, VSS,
+ 597857.900000ns, VDD,
+ 598458.300000ns, VDD,
+ 598458.400000ns, VSS,
+ 599058.800000ns, VSS,
+ 599058.900000ns, VDD,
+ 600740.200000ns, VDD,
+ 600740.300000ns, VSS,
+ 602541.700000ns, VSS,
+ 602541.800000ns, VDD,
+ 602781.900000ns, VDD,
+ 602782.000000ns, VSS,
+ 604103.000000ns, VSS,
+ 604103.100000ns, VDD,
+ 604463.300000ns, VDD,
+ 604463.400000ns, VSS,
+ 604583.400000ns, VSS,
+ 604583.500000ns, VDD,
+ 604823.600000ns, VDD,
+ 604823.700000ns, VSS,
+ 606745.200000ns, VSS,
+ 606745.300000ns, VDD,
+ 607225.600000ns, VDD,
+ 607225.700000ns, VSS,
+ 608546.700000ns, VSS,
+ 608546.800000ns, VDD,
+ 608907.000000ns, VDD,
+ 608907.100000ns, VSS,
+ 609507.500000ns, VSS,
+ 609507.600000ns, VDD,
+ 610588.400000ns, VDD,
+ 610588.500000ns, VSS,
+ 610948.700000ns, VSS,
+ 610948.800000ns, VDD,
+ 611188.900000ns, VDD,
+ 611189.000000ns, VSS,
+ 611549.200000ns, VSS,
+ 611549.300000ns, VDD,
+ 611669.300000ns, VDD,
+ 611669.400000ns, VSS,
+ 612269.800000ns, VSS,
+ 612269.900000ns, VDD,
+ 612870.300000ns, VDD,
+ 612870.400000ns, VSS,
+ 613470.800000ns, VSS,
+ 613470.900000ns, VDD,
+ 614191.400000ns, VDD,
+ 614191.500000ns, VSS,
+ 615152.200000ns, VSS,
+ 615152.300000ns, VDD,
+ 615752.700000ns, VDD,
+ 615752.800000ns, VSS,
+ 615992.900000ns, VSS,
+ 615993.000000ns, VDD,
+ 616953.700000ns, VDD,
+ 616953.800000ns, VSS,
+ 617554.200000ns, VSS,
+ 617554.300000ns, VDD,
+ 617794.400000ns, VDD,
+ 617794.500000ns, VSS,
+ 618515.000000ns, VSS,
+ 618515.100000ns, VDD,
+ 619115.500000ns, VDD,
+ 619115.600000ns, VSS,
+ 619716.000000ns, VSS,
+ 619716.100000ns, VDD,
+ 620076.300000ns, VDD,
+ 620076.400000ns, VSS,
+ 620796.900000ns, VSS,
+ 620797.000000ns, VDD,
+ 621277.300000ns, VDD,
+ 621277.400000ns, VSS,
+ 621517.500000ns, VSS,
+ 621517.600000ns, VDD,
+ 621637.600000ns, VDD,
+ 621637.700000ns, VSS,
+ 621757.700000ns, VSS,
+ 621757.800000ns, VDD,
+ 621877.800000ns, VDD,
+ 621877.900000ns, VSS,
+ 622478.300000ns, VSS,
+ 622478.400000ns, VDD,
+ 623319.000000ns, VDD,
+ 623319.100000ns, VSS,
+ 623559.200000ns, VSS,
+ 623559.300000ns, VDD,
+ 623919.500000ns, VDD,
+ 623919.600000ns, VSS,
+ 624399.900000ns, VSS,
+ 624400.000000ns, VDD,
+ 624640.100000ns, VDD,
+ 624640.200000ns, VSS,
+ 624760.200000ns, VSS,
+ 624760.300000ns, VDD,
+ 624880.300000ns, VDD,
+ 624880.400000ns, VSS,
+ 625120.500000ns, VSS,
+ 625120.600000ns, VDD,
+ 625360.700000ns, VDD,
+ 625360.800000ns, VSS,
+ 625600.900000ns, VSS,
+ 625601.000000ns, VDD,
+ 625841.100000ns, VDD,
+ 625841.200000ns, VSS,
+ 626201.400000ns, VSS,
+ 626201.500000ns, VDD,
+ 626441.600000ns, VDD,
+ 626441.700000ns, VSS,
+ 626922.000000ns, VSS,
+ 626922.100000ns, VDD,
+ 627162.200000ns, VDD,
+ 627162.300000ns, VSS,
+ 627642.600000ns, VSS,
+ 627642.700000ns, VDD,
+ 627882.800000ns, VDD,
+ 627882.900000ns, VSS,
+ 628123.000000ns, VSS,
+ 628123.100000ns, VDD,
+ 628243.100000ns, VDD,
+ 628243.200000ns, VSS,
+ 628483.300000ns, VSS,
+ 628483.400000ns, VDD,
+ 628603.400000ns, VDD,
+ 628603.500000ns, VSS,
+ 628963.700000ns, VSS,
+ 628963.800000ns, VDD,
+ 630525.000000ns, VDD,
+ 630525.100000ns, VSS,
+ 630645.100000ns, VSS,
+ 630645.200000ns, VDD,
+ 631005.400000ns, VDD,
+ 631005.500000ns, VSS,
+ 631125.500000ns, VSS,
+ 631125.600000ns, VDD,
+ 631846.100000ns, VDD,
+ 631846.200000ns, VSS,
+ 632326.500000ns, VSS,
+ 632326.600000ns, VDD,
+ 632446.600000ns, VDD,
+ 632446.700000ns, VSS,
+ 632806.900000ns, VSS,
+ 632807.000000ns, VDD,
+ 633047.100000ns, VDD,
+ 633047.200000ns, VSS,
+ 633407.400000ns, VSS,
+ 633407.500000ns, VDD,
+ 634007.900000ns, VDD,
+ 634008.000000ns, VSS,
+ 635208.900000ns, VSS,
+ 635209.000000ns, VDD,
+ 635689.300000ns, VDD,
+ 635689.400000ns, VSS,
+ 636169.700000ns, VSS,
+ 636169.800000ns, VDD,
+ 636770.200000ns, VDD,
+ 636770.300000ns, VSS,
+ 637010.400000ns, VSS,
+ 637010.500000ns, VDD,
+ 637490.800000ns, VDD,
+ 637490.900000ns, VSS,
+ 637610.900000ns, VSS,
+ 637611.000000ns, VDD,
+ 637971.200000ns, VDD,
+ 637971.300000ns, VSS,
+ 638091.300000ns, VSS,
+ 638091.400000ns, VDD,
+ 638451.600000ns, VDD,
+ 638451.700000ns, VSS,
+ 638811.900000ns, VSS,
+ 638812.000000ns, VDD,
+ 639052.100000ns, VDD,
+ 639052.200000ns, VSS,
+ 639412.400000ns, VSS,
+ 639412.500000ns, VDD,
+ 640613.400000ns, VDD,
+ 640613.500000ns, VSS,
+ 641093.800000ns, VSS,
+ 641093.900000ns, VDD,
+ 641574.200000ns, VDD,
+ 641574.300000ns, VSS,
+ 641934.500000ns, VSS,
+ 641934.600000ns, VDD,
+ 642174.700000ns, VDD,
+ 642174.800000ns, VSS,
+ 642535.000000ns, VSS,
+ 642535.100000ns, VDD,
+ 643135.500000ns, VDD,
+ 643135.600000ns, VSS,
+ 644816.900000ns, VSS,
+ 644817.000000ns, VDD,
+ 645057.100000ns, VDD,
+ 645057.200000ns, VSS,
+ 645177.200000ns, VSS,
+ 645177.300000ns, VDD,
+ 645537.500000ns, VDD,
+ 645537.600000ns, VSS,
+ 645897.800000ns, VSS,
+ 645897.900000ns, VDD,
+ 646858.600000ns, VDD,
+ 646858.700000ns, VSS,
+ 646978.700000ns, VSS,
+ 646978.800000ns, VDD,
+ 647218.900000ns, VDD,
+ 647219.000000ns, VSS,
+ 647459.100000ns, VSS,
+ 647459.200000ns, VDD,
+ 648059.600000ns, VDD,
+ 648059.700000ns, VSS,
+ 648780.200000ns, VSS,
+ 648780.300000ns, VDD,
+ 649140.500000ns, VDD,
+ 649140.600000ns, VSS,
+ 649260.600000ns, VSS,
+ 649260.700000ns, VDD,
+ 649380.700000ns, VDD,
+ 649380.800000ns, VSS,
+ 650101.300000ns, VSS,
+ 650101.400000ns, VDD,
+ 650942.000000ns, VDD,
+ 650942.100000ns, VSS,
+ 651062.100000ns, VSS,
+ 651062.200000ns, VDD,
+ 653344.000000ns, VDD,
+ 653344.100000ns, VSS,
+ 654304.800000ns, VSS,
+ 654304.900000ns, VDD,
+ 655025.400000ns, VDD,
+ 655025.500000ns, VSS,
+ 655866.100000ns, VSS,
+ 655866.200000ns, VDD,
+ 656226.400000ns, VDD,
+ 656226.500000ns, VSS,
+ 656947.000000ns, VSS,
+ 656947.100000ns, VDD,
+ 657547.500000ns, VDD,
+ 657547.600000ns, VSS,
+ 657787.700000ns, VSS,
+ 657787.800000ns, VDD,
+ 658628.400000ns, VDD,
+ 658628.500000ns, VSS,
+ 658868.600000ns, VSS,
+ 658868.700000ns, VDD,
+ 659589.200000ns, VDD,
+ 659589.300000ns, VSS,
+ 659709.300000ns, VSS,
+ 659709.400000ns, VDD,
+ 659829.400000ns, VDD,
+ 659829.500000ns, VSS,
+ 659949.500000ns, VSS,
+ 659949.600000ns, VDD,
+ 660429.900000ns, VDD,
+ 660430.000000ns, VSS,
+ 660550.000000ns, VSS,
+ 660550.100000ns, VDD,
+ 660670.100000ns, VDD,
+ 660670.200000ns, VSS,
+ 661030.400000ns, VSS,
+ 661030.500000ns, VDD,
+ 661390.700000ns, VDD,
+ 661390.800000ns, VSS,
+ 661751.000000ns, VSS,
+ 661751.100000ns, VDD,
+ 662111.300000ns, VDD,
+ 662111.400000ns, VSS,
+ 662231.400000ns, VSS,
+ 662231.500000ns, VDD,
+ 662831.900000ns, VDD,
+ 662832.000000ns, VSS,
+ 662952.000000ns, VSS,
+ 662952.100000ns, VDD,
+ 663072.100000ns, VDD,
+ 663072.200000ns, VSS,
+ 663432.400000ns, VSS,
+ 663432.500000ns, VDD,
+ 663672.600000ns, VDD,
+ 663672.700000ns, VSS,
+ 664753.500000ns, VSS,
+ 664753.600000ns, VDD,
+ 664993.700000ns, VDD,
+ 664993.800000ns, VSS,
+ 665233.900000ns, VSS,
+ 665234.000000ns, VDD,
+ 665474.100000ns, VDD,
+ 665474.200000ns, VSS,
+ 666314.800000ns, VSS,
+ 666314.900000ns, VDD,
+ 667155.500000ns, VDD,
+ 667155.600000ns, VSS,
+ 667876.100000ns, VSS,
+ 667876.200000ns, VDD,
+ 667996.200000ns, VDD,
+ 667996.300000ns, VSS,
+ 668716.800000ns, VSS,
+ 668716.900000ns, VDD,
+ 668957.000000ns, VDD,
+ 668957.100000ns, VSS,
+ 669077.100000ns, VSS,
+ 669077.200000ns, VDD,
+ 669197.200000ns, VDD,
+ 669197.300000ns, VSS,
+ 669317.300000ns, VSS,
+ 669317.400000ns, VDD,
+ 669677.600000ns, VDD,
+ 669677.700000ns, VSS,
+ 670518.300000ns, VSS,
+ 670518.400000ns, VDD,
+ 670758.500000ns, VDD,
+ 670758.600000ns, VSS,
+ 670878.600000ns, VSS,
+ 670878.700000ns, VDD,
+ 671118.800000ns, VDD,
+ 671118.900000ns, VSS,
+ 671599.200000ns, VSS,
+ 671599.300000ns, VDD,
+ 672079.600000ns, VDD,
+ 672079.700000ns, VSS,
+ 672560.000000ns, VSS,
+ 672560.100000ns, VDD,
+ 672680.100000ns, VDD,
+ 672680.200000ns, VSS,
+ 673280.600000ns, VSS,
+ 673280.700000ns, VDD,
+ 673640.900000ns, VDD,
+ 673641.000000ns, VSS,
+ 674241.400000ns, VSS,
+ 674241.500000ns, VDD,
+ 674481.600000ns, VDD,
+ 674481.700000ns, VSS,
+ 676283.100000ns, VSS,
+ 676283.200000ns, VDD,
+ 676523.300000ns, VDD,
+ 676523.400000ns, VSS,
+ 676643.400000ns, VSS,
+ 676643.500000ns, VDD,
+ 676883.600000ns, VDD,
+ 676883.700000ns, VSS,
+ 677123.800000ns, VSS,
+ 677123.900000ns, VDD,
+ 677243.900000ns, VDD,
+ 677244.000000ns, VSS,
+ 677364.000000ns, VSS,
+ 677364.100000ns, VDD,
+ 680126.300000ns, VDD,
+ 680126.400000ns, VSS,
+ 680606.700000ns, VSS,
+ 680606.800000ns, VDD,
+ 680846.900000ns, VDD,
+ 680847.000000ns, VSS,
+ 680967.000000ns, VSS,
+ 680967.100000ns, VDD,
+ 681567.500000ns, VDD,
+ 681567.600000ns, VSS,
+ 681687.600000ns, VSS,
+ 681687.700000ns, VDD,
+ 681807.700000ns, VDD,
+ 681807.800000ns, VSS,
+ 682047.900000ns, VSS,
+ 682048.000000ns, VDD,
+ 682168.000000ns, VDD,
+ 682168.100000ns, VSS,
+ 682768.500000ns, VSS,
+ 682768.600000ns, VDD,
+ 683128.800000ns, VDD,
+ 683128.900000ns, VSS,
+ 683369.000000ns, VSS,
+ 683369.100000ns, VDD,
+ 683489.100000ns, VDD,
+ 683489.200000ns, VSS,
+ 683849.400000ns, VSS,
+ 683849.500000ns, VDD,
+ 683969.500000ns, VDD,
+ 683969.600000ns, VSS,
+ 684089.600000ns, VSS,
+ 684089.700000ns, VDD,
+ 684690.100000ns, VDD,
+ 684690.200000ns, VSS,
+ 684930.300000ns, VSS,
+ 684930.400000ns, VDD,
+ 685530.800000ns, VDD,
+ 685530.900000ns, VSS,
+ 685771.000000ns, VSS,
+ 685771.100000ns, VDD,
+ 685891.100000ns, VDD,
+ 685891.200000ns, VSS,
+ 686131.300000ns, VSS,
+ 686131.400000ns, VDD,
+ 686371.500000ns, VDD,
+ 686371.600000ns, VSS,
+ 686491.600000ns, VSS,
+ 686491.700000ns, VDD,
+ 686611.700000ns, VDD,
+ 686611.800000ns, VSS,
+ 686851.900000ns, VSS,
+ 686852.000000ns, VDD,
+ 687572.500000ns, VDD,
+ 687572.600000ns, VSS,
+ 687932.800000ns, VSS,
+ 687932.900000ns, VDD,
+ 688413.200000ns, VDD,
+ 688413.300000ns, VSS,
+ 688773.500000ns, VSS,
+ 688773.600000ns, VDD,
+ 689133.800000ns, VDD,
+ 689133.900000ns, VSS,
+ 689614.200000ns, VSS,
+ 689614.300000ns, VDD,
+ 690214.700000ns, VDD,
+ 690214.800000ns, VSS,
+ 690575.000000ns, VSS,
+ 690575.100000ns, VDD,
+ 690935.300000ns, VDD,
+ 690935.400000ns, VSS,
+ 691175.500000ns, VSS,
+ 691175.600000ns, VDD,
+ 691415.700000ns, VDD,
+ 691415.800000ns, VSS,
+ 691655.900000ns, VSS,
+ 691656.000000ns, VDD,
+ 691776.000000ns, VDD,
+ 691776.100000ns, VSS,
+ 692256.400000ns, VSS,
+ 692256.500000ns, VDD,
+ 692736.800000ns, VDD,
+ 692736.900000ns, VSS,
+ 692977.000000ns, VSS,
+ 692977.100000ns, VDD,
+ 693817.700000ns, VDD,
+ 693817.800000ns, VSS,
+ 694538.300000ns, VSS,
+ 694538.400000ns, VDD,
+ 695018.700000ns, VDD,
+ 695018.800000ns, VSS,
+ 695739.300000ns, VSS,
+ 695739.400000ns, VDD,
+ 696700.100000ns, VDD,
+ 696700.200000ns, VSS,
+ 697540.800000ns, VSS,
+ 697540.900000ns, VDD,
+ 697901.100000ns, VDD,
+ 697901.200000ns, VSS,
+ 698621.700000ns, VSS,
+ 698621.800000ns, VDD,
+ 698741.800000ns, VDD,
+ 698741.900000ns, VSS,
+ 699822.700000ns, VSS,
+ 699822.800000ns, VDD,
+ 700783.500000ns, VDD,
+ 700783.600000ns, VSS,
+ 701143.800000ns, VSS,
+ 701143.900000ns, VDD,
+ 701263.900000ns, VDD,
+ 701264.000000ns, VSS,
+ 701984.500000ns, VSS,
+ 701984.600000ns, VDD,
+ 702705.100000ns, VDD,
+ 702705.200000ns, VSS,
+ 703065.400000ns, VSS,
+ 703065.500000ns, VDD,
+ 703545.800000ns, VDD,
+ 703545.900000ns, VSS,
+ 704746.800000ns, VSS,
+ 704746.900000ns, VDD,
+ 705107.100000ns, VDD,
+ 705107.200000ns, VSS,
+ 705467.400000ns, VSS,
+ 705467.500000ns, VDD,
+ 705587.500000ns, VDD,
+ 705587.600000ns, VSS,
+ 706668.400000ns, VSS,
+ 706668.500000ns, VDD,
+ 706908.600000ns, VDD,
+ 706908.700000ns, VSS,
+ 707028.700000ns, VSS,
+ 707028.800000ns, VDD,
+ 707148.800000ns, VDD,
+ 707148.900000ns, VSS,
+ 707389.000000ns, VSS,
+ 707389.100000ns, VDD,
+ 708469.900000ns, VDD,
+ 708470.000000ns, VSS,
+ 708710.100000ns, VSS,
+ 708710.200000ns, VDD,
+ 708830.200000ns, VDD,
+ 708830.300000ns, VSS,
+ 709070.400000ns, VSS,
+ 709070.500000ns, VDD,
+ 710271.400000ns, VDD,
+ 710271.500000ns, VSS,
+ 710511.600000ns, VSS,
+ 710511.700000ns, VDD,
+ 710631.700000ns, VDD,
+ 710631.800000ns, VSS,
+ 711712.600000ns, VSS,
+ 711712.700000ns, VDD,
+ 712072.900000ns, VDD,
+ 712073.000000ns, VSS,
+ 712193.000000ns, VSS,
+ 712193.100000ns, VDD,
+ 712673.400000ns, VDD,
+ 712673.500000ns, VSS,
+ 712793.500000ns, VSS,
+ 712793.600000ns, VDD,
+ 713394.000000ns, VDD,
+ 713394.100000ns, VSS,
+ 713514.100000ns, VSS,
+ 713514.200000ns, VDD,
+ 713874.400000ns, VDD,
+ 713874.500000ns, VSS,
+ 713994.500000ns, VSS,
+ 713994.600000ns, VDD,
+ 714114.600000ns, VDD,
+ 714114.700000ns, VSS,
+ 714354.800000ns, VSS,
+ 714354.900000ns, VDD,
+ 714715.100000ns, VDD,
+ 714715.200000ns, VSS,
+ 714835.200000ns, VSS,
+ 714835.300000ns, VDD,
+ 715195.500000ns, VDD,
+ 715195.600000ns, VSS,
+ 715435.700000ns, VSS,
+ 715435.800000ns, VDD,
+ 716276.400000ns, VDD,
+ 716276.500000ns, VSS,
+ 716876.900000ns, VSS,
+ 716877.000000ns, VDD,
+ 716997.000000ns, VDD,
+ 716997.100000ns, VSS,
+ 717117.100000ns, VSS,
+ 717117.200000ns, VDD,
+ 717357.300000ns, VDD,
+ 717357.400000ns, VSS,
+ 717477.400000ns, VSS,
+ 717477.500000ns, VDD,
+ 717597.500000ns, VDD,
+ 717597.600000ns, VSS,
+ 718198.000000ns, VSS,
+ 718198.100000ns, VDD,
+ 718318.100000ns, VDD,
+ 718318.200000ns, VSS,
+ 718798.500000ns, VSS,
+ 718798.600000ns, VDD,
+ 719278.900000ns, VDD,
+ 719279.000000ns, VSS,
+ 719399.000000ns, VSS,
+ 719399.100000ns, VDD,
+ 719879.400000ns, VDD,
+ 719879.500000ns, VSS,
+ 720960.300000ns, VSS,
+ 720960.400000ns, VDD,
+ 722161.300000ns, VDD,
+ 722161.400000ns, VSS,
+ 722521.600000ns, VSS,
+ 722521.700000ns, VDD,
+ 722881.900000ns, VDD,
+ 722882.000000ns, VSS,
+ 723122.100000ns, VSS,
+ 723122.200000ns, VDD,
+ 723242.200000ns, VDD,
+ 723242.300000ns, VSS,
+ 723362.300000ns, VSS,
+ 723362.400000ns, VDD,
+ 723602.500000ns, VDD,
+ 723602.600000ns, VSS,
+ 724443.200000ns, VSS,
+ 724443.300000ns, VDD,
+ 726004.500000ns, VDD,
+ 726004.600000ns, VSS,
+ 726244.700000ns, VSS,
+ 726244.800000ns, VDD,
+ 726364.800000ns, VDD,
+ 726364.900000ns, VSS,
+ 726725.100000ns, VSS,
+ 726725.200000ns, VDD,
+ 726845.200000ns, VDD,
+ 726845.300000ns, VSS,
+ 727445.700000ns, VSS,
+ 727445.800000ns, VDD,
+ 729727.600000ns, VDD,
+ 729727.700000ns, VSS,
+ 730087.900000ns, VSS,
+ 730088.000000ns, VDD,
+ 730688.400000ns, VDD,
+ 730688.500000ns, VSS,
+ 731889.400000ns, VSS,
+ 731889.500000ns, VDD,
+ 732129.600000ns, VDD,
+ 732129.700000ns, VSS,
+ 732489.900000ns, VSS,
+ 732490.000000ns, VDD,
+ 732730.100000ns, VDD,
+ 732730.200000ns, VSS,
+ 732850.200000ns, VSS,
+ 732850.300000ns, VDD,
+ 732970.300000ns, VDD,
+ 732970.400000ns, VSS,
+ 733570.800000ns, VSS,
+ 733570.900000ns, VDD,
+ 733690.900000ns, VDD,
+ 733691.000000ns, VSS,
+ 733931.100000ns, VSS,
+ 733931.200000ns, VDD,
+ 734411.500000ns, VDD,
+ 734411.600000ns, VSS,
+ 734531.600000ns, VSS,
+ 734531.700000ns, VDD,
+ 734771.800000ns, VDD,
+ 734771.900000ns, VSS,
+ 734891.900000ns, VSS,
+ 734892.000000ns, VDD,
+ 735252.200000ns, VDD,
+ 735252.300000ns, VSS,
+ 735492.400000ns, VSS,
+ 735492.500000ns, VDD,
+ 735852.700000ns, VDD,
+ 735852.800000ns, VSS,
+ 735972.800000ns, VSS,
+ 735972.900000ns, VDD,
+ 737894.400000ns, VDD,
+ 737894.500000ns, VSS,
+ 738014.500000ns, VSS,
+ 738014.600000ns, VDD,
+ 738374.800000ns, VDD,
+ 738374.900000ns, VSS,
+ 738494.900000ns, VSS,
+ 738495.000000ns, VDD,
+ 738615.000000ns, VDD,
+ 738615.100000ns, VSS,
+ 739215.500000ns, VSS,
+ 739215.600000ns, VDD,
+ 739816.000000ns, VDD,
+ 739816.100000ns, VSS,
+ 740176.300000ns, VSS,
+ 740176.400000ns, VDD,
+ 740296.400000ns, VDD,
+ 740296.500000ns, VSS,
+ 740536.600000ns, VSS,
+ 740536.700000ns, VDD,
+ 740656.700000ns, VDD,
+ 740656.800000ns, VSS,
+ 741137.100000ns, VSS,
+ 741137.200000ns, VDD,
+ 741617.500000ns, VDD,
+ 741617.600000ns, VSS,
+ 741857.700000ns, VSS,
+ 741857.800000ns, VDD,
+ 742097.900000ns, VDD,
+ 742098.000000ns, VSS,
+ 742458.200000ns, VSS,
+ 742458.300000ns, VDD,
+ 742698.400000ns, VDD,
+ 742698.500000ns, VSS,
+ 742818.500000ns, VSS,
+ 742818.600000ns, VDD,
+ 742938.600000ns, VDD,
+ 742938.700000ns, VSS,
+ 743058.700000ns, VSS,
+ 743058.800000ns, VDD,
+ 743298.900000ns, VDD,
+ 743299.000000ns, VSS,
+ 743539.100000ns, VSS,
+ 743539.200000ns, VDD,
+ 743899.400000ns, VDD,
+ 743899.500000ns, VSS,
+ 744139.600000ns, VSS,
+ 744139.700000ns, VDD,
+ 744860.200000ns, VDD,
+ 744860.300000ns, VSS,
+ 745100.400000ns, VSS,
+ 745100.500000ns, VDD,
+ 745220.500000ns, VDD,
+ 745220.600000ns, VSS,
+ 745340.600000ns, VSS,
+ 745340.700000ns, VDD,
+ 746301.400000ns, VDD,
+ 746301.500000ns, VSS,
+ 746541.600000ns, VSS,
+ 746541.700000ns, VDD,
+ 746661.700000ns, VDD,
+ 746661.800000ns, VSS,
+ 747622.500000ns, VSS,
+ 747622.600000ns, VDD,
+ 748583.300000ns, VDD,
+ 748583.400000ns, VSS,
+ 749544.100000ns, VSS,
+ 749544.200000ns, VDD,
+ 749784.300000ns, VDD,
+ 749784.400000ns, VSS,
+ 749904.400000ns, VSS,
+ 749904.500000ns, VDD,
+ 750264.700000ns, VDD,
+ 750264.800000ns, VSS,
+ 750625.000000ns, VSS,
+ 750625.100000ns, VDD,
+ 751345.600000ns, VDD,
+ 751345.700000ns, VSS,
+ 751465.700000ns, VSS,
+ 751465.800000ns, VDD,
+ 751826.000000ns, VDD,
+ 751826.100000ns, VSS,
+ 751946.100000ns, VSS,
+ 751946.200000ns, VDD,
+ 752306.400000ns, VDD,
+ 752306.500000ns, VSS,
+ 754828.500000ns, VSS,
+ 754828.600000ns, VDD,
+ 755549.100000ns, VDD,
+ 755549.200000ns, VSS,
+ 755669.200000ns, VSS,
+ 755669.300000ns, VDD,
+ 756269.700000ns, VDD,
+ 756269.800000ns, VSS,
+ 756389.800000ns, VSS,
+ 756389.900000ns, VDD,
+ 756750.100000ns, VDD,
+ 756750.200000ns, VSS,
+ 757110.400000ns, VSS,
+ 757110.500000ns, VDD,
+ 757831.000000ns, VDD,
+ 757831.100000ns, VSS,
+ 758311.400000ns, VSS,
+ 758311.500000ns, VDD,
+ 758431.500000ns, VDD,
+ 758431.600000ns, VSS,
+ 758551.600000ns, VSS,
+ 758551.700000ns, VDD,
+ 759152.100000ns, VDD,
+ 759152.200000ns, VSS,
+ 759272.200000ns, VSS,
+ 759272.300000ns, VDD,
+ 759752.600000ns, VDD,
+ 759752.700000ns, VSS,
+ 759992.800000ns, VSS,
+ 759992.900000ns, VDD,
+ 760353.100000ns, VDD,
+ 760353.200000ns, VSS,
+ 760473.200000ns, VSS,
+ 760473.300000ns, VDD,
+ 761193.800000ns, VDD,
+ 761193.900000ns, VSS,
+ 761313.900000ns, VSS,
+ 761314.000000ns, VDD,
+ 761674.200000ns, VDD,
+ 761674.300000ns, VSS,
+ 761794.300000ns, VSS,
+ 761794.400000ns, VDD,
+ 762034.500000ns, VDD,
+ 762034.600000ns, VSS,
+ 762154.600000ns, VSS,
+ 762154.700000ns, VDD,
+ 762274.700000ns, VDD,
+ 762274.800000ns, VSS,
+ 762394.800000ns, VSS,
+ 762394.900000ns, VDD,
+ 762755.100000ns, VDD,
+ 762755.200000ns, VSS,
+ 762995.300000ns, VSS,
+ 762995.400000ns, VDD,
+ 763235.500000ns, VDD,
+ 763235.600000ns, VSS,
+ 763355.600000ns, VSS,
+ 763355.700000ns, VDD,
+ 763475.700000ns, VDD,
+ 763475.800000ns, VSS,
+ 763715.900000ns, VSS,
+ 763716.000000ns, VDD,
+ 763836.000000ns, VDD,
+ 763836.100000ns, VSS,
+ 764436.500000ns, VSS,
+ 764436.600000ns, VDD,
+ 764676.700000ns, VDD,
+ 764676.800000ns, VSS,
+ 765037.000000ns, VSS,
+ 765037.100000ns, VDD,
+ 765157.100000ns, VDD,
+ 765157.200000ns, VSS,
+ 765277.200000ns, VSS,
+ 765277.300000ns, VDD,
+ 765637.500000ns, VDD,
+ 765637.600000ns, VSS,
+ 765877.700000ns, VSS,
+ 765877.800000ns, VDD,
+ 767078.700000ns, VDD,
+ 767078.800000ns, VSS,
+ 767799.300000ns, VSS,
+ 767799.400000ns, VDD,
+ 768159.600000ns, VDD,
+ 768159.700000ns, VSS,
+ 768760.100000ns, VSS,
+ 768760.200000ns, VDD,
+ 769120.400000ns, VDD,
+ 769120.500000ns, VSS,
+ 769600.800000ns, VSS,
+ 769600.900000ns, VDD,
+ 770081.200000ns, VDD,
+ 770081.300000ns, VSS,
+ 770321.400000ns, VSS,
+ 770321.500000ns, VDD,
+ 770801.800000ns, VDD,
+ 770801.900000ns, VSS,
+ 771522.400000ns, VSS,
+ 771522.500000ns, VDD,
+ 772002.800000ns, VDD,
+ 772002.900000ns, VSS,
+ 772122.900000ns, VSS,
+ 772123.000000ns, VDD,
+ 772363.100000ns, VDD,
+ 772363.200000ns, VSS,
+ 772483.200000ns, VSS,
+ 772483.300000ns, VDD,
+ 773203.800000ns, VDD,
+ 773203.900000ns, VSS,
+ 773323.900000ns, VSS,
+ 773324.000000ns, VDD,
+ 773924.400000ns, VDD,
+ 773924.500000ns, VSS,
+ 774044.500000ns, VSS,
+ 774044.600000ns, VDD,
+ 775005.300000ns, VDD,
+ 775005.400000ns, VSS,
+ 775125.400000ns, VSS,
+ 775125.500000ns, VDD,
+ 775245.500000ns, VDD,
+ 775245.600000ns, VSS,
+ 775485.700000ns, VSS,
+ 775485.800000ns, VDD,
+ 776086.200000ns, VDD,
+ 776086.300000ns, VSS,
+ 776326.400000ns, VSS,
+ 776326.500000ns, VDD,
+ 777407.300000ns, VDD,
+ 777407.400000ns, VSS,
+ 777647.500000ns, VSS,
+ 777647.600000ns, VDD,
+ 777767.600000ns, VDD,
+ 777767.700000ns, VSS,
+ 778248.000000ns, VSS,
+ 778248.100000ns, VDD,
+ 778608.300000ns, VDD,
+ 778608.400000ns, VSS,
+ 778968.600000ns, VSS,
+ 778968.700000ns, VDD,
+ 779208.800000ns, VDD,
+ 779208.900000ns, VSS,
+ 780169.600000ns, VSS,
+ 780169.700000ns, VDD,
+ 780890.200000ns, VDD,
+ 780890.300000ns, VSS,
+ 781010.300000ns, VSS,
+ 781010.400000ns, VDD,
+ 781370.600000ns, VDD,
+ 781370.700000ns, VSS,
+ 781490.700000ns, VSS,
+ 781490.800000ns, VDD,
+ 781610.800000ns, VDD,
+ 781610.900000ns, VSS,
+ 781730.900000ns, VSS,
+ 781731.000000ns, VDD,
+ 782331.400000ns, VDD,
+ 782331.500000ns, VSS,
+ 782451.500000ns, VSS,
+ 782451.600000ns, VDD,
+ 782571.600000ns, VDD,
+ 782571.700000ns, VSS,
+ 783412.300000ns, VSS,
+ 783412.400000ns, VDD,
+ 785093.700000ns, VDD,
+ 785093.800000ns, VSS,
+ 785213.800000ns, VSS,
+ 785213.900000ns, VDD,
+ 786294.700000ns, VDD,
+ 786294.800000ns, VSS,
+ 786414.800000ns, VSS,
+ 786414.900000ns, VDD,
+ 786895.200000ns, VDD,
+ 786895.300000ns, VSS,
+ 787255.500000ns, VSS,
+ 787255.600000ns, VDD,
+ 788696.700000ns, VDD,
+ 788696.800000ns, VSS,
+ 789417.300000ns, VSS,
+ 789417.400000ns, VDD,
+ 789537.400000ns, VDD,
+ 789537.500000ns, VSS,
+ 789777.600000ns, VSS,
+ 789777.700000ns, VDD,
+ 789897.700000ns, VDD,
+ 789897.800000ns, VSS,
+ 790017.800000ns, VSS,
+ 790017.900000ns, VDD,
+ 790137.900000ns, VDD,
+ 790138.000000ns, VSS,
+ 790618.300000ns, VSS,
+ 790618.400000ns, VDD,
+ 790858.500000ns, VDD,
+ 790858.600000ns, VSS,
+ 791098.700000ns, VSS,
+ 791098.800000ns, VDD,
+ 791218.800000ns, VDD,
+ 791218.900000ns, VSS,
+ 791338.900000ns, VSS,
+ 791339.000000ns, VDD,
+ 791699.200000ns, VDD,
+ 791699.300000ns, VSS,
+ 792179.600000ns, VSS,
+ 792179.700000ns, VDD,
+ 792539.900000ns, VDD,
+ 792540.000000ns, VSS,
+ 792660.000000ns, VSS,
+ 792660.100000ns, VDD,
+ 792900.200000ns, VDD,
+ 792900.300000ns, VSS,
+ 793861.000000ns, VSS,
+ 793861.100000ns, VDD,
+ 794701.700000ns, VDD,
+ 794701.800000ns, VSS,
+ 795422.300000ns, VSS,
+ 795422.400000ns, VDD,
+ 795662.500000ns, VDD,
+ 795662.600000ns, VSS,
+ 796383.100000ns, VSS,
+ 796383.200000ns, VDD,
+ 796623.300000ns, VDD,
+ 796623.400000ns, VSS,
+ 796863.500000ns, VSS,
+ 796863.600000ns, VDD,
+ 797704.200000ns, VDD,
+ 797704.300000ns, VSS,
+ 798304.700000ns, VSS,
+ 798304.800000ns, VDD,
+ 798424.800000ns, VDD,
+ 798424.900000ns, VSS,
+ 798905.200000ns, VSS,
+ 798905.300000ns, VDD,
+ 799025.300000ns, VDD,
+ 799025.400000ns, VSS,
+ 799505.700000ns, VSS,
+ 799505.800000ns, VDD,
+ 799745.900000ns, VDD,
+ 799746.000000ns, VSS,
+ 800226.300000ns, VSS,
+ 800226.400000ns, VDD,
+ 800946.900000ns, VDD,
+ 800947.000000ns, VSS,
+ 801307.200000ns, VSS,
+ 801307.300000ns, VDD,
+ 801787.600000ns, VDD,
+ 801787.700000ns, VSS,
+ 802508.200000ns, VSS,
+ 802508.300000ns, VDD,
+ 803348.900000ns, VDD,
+ 803349.000000ns, VSS,
+ 803469.000000ns, VSS,
+ 803469.100000ns, VDD,
+ 803949.400000ns, VDD,
+ 803949.500000ns, VSS,
+ 804429.800000ns, VSS,
+ 804429.900000ns, VDD,
+ 804670.000000ns, VDD,
+ 804670.100000ns, VSS,
+ 804910.200000ns, VSS,
+ 804910.300000ns, VDD,
+ 805750.900000ns, VDD,
+ 805751.000000ns, VSS,
+ 806951.900000ns, VSS,
+ 806952.000000ns, VDD,
+ 807432.300000ns, VDD,
+ 807432.400000ns, VSS,
+ 807552.400000ns, VSS,
+ 807552.500000ns, VDD,
+ 808393.100000ns, VDD,
+ 808393.200000ns, VSS,
+ 808513.200000ns, VSS,
+ 808513.300000ns, VDD,
+ 809353.900000ns, VDD,
+ 809354.000000ns, VSS,
+ 809474.000000ns, VSS,
+ 809474.100000ns, VDD,
+ 809954.400000ns, VDD,
+ 809954.500000ns, VSS,
+ 810434.800000ns, VSS,
+ 810434.900000ns, VDD,
+ 811155.400000ns, VDD,
+ 811155.500000ns, VSS,
+ 811635.800000ns, VSS,
+ 811635.900000ns, VDD,
+ 811876.000000ns, VDD,
+ 811876.100000ns, VSS,
+ 811996.100000ns, VSS,
+ 811996.200000ns, VDD,
+ 812236.300000ns, VDD,
+ 812236.400000ns, VSS,
+ 812596.600000ns, VSS,
+ 812596.700000ns, VDD,
+ 812716.700000ns, VDD,
+ 812716.800000ns, VSS,
+ 813197.100000ns, VSS,
+ 813197.200000ns, VDD,
+ 813557.400000ns, VDD,
+ 813557.500000ns, VSS,
+ 813677.500000ns, VSS,
+ 813677.600000ns, VDD,
+ 814037.800000ns, VDD,
+ 814037.900000ns, VSS,
+ 814157.900000ns, VSS,
+ 814158.000000ns, VDD,
+ 814398.100000ns, VDD,
+ 814398.200000ns, VSS,
+ 814998.600000ns, VSS,
+ 814998.700000ns, VDD,
+ 815719.200000ns, VDD,
+ 815719.300000ns, VSS,
+ 816199.600000ns, VSS,
+ 816199.700000ns, VDD,
+ 816439.800000ns, VDD,
+ 816439.900000ns, VSS,
+ 816800.100000ns, VSS,
+ 816800.200000ns, VDD,
+ 816920.200000ns, VDD,
+ 816920.300000ns, VSS,
+ 817400.600000ns, VSS,
+ 817400.700000ns, VDD,
+ 817881.000000ns, VDD,
+ 817881.100000ns, VSS,
+ 818001.100000ns, VSS,
+ 818001.200000ns, VDD,
+ 818241.300000ns, VDD,
+ 818241.400000ns, VSS,
+ 818361.400000ns, VSS,
+ 818361.500000ns, VDD,
+ 818721.700000ns, VDD,
+ 818721.800000ns, VSS,
+ 818961.900000ns, VSS,
+ 818962.000000ns, VDD,
+ 820523.200000ns, VDD,
+ 820523.300000ns, VSS,
+ 820763.400000ns, VSS,
+ 820763.500000ns, VDD,
+ 821243.800000ns, VDD,
+ 821243.900000ns, VSS,
+ 821724.200000ns, VSS,
+ 821724.300000ns, VDD,
+ 822204.600000ns, VDD,
+ 822204.700000ns, VSS,
+ 822324.700000ns, VSS,
+ 822324.800000ns, VDD,
+ 822685.000000ns, VDD,
+ 822685.100000ns, VSS,
+ 822805.100000ns, VSS,
+ 822805.200000ns, VDD,
+ 823405.600000ns, VDD,
+ 823405.700000ns, VSS,
+ 823886.000000ns, VSS,
+ 823886.100000ns, VDD,
+ 824126.200000ns, VDD,
+ 824126.300000ns, VSS,
+ 824366.400000ns, VSS,
+ 824366.500000ns, VDD,
+ 824486.500000ns, VDD,
+ 824486.600000ns, VSS,
+ 824966.900000ns, VSS,
+ 824967.000000ns, VDD,
+ 825327.200000ns, VDD,
+ 825327.300000ns, VSS,
+ 826047.800000ns, VSS,
+ 826047.900000ns, VDD,
+ 826528.200000ns, VDD,
+ 826528.300000ns, VSS,
+ 827248.800000ns, VSS,
+ 827248.900000ns, VDD,
+ 827969.400000ns, VDD,
+ 827969.500000ns, VSS,
+ 828209.600000ns, VSS,
+ 828209.700000ns, VDD,
+ 828329.700000ns, VDD,
+ 828329.800000ns, VSS,
+ 829290.500000ns, VSS,
+ 829290.600000ns, VDD,
+ 829770.900000ns, VDD,
+ 829771.000000ns, VSS,
+ 830251.300000ns, VSS,
+ 830251.400000ns, VDD,
+ 831212.100000ns, VDD,
+ 831212.200000ns, VSS,
+ 831452.300000ns, VSS,
+ 831452.400000ns, VDD,
+ 831812.600000ns, VDD,
+ 831812.700000ns, VSS,
+ 831932.700000ns, VSS,
+ 831932.800000ns, VDD,
+ 832413.100000ns, VDD,
+ 832413.200000ns, VSS,
+ 832533.200000ns, VSS,
+ 832533.300000ns, VDD,
+ 833013.600000ns, VDD,
+ 833013.700000ns, VSS,
+ 833253.800000ns, VSS,
+ 833253.900000ns, VDD,
+ 833614.100000ns, VDD,
+ 833614.200000ns, VSS,
+ 833974.400000ns, VSS,
+ 833974.500000ns, VDD,
+ 834454.800000ns, VDD,
+ 834454.900000ns, VSS,
+ 834695.000000ns, VSS,
+ 834695.100000ns, VDD,
+ 835055.300000ns, VDD,
+ 835055.400000ns, VSS,
+ 835175.400000ns, VSS,
+ 835175.500000ns, VDD,
+ 835535.700000ns, VDD,
+ 835535.800000ns, VSS,
+ 836016.100000ns, VSS,
+ 836016.200000ns, VDD,
+ 836496.500000ns, VDD,
+ 836496.600000ns, VSS,
+ 836616.600000ns, VSS,
+ 836616.700000ns, VDD,
+ 838778.400000ns, VDD,
+ 838778.500000ns, VSS,
+ 838898.500000ns, VSS,
+ 838898.600000ns, VDD,
+ 839258.800000ns, VDD,
+ 839258.900000ns, VSS,
+ 839378.900000ns, VSS,
+ 839379.000000ns, VDD,
+ 839859.300000ns, VDD,
+ 839859.400000ns, VSS,
+ 840219.600000ns, VSS,
+ 840219.700000ns, VDD,
+ 840339.700000ns, VDD,
+ 840339.800000ns, VSS,
+ 840459.800000ns, VSS,
+ 840459.900000ns, VDD,
+ 841060.300000ns, VDD,
+ 841060.400000ns, VSS,
+ 841660.800000ns, VSS,
+ 841660.900000ns, VDD,
+ 842141.200000ns, VDD,
+ 842141.300000ns, VSS,
+ 842261.300000ns, VSS,
+ 842261.400000ns, VDD,
+ 842501.500000ns, VDD,
+ 842501.600000ns, VSS,
+ 842861.800000ns, VSS,
+ 842861.900000ns, VDD,
+ 843462.300000ns, VDD,
+ 843462.400000ns, VSS,
+ 843702.500000ns, VSS,
+ 843702.600000ns, VDD,
+ 844663.300000ns, VDD,
+ 844663.400000ns, VSS,
+ 845504.000000ns, VSS,
+ 845504.100000ns, VDD,
+ 845984.400000ns, VDD,
+ 845984.500000ns, VSS,
+ 846224.600000ns, VSS,
+ 846224.700000ns, VDD,
+ 846344.700000ns, VDD,
+ 846344.800000ns, VSS,
+ 846464.800000ns, VSS,
+ 846464.900000ns, VDD,
+ 846584.900000ns, VDD,
+ 846585.000000ns, VSS,
+ 847185.400000ns, VSS,
+ 847185.500000ns, VDD,
+ 847425.600000ns, VDD,
+ 847425.700000ns, VSS,
+ 847545.700000ns, VSS,
+ 847545.800000ns, VDD,
+ 847785.900000ns, VDD,
+ 847786.000000ns, VSS,
+ 847906.000000ns, VSS,
+ 847906.100000ns, VDD,
+ 848146.200000ns, VDD,
+ 848146.300000ns, VSS,
+ 848386.400000ns, VSS,
+ 848386.500000ns, VDD,
+ 848506.500000ns, VDD,
+ 848506.600000ns, VSS,
+ 848866.800000ns, VSS,
+ 848866.900000ns, VDD,
+ 848986.900000ns, VDD,
+ 848987.000000ns, VSS,
+ 849347.200000ns, VSS,
+ 849347.300000ns, VDD,
+ 850187.900000ns, VDD,
+ 850188.000000ns, VSS,
+ 850908.500000ns, VSS,
+ 850908.600000ns, VDD,
+ 851148.700000ns, VDD,
+ 851148.800000ns, VSS,
+ 851388.900000ns, VSS,
+ 851389.000000ns, VDD,
+ 851749.200000ns, VDD,
+ 851749.300000ns, VSS,
+ 852349.700000ns, VSS,
+ 852349.800000ns, VDD,
+ 852710.000000ns, VDD,
+ 852710.100000ns, VSS,
+ 852950.200000ns, VSS,
+ 852950.300000ns, VDD,
+ 853310.500000ns, VDD,
+ 853310.600000ns, VSS,
+ 853430.600000ns, VSS,
+ 853430.700000ns, VDD,
+ 853550.700000ns, VDD,
+ 853550.800000ns, VSS,
+ 853911.000000ns, VSS,
+ 853911.100000ns, VDD,
+ 854151.200000ns, VDD,
+ 854151.300000ns, VSS,
+ 854271.300000ns, VSS,
+ 854271.400000ns, VDD,
+ 854391.400000ns, VDD,
+ 854391.500000ns, VSS,
+ 854511.500000ns, VSS,
+ 854511.600000ns, VDD,
+ 855232.100000ns, VDD,
+ 855232.200000ns, VSS,
+ 856192.900000ns, VSS,
+ 856193.000000ns, VDD,
+ 856433.100000ns, VDD,
+ 856433.200000ns, VSS,
+ 856553.200000ns, VSS,
+ 856553.300000ns, VDD,
+ 856793.400000ns, VDD,
+ 856793.500000ns, VSS,
+ 857153.700000ns, VSS,
+ 857153.800000ns, VDD,
+ 857393.900000ns, VDD,
+ 857394.000000ns, VSS,
+ 857634.100000ns, VSS,
+ 857634.200000ns, VDD,
+ 857874.300000ns, VDD,
+ 857874.400000ns, VSS,
+ 858234.600000ns, VSS,
+ 858234.700000ns, VDD,
+ 859195.400000ns, VDD,
+ 859195.500000ns, VSS,
+ 859315.500000ns, VSS,
+ 859315.600000ns, VDD,
+ 859675.800000ns, VDD,
+ 859675.900000ns, VSS,
+ 859795.900000ns, VSS,
+ 859796.000000ns, VDD,
+ 860516.500000ns, VDD,
+ 860516.600000ns, VSS,
+ 861357.200000ns, VSS,
+ 861357.300000ns, VDD,
+ 861477.300000ns, VDD,
+ 861477.400000ns, VSS,
+ 862438.100000ns, VSS,
+ 862438.200000ns, VDD,
+ 862558.200000ns, VDD,
+ 862558.300000ns, VSS,
+ 862918.500000ns, VSS,
+ 862918.600000ns, VDD,
+ 863038.600000ns, VDD,
+ 863038.700000ns, VSS,
+ 864479.800000ns, VSS,
+ 864479.900000ns, VDD,
+ 864960.200000ns, VDD,
+ 864960.300000ns, VSS,
+ 865080.300000ns, VSS,
+ 865080.400000ns, VDD,
+ 865440.600000ns, VDD,
+ 865440.700000ns, VSS,
+ 865921.000000ns, VSS,
+ 865921.100000ns, VDD,
+ 866161.200000ns, VDD,
+ 866161.300000ns, VSS,
+ 866281.300000ns, VSS,
+ 866281.400000ns, VDD,
+ 866401.400000ns, VDD,
+ 866401.500000ns, VSS,
+ 866521.500000ns, VSS,
+ 866521.600000ns, VDD,
+ 867122.000000ns, VDD,
+ 867122.100000ns, VSS,
+ 867362.200000ns, VSS,
+ 867362.300000ns, VDD,
+ 867482.300000ns, VDD,
+ 867482.400000ns, VSS,
+ 867602.400000ns, VSS,
+ 867602.500000ns, VDD,
+ 867722.500000ns, VDD,
+ 867722.600000ns, VSS,
+ 868803.400000ns, VSS,
+ 868803.500000ns, VDD,
+ 870244.600000ns, VDD,
+ 870244.700000ns, VSS,
+ 870484.800000ns, VSS,
+ 870484.900000ns, VDD,
+ 870965.200000ns, VDD,
+ 870965.300000ns, VSS,
+ 871205.400000ns, VSS,
+ 871205.500000ns, VDD,
+ 871565.700000ns, VDD,
+ 871565.800000ns, VSS,
+ 871926.000000ns, VSS,
+ 871926.100000ns, VDD,
+ 872046.100000ns, VDD,
+ 872046.200000ns, VSS,
+ 872526.500000ns, VSS,
+ 872526.600000ns, VDD,
+ 872886.800000ns, VDD,
+ 872886.900000ns, VSS,
+ 873006.900000ns, VSS,
+ 873007.000000ns, VDD,
+ 873727.500000ns, VDD,
+ 873727.600000ns, VSS,
+ 873847.600000ns, VSS,
+ 873847.700000ns, VDD,
+ 873967.700000ns, VDD,
+ 873967.800000ns, VSS,
+ 874207.900000ns, VSS,
+ 874208.000000ns, VDD,
+ 874688.300000ns, VDD,
+ 874688.400000ns, VSS,
+ 874928.500000ns, VSS,
+ 874928.600000ns, VDD,
+ 875048.600000ns, VDD,
+ 875048.700000ns, VSS,
+ 875168.700000ns, VSS,
+ 875168.800000ns, VDD,
+ 875769.200000ns, VDD,
+ 875769.300000ns, VSS,
+ 875889.300000ns, VSS,
+ 875889.400000ns, VDD,
+ 876009.400000ns, VDD,
+ 876009.500000ns, VSS,
+ 876249.600000ns, VSS,
+ 876249.700000ns, VDD,
+ 876609.900000ns, VDD,
+ 876610.000000ns, VSS,
+ 877090.300000ns, VSS,
+ 877090.400000ns, VDD,
+ 877330.500000ns, VDD,
+ 877330.600000ns, VSS,
+ 878051.100000ns, VSS,
+ 878051.200000ns, VDD,
+ 878171.200000ns, VDD,
+ 878171.300000ns, VSS,
+ 878651.600000ns, VSS,
+ 878651.700000ns, VDD,
+ 879252.100000ns, VDD,
+ 879252.200000ns, VSS,
+ 879612.400000ns, VSS,
+ 879612.500000ns, VDD,
+ 879852.600000ns, VDD,
+ 879852.700000ns, VSS,
+ 880693.300000ns, VSS,
+ 880693.400000ns, VDD,
+ 881053.600000ns, VDD,
+ 881053.700000ns, VSS,
+ 881774.200000ns, VSS,
+ 881774.300000ns, VDD,
+ 882254.600000ns, VDD,
+ 882254.700000ns, VSS,
+ 882494.800000ns, VSS,
+ 882494.900000ns, VDD,
+ 882735.000000ns, VDD,
+ 882735.100000ns, VSS,
+ 882975.200000ns, VSS,
+ 882975.300000ns, VDD,
+ 883095.300000ns, VDD,
+ 883095.400000ns, VSS,
+ 883215.400000ns, VSS,
+ 883215.500000ns, VDD,
+ 883455.600000ns, VDD,
+ 883455.700000ns, VSS,
+ 883936.000000ns, VSS,
+ 883936.100000ns, VDD,
+ 885377.200000ns, VDD,
+ 885377.300000ns, VSS,
+ 885497.300000ns, VSS,
+ 885497.400000ns, VDD,
+ 885857.600000ns, VDD,
+ 885857.700000ns, VSS,
+ 886097.800000ns, VSS,
+ 886097.900000ns, VDD,
+ 886818.400000ns, VDD,
+ 886818.500000ns, VSS,
+ 886938.500000ns, VSS,
+ 886938.600000ns, VDD,
+ 887178.700000ns, VDD,
+ 887178.800000ns, VSS,
+ 887899.300000ns, VSS,
+ 887899.400000ns, VDD,
+ 888259.600000ns, VDD,
+ 888259.700000ns, VSS,
+ 888619.900000ns, VSS,
+ 888620.000000ns, VDD,
+ 888860.100000ns, VDD,
+ 888860.200000ns, VSS,
+ 889100.300000ns, VSS,
+ 889100.400000ns, VDD,
+ 889340.500000ns, VDD,
+ 889340.600000ns, VSS,
+ 889460.600000ns, VSS,
+ 889460.700000ns, VDD,
+ 890301.300000ns, VDD,
+ 890301.400000ns, VSS,
+ 890541.500000ns, VSS,
+ 890541.600000ns, VDD,
+ 890901.800000ns, VDD,
+ 890901.900000ns, VSS,
+ 891382.200000ns, VSS,
+ 891382.300000ns, VDD,
+ 891742.500000ns, VDD,
+ 891742.600000ns, VSS,
+ 891982.700000ns, VSS,
+ 891982.800000ns, VDD,
+ 892102.800000ns, VDD,
+ 892102.900000ns, VSS,
+ 892463.100000ns, VSS,
+ 892463.200000ns, VDD,
+ 892583.200000ns, VDD,
+ 892583.300000ns, VSS,
+ 893183.700000ns, VSS,
+ 893183.800000ns, VDD,
+ 893303.800000ns, VDD,
+ 893303.900000ns, VSS,
+ 893664.100000ns, VSS,
+ 893664.200000ns, VDD,
+ 894144.500000ns, VDD,
+ 894144.600000ns, VSS,
+ 894264.600000ns, VSS,
+ 894264.700000ns, VDD,
+ 894624.900000ns, VDD,
+ 894625.000000ns, VSS,
+ 895105.300000ns, VSS,
+ 895105.400000ns, VDD,
+ 896066.100000ns, VDD,
+ 896066.200000ns, VSS,
+ 896186.200000ns, VSS,
+ 896186.300000ns, VDD,
+ 897387.200000ns, VDD,
+ 897387.300000ns, VSS,
+ 897627.400000ns, VSS,
+ 897627.500000ns, VDD,
+ 897747.500000ns, VDD,
+ 897747.600000ns, VSS,
+ 897987.700000ns, VSS,
+ 897987.800000ns, VDD,
+ 898468.100000ns, VDD,
+ 898468.200000ns, VSS,
+ 898708.300000ns, VSS,
+ 898708.400000ns, VDD,
+ 899068.600000ns, VDD,
+ 899068.700000ns, VSS,
+ 899308.800000ns, VSS,
+ 899308.900000ns, VDD,
+ 900029.400000ns, VDD,
+ 900029.500000ns, VSS,
+ 900149.500000ns, VSS,
+ 900149.600000ns, VDD,
+ 900269.600000ns, VDD,
+ 900269.700000ns, VSS,
+ 900990.200000ns, VSS,
+ 900990.300000ns, VDD,
+ 901470.600000ns, VDD,
+ 901470.700000ns, VSS,
+ 901710.800000ns, VSS,
+ 901710.900000ns, VDD,
+ 901830.900000ns, VDD,
+ 901831.000000ns, VSS,
+ 902431.400000ns, VSS,
+ 902431.500000ns, VDD,
+ 902671.600000ns, VDD,
+ 902671.700000ns, VSS,
+ 903152.000000ns, VSS,
+ 903152.100000ns, VDD,
+ 903512.300000ns, VDD,
+ 903512.400000ns, VSS,
+ 903632.400000ns, VSS,
+ 903632.500000ns, VDD,
+ 904353.000000ns, VDD,
+ 904353.100000ns, VSS,
+ 904473.100000ns, VSS,
+ 904473.200000ns, VDD,
+ 904593.200000ns, VDD,
+ 904593.300000ns, VSS,
+ 904833.400000ns, VSS,
+ 904833.500000ns, VDD,
+ 905073.600000ns, VDD,
+ 905073.700000ns, VSS,
+ 905554.000000ns, VSS,
+ 905554.100000ns, VDD,
+ 905794.200000ns, VDD,
+ 905794.300000ns, VSS,
+ 906034.400000ns, VSS,
+ 906034.500000ns, VDD,
+ 906514.800000ns, VDD,
+ 906514.900000ns, VSS,
+ 907115.300000ns, VSS,
+ 907115.400000ns, VDD,
+ 908436.400000ns, VDD,
+ 908436.500000ns, VSS,
+ 908676.600000ns, VSS,
+ 908676.700000ns, VDD,
+ 909997.700000ns, VDD,
+ 909997.800000ns, VSS,
+ 910117.800000ns, VSS,
+ 910117.900000ns, VDD,
+ 910358.000000ns, VDD,
+ 910358.100000ns, VSS,
+ 910838.400000ns, VSS,
+ 910838.500000ns, VDD,
+ 911919.300000ns, VDD,
+ 911919.400000ns, VSS,
+ 912399.700000ns, VSS,
+ 912399.800000ns, VDD,
+ 912760.000000ns, VDD,
+ 912760.100000ns, VSS,
+ 912880.100000ns, VSS,
+ 912880.200000ns, VDD,
+ 913961.000000ns, VDD,
+ 913961.100000ns, VSS,
+ 914201.200000ns, VSS,
+ 914201.300000ns, VDD,
+ 914321.300000ns, VDD,
+ 914321.400000ns, VSS,
+ 914681.600000ns, VSS,
+ 914681.700000ns, VDD,
+ 915522.300000ns, VDD,
+ 915522.400000ns, VSS,
+ 915642.400000ns, VSS,
+ 915642.500000ns, VDD,
+ 915762.500000ns, VDD,
+ 915762.600000ns, VSS,
+ 916122.800000ns, VSS,
+ 916122.900000ns, VDD,
+ 916363.000000ns, VDD,
+ 916363.100000ns, VSS,
+ 916603.200000ns, VSS,
+ 916603.300000ns, VDD,
+ 916723.300000ns, VDD,
+ 916723.400000ns, VSS,
+ 917203.700000ns, VSS,
+ 917203.800000ns, VDD,
+ 917443.900000ns, VDD,
+ 917444.000000ns, VSS,
+ 917684.100000ns, VSS,
+ 917684.200000ns, VDD,
+ 919125.300000ns, VDD,
+ 919125.400000ns, VSS,
+ 919966.000000ns, VSS,
+ 919966.100000ns, VDD,
+ 920086.100000ns, VDD,
+ 920086.200000ns, VSS,
+ 920686.600000ns, VSS,
+ 920686.700000ns, VDD,
+ 921167.000000ns, VDD,
+ 921167.100000ns, VSS,
+ 921527.300000ns, VSS,
+ 921527.400000ns, VDD,
+ 922007.700000ns, VDD,
+ 922007.800000ns, VSS,
+ 922488.100000ns, VSS,
+ 922488.200000ns, VDD,
+ 922728.300000ns, VDD,
+ 922728.400000ns, VSS,
+ 924169.500000ns, VSS,
+ 924169.600000ns, VDD,
+ 924289.600000ns, VDD,
+ 924289.700000ns, VSS,
+ 924649.900000ns, VSS,
+ 924650.000000ns, VDD,
+ 925010.200000ns, VDD,
+ 925010.300000ns, VSS,
+ 925370.500000ns, VSS,
+ 925370.600000ns, VDD,
+ 925490.600000ns, VDD,
+ 925490.700000ns, VSS,
+ 925971.000000ns, VSS,
+ 925971.100000ns, VDD,
+ 926211.200000ns, VDD,
+ 926211.300000ns, VSS,
+ 926691.600000ns, VSS,
+ 926691.700000ns, VDD,
+ 927172.000000ns, VDD,
+ 927172.100000ns, VSS,
+ 927292.100000ns, VSS,
+ 927292.200000ns, VDD,
+ 927412.200000ns, VDD,
+ 927412.300000ns, VSS,
+ 927652.400000ns, VSS,
+ 927652.500000ns, VDD,
+ 928373.000000ns, VDD,
+ 928373.100000ns, VSS,
+ 928853.400000ns, VSS,
+ 928853.500000ns, VDD,
+ 929453.900000ns, VDD,
+ 929454.000000ns, VSS,
+ 929694.100000ns, VSS,
+ 929694.200000ns, VDD,
+ 929934.300000ns, VDD,
+ 929934.400000ns, VSS,
+ 930174.500000ns, VSS,
+ 930174.600000ns, VDD,
+ 930414.700000ns, VDD,
+ 930414.800000ns, VSS,
+ 931375.500000ns, VSS,
+ 931375.600000ns, VDD,
+ 931495.600000ns, VDD,
+ 931495.700000ns, VSS,
+ 931615.700000ns, VSS,
+ 931615.800000ns, VDD,
+ 932096.100000ns, VDD,
+ 932096.200000ns, VSS,
+ 932456.400000ns, VSS,
+ 932456.500000ns, VDD,
+ 932816.700000ns, VDD,
+ 932816.800000ns, VSS,
+ 932936.800000ns, VSS,
+ 932936.900000ns, VDD,
+ 933897.600000ns, VDD,
+ 933897.700000ns, VSS,
+ 934017.700000ns, VSS,
+ 934017.800000ns, VDD,
+ 934137.800000ns, VDD,
+ 934137.900000ns, VSS,
+ 934978.500000ns, VSS,
+ 934978.600000ns, VDD,
+ 935699.100000ns, VDD,
+ 935699.200000ns, VSS,
+ 935819.200000ns, VSS,
+ 935819.300000ns, VDD,
+ 936059.400000ns, VDD,
+ 936059.500000ns, VSS,
+ 936299.600000ns, VSS,
+ 936299.700000ns, VDD,
+ 936419.700000ns, VDD,
+ 936419.800000ns, VSS,
+ 936659.900000ns, VSS,
+ 936660.000000ns, VDD,
+ 937020.200000ns, VDD,
+ 937020.300000ns, VSS,
+ 937981.000000ns, VSS,
+ 937981.100000ns, VDD,
+ 938581.500000ns, VDD,
+ 938581.600000ns, VSS,
+ 938941.800000ns, VSS,
+ 938941.900000ns, VDD,
+ 939061.900000ns, VDD,
+ 939062.000000ns, VSS,
+ 939422.200000ns, VSS,
+ 939422.300000ns, VDD,
+ 939662.400000ns, VDD,
+ 939662.500000ns, VSS,
+ 939902.600000ns, VSS,
+ 939902.700000ns, VDD,
+ 940022.700000ns, VDD,
+ 940022.800000ns, VSS,
+ 940623.200000ns, VSS,
+ 940623.300000ns, VDD,
+ 941343.800000ns, VDD,
+ 941343.900000ns, VSS,
+ 941944.300000ns, VSS,
+ 941944.400000ns, VDD,
+ 942064.400000ns, VDD,
+ 942064.500000ns, VSS,
+ 942304.600000ns, VSS,
+ 942304.700000ns, VDD,
+ 942544.800000ns, VDD,
+ 942544.900000ns, VSS,
+ 942664.900000ns, VSS,
+ 942665.000000ns, VDD,
+ 943025.200000ns, VDD,
+ 943025.300000ns, VSS,
+ 943265.400000ns, VSS,
+ 943265.500000ns, VDD,
+ 943505.600000ns, VDD,
+ 943505.700000ns, VSS,
+ 943625.700000ns, VSS,
+ 943625.800000ns, VDD,
+ 943745.800000ns, VDD,
+ 943745.900000ns, VSS,
+ 944106.100000ns, VSS,
+ 944106.200000ns, VDD,
+ 944346.300000ns, VDD,
+ 944346.400000ns, VSS,
+ 944586.500000ns, VSS,
+ 944586.600000ns, VDD,
+ 945187.000000ns, VDD,
+ 945187.100000ns, VSS,
+ 945907.600000ns, VSS,
+ 945907.700000ns, VDD,
+ 946388.000000ns, VDD,
+ 946388.100000ns, VSS,
+ 946748.300000ns, VSS,
+ 946748.400000ns, VDD,
+ 947108.600000ns, VDD,
+ 947108.700000ns, VSS,
+ 947468.900000ns, VSS,
+ 947469.000000ns, VDD,
+ 948309.600000ns, VDD,
+ 948309.700000ns, VSS,
+ 948910.100000ns, VSS,
+ 948910.200000ns, VDD,
+ 949150.300000ns, VDD,
+ 949150.400000ns, VSS,
+ 949390.500000ns, VSS,
+ 949390.600000ns, VDD,
+ 949630.700000ns, VDD,
+ 949630.800000ns, VSS,
+ 949750.800000ns, VSS,
+ 949750.900000ns, VDD,
+ 949991.000000ns, VDD,
+ 949991.100000ns, VSS,
+ 950831.700000ns, VSS,
+ 950831.800000ns, VDD,
+ 951071.900000ns, VDD,
+ 951072.000000ns, VSS,
+ 951432.200000ns, VSS,
+ 951432.300000ns, VDD,
+ 951672.400000ns, VDD,
+ 951672.500000ns, VSS,
+ 951792.500000ns, VSS,
+ 951792.600000ns, VDD,
+ 952032.700000ns, VDD,
+ 952032.800000ns, VSS,
+ 952393.000000ns, VSS,
+ 952393.100000ns, VDD,
+ 952633.200000ns, VDD,
+ 952633.300000ns, VSS,
+ 953473.900000ns, VSS,
+ 953474.000000ns, VDD,
+ 953954.300000ns, VDD,
+ 953954.400000ns, VSS,
+ 954554.800000ns, VSS,
+ 954554.900000ns, VDD,
+ 955155.300000ns, VDD,
+ 955155.400000ns, VSS,
+ 955515.600000ns, VSS,
+ 955515.700000ns, VDD,
+ 955635.700000ns, VDD,
+ 955635.800000ns, VSS,
+ 956236.200000ns, VSS,
+ 956236.300000ns, VDD,
+ 956476.400000ns, VDD,
+ 956476.500000ns, VSS,
+ 956596.500000ns, VSS,
+ 956596.600000ns, VDD,
+ 957317.100000ns, VDD,
+ 957317.200000ns, VSS,
+ 957557.300000ns, VSS,
+ 957557.400000ns, VDD,
+ 957677.400000ns, VDD,
+ 957677.500000ns, VSS,
+ 958398.000000ns, VSS,
+ 958398.100000ns, VDD,
+ 958638.200000ns, VDD,
+ 958638.300000ns, VSS,
+ 959238.700000ns, VSS,
+ 959238.800000ns, VDD,
+ 959478.900000ns, VDD,
+ 959479.000000ns, VSS,
+ 959839.200000ns, VSS,
+ 959839.300000ns, VDD,
+ 960199.500000ns, VDD,
+ 960199.600000ns, VSS,
+ 960319.600000ns, VSS,
+ 960319.700000ns, VDD,
+ 961160.300000ns, VDD,
+ 961160.400000ns, VSS,
+ 961760.800000ns, VSS,
+ 961760.900000ns, VDD,
+ 962721.600000ns, VDD,
+ 962721.700000ns, VSS,
+ 962841.700000ns, VSS,
+ 962841.800000ns, VDD,
+ 963322.100000ns, VDD,
+ 963322.200000ns, VSS,
+ 963442.200000ns, VSS,
+ 963442.300000ns, VDD,
+ 963802.500000ns, VDD,
+ 963802.600000ns, VSS,
+ 963922.600000ns, VSS,
+ 963922.700000ns, VDD,
+ 965363.800000ns, VDD,
+ 965363.900000ns, VSS,
+ 965844.200000ns, VSS,
+ 965844.300000ns, VDD,
+ 966204.500000ns, VDD,
+ 966204.600000ns, VSS,
+ 967045.200000ns, VSS,
+ 967045.300000ns, VDD,
+ 967285.400000ns, VDD,
+ 967285.500000ns, VSS,
+ 967405.500000ns, VSS,
+ 967405.600000ns, VDD,
+ 967525.600000ns, VDD,
+ 967525.700000ns, VSS,
+ 968726.600000ns, VSS,
+ 968726.700000ns, VDD,
+ 969687.400000ns, VDD,
+ 969687.500000ns, VSS,
+ 969927.600000ns, VSS,
+ 969927.700000ns, VDD,
+ 970167.800000ns, VDD,
+ 970167.900000ns, VSS,
+ 971609.000000ns, VSS,
+ 971609.100000ns, VDD,
+ 971729.100000ns, VDD,
+ 971729.200000ns, VSS,
+ 972089.400000ns, VSS,
+ 972089.500000ns, VDD,
+ 972329.600000ns, VDD,
+ 972329.700000ns, VSS,
+ 972569.800000ns, VSS,
+ 972569.900000ns, VDD,
+ 972689.900000ns, VDD,
+ 972690.000000ns, VSS,
+ 973050.200000ns, VSS,
+ 973050.300000ns, VDD,
+ 973290.400000ns, VDD,
+ 973290.500000ns, VSS,
+ 973770.800000ns, VSS,
+ 973770.900000ns, VDD,
+ 974611.500000ns, VDD,
+ 974611.600000ns, VSS,
+ 976172.800000ns, VSS,
+ 976172.900000ns, VDD,
+ 976413.000000ns, VDD,
+ 976413.100000ns, VSS,
+ 976773.300000ns, VSS,
+ 976773.400000ns, VDD,
+ 977493.900000ns, VDD,
+ 977494.000000ns, VSS,
+ 977974.300000ns, VSS,
+ 977974.400000ns, VDD,
+ 978214.500000ns, VDD,
+ 978214.600000ns, VSS,
+ 978454.700000ns, VSS,
+ 978454.800000ns, VDD,
+ 978574.800000ns, VDD,
+ 978574.900000ns, VSS,
+ 979055.200000ns, VSS,
+ 979055.300000ns, VDD,
+ 979415.500000ns, VDD,
+ 979415.600000ns, VSS,
+ 979775.800000ns, VSS,
+ 979775.900000ns, VDD,
+ 980016.000000ns, VDD,
+ 980016.100000ns, VSS,
+ 980496.400000ns, VSS,
+ 980496.500000ns, VDD,
+ 980736.600000ns, VDD,
+ 980736.700000ns, VSS,
+ 980856.700000ns, VSS,
+ 980856.800000ns, VDD,
+ 981096.900000ns, VDD,
+ 981097.000000ns, VSS,
+ 981697.400000ns, VSS,
+ 981697.500000ns, VDD,
+ 981817.500000ns, VDD,
+ 981817.600000ns, VSS,
+ 981937.600000ns, VSS,
+ 981937.700000ns, VDD,
+ 982297.900000ns, VDD,
+ 982298.000000ns, VSS,
+ 982418.000000ns, VSS,
+ 982418.100000ns, VDD,
+ 982658.200000ns, VDD,
+ 982658.300000ns, VSS,
+ 982778.300000ns, VSS,
+ 982778.400000ns, VDD,
+ 983378.800000ns, VDD,
+ 983378.900000ns, VSS,
+ 983498.900000ns, VSS,
+ 983499.000000ns, VDD,
+ 983739.100000ns, VDD,
+ 983739.200000ns, VSS,
+ 984339.600000ns, VSS,
+ 984339.700000ns, VDD,
+ 985060.200000ns, VDD,
+ 985060.300000ns, VSS,
+ 985420.500000ns, VSS,
+ 985420.600000ns, VDD,
+ 985660.700000ns, VDD,
+ 985660.800000ns, VSS,
+ 986021.000000ns, VSS,
+ 986021.100000ns, VDD,
+ 986621.500000ns, VDD,
+ 986621.600000ns, VSS,
+ 987342.100000ns, VSS,
+ 987342.200000ns, VDD,
+ 987702.400000ns, VDD,
+ 987702.500000ns, VSS,
+ 987822.500000ns, VSS,
+ 987822.600000ns, VDD,
+ 988182.800000ns, VDD,
+ 988182.900000ns, VSS,
+ 988543.100000ns, VSS,
+ 988543.200000ns, VDD,
+ 988663.200000ns, VDD,
+ 988663.300000ns, VSS,
+ 989263.700000ns, VSS,
+ 989263.800000ns, VDD,
+ 989624.000000ns, VDD,
+ 989624.100000ns, VSS,
+ 989984.300000ns, VSS,
+ 989984.400000ns, VDD,
+ 990464.700000ns, VDD,
+ 990464.800000ns, VSS,
+ 990945.100000ns, VSS,
+ 990945.200000ns, VDD,
+ 991425.500000ns, VDD,
+ 991425.600000ns, VSS,
+ 991665.700000ns, VSS,
+ 991665.800000ns, VDD,
+ 991785.800000ns, VDD,
+ 991785.900000ns, VSS,
+ 992506.400000ns, VSS,
+ 992506.500000ns, VDD,
+ 992746.600000ns, VDD,
+ 992746.700000ns, VSS,
+ 992866.700000ns, VSS,
+ 992866.800000ns, VDD,
+ 993227.000000ns, VDD,
+ 993227.100000ns, VSS,
+ 993947.600000ns, VSS,
+ 993947.700000ns, VDD,
+ 994187.800000ns, VDD,
+ 994187.900000ns, VSS,
+ 994548.100000ns, VSS,
+ 994548.200000ns, VDD,
+ 995028.500000ns, VDD,
+ 995028.600000ns, VSS,
+ 995148.600000ns, VSS,
+ 995148.700000ns, VDD,
+ 995388.800000ns, VDD,
+ 995388.900000ns, VSS,
+ 995508.900000ns, VSS,
+ 995509.000000ns, VDD,
+ 995869.200000ns, VDD,
+ 995869.300000ns, VSS,
+ 995989.300000ns, VSS,
+ 995989.400000ns, VDD,
+ 996109.400000ns, VDD,
+ 996109.500000ns, VSS,
+ 996589.800000ns, VSS,
+ 996589.900000ns, VDD,
+ 998031.000000ns, VDD,
+ 998031.100000ns, VSS,
+ 998151.100000ns, VSS,
+ 998151.200000ns, VDD,
+ 998631.500000ns, VDD,
+ 998631.600000ns, VSS,
+ 1000553.100000ns, VSS,
+ 1000553.200000ns, VDD,
+ 1001273.700000ns, VDD,
+ 1001273.800000ns, VSS,
+ 1001393.800000ns, VSS,
+ 1001393.900000ns, VDD,
+ 1001754.100000ns, VDD,
+ 1001754.200000ns, VSS,
+ 1002234.500000ns, VSS,
+ 1002234.600000ns, VDD,
+ 1002955.100000ns, VDD,
+ 1002955.200000ns, VSS,
+ 1003435.500000ns, VSS,
+ 1003435.600000ns, VDD,
+ 1004156.100000ns, VDD,
+ 1004156.200000ns, VSS,
+ 1004876.700000ns, VSS,
+ 1004876.800000ns, VDD,
+ 1006077.700000ns, VDD,
+ 1006077.800000ns, VSS,
+ 1006197.800000ns, VSS,
+ 1006197.900000ns, VDD,
+ 1006678.200000ns, VDD,
+ 1006678.300000ns, VSS,
+ 1006798.300000ns, VSS,
+ 1006798.400000ns, VDD,
+ 1007398.800000ns, VDD,
+ 1007398.900000ns, VSS,
+ 1007518.900000ns, VSS,
+ 1007519.000000ns, VDD,
+ 1008119.400000ns, VDD,
+ 1008119.500000ns, VSS,
+ 1008599.800000ns, VSS,
+ 1008599.900000ns, VDD,
+ 1009080.200000ns, VDD,
+ 1009080.300000ns, VSS,
+ 1010521.400000ns, VSS,
+ 1010521.500000ns, VDD,
+ 1010641.500000ns, VDD,
+ 1010641.600000ns, VSS,
+ 1010761.600000ns, VSS,
+ 1010761.700000ns, VDD,
+ 1011121.900000ns, VDD,
+ 1011122.000000ns, VSS,
+ 1011602.300000ns, VSS,
+ 1011602.400000ns, VDD,
+ 1011842.500000ns, VDD,
+ 1011842.600000ns, VSS,
+ 1012322.900000ns, VSS,
+ 1012323.000000ns, VDD,
+ 1012443.000000ns, VDD,
+ 1012443.100000ns, VSS,
+ 1012683.200000ns, VSS,
+ 1012683.300000ns, VDD,
+ 1013043.500000ns, VDD,
+ 1013043.600000ns, VSS,
+ 1013163.600000ns, VSS,
+ 1013163.700000ns, VDD,
+ 1013283.700000ns, VDD,
+ 1013283.800000ns, VSS,
+ 1013644.000000ns, VSS,
+ 1013644.100000ns, VDD,
+ 1013884.200000ns, VDD,
+ 1013884.300000ns, VSS,
+ 1014124.400000ns, VSS,
+ 1014124.500000ns, VDD,
+ 1014244.500000ns, VDD,
+ 1014244.600000ns, VSS,
+ 1014724.900000ns, VSS,
+ 1014725.000000ns, VDD,
+ 1015805.800000ns, VDD,
+ 1015805.900000ns, VSS,
+ 1016046.000000ns, VSS,
+ 1016046.100000ns, VDD,
+ 1016166.100000ns, VDD,
+ 1016166.200000ns, VSS,
+ 1016766.600000ns, VSS,
+ 1016766.700000ns, VDD,
+ 1017367.100000ns, VDD,
+ 1017367.200000ns, VSS,
+ 1017487.200000ns, VSS,
+ 1017487.300000ns, VDD,
+ 1017607.300000ns, VDD,
+ 1017607.400000ns, VSS,
+ 1017727.400000ns, VSS,
+ 1017727.500000ns, VDD,
+ 1018087.700000ns, VDD,
+ 1018087.800000ns, VSS,
+ 1018568.100000ns, VSS,
+ 1018568.200000ns, VDD,
+ 1019048.500000ns, VDD,
+ 1019048.600000ns, VSS,
+ 1019408.800000ns, VSS,
+ 1019408.900000ns, VDD,
+ 1020249.500000ns, VDD,
+ 1020249.600000ns, VSS,
+ 1020489.700000ns, VSS,
+ 1020489.800000ns, VDD,
+ 1020970.100000ns, VDD,
+ 1020970.200000ns, VSS,
+ 1021210.300000ns, VSS,
+ 1021210.400000ns, VDD,
+ 1021810.800000ns, VDD,
+ 1021810.900000ns, VSS,
+ 1022171.100000ns, VSS,
+ 1022171.200000ns, VDD,
+ 1022771.600000ns, VDD,
+ 1022771.700000ns, VSS,
+ 1022891.700000ns, VSS,
+ 1022891.800000ns, VDD,
+ 1024693.200000ns, VDD,
+ 1024693.300000ns, VSS,
+ 1024813.300000ns, VSS,
+ 1024813.400000ns, VDD,
+ 1024933.400000ns, VDD,
+ 1024933.500000ns, VSS,
+ 1025053.500000ns, VSS,
+ 1025053.600000ns, VDD,
+ 1025293.700000ns, VDD,
+ 1025293.800000ns, VSS,
+ 1026134.400000ns, VSS,
+ 1026134.500000ns, VDD,
+ 1026494.700000ns, VDD,
+ 1026494.800000ns, VSS,
+ 1026614.800000ns, VSS,
+ 1026614.900000ns, VDD,
+ 1027095.200000ns, VDD,
+ 1027095.300000ns, VSS,
+ 1028296.200000ns, VSS,
+ 1028296.300000ns, VDD,
+ 1029377.100000ns, VDD,
+ 1029377.200000ns, VSS,
+ 1029857.500000ns, VSS,
+ 1029857.600000ns, VDD,
+ 1030097.700000ns, VDD,
+ 1030097.800000ns, VSS,
+ 1030337.900000ns, VSS,
+ 1030338.000000ns, VDD,
+ 1030458.000000ns, VDD,
+ 1030458.100000ns, VSS,
+ 1031298.700000ns, VSS,
+ 1031298.800000ns, VDD,
+ 1031779.100000ns, VDD,
+ 1031779.200000ns, VSS,
+ 1031899.200000ns, VSS,
+ 1031899.300000ns, VDD,
+ 1032139.400000ns, VDD,
+ 1032139.500000ns, VSS,
+ 1033100.200000ns, VSS,
+ 1033100.300000ns, VDD,
+ 1033580.600000ns, VDD,
+ 1033580.700000ns, VSS,
+ 1033820.800000ns, VSS,
+ 1033820.900000ns, VDD,
+ 1035382.100000ns, VDD,
+ 1035382.200000ns, VSS,
+ 1036463.000000ns, VSS,
+ 1036463.100000ns, VDD,
+ 1037183.600000ns, VDD,
+ 1037183.700000ns, VSS,
+ 1037303.700000ns, VSS,
+ 1037303.800000ns, VDD,
+ 1037904.200000ns, VDD,
+ 1037904.300000ns, VSS,
+ 1038024.300000ns, VSS,
+ 1038024.400000ns, VDD,
+ 1038144.400000ns, VDD,
+ 1038144.500000ns, VSS,
+ 1038264.500000ns, VSS,
+ 1038264.600000ns, VDD,
+ 1038865.000000ns, VDD,
+ 1038865.100000ns, VSS,
+ 1039225.300000ns, VSS,
+ 1039225.400000ns, VDD,
+ 1039465.500000ns, VDD,
+ 1039465.600000ns, VSS,
+ 1040426.300000ns, VSS,
+ 1040426.400000ns, VDD,
+ 1041387.100000ns, VDD,
+ 1041387.200000ns, VSS,
+ 1042107.700000ns, VSS,
+ 1042107.800000ns, VDD,
+ 1042347.900000ns, VDD,
+ 1042348.000000ns, VSS,
+ 1043548.900000ns, VSS,
+ 1043549.000000ns, VDD,
+ 1044029.300000ns, VDD,
+ 1044029.400000ns, VSS,
+ 1044629.800000ns, VSS,
+ 1044629.900000ns, VDD,
+ 1044990.100000ns, VDD,
+ 1044990.200000ns, VSS,
+ 1045590.600000ns, VSS,
+ 1045590.700000ns, VDD,
+ 1046191.100000ns, VDD,
+ 1046191.200000ns, VSS,
+ 1046671.500000ns, VSS,
+ 1046671.600000ns, VDD,
+ 1047151.900000ns, VDD,
+ 1047152.000000ns, VSS,
+ 1048713.200000ns, VSS,
+ 1048713.300000ns, VDD,
+ 1049193.600000ns, VDD,
+ 1049193.700000ns, VSS,
+ 1049794.100000ns, VSS,
+ 1049794.200000ns, VDD,
+ 1050154.400000ns, VDD,
+ 1050154.500000ns, VSS,
+ 1050274.500000ns, VSS,
+ 1050274.600000ns, VDD,
+ 1050875.000000ns, VDD,
+ 1050875.100000ns, VSS,
+ 1051115.200000ns, VSS,
+ 1051115.300000ns, VDD,
+ 1051715.700000ns, VDD,
+ 1051715.800000ns, VSS,
+ 1051835.800000ns, VSS,
+ 1051835.900000ns, VDD,
+ 1052196.100000ns, VDD,
+ 1052196.200000ns, VSS,
+ 1052316.200000ns, VSS,
+ 1052316.300000ns, VDD,
+ 1052916.700000ns, VDD,
+ 1052916.800000ns, VSS,
+ 1053277.000000ns, VSS,
+ 1053277.100000ns, VDD,
+ 1053397.100000ns, VDD,
+ 1053397.200000ns, VSS,
+ 1053877.500000ns, VSS,
+ 1053877.600000ns, VDD,
+ 1053997.600000ns, VDD,
+ 1053997.700000ns, VSS,
+ 1054237.800000ns, VSS,
+ 1054237.900000ns, VDD,
+ 1055558.900000ns, VDD,
+ 1055559.000000ns, VSS,
+ 1055679.000000ns, VSS,
+ 1055679.100000ns, VDD,
+ 1055919.200000ns, VDD,
+ 1055919.300000ns, VSS,
+ 1056880.000000ns, VSS,
+ 1056880.100000ns, VDD,
+ 1057360.400000ns, VDD,
+ 1057360.500000ns, VSS,
+ 1057480.500000ns, VSS,
+ 1057480.600000ns, VDD,
+ 1057720.700000ns, VDD,
+ 1057720.800000ns, VSS,
+ 1057960.900000ns, VSS,
+ 1057961.000000ns, VDD,
+ 1058441.300000ns, VDD,
+ 1058441.400000ns, VSS,
+ 1058801.600000ns, VSS,
+ 1058801.700000ns, VDD,
+ 1058921.700000ns, VDD,
+ 1058921.800000ns, VSS,
+ 1059161.900000ns, VSS,
+ 1059162.000000ns, VDD,
+ 1059522.200000ns, VDD,
+ 1059522.300000ns, VSS,
+ 1059642.300000ns, VSS,
+ 1059642.400000ns, VDD,
+ 1059882.500000ns, VDD,
+ 1059882.600000ns, VSS,
+ 1060242.800000ns, VSS,
+ 1060242.900000ns, VDD,
+ 1060483.000000ns, VDD,
+ 1060483.100000ns, VSS,
+ 1060603.100000ns, VSS,
+ 1060603.200000ns, VDD,
+ 1060723.200000ns, VDD,
+ 1060723.300000ns, VSS,
+ 1060963.400000ns, VSS,
+ 1060963.500000ns, VDD,
+ 1061323.700000ns, VDD,
+ 1061323.800000ns, VSS,
+ 1061563.900000ns, VSS,
+ 1061564.000000ns, VDD,
+ 1062044.300000ns, VDD,
+ 1062044.400000ns, VSS,
+ 1062404.600000ns, VSS,
+ 1062404.700000ns, VDD,
+ 1062524.700000ns, VDD,
+ 1062524.800000ns, VSS,
+ 1062644.800000ns, VSS,
+ 1062644.900000ns, VDD,
+ 1063125.200000ns, VDD,
+ 1063125.300000ns, VSS,
+ 1063245.300000ns, VSS,
+ 1063245.400000ns, VDD,
+ 1063605.600000ns, VDD,
+ 1063605.700000ns, VSS,
+ 1063725.700000ns, VSS,
+ 1063725.800000ns, VDD,
+ 1064206.100000ns, VDD,
+ 1064206.200000ns, VSS,
+ 1064446.300000ns, VSS,
+ 1064446.400000ns, VDD,
+ 1064566.400000ns, VDD,
+ 1064566.500000ns, VSS,
+ 1064686.500000ns, VSS,
+ 1064686.600000ns, VDD,
+ 1065407.100000ns, VDD,
+ 1065407.200000ns, VSS,
+ 1066247.800000ns, VSS,
+ 1066247.900000ns, VDD,
+ 1066608.100000ns, VDD,
+ 1066608.200000ns, VSS,
+ 1066848.300000ns, VSS,
+ 1066848.400000ns, VDD,
+ 1067208.600000ns, VDD,
+ 1067208.700000ns, VSS,
+ 1067568.900000ns, VSS,
+ 1067569.000000ns, VDD,
+ 1068289.500000ns, VDD,
+ 1068289.600000ns, VSS,
+ 1068649.800000ns, VSS,
+ 1068649.900000ns, VDD,
+ 1069130.200000ns, VDD,
+ 1069130.300000ns, VSS,
+ 1069850.800000ns, VSS,
+ 1069850.900000ns, VDD,
+ 1070451.300000ns, VDD,
+ 1070451.400000ns, VSS,
+ 1070691.500000ns, VSS,
+ 1070691.600000ns, VDD,
+ 1071171.900000ns, VDD,
+ 1071172.000000ns, VSS,
+ 1071892.500000ns, VSS,
+ 1071892.600000ns, VDD,
+ 1072012.600000ns, VDD,
+ 1072012.700000ns, VSS,
+ 1072372.900000ns, VSS,
+ 1072373.000000ns, VDD,
+ 1072493.000000ns, VDD,
+ 1072493.100000ns, VSS,
+ 1073093.500000ns, VSS,
+ 1073093.600000ns, VDD,
+ 1073333.700000ns, VDD,
+ 1073333.800000ns, VSS,
+ 1073453.800000ns, VSS,
+ 1073453.900000ns, VDD,
+ 1074054.300000ns, VDD,
+ 1074054.400000ns, VSS,
+ 1075255.300000ns, VSS,
+ 1075255.400000ns, VDD,
+ 1075855.800000ns, VDD,
+ 1075855.900000ns, VSS,
+ 1076096.000000ns, VSS,
+ 1076096.100000ns, VDD,
+ 1076216.100000ns, VDD,
+ 1076216.200000ns, VSS,
+ 1076336.200000ns, VSS,
+ 1076336.300000ns, VDD,
+ 1077537.200000ns, VDD,
+ 1077537.300000ns, VSS,
+ 1077657.300000ns, VSS,
+ 1077657.400000ns, VDD,
+ 1078017.600000ns, VDD,
+ 1078017.700000ns, VSS,
+ 1078137.700000ns, VSS,
+ 1078137.800000ns, VDD,
+ 1078257.800000ns, VDD,
+ 1078257.900000ns, VSS,
+ 1078498.000000ns, VSS,
+ 1078498.100000ns, VDD,
+ 1078978.400000ns, VDD,
+ 1078978.500000ns, VSS,
+ 1079098.500000ns, VSS,
+ 1079098.600000ns, VDD,
+ 1079218.600000ns, VDD,
+ 1079218.700000ns, VSS,
+ 1079338.700000ns, VSS,
+ 1079338.800000ns, VDD,
+ 1079699.000000ns, VDD,
+ 1079699.100000ns, VSS,
+ 1080059.300000ns, VSS,
+ 1080059.400000ns, VDD,
+ 1080419.600000ns, VDD,
+ 1080419.700000ns, VSS,
+ 1080659.800000ns, VSS,
+ 1080659.900000ns, VDD,
+ 1081140.200000ns, VDD,
+ 1081140.300000ns, VSS,
+ 1082821.600000ns, VSS,
+ 1082821.700000ns, VDD,
+ 1083061.800000ns, VDD,
+ 1083061.900000ns, VSS,
+ 1083181.900000ns, VSS,
+ 1083182.000000ns, VDD,
+ 1083302.000000ns, VDD,
+ 1083302.100000ns, VSS,
+ 1083782.400000ns, VSS,
+ 1083782.500000ns, VDD,
+ 1084262.800000ns, VDD,
+ 1084262.900000ns, VSS,
+ 1084503.000000ns, VSS,
+ 1084503.100000ns, VDD,
+ 1084983.400000ns, VDD,
+ 1084983.500000ns, VSS,
+ 1085223.600000ns, VSS,
+ 1085223.700000ns, VDD,
+ 1085704.000000ns, VDD,
+ 1085704.100000ns, VSS,
+ 1085944.200000ns, VSS,
+ 1085944.300000ns, VDD,
+ 1086184.400000ns, VDD,
+ 1086184.500000ns, VSS,
+ 1086304.500000ns, VSS,
+ 1086304.600000ns, VDD,
+ 1086424.600000ns, VDD,
+ 1086424.700000ns, VSS,
+ 1086544.700000ns, VSS,
+ 1086544.800000ns, VDD,
+ 1086905.000000ns, VDD,
+ 1086905.100000ns, VSS,
+ 1087385.400000ns, VSS,
+ 1087385.500000ns, VDD,
+ 1088586.400000ns, VDD,
+ 1088586.500000ns, VSS,
+ 1088706.500000ns, VSS,
+ 1088706.600000ns, VDD,
+ 1088826.600000ns, VDD,
+ 1088826.700000ns, VSS,
+ 1089066.800000ns, VSS,
+ 1089066.900000ns, VDD,
+ 1089186.900000ns, VDD,
+ 1089187.000000ns, VSS,
+ 1089307.000000ns, VSS,
+ 1089307.100000ns, VDD,
+ 1089427.100000ns, VDD,
+ 1089427.200000ns, VSS,
+ 1090748.200000ns, VSS,
+ 1090748.300000ns, VDD,
+ 1090868.300000ns, VDD,
+ 1090868.400000ns, VSS,
+ 1090988.400000ns, VSS,
+ 1090988.500000ns, VDD,
+ 1091228.600000ns, VDD,
+ 1091228.700000ns, VSS,
+ 1091348.700000ns, VSS,
+ 1091348.800000ns, VDD,
+ 1091709.000000ns, VDD,
+ 1091709.100000ns, VSS,
+ 1091949.200000ns, VSS,
+ 1091949.300000ns, VDD,
+ 1092189.400000ns, VDD,
+ 1092189.500000ns, VSS,
+ 1092309.500000ns, VSS,
+ 1092309.600000ns, VDD,
+ 1092669.800000ns, VDD,
+ 1092669.900000ns, VSS,
+ 1093150.200000ns, VSS,
+ 1093150.300000ns, VDD,
+ 1094111.000000ns, VDD,
+ 1094111.100000ns, VSS,
+ 1094471.300000ns, VSS,
+ 1094471.400000ns, VDD,
+ 1094831.600000ns, VDD,
+ 1094831.700000ns, VSS,
+ 1095071.800000ns, VSS,
+ 1095071.900000ns, VDD,
+ 1095552.200000ns, VDD,
+ 1095552.300000ns, VSS,
+ 1095672.300000ns, VSS,
+ 1095672.400000ns, VDD,
+ 1096753.200000ns, VDD,
+ 1096753.300000ns, VSS,
+ 1096993.400000ns, VSS,
+ 1096993.500000ns, VDD,
+ 1097714.000000ns, VDD,
+ 1097714.100000ns, VSS,
+ 1098194.400000ns, VSS,
+ 1098194.500000ns, VDD,
+ 1098434.600000ns, VDD,
+ 1098434.700000ns, VSS,
+ 1098554.700000ns, VSS,
+ 1098554.800000ns, VDD,
+ 1098674.800000ns, VDD,
+ 1098674.900000ns, VSS,
+ 1098915.000000ns, VSS,
+ 1098915.100000ns, VDD,
+ 1099035.100000ns, VDD,
+ 1099035.200000ns, VSS,
+ 1099155.200000ns, VSS,
+ 1099155.300000ns, VDD,
+ 1099635.600000ns, VDD,
+ 1099635.700000ns, VSS,
+ 1099995.900000ns, VSS,
+ 1099996.000000ns, VDD,
+ 1100236.100000ns, VDD,
+ 1100236.200000ns, VSS,
+ 1100356.200000ns, VSS,
+ 1100356.300000ns, VDD,
+ 1100716.500000ns, VDD,
+ 1100716.600000ns, VSS,
+ 1101196.900000ns, VSS,
+ 1101197.000000ns, VDD,
+ 1101317.000000ns, VDD,
+ 1101317.100000ns, VSS,
+ 1101677.300000ns, VSS,
+ 1101677.400000ns, VDD,
+ 1103118.500000ns, VDD,
+ 1103118.600000ns, VSS,
+ 1103238.600000ns, VSS,
+ 1103238.700000ns, VDD,
+ 1103598.900000ns, VDD,
+ 1103599.000000ns, VSS,
+ 1104079.300000ns, VSS,
+ 1104079.400000ns, VDD,
+ 1104199.400000ns, VDD,
+ 1104199.500000ns, VSS,
+ 1104559.700000ns, VSS,
+ 1104559.800000ns, VDD,
+ 1104679.800000ns, VDD,
+ 1104679.900000ns, VSS,
+ 1104920.000000ns, VSS,
+ 1104920.100000ns, VDD,
+ 1106241.100000ns, VDD,
+ 1106241.200000ns, VSS,
+ 1106481.300000ns, VSS,
+ 1106481.400000ns, VDD,
+ 1106601.400000ns, VDD,
+ 1106601.500000ns, VSS,
+ 1106721.500000ns, VSS,
+ 1106721.600000ns, VDD,
+ 1107322.000000ns, VDD,
+ 1107322.100000ns, VSS,
+ 1107442.100000ns, VSS,
+ 1107442.200000ns, VDD,
+ 1107922.500000ns, VDD,
+ 1107922.600000ns, VSS,
+ 1108282.800000ns, VSS,
+ 1108282.900000ns, VDD,
+ 1108643.100000ns, VDD,
+ 1108643.200000ns, VSS,
+ 1108763.200000ns, VSS,
+ 1108763.300000ns, VDD,
+ 1110204.400000ns, VDD,
+ 1110204.500000ns, VSS,
+ 1110684.800000ns, VSS,
+ 1110684.900000ns, VDD,
+ 1111405.400000ns, VDD,
+ 1111405.500000ns, VSS,
+ 1112126.000000ns, VSS,
+ 1112126.100000ns, VDD,
+ 1113206.900000ns, VDD,
+ 1113207.000000ns, VSS,
+ 1113687.300000ns, VSS,
+ 1113687.400000ns, VDD,
+ 1114047.600000ns, VDD,
+ 1114047.700000ns, VSS,
+ 1114167.700000ns, VSS,
+ 1114167.800000ns, VDD,
+ 1114407.900000ns, VDD,
+ 1114408.000000ns, VSS,
+ 1114528.000000ns, VSS,
+ 1114528.100000ns, VDD,
+ 1114888.300000ns, VDD,
+ 1114888.400000ns, VSS,
+ 1115008.400000ns, VSS,
+ 1115008.500000ns, VDD,
+ 1115368.700000ns, VDD,
+ 1115368.800000ns, VSS,
+ 1116089.300000ns, VSS,
+ 1116089.400000ns, VDD,
+ 1116689.800000ns, VDD,
+ 1116689.900000ns, VSS,
+ 1116930.000000ns, VSS,
+ 1116930.100000ns, VDD,
+ 1117530.500000ns, VDD,
+ 1117530.600000ns, VSS,
+ 1117650.600000ns, VSS,
+ 1117650.700000ns, VDD,
+ 1118010.900000ns, VDD,
+ 1118011.000000ns, VSS,
+ 1118611.400000ns, VSS,
+ 1118611.500000ns, VDD,
+ 1118731.500000ns, VDD,
+ 1118731.600000ns, VSS,
+ 1118971.700000ns, VSS,
+ 1118971.800000ns, VDD,
+ 1119572.200000ns, VDD,
+ 1119572.300000ns, VSS,
+ 1119692.300000ns, VSS,
+ 1119692.400000ns, VDD,
+ 1120052.600000ns, VDD,
+ 1120052.700000ns, VSS,
+ 1120172.700000ns, VSS,
+ 1120172.800000ns, VDD,
+ 1120653.100000ns, VDD,
+ 1120653.200000ns, VSS,
+ 1121133.500000ns, VSS,
+ 1121133.600000ns, VDD,
+ 1121734.000000ns, VDD,
+ 1121734.100000ns, VSS,
+ 1122094.300000ns, VSS,
+ 1122094.400000ns, VDD,
+ 1122334.500000ns, VDD,
+ 1122334.600000ns, VSS,
+ 1122454.600000ns, VSS,
+ 1122454.700000ns, VDD,
+ 1122574.700000ns, VDD,
+ 1122574.800000ns, VSS,
+ 1122814.900000ns, VSS,
+ 1122815.000000ns, VDD,
+ 1123175.200000ns, VDD,
+ 1123175.300000ns, VSS,
+ 1123775.700000ns, VSS,
+ 1123775.800000ns, VDD,
+ 1124376.200000ns, VDD,
+ 1124376.300000ns, VSS,
+ 1124736.500000ns, VSS,
+ 1124736.600000ns, VDD,
+ 1124976.700000ns, VDD,
+ 1124976.800000ns, VSS,
+ 1125096.800000ns, VSS,
+ 1125096.900000ns, VDD,
+ 1125216.900000ns, VDD,
+ 1125217.000000ns, VSS,
+ 1125337.000000ns, VSS,
+ 1125337.100000ns, VDD,
+ 1125937.500000ns, VDD,
+ 1125937.600000ns, VSS,
+ 1126177.700000ns, VSS,
+ 1126177.800000ns, VDD,
+ 1126417.900000ns, VDD,
+ 1126418.000000ns, VSS,
+ 1126778.200000ns, VSS,
+ 1126778.300000ns, VDD,
+ 1127378.700000ns, VDD,
+ 1127378.800000ns, VSS,
+ 1128819.900000ns, VSS,
+ 1128820.000000ns, VDD,
+ 1129780.700000ns, VDD,
+ 1129780.800000ns, VSS,
+ 1130621.400000ns, VSS,
+ 1130621.500000ns, VDD,
+ 1130861.600000ns, VDD,
+ 1130861.700000ns, VSS,
+ 1131221.900000ns, VSS,
+ 1131222.000000ns, VDD,
+ 1131462.100000ns, VDD,
+ 1131462.200000ns, VSS,
+ 1131942.500000ns, VSS,
+ 1131942.600000ns, VDD,
+ 1132182.700000ns, VDD,
+ 1132182.800000ns, VSS,
+ 1133143.500000ns, VSS,
+ 1133143.600000ns, VDD,
+ 1133263.600000ns, VDD,
+ 1133263.700000ns, VSS,
+ 1133864.100000ns, VSS,
+ 1133864.200000ns, VDD,
+ 1134464.600000ns, VDD,
+ 1134464.700000ns, VSS,
+ 1134704.800000ns, VSS,
+ 1134704.900000ns, VDD,
+ 1134824.900000ns, VDD,
+ 1134825.000000ns, VSS,
+ 1135305.300000ns, VSS,
+ 1135305.400000ns, VDD,
+ 1135665.600000ns, VDD,
+ 1135665.700000ns, VSS,
+ 1136025.900000ns, VSS,
+ 1136026.000000ns, VDD,
+ 1136146.000000ns, VDD,
+ 1136146.100000ns, VSS,
+ 1136386.200000ns, VSS,
+ 1136386.300000ns, VDD,
+ 1136626.400000ns, VDD,
+ 1136626.500000ns, VSS,
+ 1136746.500000ns, VSS,
+ 1136746.600000ns, VDD,
+ 1136866.600000ns, VDD,
+ 1136866.700000ns, VSS,
+ 1138307.800000ns, VSS,
+ 1138307.900000ns, VDD,
+ 1138427.900000ns, VDD,
+ 1138428.000000ns, VSS,
+ 1138788.200000ns, VSS,
+ 1138788.300000ns, VDD,
+ 1139628.900000ns, VDD,
+ 1139629.000000ns, VSS,
+ 1139869.100000ns, VSS,
+ 1139869.200000ns, VDD,
+ 1140349.500000ns, VDD,
+ 1140349.600000ns, VSS,
+ 1140589.700000ns, VSS,
+ 1140589.800000ns, VDD,
+ 1140709.800000ns, VDD,
+ 1140709.900000ns, VSS,
+ 1140829.900000ns, VSS,
+ 1140830.000000ns, VDD,
+ 1141310.300000ns, VDD,
+ 1141310.400000ns, VSS,
+ 1141430.400000ns, VSS,
+ 1141430.500000ns, VDD,
+ 1141790.700000ns, VDD,
+ 1141790.800000ns, VSS,
+ 1141910.800000ns, VSS,
+ 1141910.900000ns, VDD,
+ 1143352.000000ns, VDD,
+ 1143352.100000ns, VSS,
+ 1143712.300000ns, VSS,
+ 1143712.400000ns, VDD,
+ 1144312.800000ns, VDD,
+ 1144312.900000ns, VSS,
+ 1144432.900000ns, VSS,
+ 1144433.000000ns, VDD,
+ 1144793.200000ns, VDD,
+ 1144793.300000ns, VSS,
+ 1144913.300000ns, VSS,
+ 1144913.400000ns, VDD,
+ 1145273.600000ns, VDD,
+ 1145273.700000ns, VSS,
+ 1145994.200000ns, VSS,
+ 1145994.300000ns, VDD,
+ 1146114.300000ns, VDD,
+ 1146114.400000ns, VSS,
+ 1147195.200000ns, VSS,
+ 1147195.300000ns, VDD,
+ 1147435.400000ns, VDD,
+ 1147435.500000ns, VSS,
+ 1147675.600000ns, VSS,
+ 1147675.700000ns, VDD,
+ 1148396.200000ns, VDD,
+ 1148396.300000ns, VSS,
+ 1148516.300000ns, VSS,
+ 1148516.400000ns, VDD,
+ 1150317.800000ns, VDD,
+ 1150317.900000ns, VSS,
+ 1151158.500000ns, VSS,
+ 1151158.600000ns, VDD,
+ 1151398.700000ns, VDD,
+ 1151398.800000ns, VSS,
+ 1151999.200000ns, VSS,
+ 1151999.300000ns, VDD,
+ 1152119.300000ns, VDD,
+ 1152119.400000ns, VSS,
+ 1152239.400000ns, VSS,
+ 1152239.500000ns, VDD,
+ 1152479.600000ns, VDD,
+ 1152479.700000ns, VSS,
+ 1152839.900000ns, VSS,
+ 1152840.000000ns, VDD,
+ 1153440.400000ns, VDD,
+ 1153440.500000ns, VSS,
+ 1153920.800000ns, VSS,
+ 1153920.900000ns, VDD,
+ 1155241.900000ns, VDD,
+ 1155242.000000ns, VSS,
+ 1155362.000000ns, VSS,
+ 1155362.100000ns, VDD,
+ 1155602.200000ns, VDD,
+ 1155602.300000ns, VSS,
+ 1155722.300000ns, VSS,
+ 1155722.400000ns, VDD,
+ 1156082.600000ns, VDD,
+ 1156082.700000ns, VSS,
+ 1157163.500000ns, VSS,
+ 1157163.600000ns, VDD,
+ 1157283.600000ns, VDD,
+ 1157283.700000ns, VSS,
+ 1158124.300000ns, VSS,
+ 1158124.400000ns, VDD,
+ 1158364.500000ns, VDD,
+ 1158364.600000ns, VSS,
+ 1158484.600000ns, VSS,
+ 1158484.700000ns, VDD,
+ 1158724.800000ns, VDD,
+ 1158724.900000ns, VSS,
+ 1158965.000000ns, VSS,
+ 1158965.100000ns, VDD,
+ 1159325.300000ns, VDD,
+ 1159325.400000ns, VSS,
+ 1160406.200000ns, VSS,
+ 1160406.300000ns, VDD,
+ 1160646.400000ns, VDD,
+ 1160646.500000ns, VSS,
+ 1161126.800000ns, VSS,
+ 1161126.900000ns, VDD,
+ 1161607.200000ns, VDD,
+ 1161607.300000ns, VSS,
+ 1161967.500000ns, VSS,
+ 1161967.600000ns, VDD,
+ 1162808.200000ns, VDD,
+ 1162808.300000ns, VSS,
+ 1163288.600000ns, VSS,
+ 1163288.700000ns, VDD,
+ 1163528.800000ns, VDD,
+ 1163528.900000ns, VSS,
+ 1163648.900000ns, VSS,
+ 1163649.000000ns, VDD,
+ 1163769.000000ns, VDD,
+ 1163769.100000ns, VSS,
+ 1163889.100000ns, VSS,
+ 1163889.200000ns, VDD,
+ 1164609.700000ns, VDD,
+ 1164609.800000ns, VSS,
+ 1165330.300000ns, VSS,
+ 1165330.400000ns, VDD,
+ 1165450.400000ns, VDD,
+ 1165450.500000ns, VSS,
+ 1165810.700000ns, VSS,
+ 1165810.800000ns, VDD,
+ 1167251.900000ns, VDD,
+ 1167252.000000ns, VSS,
+ 1167612.200000ns, VSS,
+ 1167612.300000ns, VDD,
+ 1168573.000000ns, VDD,
+ 1168573.100000ns, VSS,
+ 1168693.100000ns, VSS,
+ 1168693.200000ns, VDD,
+ 1169053.400000ns, VDD,
+ 1169053.500000ns, VSS,
+ 1169293.600000ns, VSS,
+ 1169293.700000ns, VDD,
+ 1169413.700000ns, VDD,
+ 1169413.800000ns, VSS,
+ 1169653.900000ns, VSS,
+ 1169654.000000ns, VDD,
+ 1170014.200000ns, VDD,
+ 1170014.300000ns, VSS,
+ 1170134.300000ns, VSS,
+ 1170134.400000ns, VDD,
+ 1170254.400000ns, VDD,
+ 1170254.500000ns, VSS,
+ 1170614.700000ns, VSS,
+ 1170614.800000ns, VDD,
+ 1171095.100000ns, VDD,
+ 1171095.200000ns, VSS,
+ 1171695.600000ns, VSS,
+ 1171695.700000ns, VDD,
+ 1173016.700000ns, VDD,
+ 1173016.800000ns, VSS,
+ 1173737.300000ns, VSS,
+ 1173737.400000ns, VDD,
+ 1174097.600000ns, VDD,
+ 1174097.700000ns, VSS,
+ 1174818.200000ns, VSS,
+ 1174818.300000ns, VDD,
+ 1176019.200000ns, VDD,
+ 1176019.300000ns, VSS,
+ 1176259.400000ns, VSS,
+ 1176259.500000ns, VDD,
+ 1176739.800000ns, VDD,
+ 1176739.900000ns, VSS,
+ 1176859.900000ns, VSS,
+ 1176860.000000ns, VDD,
+ 1177580.500000ns, VDD,
+ 1177580.600000ns, VSS,
+ 1177820.700000ns, VSS,
+ 1177820.800000ns, VDD,
+ 1177940.800000ns, VDD,
+ 1177940.900000ns, VSS,
+ 1178421.200000ns, VSS,
+ 1178421.300000ns, VDD,
+ 1179141.800000ns, VDD,
+ 1179141.900000ns, VSS,
+ 1179742.300000ns, VSS,
+ 1179742.400000ns, VDD,
+ 1179862.400000ns, VDD,
+ 1179862.500000ns, VSS,
+ 1180222.700000ns, VSS,
+ 1180222.800000ns, VDD,
+ 1180342.800000ns, VDD,
+ 1180342.900000ns, VSS,
+ 1181063.400000ns, VSS,
+ 1181063.500000ns, VDD,
+ 1181183.500000ns, VDD,
+ 1181183.600000ns, VSS,
+ 1181303.600000ns, VSS,
+ 1181303.700000ns, VDD,
+ 1181543.800000ns, VDD,
+ 1181543.900000ns, VSS,
+ 1182024.200000ns, VSS,
+ 1182024.300000ns, VDD,
+ 1183705.600000ns, VDD,
+ 1183705.700000ns, VSS,
+ 1184666.400000ns, VSS,
+ 1184666.500000ns, VDD,
+ 1184906.600000ns, VDD,
+ 1184906.700000ns, VSS,
+ 1185266.900000ns, VSS,
+ 1185267.000000ns, VDD,
+ 1185747.300000ns, VDD,
+ 1185747.400000ns, VSS,
+ 1185867.400000ns, VSS,
+ 1185867.500000ns, VDD,
+ 1186227.700000ns, VDD,
+ 1186227.800000ns, VSS,
+ 1186347.800000ns, VSS,
+ 1186347.900000ns, VDD,
+ 1187789.000000ns, VDD,
+ 1187789.100000ns, VSS,
+ 1188029.200000ns, VSS,
+ 1188029.300000ns, VDD,
+ 1188509.600000ns, VDD,
+ 1188509.700000ns, VSS,
+ 1188749.800000ns, VSS,
+ 1188749.900000ns, VDD,
+ 1188869.900000ns, VDD,
+ 1188870.000000ns, VSS,
+ 1189590.500000ns, VSS,
+ 1189590.600000ns, VDD,
+ 1189830.700000ns, VDD,
+ 1189830.800000ns, VSS,
+ 1189950.800000ns, VSS,
+ 1189950.900000ns, VDD,
+ 1190671.400000ns, VDD,
+ 1190671.500000ns, VSS,
+ 1191031.700000ns, VSS,
+ 1191031.800000ns, VDD,
+ 1191512.100000ns, VDD,
+ 1191512.200000ns, VSS,
+ 1191872.400000ns, VSS,
+ 1191872.500000ns, VDD,
+ 1192232.700000ns, VDD,
+ 1192232.800000ns, VSS,
+ 1192352.800000ns, VSS,
+ 1192352.900000ns, VDD,
+ 1193193.500000ns, VDD,
+ 1193193.600000ns, VSS,
+ 1193313.600000ns, VSS,
+ 1193313.700000ns, VDD,
+ 1193914.100000ns, VDD,
+ 1193914.200000ns, VSS,
+ 1194154.300000ns, VSS,
+ 1194154.400000ns, VDD,
+ 1194394.500000ns, VDD,
+ 1194394.600000ns, VSS,
+ 1194634.700000ns, VSS,
+ 1194634.800000ns, VDD,
+ 1194995.000000ns, VDD,
+ 1194995.100000ns, VSS,
+ 1195235.200000ns, VSS,
+ 1195235.300000ns, VDD,
+ 1196556.300000ns, VDD,
+ 1196556.400000ns, VSS,
+ 1196676.400000ns, VSS,
+ 1196676.500000ns, VDD,
+ 1196916.600000ns, VDD,
+ 1196916.700000ns, VSS,
+ 1197397.000000ns, VSS,
+ 1197397.100000ns, VDD,
+ 1197637.200000ns, VDD,
+ 1197637.300000ns, VSS,
+ 1197757.300000ns, VSS,
+ 1197757.400000ns, VDD,
+ 1198718.100000ns, VDD,
+ 1198718.200000ns, VSS,
+ 1198838.200000ns, VSS,
+ 1198838.300000ns, VDD,
+ 1199318.600000ns, VDD,
+ 1199318.700000ns, VSS,
+ 1199438.700000ns, VSS,
+ 1199438.800000ns, VDD,
+ 1199678.900000ns, VDD,
+ 1199679.000000ns, VSS,
+ 1199919.100000ns, VSS,
+ 1199919.200000ns, VDD,
+ 1200039.200000ns, VDD,
+ 1200039.300000ns, VSS,
+ 1200279.400000ns, VSS,
+ 1200279.500000ns, VDD,
+ 1200639.700000ns, VDD,
+ 1200639.800000ns, VSS,
+ 1201000.000000ns, VSS,
+ 1201000.100000ns, VDD,
+ 1201720.600000ns, VDD,
+ 1201720.700000ns, VSS,
+ 1202201.000000ns, VSS,
+ 1202201.100000ns, VDD,
+ 1203161.800000ns, VDD,
+ 1203161.900000ns, VSS,
+ 1203402.000000ns, VSS,
+ 1203402.100000ns, VDD,
+ 1203642.200000ns, VDD,
+ 1203642.300000ns, VSS,
+ 1203762.300000ns, VSS,
+ 1203762.400000ns, VDD,
+ 1203882.400000ns, VDD,
+ 1203882.500000ns, VSS,
+ 1204122.600000ns, VSS,
+ 1204122.700000ns, VDD,
+ 1204362.800000ns, VDD,
+ 1204362.900000ns, VSS,
+ 1204482.900000ns, VSS,
+ 1204483.000000ns, VDD,
+ 1204843.200000ns, VDD,
+ 1204843.300000ns, VSS,
+ 1204963.300000ns, VSS,
+ 1204963.400000ns, VDD,
+ 1205323.600000ns, VDD,
+ 1205323.700000ns, VSS,
+ 1205443.700000ns, VSS,
+ 1205443.800000ns, VDD,
+ 1206044.200000ns, VDD,
+ 1206044.300000ns, VSS,
+ 1206644.700000ns, VSS,
+ 1206644.800000ns, VDD,
+ 1207125.100000ns, VDD,
+ 1207125.200000ns, VSS,
+ 1207365.300000ns, VSS,
+ 1207365.400000ns, VDD,
+ 1207605.500000ns, VDD,
+ 1207605.600000ns, VSS,
+ 1208326.100000ns, VSS,
+ 1208326.200000ns, VDD,
+ 1208686.400000ns, VDD,
+ 1208686.500000ns, VSS,
+ 1209647.200000ns, VSS,
+ 1209647.300000ns, VDD,
+ 1210247.700000ns, VDD,
+ 1210247.800000ns, VSS,
+ 1210367.800000ns, VSS,
+ 1210367.900000ns, VDD,
+ 1210487.900000ns, VDD,
+ 1210488.000000ns, VSS,
+ 1210608.000000ns, VSS,
+ 1210608.100000ns, VDD,
+ 1210728.100000ns, VDD,
+ 1210728.200000ns, VSS,
+ 1211088.400000ns, VSS,
+ 1211088.500000ns, VDD,
+ 1212169.300000ns, VDD,
+ 1212169.400000ns, VSS,
+ 1212409.500000ns, VSS,
+ 1212409.600000ns, VDD,
+ 1212649.700000ns, VDD,
+ 1212649.800000ns, VSS,
+ 1212769.800000ns, VSS,
+ 1212769.900000ns, VDD,
+ 1212889.900000ns, VDD,
+ 1212890.000000ns, VSS,
+ 1213010.000000ns, VSS,
+ 1213010.100000ns, VDD,
+ 1213730.600000ns, VDD,
+ 1213730.700000ns, VSS,
+ 1213850.700000ns, VSS,
+ 1213850.800000ns, VDD,
+ 1215171.800000ns, VDD,
+ 1215171.900000ns, VSS,
+ 1215291.900000ns, VSS,
+ 1215292.000000ns, VDD,
+ 1215412.000000ns, VDD,
+ 1215412.100000ns, VSS,
+ 1215532.100000ns, VSS,
+ 1215532.200000ns, VDD,
+ 1215892.400000ns, VDD,
+ 1215892.500000ns, VSS,
+ 1216733.100000ns, VSS,
+ 1216733.200000ns, VDD,
+ 1218294.400000ns, VDD,
+ 1218294.500000ns, VSS,
+ 1218414.500000ns, VSS,
+ 1218414.600000ns, VDD,
+ 1219015.000000ns, VDD,
+ 1219015.100000ns, VSS,
+ 1219135.100000ns, VSS,
+ 1219135.200000ns, VDD,
+ 1219255.200000ns, VDD,
+ 1219255.300000ns, VSS,
+ 1219375.300000ns, VSS,
+ 1219375.400000ns, VDD,
+ 1219975.800000ns, VDD,
+ 1219975.900000ns, VSS,
+ 1220095.900000ns, VSS,
+ 1220096.000000ns, VDD,
+ 1220216.000000ns, VDD,
+ 1220216.100000ns, VSS,
+ 1220336.100000ns, VSS,
+ 1220336.200000ns, VDD,
+ 1220816.500000ns, VDD,
+ 1220816.600000ns, VSS,
+ 1221176.800000ns, VSS,
+ 1221176.900000ns, VDD,
+ 1221657.200000ns, VDD,
+ 1221657.300000ns, VSS,
+ 1221897.400000ns, VSS,
+ 1221897.500000ns, VDD,
+ 1222257.700000ns, VDD,
+ 1222257.800000ns, VSS,
+ 1222738.100000ns, VSS,
+ 1222738.200000ns, VDD,
+ 1224059.200000ns, VDD,
+ 1224059.300000ns, VSS,
+ 1224539.600000ns, VSS,
+ 1224539.700000ns, VDD,
+ 1224899.900000ns, VDD,
+ 1224900.000000ns, VSS,
+ 1225140.100000ns, VSS,
+ 1225140.200000ns, VDD,
+ 1225260.200000ns, VDD,
+ 1225260.300000ns, VSS,
+ 1225500.400000ns, VSS,
+ 1225500.500000ns, VDD,
+ 1225860.700000ns, VDD,
+ 1225860.800000ns, VSS,
+ 1226100.900000ns, VSS,
+ 1226101.000000ns, VDD,
+ 1226341.100000ns, VDD,
+ 1226341.200000ns, VSS,
+ 1226581.300000ns, VSS,
+ 1226581.400000ns, VDD,
+ 1226701.400000ns, VDD,
+ 1226701.500000ns, VSS,
+ 1227301.900000ns, VSS,
+ 1227302.000000ns, VDD,
+ 1227542.100000ns, VDD,
+ 1227542.200000ns, VSS,
+ 1228022.500000ns, VSS,
+ 1228022.600000ns, VDD,
+ 1228983.300000ns, VDD,
+ 1228983.400000ns, VSS,
+ 1229463.700000ns, VSS,
+ 1229463.800000ns, VDD,
+ 1231025.000000ns, VDD,
+ 1231025.100000ns, VSS,
+ 1231265.200000ns, VSS,
+ 1231265.300000ns, VDD,
+ 1231385.300000ns, VDD,
+ 1231385.400000ns, VSS,
+ 1232226.000000ns, VSS,
+ 1232226.100000ns, VDD,
+ 1232946.600000ns, VDD,
+ 1232946.700000ns, VSS,
+ 1233306.900000ns, VSS,
+ 1233307.000000ns, VDD,
+ 1233787.300000ns, VDD,
+ 1233787.400000ns, VSS,
+ 1234027.500000ns, VSS,
+ 1234027.600000ns, VDD,
+ 1234387.800000ns, VDD,
+ 1234387.900000ns, VSS,
+ 1234868.200000ns, VSS,
+ 1234868.300000ns, VDD,
+ 1235228.500000ns, VDD,
+ 1235228.600000ns, VSS,
+ 1236549.600000ns, VSS,
+ 1236549.700000ns, VDD,
+ 1236789.800000ns, VDD,
+ 1236789.900000ns, VSS,
+ 1237390.300000ns, VSS,
+ 1237390.400000ns, VDD,
+ 1237750.600000ns, VDD,
+ 1237750.700000ns, VSS,
+ 1238231.000000ns, VSS,
+ 1238231.100000ns, VDD,
+ 1239071.700000ns, VDD,
+ 1239071.800000ns, VSS,
+ 1239191.800000ns, VSS,
+ 1239191.900000ns, VDD,
+ 1239792.300000ns, VDD,
+ 1239792.400000ns, VSS,
+ 1240272.700000ns, VSS,
+ 1240272.800000ns, VDD,
+ 1241233.500000ns, VDD,
+ 1241233.600000ns, VSS,
+ 1241353.600000ns, VSS,
+ 1241353.700000ns, VDD,
+ 1241593.800000ns, VDD,
+ 1241593.900000ns, VSS,
+ 1242314.400000ns, VSS,
+ 1242314.500000ns, VDD,
+ 1242434.500000ns, VDD,
+ 1242434.600000ns, VSS,
+ 1242794.800000ns, VSS,
+ 1242794.900000ns, VDD,
+ 1243035.000000ns, VDD,
+ 1243035.100000ns, VSS,
+ 1243515.400000ns, VSS,
+ 1243515.500000ns, VDD,
+ 1243755.600000ns, VDD,
+ 1243755.700000ns, VSS,
+ 1244356.100000ns, VSS,
+ 1244356.200000ns, VDD,
+ 1244476.200000ns, VDD,
+ 1244476.300000ns, VSS,
+ 1244956.600000ns, VSS,
+ 1244956.700000ns, VDD,
+ 1245076.700000ns, VDD,
+ 1245076.800000ns, VSS,
+ 1245196.800000ns, VSS,
+ 1245196.900000ns, VDD,
+ 1245557.100000ns, VDD,
+ 1245557.200000ns, VSS,
+ 1245677.200000ns, VSS,
+ 1245677.300000ns, VDD,
+ 1246277.700000ns, VDD,
+ 1246277.800000ns, VSS,
+ 1246758.100000ns, VSS,
+ 1246758.200000ns, VDD,
+ 1247358.600000ns, VDD,
+ 1247358.700000ns, VSS,
+ 1247598.800000ns, VSS,
+ 1247598.900000ns, VDD,
+ 1247718.900000ns, VDD,
+ 1247719.000000ns, VSS,
+ 1247839.000000ns, VSS,
+ 1247839.100000ns, VDD,
+ 1248079.200000ns, VDD,
+ 1248079.300000ns, VSS,
+ 1248679.700000ns, VSS,
+ 1248679.800000ns, VDD,
+ 1249160.100000ns, VDD,
+ 1249160.200000ns, VSS,
+ 1249400.300000ns, VSS,
+ 1249400.400000ns, VDD,
+ 1249640.500000ns, VDD,
+ 1249640.600000ns, VSS,
+ 1249760.600000ns, VSS,
+ 1249760.700000ns, VDD,
+ 1249880.700000ns, VDD,
+ 1249880.800000ns, VSS,
+ 1250120.900000ns, VSS,
+ 1250121.000000ns, VDD,
+ 1250361.100000ns, VDD,
+ 1250361.200000ns, VSS,
+ 1250721.400000ns, VSS,
+ 1250721.500000ns, VDD,
+ 1251922.400000ns, VDD,
+ 1251922.500000ns, VSS,
+ 1252162.600000ns, VSS,
+ 1252162.700000ns, VDD,
+ 1252282.700000ns, VDD,
+ 1252282.800000ns, VSS,
+ 1252763.100000ns, VSS,
+ 1252763.200000ns, VDD,
+ 1253363.600000ns, VDD,
+ 1253363.700000ns, VSS,
+ 1253844.000000ns, VSS,
+ 1253844.100000ns, VDD,
+ 1254204.300000ns, VDD,
+ 1254204.400000ns, VSS,
+ 1254444.500000ns, VSS,
+ 1254444.600000ns, VDD,
+ 1254804.800000ns, VDD,
+ 1254804.900000ns, VSS,
+ 1254924.900000ns, VSS,
+ 1254925.000000ns, VDD,
+ 1255765.600000ns, VDD,
+ 1255765.700000ns, VSS,
+ 1255885.700000ns, VSS,
+ 1255885.800000ns, VDD,
+ 1256125.900000ns, VDD,
+ 1256126.000000ns, VSS,
+ 1256366.100000ns, VSS,
+ 1256366.200000ns, VDD,
+ 1256726.400000ns, VDD,
+ 1256726.500000ns, VSS,
+ 1256846.500000ns, VSS,
+ 1256846.600000ns, VDD,
+ 1257086.700000ns, VDD,
+ 1257086.800000ns, VSS,
+ 1257447.000000ns, VSS,
+ 1257447.100000ns, VDD,
+ 1257927.400000ns, VDD,
+ 1257927.500000ns, VSS,
+ 1258167.600000ns, VSS,
+ 1258167.700000ns, VDD,
+ 1258287.700000ns, VDD,
+ 1258287.800000ns, VSS,
+ 1258648.000000ns, VSS,
+ 1258648.100000ns, VDD,
+ 1258888.200000ns, VDD,
+ 1258888.300000ns, VSS,
+ 1259128.400000ns, VSS,
+ 1259128.500000ns, VDD,
+ 1259608.800000ns, VDD,
+ 1259608.900000ns, VSS,
+ 1259969.100000ns, VSS,
+ 1259969.200000ns, VDD,
+ 1260089.200000ns, VDD,
+ 1260089.300000ns, VSS,
+ 1260209.300000ns, VSS,
+ 1260209.400000ns, VDD,
+ 1260329.400000ns, VDD,
+ 1260329.500000ns, VSS,
+ 1261170.100000ns, VSS,
+ 1261170.200000ns, VDD,
+ 1261410.300000ns, VDD,
+ 1261410.400000ns, VSS,
+ 1262251.000000ns, VSS,
+ 1262251.100000ns, VDD,
+ 1262731.400000ns, VDD,
+ 1262731.500000ns, VSS,
+ 1262971.600000ns, VSS,
+ 1262971.700000ns, VDD,
+ 1263452.000000ns, VDD,
+ 1263452.100000ns, VSS,
+ 1263572.100000ns, VSS,
+ 1263572.200000ns, VDD,
+ 1263692.200000ns, VDD,
+ 1263692.300000ns, VSS,
+ 1265133.400000ns, VSS,
+ 1265133.500000ns, VDD,
+ 1265373.600000ns, VDD,
+ 1265373.700000ns, VSS,
+ 1265493.700000ns, VSS,
+ 1265493.800000ns, VDD,
+ 1265974.100000ns, VDD,
+ 1265974.200000ns, VSS,
+ 1266214.300000ns, VSS,
+ 1266214.400000ns, VDD,
+ 1266574.600000ns, VDD,
+ 1266574.700000ns, VSS,
+ 1267655.500000ns, VSS,
+ 1267655.600000ns, VDD,
+ 1268135.900000ns, VDD,
+ 1268136.000000ns, VSS,
+ 1268496.200000ns, VSS,
+ 1268496.300000ns, VDD,
+ 1268616.300000ns, VDD,
+ 1268616.400000ns, VSS,
+ 1268736.400000ns, VSS,
+ 1268736.500000ns, VDD,
+ 1269457.000000ns, VDD,
+ 1269457.100000ns, VSS,
+ 1269817.300000ns, VSS,
+ 1269817.400000ns, VDD,
+ 1270297.700000ns, VDD,
+ 1270297.800000ns, VSS,
+ 1270417.800000ns, VSS,
+ 1270417.900000ns, VDD,
+ 1270658.000000ns, VDD,
+ 1270658.100000ns, VSS,
+ 1271138.400000ns, VSS,
+ 1271138.500000ns, VDD,
+ 1272819.800000ns, VDD,
+ 1272819.900000ns, VSS,
+ 1274381.100000ns, VSS,
+ 1274381.200000ns, VDD,
+ 1274861.500000ns, VDD,
+ 1274861.600000ns, VSS,
+ 1275582.100000ns, VSS,
+ 1275582.200000ns, VDD,
+ 1275822.300000ns, VDD,
+ 1275822.400000ns, VSS,
+ 1276062.500000ns, VSS,
+ 1276062.600000ns, VDD,
+ 1277503.700000ns, VDD,
+ 1277503.800000ns, VSS,
+ 1277743.900000ns, VSS,
+ 1277744.000000ns, VDD,
+ 1278104.200000ns, VDD,
+ 1278104.300000ns, VSS,
+ 1278704.700000ns, VSS,
+ 1278704.800000ns, VDD,
+ 1279305.200000ns, VDD,
+ 1279305.300000ns, VSS,
+ 1279545.400000ns, VSS,
+ 1279545.500000ns, VDD,
+ 1280506.200000ns, VDD,
+ 1280506.300000ns, VSS,
+ 1281106.700000ns, VSS,
+ 1281106.800000ns, VDD,
+ 1281587.100000ns, VDD,
+ 1281587.200000ns, VSS,
+ 1281707.200000ns, VSS,
+ 1281707.300000ns, VDD,
+ 1282187.600000ns, VDD,
+ 1282187.700000ns, VSS,
+ 1282547.900000ns, VSS,
+ 1282548.000000ns, VDD,
+ 1283989.100000ns, VDD,
+ 1283989.200000ns, VSS,
+ 1284109.200000ns, VSS,
+ 1284109.300000ns, VDD,
+ 1284469.500000ns, VDD,
+ 1284469.600000ns, VSS,
+ 1284829.800000ns, VSS,
+ 1284829.900000ns, VDD,
+ 1284949.900000ns, VDD,
+ 1284950.000000ns, VSS,
+ 1285670.500000ns, VSS,
+ 1285670.600000ns, VDD,
+ 1285790.600000ns, VDD,
+ 1285790.700000ns, VSS,
+ 1285910.700000ns, VSS,
+ 1285910.800000ns, VDD,
+ 1286271.000000ns, VDD,
+ 1286271.100000ns, VSS,
+ 1286631.300000ns, VSS,
+ 1286631.400000ns, VDD,
+ 1286871.500000ns, VDD,
+ 1286871.600000ns, VSS,
+ 1287111.700000ns, VSS,
+ 1287111.800000ns, VDD,
+ 1287592.100000ns, VDD,
+ 1287592.200000ns, VSS,
+ 1287712.200000ns, VSS,
+ 1287712.300000ns, VDD,
+ 1289393.600000ns, VDD,
+ 1289393.700000ns, VSS,
+ 1289513.700000ns, VSS,
+ 1289513.800000ns, VDD,
+ 1289994.100000ns, VDD,
+ 1289994.200000ns, VSS,
+ 1290354.400000ns, VSS,
+ 1290354.500000ns, VDD,
+ 1291075.000000ns, VDD,
+ 1291075.100000ns, VSS,
+ 1291315.200000ns, VSS,
+ 1291315.300000ns, VDD,
+ 1291795.600000ns, VDD,
+ 1291795.700000ns, VSS,
+ 1292276.000000ns, VSS,
+ 1292276.100000ns, VDD,
+ 1293116.700000ns, VDD,
+ 1293116.800000ns, VSS,
+ 1293236.800000ns, VSS,
+ 1293236.900000ns, VDD,
+ 1293356.900000ns, VDD,
+ 1293357.000000ns, VSS,
+ 1293477.000000ns, VSS,
+ 1293477.100000ns, VDD,
+ 1293837.300000ns, VDD,
+ 1293837.400000ns, VSS,
+ 1293957.400000ns, VSS,
+ 1293957.500000ns, VDD,
+ 1294317.700000ns, VDD,
+ 1294317.800000ns, VSS,
+ 1294678.000000ns, VSS,
+ 1294678.100000ns, VDD,
+ 1295278.500000ns, VDD,
+ 1295278.600000ns, VSS,
+ 1295879.000000ns, VSS,
+ 1295879.100000ns, VDD,
+ 1296959.900000ns, VDD,
+ 1296960.000000ns, VSS,
+ 1297080.000000ns, VSS,
+ 1297080.100000ns, VDD,
+ 1297200.100000ns, VDD,
+ 1297200.200000ns, VSS,
+ 1298040.800000ns, VSS,
+ 1298040.900000ns, VDD,
+ 1298641.300000ns, VDD,
+ 1298641.400000ns, VSS,
+ 1299241.800000ns, VSS,
+ 1299241.900000ns, VDD,
+ 1299722.200000ns, VDD,
+ 1299722.300000ns, VSS,
+ 1299962.400000ns, VSS,
+ 1299962.500000ns, VDD,
+ 1300082.500000ns, VDD,
+ 1300082.600000ns, VSS,
+ 1301043.300000ns, VSS,
+ 1301043.400000ns, VDD,
+ 1301283.500000ns, VDD,
+ 1301283.600000ns, VSS,
+ 1301403.600000ns, VSS,
+ 1301403.700000ns, VDD,
+ 1301523.700000ns, VDD,
+ 1301523.800000ns, VSS,
+ 1302364.400000ns, VSS,
+ 1302364.500000ns, VDD,
+ 1302484.500000ns, VDD,
+ 1302484.600000ns, VSS,
+ 1303085.000000ns, VSS,
+ 1303085.100000ns, VDD,
+ 1303565.400000ns, VDD,
+ 1303565.500000ns, VSS,
+ 1303805.600000ns, VSS,
+ 1303805.700000ns, VDD,
+ 1304045.800000ns, VDD,
+ 1304045.900000ns, VSS,
+ 1304406.100000ns, VSS,
+ 1304406.200000ns, VDD,
+ 1305006.600000ns, VDD,
+ 1305006.700000ns, VSS,
+ 1305727.200000ns, VSS,
+ 1305727.300000ns, VDD,
+ 1306087.500000ns, VDD,
+ 1306087.600000ns, VSS,
+ 1306567.900000ns, VSS,
+ 1306568.000000ns, VDD,
+ 1307168.400000ns, VDD,
+ 1307168.500000ns, VSS,
+ 1307408.600000ns, VSS,
+ 1307408.700000ns, VDD,
+ 1307528.700000ns, VDD,
+ 1307528.800000ns, VSS,
+ 1307648.800000ns, VSS,
+ 1307648.900000ns, VDD,
+ 1308969.900000ns, VDD,
+ 1308970.000000ns, VSS,
+ 1309090.000000ns, VSS,
+ 1309090.100000ns, VDD,
+ 1309570.400000ns, VDD,
+ 1309570.500000ns, VSS,
+ 1310411.100000ns, VSS,
+ 1310411.200000ns, VDD,
+ 1311131.700000ns, VDD,
+ 1311131.800000ns, VSS,
+ 1311732.200000ns, VSS,
+ 1311732.300000ns, VDD,
+ 1311852.300000ns, VDD,
+ 1311852.400000ns, VSS,
+ 1312452.800000ns, VSS,
+ 1312452.900000ns, VDD,
+ 1312572.900000ns, VDD,
+ 1312573.000000ns, VSS,
+ 1312813.100000ns, VSS,
+ 1312813.200000ns, VDD,
+ 1313173.400000ns, VDD,
+ 1313173.500000ns, VSS,
+ 1313653.800000ns, VSS,
+ 1313653.900000ns, VDD,
+ 1314854.800000ns, VDD,
+ 1314854.900000ns, VSS,
+ 1315935.700000ns, VSS,
+ 1315935.800000ns, VDD,
+ 1316296.000000ns, VDD,
+ 1316296.100000ns, VSS,
+ 1316416.100000ns, VSS,
+ 1316416.200000ns, VDD,
+ 1316776.400000ns, VDD,
+ 1316776.500000ns, VSS,
+ 1317016.600000ns, VSS,
+ 1317016.700000ns, VDD,
+ 1317136.700000ns, VDD,
+ 1317136.800000ns, VSS,
+ 1317497.000000ns, VSS,
+ 1317497.100000ns, VDD,
+ 1317737.200000ns, VDD,
+ 1317737.300000ns, VSS,
+ 1317857.300000ns, VSS,
+ 1317857.400000ns, VDD,
+ 1317977.400000ns, VDD,
+ 1317977.500000ns, VSS,
+ 1318457.800000ns, VSS,
+ 1318457.900000ns, VDD,
+ 1318698.000000ns, VDD,
+ 1318698.100000ns, VSS,
+ 1319058.300000ns, VSS,
+ 1319058.400000ns, VDD,
+ 1319298.500000ns, VDD,
+ 1319298.600000ns, VSS,
+ 1320019.100000ns, VSS,
+ 1320019.200000ns, VDD,
+ 1320259.300000ns, VDD,
+ 1320259.400000ns, VSS,
+ 1320379.400000ns, VSS,
+ 1320379.500000ns, VDD,
+ 1320499.500000ns, VDD,
+ 1320499.600000ns, VSS,
+ 1320619.600000ns, VSS,
+ 1320619.700000ns, VDD,
+ 1321220.100000ns, VDD,
+ 1321220.200000ns, VSS,
+ 1321580.400000ns, VSS,
+ 1321580.500000ns, VDD,
+ 1322060.800000ns, VDD,
+ 1322060.900000ns, VSS,
+ 1322541.200000ns, VSS,
+ 1322541.300000ns, VDD,
+ 1322901.500000ns, VDD,
+ 1322901.600000ns, VSS,
+ 1323021.600000ns, VSS,
+ 1323021.700000ns, VDD,
+ 1323622.100000ns, VDD,
+ 1323622.200000ns, VSS,
+ 1324102.500000ns, VSS,
+ 1324102.600000ns, VDD,
+ 1324703.000000ns, VDD,
+ 1324703.100000ns, VSS,
+ 1324823.100000ns, VSS,
+ 1324823.200000ns, VDD,
+ 1325183.400000ns, VDD,
+ 1325183.500000ns, VSS,
+ 1325423.600000ns, VSS,
+ 1325423.700000ns, VDD,
+ 1325543.700000ns, VDD,
+ 1325543.800000ns, VSS,
+ 1326984.900000ns, VSS,
+ 1326985.000000ns, VDD,
+ 1327465.300000ns, VDD,
+ 1327465.400000ns, VSS,
+ 1327825.600000ns, VSS,
+ 1327825.700000ns, VDD,
+ 1328185.900000ns, VDD,
+ 1328186.000000ns, VSS,
+ 1329026.600000ns, VSS,
+ 1329026.700000ns, VDD,
+ 1329507.000000ns, VDD,
+ 1329507.100000ns, VSS,
+ 1329747.200000ns, VSS,
+ 1329747.300000ns, VDD,
+ 1329867.300000ns, VDD,
+ 1329867.400000ns, VSS,
+ 1330708.000000ns, VSS,
+ 1330708.100000ns, VDD,
+ 1330948.200000ns, VDD,
+ 1330948.300000ns, VSS,
+ 1331668.800000ns, VSS,
+ 1331668.900000ns, VDD,
+ 1332029.100000ns, VDD,
+ 1332029.200000ns, VSS,
+ 1332149.200000ns, VSS,
+ 1332149.300000ns, VDD,
+ 1332269.300000ns, VDD,
+ 1332269.400000ns, VSS,
+ 1333710.500000ns, VSS,
+ 1333710.600000ns, VDD,
+ 1334070.800000ns, VDD,
+ 1334070.900000ns, VSS,
+ 1334190.900000ns, VSS,
+ 1334191.000000ns, VDD,
+ 1335031.600000ns, VDD,
+ 1335031.700000ns, VSS,
+ 1335271.800000ns, VSS,
+ 1335271.900000ns, VDD,
+ 1335632.100000ns, VDD,
+ 1335632.200000ns, VSS,
+ 1335872.300000ns, VSS,
+ 1335872.400000ns, VDD,
+ 1336472.800000ns, VDD,
+ 1336472.900000ns, VSS,
+ 1336713.000000ns, VSS,
+ 1336713.100000ns, VDD,
+ 1336833.100000ns, VDD,
+ 1336833.200000ns, VSS,
+ 1337793.900000ns, VSS,
+ 1337794.000000ns, VDD,
+ 1338154.200000ns, VDD,
+ 1338154.300000ns, VSS,
+ 1338394.400000ns, VSS,
+ 1338394.500000ns, VDD,
+ 1338754.700000ns, VDD,
+ 1338754.800000ns, VSS,
+ 1339115.000000ns, VSS,
+ 1339115.100000ns, VDD,
+ 1339835.600000ns, VDD,
+ 1339835.700000ns, VSS,
+ 1339955.700000ns, VSS,
+ 1339955.800000ns, VDD,
+ 1340916.500000ns, VDD,
+ 1340916.600000ns, VSS,
+ 1341517.000000ns, VSS,
+ 1341517.100000ns, VDD,
+ 1341637.100000ns, VDD,
+ 1341637.200000ns, VSS,
+ 1341997.400000ns, VSS,
+ 1341997.500000ns, VDD,
+ 1342958.200000ns, VDD,
+ 1342958.300000ns, VSS,
+ 1343558.700000ns, VSS,
+ 1343558.800000ns, VDD,
+ 1343919.000000ns, VDD,
+ 1343919.100000ns, VSS,
+ 1344279.300000ns, VSS,
+ 1344279.400000ns, VDD,
+ 1344639.600000ns, VDD,
+ 1344639.700000ns, VSS,
+ 1344759.700000ns, VSS,
+ 1344759.800000ns, VDD,
+ 1344879.800000ns, VDD,
+ 1344879.900000ns, VSS,
+ 1345120.000000ns, VSS,
+ 1345120.100000ns, VDD,
+ 1345240.100000ns, VDD,
+ 1345240.200000ns, VSS,
+ 1345840.600000ns, VSS,
+ 1345840.700000ns, VDD,
+ 1346321.000000ns, VDD,
+ 1346321.100000ns, VSS,
+ 1346561.200000ns, VSS,
+ 1346561.300000ns, VDD,
+ 1347041.600000ns, VDD,
+ 1347041.700000ns, VSS,
+ 1347161.700000ns, VSS,
+ 1347161.800000ns, VDD,
+ 1347642.100000ns, VDD,
+ 1347642.200000ns, VSS,
+ 1348002.400000ns, VSS,
+ 1348002.500000ns, VDD,
+ 1348723.000000ns, VDD,
+ 1348723.100000ns, VSS,
+ 1349083.300000ns, VSS,
+ 1349083.400000ns, VDD,
+ 1349683.800000ns, VDD,
+ 1349683.900000ns, VSS,
+ 1350164.200000ns, VSS,
+ 1350164.300000ns, VDD,
+ 1350284.300000ns, VDD,
+ 1350284.400000ns, VSS,
+ 1350524.500000ns, VSS,
+ 1350524.600000ns, VDD,
+ 1350764.700000ns, VDD,
+ 1350764.800000ns, VSS,
+ 1351004.900000ns, VSS,
+ 1351005.000000ns, VDD,
+ 1351605.400000ns, VDD,
+ 1351605.500000ns, VSS,
+ 1351725.500000ns, VSS,
+ 1351725.600000ns, VDD,
+ 1351965.700000ns, VDD,
+ 1351965.800000ns, VSS,
+ 1352085.800000ns, VSS,
+ 1352085.900000ns, VDD,
+ 1352686.300000ns, VDD,
+ 1352686.400000ns, VSS,
+ 1352806.400000ns, VSS,
+ 1352806.500000ns, VDD,
+ 1353166.700000ns, VDD,
+ 1353166.800000ns, VSS,
+ 1353406.900000ns, VSS,
+ 1353407.000000ns, VDD,
+ 1353767.200000ns, VDD,
+ 1353767.300000ns, VSS,
+ 1354127.500000ns, VSS,
+ 1354127.600000ns, VDD,
+ 1354247.600000ns, VDD,
+ 1354247.700000ns, VSS,
+ 1354367.700000ns, VSS,
+ 1354367.800000ns, VDD,
+ 1355088.300000ns, VDD,
+ 1355088.400000ns, VSS,
+ 1355448.600000ns, VSS,
+ 1355448.700000ns, VDD,
+ 1355929.000000ns, VDD,
+ 1355929.100000ns, VSS,
+ 1356289.300000ns, VSS,
+ 1356289.400000ns, VDD,
+ 1356529.500000ns, VDD,
+ 1356529.600000ns, VSS,
+ 1357490.300000ns, VSS,
+ 1357490.400000ns, VDD,
+ 1357970.700000ns, VDD,
+ 1357970.800000ns, VSS,
+ 1358451.100000ns, VSS,
+ 1358451.200000ns, VDD,
+ 1358571.200000ns, VDD,
+ 1358571.300000ns, VSS,
+ 1359051.600000ns, VSS,
+ 1359051.700000ns, VDD,
+ 1360252.600000ns, VDD,
+ 1360252.700000ns, VSS,
+ 1360733.000000ns, VSS,
+ 1360733.100000ns, VDD,
+ 1360853.100000ns, VDD,
+ 1360853.200000ns, VSS,
+ 1361213.400000ns, VSS,
+ 1361213.500000ns, VDD,
+ 1362054.100000ns, VDD,
+ 1362054.200000ns, VSS,
+ 1362174.200000ns, VSS,
+ 1362174.300000ns, VDD,
+ 1362534.500000ns, VDD,
+ 1362534.600000ns, VSS,
+ 1362654.600000ns, VSS,
+ 1362654.700000ns, VDD,
+ 1362894.800000ns, VDD,
+ 1362894.900000ns, VSS,
+ 1363135.000000ns, VSS,
+ 1363135.100000ns, VDD,
+ 1363255.100000ns, VDD,
+ 1363255.200000ns, VSS,
+ 1363495.300000ns, VSS,
+ 1363495.400000ns, VDD,
+ 1363975.700000ns, VDD,
+ 1363975.800000ns, VSS,
+ 1365176.700000ns, VSS,
+ 1365176.800000ns, VDD,
+ 1365537.000000ns, VDD,
+ 1365537.100000ns, VSS,
+ 1365777.200000ns, VSS,
+ 1365777.300000ns, VDD,
+ 1365897.300000ns, VDD,
+ 1365897.400000ns, VSS,
+ 1366137.500000ns, VSS,
+ 1366137.600000ns, VDD,
+ 1366257.600000ns, VDD,
+ 1366257.700000ns, VSS,
+ 1366978.200000ns, VSS,
+ 1366978.300000ns, VDD,
+ 1367218.400000ns, VDD,
+ 1367218.500000ns, VSS,
+ 1367939.000000ns, VSS,
+ 1367939.100000ns, VDD,
+ 1368179.200000ns, VDD,
+ 1368179.300000ns, VSS,
+ 1368299.300000ns, VSS,
+ 1368299.400000ns, VDD,
+ 1368659.600000ns, VDD,
+ 1368659.700000ns, VSS,
+ 1369140.000000ns, VSS,
+ 1369140.100000ns, VDD,
+ 1369500.300000ns, VDD,
+ 1369500.400000ns, VSS,
+ 1369620.400000ns, VSS,
+ 1369620.500000ns, VDD,
+ 1369980.700000ns, VDD,
+ 1369980.800000ns, VSS,
+ 1370220.900000ns, VSS,
+ 1370221.000000ns, VDD,
+ 1370581.200000ns, VDD,
+ 1370581.300000ns, VSS,
+ 1371061.600000ns, VSS,
+ 1371061.700000ns, VDD,
+ 1371421.900000ns, VDD,
+ 1371422.000000ns, VSS,
+ 1371662.100000ns, VSS,
+ 1371662.200000ns, VDD,
+ 1372022.400000ns, VDD,
+ 1372022.500000ns, VSS,
+ 1372142.500000ns, VSS,
+ 1372142.600000ns, VDD,
+ 1372262.600000ns, VDD,
+ 1372262.700000ns, VSS,
+ 1372622.900000ns, VSS,
+ 1372623.000000ns, VDD,
+ 1373103.300000ns, VDD,
+ 1373103.400000ns, VSS,
+ 1373343.500000ns, VSS,
+ 1373343.600000ns, VDD,
+ 1373463.600000ns, VDD,
+ 1373463.700000ns, VSS,
+ 1373823.900000ns, VSS,
+ 1373824.000000ns, VDD,
+ 1374184.200000ns, VDD,
+ 1374184.300000ns, VSS,
+ 1374544.500000ns, VSS,
+ 1374544.600000ns, VDD,
+ 1374904.800000ns, VDD,
+ 1374904.900000ns, VSS,
+ 1375024.900000ns, VSS,
+ 1375025.000000ns, VDD,
+ 1375265.100000ns, VDD,
+ 1375265.200000ns, VSS,
+ 1375385.200000ns, VSS,
+ 1375385.300000ns, VDD,
+ 1375865.600000ns, VDD,
+ 1375865.700000ns, VSS,
+ 1376346.000000ns, VSS,
+ 1376346.100000ns, VDD,
+ 1376946.500000ns, VDD,
+ 1376946.600000ns, VSS,
+ 1377066.600000ns, VSS,
+ 1377066.700000ns, VDD,
+ 1377547.000000ns, VDD,
+ 1377547.100000ns, VSS,
+ 1377667.100000ns, VSS,
+ 1377667.200000ns, VDD,
+ 1378627.900000ns, VDD,
+ 1378628.000000ns, VSS,
+ 1378748.000000ns, VSS,
+ 1378748.100000ns, VDD,
+ 1379108.300000ns, VDD,
+ 1379108.400000ns, VSS,
+ 1379228.400000ns, VSS,
+ 1379228.500000ns, VDD,
+ 1379468.600000ns, VDD,
+ 1379468.700000ns, VSS,
+ 1379588.700000ns, VSS,
+ 1379588.800000ns, VDD,
+ 1379708.800000ns, VDD,
+ 1379708.900000ns, VSS,
+ 1379828.900000ns, VSS,
+ 1379829.000000ns, VDD,
+ 1380189.200000ns, VDD,
+ 1380189.300000ns, VSS,
+ 1380309.300000ns, VSS,
+ 1380309.400000ns, VDD,
+ 1380429.400000ns, VDD,
+ 1380429.500000ns, VSS,
+ 1381270.100000ns, VSS,
+ 1381270.200000ns, VDD,
+ 1381870.600000ns, VDD,
+ 1381870.700000ns, VSS,
+ 1382351.000000ns, VSS,
+ 1382351.100000ns, VDD,
+ 1383191.700000ns, VDD,
+ 1383191.800000ns, VSS,
+ 1383431.900000ns, VSS,
+ 1383432.000000ns, VDD,
+ 1383672.100000ns, VDD,
+ 1383672.200000ns, VSS,
+ 1384152.500000ns, VSS,
+ 1384152.600000ns, VDD,
+ 1384392.700000ns, VDD,
+ 1384392.800000ns, VSS,
+ 1384632.900000ns, VSS,
+ 1384633.000000ns, VDD,
+ 1384753.000000ns, VDD,
+ 1384753.100000ns, VSS,
+ 1384873.100000ns, VSS,
+ 1384873.200000ns, VDD,
+ 1385233.400000ns, VDD,
+ 1385233.500000ns, VSS,
+ 1385713.800000ns, VSS,
+ 1385713.900000ns, VDD,
+ 1386554.500000ns, VDD,
+ 1386554.600000ns, VSS,
+ 1386794.700000ns, VSS,
+ 1386794.800000ns, VDD,
+ 1386914.800000ns, VDD,
+ 1386914.900000ns, VSS,
+ 1387155.000000ns, VSS,
+ 1387155.100000ns, VDD,
+ 1387515.300000ns, VDD,
+ 1387515.400000ns, VSS,
+ 1387755.500000ns, VSS,
+ 1387755.600000ns, VDD,
+ 1387995.700000ns, VDD,
+ 1387995.800000ns, VSS,
+ 1388235.900000ns, VSS,
+ 1388236.000000ns, VDD,
+ 1388716.300000ns, VDD,
+ 1388716.400000ns, VSS,
+ 1389196.700000ns, VSS,
+ 1389196.800000ns, VDD,
+ 1389316.800000ns, VDD,
+ 1389316.900000ns, VSS,
+ 1389797.200000ns, VSS,
+ 1389797.300000ns, VDD,
+ 1390157.500000ns, VDD,
+ 1390157.600000ns, VSS,
+ 1390277.600000ns, VSS,
+ 1390277.700000ns, VDD,
+ 1390758.000000ns, VDD,
+ 1390758.100000ns, VSS,
+ 1390878.100000ns, VSS,
+ 1390878.200000ns, VDD,
+ 1390998.200000ns, VDD,
+ 1390998.300000ns, VSS,
+ 1391478.600000ns, VSS,
+ 1391478.700000ns, VDD,
+ 1391959.000000ns, VDD,
+ 1391959.100000ns, VSS,
+ 1392079.100000ns, VSS,
+ 1392079.200000ns, VDD,
+ 1392559.500000ns, VDD,
+ 1392559.600000ns, VSS,
+ 1392919.800000ns, VSS,
+ 1392919.900000ns, VDD,
+ 1393400.200000ns, VDD,
+ 1393400.300000ns, VSS,
+ 1393640.400000ns, VSS,
+ 1393640.500000ns, VDD,
+ 1393880.600000ns, VDD,
+ 1393880.700000ns, VSS,
+ 1394240.900000ns, VSS,
+ 1394241.000000ns, VDD,
+ 1394361.000000ns, VDD,
+ 1394361.100000ns, VSS,
+ 1394481.100000ns, VSS,
+ 1394481.200000ns, VDD,
+ 1394841.400000ns, VDD,
+ 1394841.500000ns, VSS,
+ 1395081.600000ns, VSS,
+ 1395081.700000ns, VDD,
+ 1395562.000000ns, VDD,
+ 1395562.100000ns, VSS,
+ 1395922.300000ns, VSS,
+ 1395922.400000ns, VDD,
+ 1396282.600000ns, VDD,
+ 1396282.700000ns, VSS,
+ 1396402.700000ns, VSS,
+ 1396402.800000ns, VDD,
+ 1397003.200000ns, VDD,
+ 1397003.300000ns, VSS,
+ 1397123.300000ns, VSS,
+ 1397123.400000ns, VDD,
+ 1397483.600000ns, VDD,
+ 1397483.700000ns, VSS,
+ 1399165.000000ns, VSS,
+ 1399165.100000ns, VDD,
+ 1399405.200000ns, VDD,
+ 1399405.300000ns, VSS,
+ 1399885.600000ns, VSS,
+ 1399885.700000ns, VDD,
+ 1400245.900000ns, VDD,
+ 1400246.000000ns, VSS,
+ 1400486.100000ns, VSS,
+ 1400486.200000ns, VDD,
+ 1400846.400000ns, VDD,
+ 1400846.500000ns, VSS,
+ 1401206.700000ns, VSS,
+ 1401206.800000ns, VDD,
+ 1401446.900000ns, VDD,
+ 1401447.000000ns, VSS,
+ 1401567.000000ns, VSS,
+ 1401567.100000ns, VDD,
+ 1402047.400000ns, VDD,
+ 1402047.500000ns, VSS,
+ 1402167.500000ns, VSS,
+ 1402167.600000ns, VDD,
+ 1402527.800000ns, VDD,
+ 1402527.900000ns, VSS,
+ 1402768.000000ns, VSS,
+ 1402768.100000ns, VDD,
+ 1403248.400000ns, VDD,
+ 1403248.500000ns, VSS,
+ 1403368.500000ns, VSS,
+ 1403368.600000ns, VDD,
+ 1405410.200000ns, VDD,
+ 1405410.300000ns, VSS,
+ 1405650.400000ns, VSS,
+ 1405650.500000ns, VDD,
+ 1405890.600000ns, VDD,
+ 1405890.700000ns, VSS,
+ 1406250.900000ns, VSS,
+ 1406251.000000ns, VDD,
+ 1406611.200000ns, VDD,
+ 1406611.300000ns, VSS,
+ 1406731.300000ns, VSS,
+ 1406731.400000ns, VDD,
+ 1407091.600000ns, VDD,
+ 1407091.700000ns, VSS,
+ 1407451.900000ns, VSS,
+ 1407452.000000ns, VDD,
+ 1407692.100000ns, VDD,
+ 1407692.200000ns, VSS,
+ 1408172.500000ns, VSS,
+ 1408172.600000ns, VDD,
+ 1408412.700000ns, VDD,
+ 1408412.800000ns, VSS,
+ 1408893.100000ns, VSS,
+ 1408893.200000ns, VDD,
+ 1409373.500000ns, VDD,
+ 1409373.600000ns, VSS,
+ 1409493.600000ns, VSS,
+ 1409493.700000ns, VDD,
+ 1409613.700000ns, VDD,
+ 1409613.800000ns, VSS,
+ 1409733.800000ns, VSS,
+ 1409733.900000ns, VDD,
+ 1410214.200000ns, VDD,
+ 1410214.300000ns, VSS,
+ 1410334.300000ns, VSS,
+ 1410334.400000ns, VDD,
+ 1412616.200000ns, VDD,
+ 1412616.300000ns, VSS,
+ 1412976.500000ns, VSS,
+ 1412976.600000ns, VDD,
+ 1413697.100000ns, VDD,
+ 1413697.200000ns, VSS,
+ 1414057.400000ns, VSS,
+ 1414057.500000ns, VDD,
+ 1414177.500000ns, VDD,
+ 1414177.600000ns, VSS,
+ 1414537.800000ns, VSS,
+ 1414537.900000ns, VDD,
+ 1414657.900000ns, VDD,
+ 1414658.000000ns, VSS,
+ 1415018.200000ns, VSS,
+ 1415018.300000ns, VDD,
+ 1415378.500000ns, VDD,
+ 1415378.600000ns, VSS,
+ 1416219.200000ns, VSS,
+ 1416219.300000ns, VDD,
+ 1416939.800000ns, VDD,
+ 1416939.900000ns, VSS,
+ 1417180.000000ns, VSS,
+ 1417180.100000ns, VDD,
+ 1417300.100000ns, VDD,
+ 1417300.200000ns, VSS,
+ 1417660.400000ns, VSS,
+ 1417660.500000ns, VDD,
+ 1418020.700000ns, VDD,
+ 1418020.800000ns, VSS,
+ 1418140.800000ns, VSS,
+ 1418140.900000ns, VDD,
+ 1418381.000000ns, VDD,
+ 1418381.100000ns, VSS,
+ 1418501.100000ns, VSS,
+ 1418501.200000ns, VDD,
+ 1418621.200000ns, VDD,
+ 1418621.300000ns, VSS,
+ 1418741.300000ns, VSS,
+ 1418741.400000ns, VDD,
+ 1419341.800000ns, VDD,
+ 1419341.900000ns, VSS,
+ 1420182.500000ns, VSS,
+ 1420182.600000ns, VDD,
+ 1420662.900000ns, VDD,
+ 1420663.000000ns, VSS,
+ 1420903.100000ns, VSS,
+ 1420903.200000ns, VDD,
+ 1421743.800000ns, VDD,
+ 1421743.900000ns, VSS,
+ 1421863.900000ns, VSS,
+ 1421864.000000ns, VDD,
+ 1422344.300000ns, VDD,
+ 1422344.400000ns, VSS,
+ 1422464.400000ns, VSS,
+ 1422464.500000ns, VDD,
+ 1422704.600000ns, VDD,
+ 1422704.700000ns, VSS,
+ 1423064.900000ns, VSS,
+ 1423065.000000ns, VDD,
+ 1423185.000000ns, VDD,
+ 1423185.100000ns, VSS,
+ 1423665.400000ns, VSS,
+ 1423665.500000ns, VDD,
+ 1424025.700000ns, VDD,
+ 1424025.800000ns, VSS,
+ 1424506.100000ns, VSS,
+ 1424506.200000ns, VDD,
+ 1424746.300000ns, VDD,
+ 1424746.400000ns, VSS,
+ 1424986.500000ns, VSS,
+ 1424986.600000ns, VDD,
+ 1425226.700000ns, VDD,
+ 1425226.800000ns, VSS,
+ 1425707.100000ns, VSS,
+ 1425707.200000ns, VDD,
+ 1426307.600000ns, VDD,
+ 1426307.700000ns, VSS,
+ 1427628.700000ns, VSS,
+ 1427628.800000ns, VDD,
+ 1428229.200000ns, VDD,
+ 1428229.300000ns, VSS,
+ 1428349.300000ns, VSS,
+ 1428349.400000ns, VDD,
+ 1428829.700000ns, VDD,
+ 1428829.800000ns, VSS,
+ 1429190.000000ns, VSS,
+ 1429190.100000ns, VDD,
+ 1429310.100000ns, VDD,
+ 1429310.200000ns, VSS,
+ 1429550.300000ns, VSS,
+ 1429550.400000ns, VDD,
+ 1429670.400000ns, VDD,
+ 1429670.500000ns, VSS,
+ 1429790.500000ns, VSS,
+ 1429790.600000ns, VDD,
+ 1430511.100000ns, VDD,
+ 1430511.200000ns, VSS,
+ 1431111.600000ns, VSS,
+ 1431111.700000ns, VDD,
+ 1431351.800000ns, VDD,
+ 1431351.900000ns, VSS,
+ 1431592.000000ns, VSS,
+ 1431592.100000ns, VDD,
+ 1431712.100000ns, VDD,
+ 1431712.200000ns, VSS,
+ 1431952.300000ns, VSS,
+ 1431952.400000ns, VDD,
+ 1432312.600000ns, VDD,
+ 1432312.700000ns, VSS,
+ 1432432.700000ns, VSS,
+ 1432432.800000ns, VDD,
+ 1432913.100000ns, VDD,
+ 1432913.200000ns, VSS,
+ 1433753.800000ns, VSS,
+ 1433753.900000ns, VDD,
+ 1433873.900000ns, VDD,
+ 1433874.000000ns, VSS,
+ 1434234.200000ns, VSS,
+ 1434234.300000ns, VDD,
+ 1435315.100000ns, VDD,
+ 1435315.200000ns, VSS,
+ 1436275.900000ns, VSS,
+ 1436276.000000ns, VDD,
+ 1436396.000000ns, VDD,
+ 1436396.100000ns, VSS,
+ 1436756.300000ns, VSS,
+ 1436756.400000ns, VDD,
+ 1436876.400000ns, VDD,
+ 1436876.500000ns, VSS,
+ 1437476.900000ns, VSS,
+ 1437477.000000ns, VDD,
+ 1438918.100000ns, VDD,
+ 1438918.200000ns, VSS,
+ 1439038.200000ns, VSS,
+ 1439038.300000ns, VDD,
+ 1439278.400000ns, VDD,
+ 1439278.500000ns, VSS,
+ 1439398.500000ns, VSS,
+ 1439398.600000ns, VDD,
+ 1439518.600000ns, VDD,
+ 1439518.700000ns, VSS,
+ 1439758.800000ns, VSS,
+ 1439758.900000ns, VDD,
+ 1439878.900000ns, VDD,
+ 1439879.000000ns, VSS,
+ 1440359.300000ns, VSS,
+ 1440359.400000ns, VDD,
+ 1440479.400000ns, VDD,
+ 1440479.500000ns, VSS,
+ 1440959.800000ns, VSS,
+ 1440959.900000ns, VDD,
+ 1441680.400000ns, VDD,
+ 1441680.500000ns, VSS,
+ 1441800.500000ns, VSS,
+ 1441800.600000ns, VDD,
+ 1443121.600000ns, VDD,
+ 1443121.700000ns, VSS,
+ 1443361.800000ns, VSS,
+ 1443361.900000ns, VDD,
+ 1444322.600000ns, VDD,
+ 1444322.700000ns, VSS,
+ 1444682.900000ns, VSS,
+ 1444683.000000ns, VDD,
+ 1445883.900000ns, VDD,
+ 1445884.000000ns, VSS,
+ 1446004.000000ns, VSS,
+ 1446004.100000ns, VDD,
+ 1446364.300000ns, VDD,
+ 1446364.400000ns, VSS,
+ 1446604.500000ns, VSS,
+ 1446604.600000ns, VDD,
+ 1446844.700000ns, VDD,
+ 1446844.800000ns, VSS,
+ 1447205.000000ns, VSS,
+ 1447205.100000ns, VDD,
+ 1448285.900000ns, VDD,
+ 1448286.000000ns, VSS,
+ 1448766.300000ns, VSS,
+ 1448766.400000ns, VDD,
+ 1449486.900000ns, VDD,
+ 1449487.000000ns, VSS,
+ 1449847.200000ns, VSS,
+ 1449847.300000ns, VDD,
+ 1450327.600000ns, VDD,
+ 1450327.700000ns, VSS,
+ 1450567.800000ns, VSS,
+ 1450567.900000ns, VDD,
+ 1451048.200000ns, VDD,
+ 1451048.300000ns, VSS,
+ 1451168.300000ns, VSS,
+ 1451168.400000ns, VDD,
+ 1451528.600000ns, VDD,
+ 1451528.700000ns, VSS,
+ 1451768.800000ns, VSS,
+ 1451768.900000ns, VDD,
+ 1452009.000000ns, VDD,
+ 1452009.100000ns, VSS,
+ 1452249.200000ns, VSS,
+ 1452249.300000ns, VDD,
+ 1452849.700000ns, VDD,
+ 1452849.800000ns, VSS,
+ 1452969.800000ns, VSS,
+ 1452969.900000ns, VDD,
+ 1453210.000000ns, VDD,
+ 1453210.100000ns, VSS,
+ 1453690.400000ns, VSS,
+ 1453690.500000ns, VDD,
+ 1453930.600000ns, VDD,
+ 1453930.700000ns, VSS,
+ 1454771.300000ns, VSS,
+ 1454771.400000ns, VDD,
+ 1455131.600000ns, VDD,
+ 1455131.700000ns, VSS,
+ 1455612.000000ns, VSS,
+ 1455612.100000ns, VDD,
+ 1455972.300000ns, VDD,
+ 1455972.400000ns, VSS,
+ 1456813.000000ns, VSS,
+ 1456813.100000ns, VDD,
+ 1458014.000000ns, VDD,
+ 1458014.100000ns, VSS,
+ 1458134.100000ns, VSS,
+ 1458134.200000ns, VDD,
+ 1458254.200000ns, VDD,
+ 1458254.300000ns, VSS,
+ 1458614.500000ns, VSS,
+ 1458614.600000ns, VDD,
+ 1458854.700000ns, VDD,
+ 1458854.800000ns, VSS,
+ 1459215.000000ns, VSS,
+ 1459215.100000ns, VDD,
+ 1459695.400000ns, VDD,
+ 1459695.500000ns, VSS,
+ 1459815.500000ns, VSS,
+ 1459815.600000ns, VDD,
+ 1460536.100000ns, VDD,
+ 1460536.200000ns, VSS,
+ 1460776.300000ns, VSS,
+ 1460776.400000ns, VDD,
+ 1461016.500000ns, VDD,
+ 1461016.600000ns, VSS,
+ 1461376.800000ns, VSS,
+ 1461376.900000ns, VDD,
+ 1461617.000000ns, VDD,
+ 1461617.100000ns, VSS,
+ 1461737.100000ns, VSS,
+ 1461737.200000ns, VDD,
+ 1461857.200000ns, VDD,
+ 1461857.300000ns, VSS,
+ 1463058.200000ns, VSS,
+ 1463058.300000ns, VDD,
+ 1463418.500000ns, VDD,
+ 1463418.600000ns, VSS,
+ 1463538.600000ns, VSS,
+ 1463538.700000ns, VDD,
+ 1463658.700000ns, VDD,
+ 1463658.800000ns, VSS,
+ 1463778.800000ns, VSS,
+ 1463778.900000ns, VDD,
+ 1464619.500000ns, VDD,
+ 1464619.600000ns, VSS,
+ 1465099.900000ns, VSS,
+ 1465100.000000ns, VDD,
+ 1465340.100000ns, VDD,
+ 1465340.200000ns, VSS,
+ 1465580.300000ns, VSS,
+ 1465580.400000ns, VDD,
+ 1465940.600000ns, VDD,
+ 1465940.700000ns, VSS,
+ 1466300.900000ns, VSS,
+ 1466301.000000ns, VDD,
+ 1466541.100000ns, VDD,
+ 1466541.200000ns, VSS,
+ 1466661.200000ns, VSS,
+ 1466661.300000ns, VDD,
+ 1466901.400000ns, VDD,
+ 1466901.500000ns, VSS,
+ 1467021.500000ns, VSS,
+ 1467021.600000ns, VDD,
+ 1467141.600000ns, VDD,
+ 1467141.700000ns, VSS,
+ 1467381.800000ns, VSS,
+ 1467381.900000ns, VDD,
+ 1467742.100000ns, VDD,
+ 1467742.200000ns, VSS,
+ 1468342.600000ns, VSS,
+ 1468342.700000ns, VDD,
+ 1468702.900000ns, VDD,
+ 1468703.000000ns, VSS,
+ 1469663.700000ns, VSS,
+ 1469663.800000ns, VDD,
+ 1470264.200000ns, VDD,
+ 1470264.300000ns, VSS,
+ 1470744.600000ns, VSS,
+ 1470744.700000ns, VDD,
+ 1470984.800000ns, VDD,
+ 1470984.900000ns, VSS,
+ 1471104.900000ns, VSS,
+ 1471105.000000ns, VDD,
+ 1471225.000000ns, VDD,
+ 1471225.100000ns, VSS,
+ 1471945.600000ns, VSS,
+ 1471945.700000ns, VDD,
+ 1472666.200000ns, VDD,
+ 1472666.300000ns, VSS,
+ 1472786.300000ns, VSS,
+ 1472786.400000ns, VDD,
+ 1473386.800000ns, VDD,
+ 1473386.900000ns, VSS,
+ 1473506.900000ns, VSS,
+ 1473507.000000ns, VDD,
+ 1473627.000000ns, VDD,
+ 1473627.100000ns, VSS,
+ 1473747.100000ns, VSS,
+ 1473747.200000ns, VDD,
+ 1473987.300000ns, VDD,
+ 1473987.400000ns, VSS,
+ 1474107.400000ns, VSS,
+ 1474107.500000ns, VDD,
+ 1474587.800000ns, VDD,
+ 1474587.900000ns, VSS,
+ 1474707.900000ns, VSS,
+ 1474708.000000ns, VDD,
+ 1474948.100000ns, VDD,
+ 1474948.200000ns, VSS,
+ 1475428.500000ns, VSS,
+ 1475428.600000ns, VDD,
+ 1475908.900000ns, VDD,
+ 1475909.000000ns, VSS,
+ 1476029.000000ns, VSS,
+ 1476029.100000ns, VDD,
+ 1476149.100000ns, VDD,
+ 1476149.200000ns, VSS,
+ 1476629.500000ns, VSS,
+ 1476629.600000ns, VDD,
+ 1477590.300000ns, VDD,
+ 1477590.400000ns, VSS,
+ 1478190.800000ns, VSS,
+ 1478190.900000ns, VDD,
+ 1478551.100000ns, VDD,
+ 1478551.200000ns, VSS,
+ 1478671.200000ns, VSS,
+ 1478671.300000ns, VDD,
+ 1478791.300000ns, VDD,
+ 1478791.400000ns, VSS,
+ 1479031.500000ns, VSS,
+ 1479031.600000ns, VDD,
+ 1479872.200000ns, VDD,
+ 1479872.300000ns, VSS,
+ 1480112.400000ns, VSS,
+ 1480112.500000ns, VDD,
+ 1480712.900000ns, VDD,
+ 1480713.000000ns, VSS,
+ 1480833.000000ns, VSS,
+ 1480833.100000ns, VDD,
+ 1481433.500000ns, VDD,
+ 1481433.600000ns, VSS,
+ 1481913.900000ns, VSS,
+ 1481914.000000ns, VDD,
+ 1482034.000000ns, VDD,
+ 1482034.100000ns, VSS,
+ 1482634.500000ns, VSS,
+ 1482634.600000ns, VDD,
+ 1482874.700000ns, VDD,
+ 1482874.800000ns, VSS,
+ 1483595.300000ns, VSS,
+ 1483595.400000ns, VDD,
+ 1483955.600000ns, VDD,
+ 1483955.700000ns, VSS,
+ 1484436.000000ns, VSS,
+ 1484436.100000ns, VDD,
+ 1485396.800000ns, VDD,
+ 1485396.900000ns, VSS,
+ 1485997.300000ns, VSS,
+ 1485997.400000ns, VDD,
+ 1486477.700000ns, VDD,
+ 1486477.800000ns, VSS,
+ 1487198.300000ns, VSS,
+ 1487198.400000ns, VDD,
+ 1487558.600000ns, VDD,
+ 1487558.700000ns, VSS,
+ 1487678.700000ns, VSS,
+ 1487678.800000ns, VDD,
+ 1487918.900000ns, VDD,
+ 1487919.000000ns, VSS,
+ 1488399.300000ns, VSS,
+ 1488399.400000ns, VDD,
+ 1488519.400000ns, VDD,
+ 1488519.500000ns, VSS,
+ 1488999.800000ns, VSS,
+ 1488999.900000ns, VDD,
+ 1489840.500000ns, VDD,
+ 1489840.600000ns, VSS,
+ 1490080.700000ns, VSS,
+ 1490080.800000ns, VDD,
+ 1490561.100000ns, VDD,
+ 1490561.200000ns, VSS,
+ 1490681.200000ns, VSS,
+ 1490681.300000ns, VDD,
+ 1491281.700000ns, VDD,
+ 1491281.800000ns, VSS,
+ 1491762.100000ns, VSS,
+ 1491762.200000ns, VDD,
+ 1492002.300000ns, VDD,
+ 1492002.400000ns, VSS,
+ 1492242.500000ns, VSS,
+ 1492242.600000ns, VDD,
+ 1492362.600000ns, VDD,
+ 1492362.700000ns, VSS,
+ 1492843.000000ns, VSS,
+ 1492843.100000ns, VDD,
+ 1493203.300000ns, VDD,
+ 1493203.400000ns, VSS,
+ 1493563.600000ns, VSS,
+ 1493563.700000ns, VDD,
+ 1494524.400000ns, VDD,
+ 1494524.500000ns, VSS,
+ 1495365.100000ns, VSS,
+ 1495365.200000ns, VDD,
+ 1495485.200000ns, VDD,
+ 1495485.300000ns, VSS,
+ 1496446.000000ns, VSS,
+ 1496446.100000ns, VDD,
+ 1497046.500000ns, VDD,
+ 1497046.600000ns, VSS,
+ 1497286.700000ns, VSS,
+ 1497286.800000ns, VDD,
+ 1497406.800000ns, VDD,
+ 1497406.900000ns, VSS,
+ 1497526.900000ns, VSS,
+ 1497527.000000ns, VDD,
+ 1497887.200000ns, VDD,
+ 1497887.300000ns, VSS,
+ 1498127.400000ns, VSS,
+ 1498127.500000ns, VDD,
+ 1498848.000000ns, VDD,
+ 1498848.100000ns, VSS,
+ 1498968.100000ns, VSS,
+ 1498968.200000ns, VDD,
+ 1499208.300000ns, VDD,
+ 1499208.400000ns, VSS,
+ 1500049.000000ns, VSS,
+ 1500049.100000ns, VDD,
+ 1500289.200000ns, VDD,
+ 1500289.300000ns, VSS,
+ 1500769.600000ns, VSS,
+ 1500769.700000ns, VDD,
+ 1501370.100000ns, VDD,
+ 1501370.200000ns, VSS,
+ 1501850.500000ns, VSS,
+ 1501850.600000ns, VDD,
+ 1502090.700000ns, VDD,
+ 1502090.800000ns, VSS,
+ 1502210.800000ns, VSS,
+ 1502210.900000ns, VDD,
+ 1502811.300000ns, VDD,
+ 1502811.400000ns, VSS,
+ 1502931.400000ns, VSS,
+ 1502931.500000ns, VDD,
+ 1503291.700000ns, VDD,
+ 1503291.800000ns, VSS,
+ 1503531.900000ns, VSS,
+ 1503532.000000ns, VDD,
+ 1503652.000000ns, VDD,
+ 1503652.100000ns, VSS,
+ 1503892.200000ns, VSS,
+ 1503892.300000ns, VDD,
+ 1504252.500000ns, VDD,
+ 1504252.600000ns, VSS,
+ 1504612.800000ns, VSS,
+ 1504612.900000ns, VDD,
+ 1504973.100000ns, VDD,
+ 1504973.200000ns, VSS,
+ 1505213.300000ns, VSS,
+ 1505213.400000ns, VDD,
+ 1505693.700000ns, VDD,
+ 1505693.800000ns, VSS,
+ 1505933.900000ns, VSS,
+ 1505934.000000ns, VDD,
+ 1506054.000000ns, VDD,
+ 1506054.100000ns, VSS,
+ 1506174.100000ns, VSS,
+ 1506174.200000ns, VDD,
+ 1506894.700000ns, VDD,
+ 1506894.800000ns, VSS,
+ 1507375.100000ns, VSS,
+ 1507375.200000ns, VDD,
+ 1507615.300000ns, VDD,
+ 1507615.400000ns, VSS,
+ 1507975.600000ns, VSS,
+ 1507975.700000ns, VDD,
+ 1508215.800000ns, VDD,
+ 1508215.900000ns, VSS,
+ 1508696.200000ns, VSS,
+ 1508696.300000ns, VDD,
+ 1508936.400000ns, VDD,
+ 1508936.500000ns, VSS,
+ 1509056.500000ns, VSS,
+ 1509056.600000ns, VDD,
+ 1509416.800000ns, VDD,
+ 1509416.900000ns, VSS,
+ 1509777.100000ns, VSS,
+ 1509777.200000ns, VDD,
+ 1510137.400000ns, VDD,
+ 1510137.500000ns, VSS,
+ 1510497.700000ns, VSS,
+ 1510497.800000ns, VDD,
+ 1511338.400000ns, VDD,
+ 1511338.500000ns, VSS,
+ 1511578.600000ns, VSS,
+ 1511578.700000ns, VDD,
+ 1512419.300000ns, VDD,
+ 1512419.400000ns, VSS,
+ 1512539.400000ns, VSS,
+ 1512539.500000ns, VDD,
+ 1512899.700000ns, VDD,
+ 1512899.800000ns, VSS,
+ 1513139.900000ns, VSS,
+ 1513140.000000ns, VDD,
+ 1513620.300000ns, VDD,
+ 1513620.400000ns, VSS,
+ 1513740.400000ns, VSS,
+ 1513740.500000ns, VDD,
+ 1514100.700000ns, VDD,
+ 1514100.800000ns, VSS,
+ 1514701.200000ns, VSS,
+ 1514701.300000ns, VDD,
+ 1515061.500000ns, VDD,
+ 1515061.600000ns, VSS,
+ 1515421.800000ns, VSS,
+ 1515421.900000ns, VDD,
+ 1515782.100000ns, VDD,
+ 1515782.200000ns, VSS,
+ 1516022.300000ns, VSS,
+ 1516022.400000ns, VDD,
+ 1516502.700000ns, VDD,
+ 1516502.800000ns, VSS,
+ 1516983.100000ns, VSS,
+ 1516983.200000ns, VDD,
+ 1517583.600000ns, VDD,
+ 1517583.700000ns, VSS,
+ 1517823.800000ns, VSS,
+ 1517823.900000ns, VDD,
+ 1517943.900000ns, VDD,
+ 1517944.000000ns, VSS,
+ 1518064.000000ns, VSS,
+ 1518064.100000ns, VDD,
+ 1518544.400000ns, VDD,
+ 1518544.500000ns, VSS,
+ 1519385.100000ns, VSS,
+ 1519385.200000ns, VDD,
+ 1519745.400000ns, VDD,
+ 1519745.500000ns, VSS,
+ 1520105.700000ns, VSS,
+ 1520105.800000ns, VDD,
+ 1520946.400000ns, VDD,
+ 1520946.500000ns, VSS,
+ 1521426.800000ns, VSS,
+ 1521426.900000ns, VDD,
+ 1521907.200000ns, VDD,
+ 1521907.300000ns, VSS,
+ 1522027.300000ns, VSS,
+ 1522027.400000ns, VDD,
+ 1522147.400000ns, VDD,
+ 1522147.500000ns, VSS,
+ 1522868.000000ns, VSS,
+ 1522868.100000ns, VDD,
+ 1523228.300000ns, VDD,
+ 1523228.400000ns, VSS,
+ 1523468.500000ns, VSS,
+ 1523468.600000ns, VDD,
+ 1523948.900000ns, VDD,
+ 1523949.000000ns, VSS,
+ 1524069.000000ns, VSS,
+ 1524069.100000ns, VDD,
+ 1524189.100000ns, VDD,
+ 1524189.200000ns, VSS,
+ 1524309.200000ns, VSS,
+ 1524309.300000ns, VDD,
+ 1524669.500000ns, VDD,
+ 1524669.600000ns, VSS,
+ 1525149.900000ns, VSS,
+ 1525150.000000ns, VDD,
+ 1525870.500000ns, VDD,
+ 1525870.600000ns, VSS,
+ 1526350.900000ns, VSS,
+ 1526351.000000ns, VDD,
+ 1527551.900000ns, VDD,
+ 1527552.000000ns, VSS,
+ 1527912.200000ns, VSS,
+ 1527912.300000ns, VDD,
+ 1528152.400000ns, VDD,
+ 1528152.500000ns, VSS,
+ 1528272.500000ns, VSS,
+ 1528272.600000ns, VDD,
+ 1528512.700000ns, VDD,
+ 1528512.800000ns, VSS,
+ 1530314.200000ns, VSS,
+ 1530314.300000ns, VDD,
+ 1530674.500000ns, VDD,
+ 1530674.600000ns, VSS,
+ 1530914.700000ns, VSS,
+ 1530914.800000ns, VDD,
+ 1531154.900000ns, VDD,
+ 1531155.000000ns, VSS,
+ 1531275.000000ns, VSS,
+ 1531275.100000ns, VDD,
+ 1531395.100000ns, VDD,
+ 1531395.200000ns, VSS,
+ 1531755.400000ns, VSS,
+ 1531755.500000ns, VDD,
+ 1533196.600000ns, VDD,
+ 1533196.700000ns, VSS,
+ 1533917.200000ns, VSS,
+ 1533917.300000ns, VDD,
+ 1534037.300000ns, VDD,
+ 1534037.400000ns, VSS,
+ 1534637.800000ns, VSS,
+ 1534637.900000ns, VDD,
+ 1534878.000000ns, VDD,
+ 1534878.100000ns, VSS,
+ 1535238.300000ns, VSS,
+ 1535238.400000ns, VDD,
+ 1535598.600000ns, VDD,
+ 1535598.700000ns, VSS,
+ 1536319.200000ns, VSS,
+ 1536319.300000ns, VDD,
+ 1536439.300000ns, VDD,
+ 1536439.400000ns, VSS,
+ 1536679.500000ns, VSS,
+ 1536679.600000ns, VDD,
+ 1538481.000000ns, VDD,
+ 1538481.100000ns, VSS,
+ 1538841.300000ns, VSS,
+ 1538841.400000ns, VDD,
+ 1539201.600000ns, VDD,
+ 1539201.700000ns, VSS,
+ 1539321.700000ns, VSS,
+ 1539321.800000ns, VDD,
+ 1539682.000000ns, VDD,
+ 1539682.100000ns, VSS,
+ 1539922.200000ns, VSS,
+ 1539922.300000ns, VDD,
+ 1540282.500000ns, VDD,
+ 1540282.600000ns, VSS,
+ 1540402.600000ns, VSS,
+ 1540402.700000ns, VDD,
+ 1540522.700000ns, VDD,
+ 1540522.800000ns, VSS,
+ 1540883.000000ns, VSS,
+ 1540883.100000ns, VDD,
+ 1541363.400000ns, VDD,
+ 1541363.500000ns, VSS,
+ 1541843.800000ns, VSS,
+ 1541843.900000ns, VDD,
+ 1543164.900000ns, VDD,
+ 1543165.000000ns, VSS,
+ 1543765.400000ns, VSS,
+ 1543765.500000ns, VDD,
+ 1544005.600000ns, VDD,
+ 1544005.700000ns, VSS,
+ 1544125.700000ns, VSS,
+ 1544125.800000ns, VDD,
+ 1544486.000000ns, VDD,
+ 1544486.100000ns, VSS,
+ 1544726.200000ns, VSS,
+ 1544726.300000ns, VDD,
+ 1544966.400000ns, VDD,
+ 1544966.500000ns, VSS,
+ 1545326.700000ns, VSS,
+ 1545326.800000ns, VDD,
+ 1546767.900000ns, VDD,
+ 1546768.000000ns, VSS,
+ 1546888.000000ns, VSS,
+ 1546888.100000ns, VDD,
+ 1547488.500000ns, VDD,
+ 1547488.600000ns, VSS,
+ 1547608.600000ns, VSS,
+ 1547608.700000ns, VDD,
+ 1547848.800000ns, VDD,
+ 1547848.900000ns, VSS,
+ 1548209.100000ns, VSS,
+ 1548209.200000ns, VDD,
+ 1549049.800000ns, VDD,
+ 1549049.900000ns, VSS,
+ 1549290.000000ns, VSS,
+ 1549290.100000ns, VDD,
+ 1549890.500000ns, VDD,
+ 1549890.600000ns, VSS,
+ 1550010.600000ns, VSS,
+ 1550010.700000ns, VDD
+)}


RSD in_SD 0 1.0
BSD in_SD 0 V={table(time,
+ 0.100000ns, VSS,
+ 240.200000ns, VSS,
+ 240.300000ns, VDD,
+ 720.600000ns, VDD,
+ 720.700000ns, VSS,
+ 960.800000ns, VSS,
+ 960.900000ns, VDD,
+ 1201.000000ns, VDD,
+ 1201.100000ns, VSS,
+ 1321.100000ns, VSS,
+ 1321.200000ns, VDD,
+ 1441.200000ns, VDD,
+ 1441.300000ns, VSS,
+ 1681.400000ns, VSS,
+ 1681.500000ns, VDD,
+ 1801.500000ns, VDD,
+ 1801.600000ns, VSS,
+ 1921.600000ns, VSS,
+ 1921.700000ns, VDD,
+ 2402.000000ns, VDD,
+ 2402.100000ns, VSS,
+ 3362.800000ns, VSS,
+ 3362.900000ns, VDD,
+ 3603.000000ns, VDD,
+ 3603.100000ns, VSS,
+ 3723.100000ns, VSS,
+ 3723.200000ns, VDD,
+ 3843.200000ns, VDD,
+ 3843.300000ns, VSS,
+ 5524.600000ns, VSS,
+ 5524.700000ns, VDD,
+ 7926.600000ns, VDD,
+ 7926.700000ns, VSS,
+ 8166.800000ns, VSS,
+ 8166.900000ns, VDD,
+ 8286.900000ns, VDD,
+ 8287.000000ns, VSS,
+ 9007.500000ns, VSS,
+ 9007.600000ns, VDD,
+ 9247.700000ns, VDD,
+ 9247.800000ns, VSS,
+ 9728.100000ns, VSS,
+ 9728.200000ns, VDD,
+ 10929.100000ns, VDD,
+ 10929.200000ns, VSS,
+ 11649.700000ns, VSS,
+ 11649.800000ns, VDD,
+ 12370.300000ns, VDD,
+ 12370.400000ns, VSS,
+ 12490.400000ns, VSS,
+ 12490.500000ns, VDD,
+ 12850.700000ns, VDD,
+ 12850.800000ns, VSS,
+ 13090.900000ns, VSS,
+ 13091.000000ns, VDD,
+ 13811.500000ns, VDD,
+ 13811.600000ns, VSS,
+ 15613.000000ns, VSS,
+ 15613.100000ns, VDD,
+ 16093.400000ns, VDD,
+ 16093.500000ns, VSS,
+ 19576.300000ns, VSS,
+ 19576.400000ns, VDD,
+ 19696.400000ns, VDD,
+ 19696.500000ns, VSS,
+ 20176.800000ns, VSS,
+ 20176.900000ns, VDD,
+ 20417.000000ns, VDD,
+ 20417.100000ns, VSS,
+ 20537.100000ns, VSS,
+ 20537.200000ns, VDD,
+ 20657.200000ns, VDD,
+ 20657.300000ns, VSS,
+ 21137.600000ns, VSS,
+ 21137.700000ns, VDD,
+ 21618.000000ns, VDD,
+ 21618.100000ns, VSS,
+ 22338.600000ns, VSS,
+ 22338.700000ns, VDD,
+ 22819.000000ns, VDD,
+ 22819.100000ns, VSS,
+ 23299.400000ns, VSS,
+ 23299.500000ns, VDD,
+ 23779.800000ns, VDD,
+ 23779.900000ns, VSS,
+ 24380.300000ns, VSS,
+ 24380.400000ns, VDD,
+ 24740.600000ns, VDD,
+ 24740.700000ns, VSS,
+ 26181.800000ns, VSS,
+ 26181.900000ns, VDD,
+ 26301.900000ns, VDD,
+ 26302.000000ns, VSS,
+ 26422.000000ns, VSS,
+ 26422.100000ns, VDD,
+ 26662.200000ns, VDD,
+ 26662.300000ns, VSS,
+ 26782.300000ns, VSS,
+ 26782.400000ns, VDD,
+ 27262.700000ns, VDD,
+ 27262.800000ns, VSS,
+ 28343.600000ns, VSS,
+ 28343.700000ns, VDD,
+ 29664.700000ns, VDD,
+ 29664.800000ns, VSS,
+ 30265.200000ns, VSS,
+ 30265.300000ns, VDD,
+ 30505.400000ns, VDD,
+ 30505.500000ns, VSS,
+ 30985.800000ns, VSS,
+ 30985.900000ns, VDD,
+ 31466.200000ns, VDD,
+ 31466.300000ns, VSS,
+ 31826.500000ns, VSS,
+ 31826.600000ns, VDD,
+ 32547.100000ns, VDD,
+ 32547.200000ns, VSS,
+ 33147.600000ns, VSS,
+ 33147.700000ns, VDD,
+ 33267.700000ns, VDD,
+ 33267.800000ns, VSS,
+ 33628.000000ns, VSS,
+ 33628.100000ns, VDD,
+ 33748.100000ns, VDD,
+ 33748.200000ns, VSS,
+ 34228.500000ns, VSS,
+ 34228.600000ns, VDD,
+ 34708.900000ns, VDD,
+ 34709.000000ns, VSS,
+ 35429.500000ns, VSS,
+ 35429.600000ns, VDD,
+ 35909.900000ns, VDD,
+ 35910.000000ns, VSS,
+ 36390.300000ns, VSS,
+ 36390.400000ns, VDD,
+ 38792.300000ns, VDD,
+ 38792.400000ns, VSS,
+ 39873.200000ns, VSS,
+ 39873.300000ns, VDD,
+ 39993.300000ns, VDD,
+ 39993.400000ns, VSS,
+ 40834.000000ns, VSS,
+ 40834.100000ns, VDD,
+ 41074.200000ns, VDD,
+ 41074.300000ns, VSS,
+ 41434.500000ns, VSS,
+ 41434.600000ns, VDD,
+ 41674.700000ns, VDD,
+ 41674.800000ns, VSS,
+ 42515.400000ns, VSS,
+ 42515.500000ns, VDD,
+ 42755.600000ns, VDD,
+ 42755.700000ns, VSS,
+ 42875.700000ns, VSS,
+ 42875.800000ns, VDD,
+ 44557.100000ns, VDD,
+ 44557.200000ns, VSS,
+ 45037.500000ns, VSS,
+ 45037.600000ns, VDD,
+ 46238.500000ns, VDD,
+ 46238.600000ns, VSS,
+ 46358.600000ns, VSS,
+ 46358.700000ns, VDD,
+ 46478.700000ns, VDD,
+ 46478.800000ns, VSS,
+ 46718.900000ns, VSS,
+ 46719.000000ns, VDD,
+ 47319.400000ns, VDD,
+ 47319.500000ns, VSS,
+ 48400.300000ns, VSS,
+ 48400.400000ns, VDD,
+ 48640.500000ns, VDD,
+ 48640.600000ns, VSS,
+ 51042.500000ns, VSS,
+ 51042.600000ns, VDD,
+ 51643.000000ns, VDD,
+ 51643.100000ns, VSS,
+ 52483.700000ns, VSS,
+ 52483.800000ns, VDD,
+ 53084.200000ns, VDD,
+ 53084.300000ns, VSS,
+ 53204.300000ns, VSS,
+ 53204.400000ns, VDD,
+ 53324.400000ns, VDD,
+ 53324.500000ns, VSS,
+ 54405.300000ns, VSS,
+ 54405.400000ns, VDD,
+ 54765.600000ns, VDD,
+ 54765.700000ns, VSS,
+ 55726.400000ns, VSS,
+ 55726.500000ns, VDD,
+ 57527.900000ns, VDD,
+ 57528.000000ns, VSS,
+ 58008.300000ns, VSS,
+ 58008.400000ns, VDD,
+ 59209.300000ns, VDD,
+ 59209.400000ns, VSS,
+ 59449.500000ns, VSS,
+ 59449.600000ns, VDD,
+ 59569.600000ns, VDD,
+ 59569.700000ns, VSS,
+ 60290.200000ns, VSS,
+ 60290.300000ns, VDD,
+ 60650.500000ns, VDD,
+ 60650.600000ns, VSS,
+ 61611.300000ns, VSS,
+ 61611.400000ns, VDD,
+ 61731.400000ns, VDD,
+ 61731.500000ns, VSS,
+ 62211.800000ns, VSS,
+ 62211.900000ns, VDD,
+ 62452.000000ns, VDD,
+ 62452.100000ns, VSS,
+ 62572.100000ns, VSS,
+ 62572.200000ns, VDD,
+ 63172.600000ns, VDD,
+ 63172.700000ns, VSS,
+ 65814.800000ns, VSS,
+ 65814.900000ns, VDD,
+ 66175.100000ns, VDD,
+ 66175.200000ns, VSS,
+ 69177.600000ns, VSS,
+ 69177.700000ns, VDD,
+ 69898.200000ns, VDD,
+ 69898.300000ns, VSS,
+ 70979.100000ns, VSS,
+ 70979.200000ns, VDD,
+ 71459.500000ns, VDD,
+ 71459.600000ns, VSS,
+ 72060.000000ns, VSS,
+ 72060.100000ns, VDD,
+ 72300.200000ns, VDD,
+ 72300.300000ns, VSS,
+ 73140.900000ns, VSS,
+ 73141.000000ns, VDD,
+ 74221.800000ns, VDD,
+ 74221.900000ns, VSS,
+ 75302.700000ns, VSS,
+ 75302.800000ns, VDD,
+ 75542.900000ns, VDD,
+ 75543.000000ns, VSS,
+ 78305.200000ns, VSS,
+ 78305.300000ns, VDD,
+ 79266.000000ns, VDD,
+ 79266.100000ns, VSS,
+ 80106.700000ns, VSS,
+ 80106.800000ns, VDD,
+ 80587.100000ns, VDD,
+ 80587.200000ns, VSS,
+ 81908.200000ns, VSS,
+ 81908.300000ns, VDD,
+ 83229.300000ns, VDD,
+ 83229.400000ns, VSS,
+ 83349.400000ns, VSS,
+ 83349.500000ns, VDD,
+ 83469.500000ns, VDD,
+ 83469.600000ns, VSS,
+ 83709.700000ns, VSS,
+ 83709.800000ns, VDD,
+ 84550.400000ns, VDD,
+ 84550.500000ns, VSS,
+ 84670.500000ns, VSS,
+ 84670.600000ns, VDD,
+ 84790.600000ns, VDD,
+ 84790.700000ns, VSS,
+ 86111.700000ns, VSS,
+ 86111.800000ns, VDD,
+ 86832.300000ns, VDD,
+ 86832.400000ns, VSS,
+ 87192.600000ns, VSS,
+ 87192.700000ns, VDD,
+ 88033.300000ns, VDD,
+ 88033.400000ns, VSS,
+ 88513.700000ns, VSS,
+ 88513.800000ns, VDD,
+ 89234.300000ns, VDD,
+ 89234.400000ns, VSS,
+ 90195.100000ns, VSS,
+ 90195.200000ns, VDD,
+ 90555.400000ns, VDD,
+ 90555.500000ns, VSS,
+ 90915.700000ns, VSS,
+ 90915.800000ns, VDD,
+ 91636.300000ns, VDD,
+ 91636.400000ns, VSS,
+ 91876.500000ns, VSS,
+ 91876.600000ns, VDD,
+ 92356.900000ns, VDD,
+ 92357.000000ns, VSS,
+ 92717.200000ns, VSS,
+ 92717.300000ns, VDD,
+ 92837.300000ns, VDD,
+ 92837.400000ns, VSS,
+ 92957.400000ns, VSS,
+ 92957.500000ns, VDD,
+ 94158.400000ns, VDD,
+ 94158.500000ns, VSS,
+ 95719.700000ns, VSS,
+ 95719.800000ns, VDD,
+ 96440.300000ns, VDD,
+ 96440.400000ns, VSS,
+ 97040.800000ns, VSS,
+ 97040.900000ns, VDD,
+ 98241.800000ns, VDD,
+ 98241.900000ns, VSS,
+ 98962.400000ns, VSS,
+ 98962.500000ns, VDD,
+ 99202.600000ns, VDD,
+ 99202.700000ns, VSS,
+ 99683.000000ns, VSS,
+ 99683.100000ns, VDD,
+ 99923.200000ns, VDD,
+ 99923.300000ns, VSS,
+ 100043.300000ns, VSS,
+ 100043.400000ns, VDD,
+ 100643.800000ns, VDD,
+ 100643.900000ns, VSS,
+ 102685.500000ns, VSS,
+ 102685.600000ns, VDD,
+ 102925.700000ns, VDD,
+ 102925.800000ns, VSS,
+ 103646.300000ns, VSS,
+ 103646.400000ns, VDD,
+ 104006.600000ns, VDD,
+ 104006.700000ns, VSS,
+ 105928.200000ns, VSS,
+ 105928.300000ns, VDD,
+ 106528.700000ns, VDD,
+ 106528.800000ns, VSS,
+ 107489.500000ns, VSS,
+ 107489.600000ns, VDD,
+ 108450.300000ns, VDD,
+ 108450.400000ns, VSS,
+ 108810.600000ns, VSS,
+ 108810.700000ns, VDD,
+ 109050.800000ns, VDD,
+ 109050.900000ns, VSS,
+ 109891.500000ns, VSS,
+ 109891.600000ns, VDD,
+ 110011.600000ns, VDD,
+ 110011.700000ns, VSS,
+ 110492.000000ns, VSS,
+ 110492.100000ns, VDD,
+ 110612.100000ns, VDD,
+ 110612.200000ns, VSS,
+ 110732.200000ns, VSS,
+ 110732.300000ns, VDD,
+ 111092.500000ns, VDD,
+ 111092.600000ns, VSS,
+ 111572.900000ns, VSS,
+ 111573.000000ns, VDD,
+ 112293.500000ns, VDD,
+ 112293.600000ns, VSS,
+ 112413.600000ns, VSS,
+ 112413.700000ns, VDD,
+ 113014.100000ns, VDD,
+ 113014.200000ns, VSS,
+ 113374.400000ns, VSS,
+ 113374.500000ns, VDD,
+ 113494.500000ns, VDD,
+ 113494.600000ns, VSS,
+ 113614.600000ns, VSS,
+ 113614.700000ns, VDD,
+ 114935.700000ns, VDD,
+ 114935.800000ns, VSS,
+ 115175.900000ns, VSS,
+ 115176.000000ns, VDD,
+ 116737.200000ns, VDD,
+ 116737.300000ns, VSS,
+ 117577.900000ns, VSS,
+ 117578.000000ns, VDD,
+ 117698.000000ns, VDD,
+ 117698.100000ns, VSS,
+ 118899.000000ns, VSS,
+ 118899.100000ns, VDD,
+ 119139.200000ns, VDD,
+ 119139.300000ns, VSS,
+ 119259.300000ns, VSS,
+ 119259.400000ns, VDD,
+ 119379.400000ns, VDD,
+ 119379.500000ns, VSS,
+ 120100.000000ns, VSS,
+ 120100.100000ns, VDD,
+ 121301.000000ns, VDD,
+ 121301.100000ns, VSS,
+ 122021.600000ns, VSS,
+ 122021.700000ns, VDD,
+ 123342.700000ns, VDD,
+ 123342.800000ns, VSS,
+ 123582.900000ns, VSS,
+ 123583.000000ns, VDD,
+ 123703.000000ns, VDD,
+ 123703.100000ns, VSS,
+ 125384.400000ns, VSS,
+ 125384.500000ns, VDD,
+ 125504.500000ns, VDD,
+ 125504.600000ns, VSS,
+ 125744.700000ns, VSS,
+ 125744.800000ns, VDD,
+ 125864.800000ns, VDD,
+ 125864.900000ns, VSS,
+ 125984.900000ns, VSS,
+ 125985.000000ns, VDD,
+ 127786.400000ns, VDD,
+ 127786.500000ns, VSS,
+ 128386.900000ns, VSS,
+ 128387.000000ns, VDD,
+ 129347.700000ns, VDD,
+ 129347.800000ns, VSS,
+ 129467.800000ns, VSS,
+ 129467.900000ns, VDD,
+ 131869.800000ns, VDD,
+ 131869.900000ns, VSS,
+ 132710.500000ns, VSS,
+ 132710.600000ns, VDD,
+ 133311.000000ns, VDD,
+ 133311.100000ns, VSS,
+ 133671.300000ns, VSS,
+ 133671.400000ns, VDD,
+ 134031.600000ns, VDD,
+ 134031.700000ns, VSS,
+ 134151.700000ns, VSS,
+ 134151.800000ns, VDD,
+ 134992.400000ns, VDD,
+ 134992.500000ns, VSS,
+ 135352.700000ns, VSS,
+ 135352.800000ns, VDD,
+ 136914.000000ns, VDD,
+ 136914.100000ns, VSS,
+ 137274.300000ns, VSS,
+ 137274.400000ns, VDD,
+ 137634.600000ns, VDD,
+ 137634.700000ns, VSS,
+ 138595.400000ns, VSS,
+ 138595.500000ns, VDD,
+ 139556.200000ns, VDD,
+ 139556.300000ns, VSS,
+ 140036.600000ns, VSS,
+ 140036.700000ns, VDD,
+ 140156.700000ns, VDD,
+ 140156.800000ns, VSS,
+ 141597.900000ns, VSS,
+ 141598.000000ns, VDD,
+ 142318.500000ns, VDD,
+ 142318.600000ns, VSS,
+ 143399.400000ns, VSS,
+ 143399.500000ns, VDD,
+ 143519.500000ns, VDD,
+ 143519.600000ns, VSS,
+ 143639.600000ns, VSS,
+ 143639.700000ns, VDD,
+ 144480.300000ns, VDD,
+ 144480.400000ns, VSS,
+ 144600.400000ns, VSS,
+ 144600.500000ns, VDD,
+ 144960.700000ns, VDD,
+ 144960.800000ns, VSS,
+ 146041.600000ns, VSS,
+ 146041.700000ns, VDD,
+ 146762.200000ns, VDD,
+ 146762.300000ns, VSS,
+ 147362.700000ns, VSS,
+ 147362.800000ns, VDD,
+ 148443.600000ns, VDD,
+ 148443.700000ns, VSS,
+ 148924.000000ns, VSS,
+ 148924.100000ns, VDD,
+ 149284.300000ns, VDD,
+ 149284.400000ns, VSS,
+ 149884.800000ns, VSS,
+ 149884.900000ns, VDD,
+ 150485.300000ns, VDD,
+ 150485.400000ns, VSS,
+ 151446.100000ns, VSS,
+ 151446.200000ns, VDD,
+ 151926.500000ns, VDD,
+ 151926.600000ns, VSS,
+ 152046.600000ns, VSS,
+ 152046.700000ns, VDD,
+ 152767.200000ns, VDD,
+ 152767.300000ns, VSS,
+ 153367.700000ns, VSS,
+ 153367.800000ns, VDD,
+ 153728.000000ns, VDD,
+ 153728.100000ns, VSS,
+ 155049.100000ns, VSS,
+ 155049.200000ns, VDD,
+ 155529.500000ns, VDD,
+ 155529.600000ns, VSS,
+ 155769.700000ns, VSS,
+ 155769.800000ns, VDD,
+ 156730.500000ns, VDD,
+ 156730.600000ns, VSS,
+ 159492.800000ns, VSS,
+ 159492.900000ns, VDD,
+ 159973.200000ns, VDD,
+ 159973.300000ns, VSS,
+ 162135.000000ns, VSS,
+ 162135.100000ns, VDD,
+ 162975.700000ns, VDD,
+ 162975.800000ns, VSS,
+ 163095.800000ns, VSS,
+ 163095.900000ns, VDD,
+ 164657.100000ns, VDD,
+ 164657.200000ns, VSS,
+ 165137.500000ns, VSS,
+ 165137.600000ns, VDD,
+ 165738.000000ns, VDD,
+ 165738.100000ns, VSS,
+ 166458.600000ns, VSS,
+ 166458.700000ns, VDD,
+ 166698.800000ns, VDD,
+ 166698.900000ns, VSS,
+ 166939.000000ns, VSS,
+ 166939.100000ns, VDD,
+ 167179.200000ns, VDD,
+ 167179.300000ns, VSS,
+ 167299.300000ns, VSS,
+ 167299.400000ns, VDD,
+ 167419.400000ns, VDD,
+ 167419.500000ns, VSS,
+ 167779.700000ns, VSS,
+ 167779.800000ns, VDD,
+ 168019.900000ns, VDD,
+ 168020.000000ns, VSS,
+ 168500.300000ns, VSS,
+ 168500.400000ns, VDD,
+ 170061.600000ns, VDD,
+ 170061.700000ns, VSS,
+ 170301.800000ns, VSS,
+ 170301.900000ns, VDD,
+ 170542.000000ns, VDD,
+ 170542.100000ns, VSS,
+ 171022.400000ns, VSS,
+ 171022.500000ns, VDD,
+ 171502.800000ns, VDD,
+ 171502.900000ns, VSS,
+ 172703.800000ns, VSS,
+ 172703.900000ns, VDD,
+ 172944.000000ns, VDD,
+ 172944.100000ns, VSS,
+ 173184.200000ns, VSS,
+ 173184.300000ns, VDD,
+ 174024.900000ns, VDD,
+ 174025.000000ns, VSS,
+ 174265.100000ns, VSS,
+ 174265.200000ns, VDD,
+ 175225.900000ns, VDD,
+ 175226.000000ns, VSS,
+ 176186.700000ns, VSS,
+ 176186.800000ns, VDD,
+ 176306.800000ns, VDD,
+ 176306.900000ns, VSS,
+ 177748.000000ns, VSS,
+ 177748.100000ns, VDD,
+ 178348.500000ns, VDD,
+ 178348.600000ns, VSS,
+ 178708.800000ns, VSS,
+ 178708.900000ns, VDD,
+ 179189.200000ns, VDD,
+ 179189.300000ns, VSS,
+ 179549.500000ns, VSS,
+ 179549.600000ns, VDD,
+ 180029.900000ns, VDD,
+ 180030.000000ns, VSS,
+ 181110.800000ns, VSS,
+ 181110.900000ns, VDD,
+ 181591.200000ns, VDD,
+ 181591.300000ns, VSS,
+ 181831.400000ns, VSS,
+ 181831.500000ns, VDD,
+ 182071.600000ns, VDD,
+ 182071.700000ns, VSS,
+ 182191.700000ns, VSS,
+ 182191.800000ns, VDD,
+ 182311.800000ns, VDD,
+ 182311.900000ns, VSS,
+ 184233.400000ns, VSS,
+ 184233.500000ns, VDD,
+ 185314.300000ns, VDD,
+ 185314.400000ns, VSS,
+ 185674.600000ns, VSS,
+ 185674.700000ns, VDD,
+ 186635.400000ns, VDD,
+ 186635.500000ns, VSS,
+ 186995.700000ns, VSS,
+ 186995.800000ns, VDD,
+ 187115.800000ns, VDD,
+ 187115.900000ns, VSS,
+ 187356.000000ns, VSS,
+ 187356.100000ns, VDD,
+ 187476.100000ns, VDD,
+ 187476.200000ns, VSS,
+ 188557.000000ns, VSS,
+ 188557.100000ns, VDD,
+ 190238.400000ns, VDD,
+ 190238.500000ns, VSS,
+ 190598.700000ns, VSS,
+ 190598.800000ns, VDD,
+ 191799.700000ns, VDD,
+ 191799.800000ns, VSS,
+ 192520.300000ns, VSS,
+ 192520.400000ns, VDD,
+ 192880.600000ns, VDD,
+ 192880.700000ns, VSS,
+ 193841.400000ns, VSS,
+ 193841.500000ns, VDD,
+ 194802.200000ns, VDD,
+ 194802.300000ns, VSS,
+ 195402.700000ns, VSS,
+ 195402.800000ns, VDD,
+ 195522.800000ns, VDD,
+ 195522.900000ns, VSS,
+ 195642.900000ns, VSS,
+ 195643.000000ns, VDD,
+ 196843.900000ns, VDD,
+ 196844.000000ns, VSS,
+ 199245.900000ns, VSS,
+ 199246.000000ns, VDD,
+ 199486.100000ns, VDD,
+ 199486.200000ns, VSS,
+ 199966.500000ns, VSS,
+ 199966.600000ns, VDD,
+ 200446.900000ns, VDD,
+ 200447.000000ns, VSS,
+ 200567.000000ns, VSS,
+ 200567.100000ns, VDD,
+ 200687.100000ns, VDD,
+ 200687.200000ns, VSS,
+ 201768.000000ns, VSS,
+ 201768.100000ns, VDD,
+ 202368.500000ns, VDD,
+ 202368.600000ns, VSS,
+ 203209.200000ns, VSS,
+ 203209.300000ns, VDD,
+ 204890.600000ns, VDD,
+ 204890.700000ns, VSS,
+ 205851.400000ns, VSS,
+ 205851.500000ns, VDD,
+ 206091.600000ns, VDD,
+ 206091.700000ns, VSS,
+ 206331.800000ns, VSS,
+ 206331.900000ns, VDD,
+ 206692.100000ns, VDD,
+ 206692.200000ns, VSS,
+ 206812.200000ns, VSS,
+ 206812.300000ns, VDD,
+ 208253.400000ns, VDD,
+ 208253.500000ns, VSS,
+ 208853.900000ns, VSS,
+ 208854.000000ns, VDD,
+ 208974.000000ns, VDD,
+ 208974.100000ns, VSS,
+ 210295.100000ns, VSS,
+ 210295.200000ns, VDD,
+ 210655.400000ns, VDD,
+ 210655.500000ns, VSS,
+ 211496.100000ns, VSS,
+ 211496.200000ns, VDD,
+ 212456.900000ns, VDD,
+ 212457.000000ns, VSS,
+ 214378.500000ns, VSS,
+ 214378.600000ns, VDD,
+ 216059.900000ns, VDD,
+ 216060.000000ns, VSS,
+ 216300.100000ns, VSS,
+ 216300.200000ns, VDD,
+ 217260.900000ns, VDD,
+ 217261.000000ns, VSS,
+ 219662.900000ns, VSS,
+ 219663.000000ns, VDD,
+ 220503.600000ns, VDD,
+ 220503.700000ns, VSS,
+ 220743.800000ns, VSS,
+ 220743.900000ns, VDD,
+ 221224.200000ns, VDD,
+ 221224.300000ns, VSS,
+ 223025.700000ns, VSS,
+ 223025.800000ns, VDD,
+ 223626.200000ns, VDD,
+ 223626.300000ns, VSS,
+ 223746.300000ns, VSS,
+ 223746.400000ns, VDD,
+ 223986.500000ns, VDD,
+ 223986.600000ns, VSS,
+ 224226.700000ns, VSS,
+ 224226.800000ns, VDD,
+ 224466.900000ns, VDD,
+ 224467.000000ns, VSS,
+ 225187.500000ns, VSS,
+ 225187.600000ns, VDD,
+ 225307.600000ns, VDD,
+ 225307.700000ns, VSS,
+ 225547.800000ns, VSS,
+ 225547.900000ns, VDD,
+ 225667.900000ns, VDD,
+ 225668.000000ns, VSS,
+ 226148.300000ns, VSS,
+ 226148.400000ns, VDD,
+ 226628.700000ns, VDD,
+ 226628.800000ns, VSS,
+ 227469.400000ns, VSS,
+ 227469.500000ns, VDD,
+ 228190.000000ns, VDD,
+ 228190.100000ns, VSS,
+ 228310.100000ns, VSS,
+ 228310.200000ns, VDD,
+ 228550.300000ns, VDD,
+ 228550.400000ns, VSS,
+ 230111.600000ns, VSS,
+ 230111.700000ns, VDD,
+ 230351.800000ns, VDD,
+ 230351.900000ns, VSS,
+ 231072.400000ns, VSS,
+ 231072.500000ns, VDD,
+ 231552.800000ns, VDD,
+ 231552.900000ns, VSS,
+ 232513.600000ns, VSS,
+ 232513.700000ns, VDD,
+ 233114.100000ns, VDD,
+ 233114.200000ns, VSS,
+ 233234.200000ns, VSS,
+ 233234.300000ns, VDD,
+ 234074.900000ns, VDD,
+ 234075.000000ns, VSS,
+ 234315.100000ns, VSS,
+ 234315.200000ns, VDD,
+ 234795.500000ns, VDD,
+ 234795.600000ns, VSS,
+ 235275.900000ns, VSS,
+ 235276.000000ns, VDD,
+ 236957.300000ns, VDD,
+ 236957.400000ns, VSS,
+ 237557.800000ns, VSS,
+ 237557.900000ns, VDD,
+ 238038.200000ns, VDD,
+ 238038.300000ns, VSS,
+ 238638.700000ns, VSS,
+ 238638.800000ns, VDD,
+ 238758.800000ns, VDD,
+ 238758.900000ns, VSS,
+ 239839.700000ns, VSS,
+ 239839.800000ns, VDD,
+ 242121.600000ns, VDD,
+ 242121.700000ns, VSS,
+ 243082.400000ns, VSS,
+ 243082.500000ns, VDD,
+ 244643.700000ns, VDD,
+ 244643.800000ns, VSS,
+ 245124.100000ns, VSS,
+ 245124.200000ns, VDD,
+ 246925.600000ns, VDD,
+ 246925.700000ns, VSS,
+ 248126.600000ns, VSS,
+ 248126.700000ns, VDD,
+ 248486.900000ns, VDD,
+ 248487.000000ns, VSS,
+ 249687.900000ns, VSS,
+ 249688.000000ns, VDD,
+ 249928.100000ns, VDD,
+ 249928.200000ns, VSS,
+ 250048.200000ns, VSS,
+ 250048.300000ns, VDD,
+ 251009.000000ns, VDD,
+ 251009.100000ns, VSS,
+ 251969.800000ns, VSS,
+ 251969.900000ns, VDD,
+ 252450.200000ns, VDD,
+ 252450.300000ns, VSS,
+ 253891.400000ns, VSS,
+ 253891.500000ns, VDD,
+ 254131.600000ns, VDD,
+ 254131.700000ns, VSS,
+ 254732.100000ns, VSS,
+ 254732.200000ns, VDD,
+ 255813.000000ns, VDD,
+ 255813.100000ns, VSS,
+ 256413.500000ns, VSS,
+ 256413.600000ns, VDD,
+ 258094.900000ns, VDD,
+ 258095.000000ns, VSS,
+ 258335.100000ns, VSS,
+ 258335.200000ns, VDD,
+ 258575.300000ns, VDD,
+ 258575.400000ns, VSS,
+ 258815.500000ns, VSS,
+ 258815.600000ns, VDD,
+ 259295.900000ns, VDD,
+ 259296.000000ns, VSS,
+ 260136.600000ns, VSS,
+ 260136.700000ns, VDD,
+ 260857.200000ns, VDD,
+ 260857.300000ns, VSS,
+ 261457.700000ns, VSS,
+ 261457.800000ns, VDD,
+ 261938.100000ns, VDD,
+ 261938.200000ns, VSS,
+ 262298.400000ns, VSS,
+ 262298.500000ns, VDD,
+ 262418.500000ns, VDD,
+ 262418.600000ns, VSS,
+ 262778.800000ns, VSS,
+ 262778.900000ns, VDD,
+ 262898.900000ns, VDD,
+ 262899.000000ns, VSS,
+ 263379.300000ns, VSS,
+ 263379.400000ns, VDD,
+ 264220.000000ns, VDD,
+ 264220.100000ns, VSS,
+ 265060.700000ns, VSS,
+ 265060.800000ns, VDD,
+ 265541.100000ns, VDD,
+ 265541.200000ns, VSS,
+ 266501.900000ns, VSS,
+ 266502.000000ns, VDD,
+ 267342.600000ns, VDD,
+ 267342.700000ns, VSS,
+ 268063.200000ns, VSS,
+ 268063.300000ns, VDD,
+ 268543.600000ns, VDD,
+ 268543.700000ns, VSS,
+ 269144.100000ns, VSS,
+ 269144.200000ns, VDD,
+ 270104.900000ns, VDD,
+ 270105.000000ns, VSS,
+ 270345.100000ns, VSS,
+ 270345.200000ns, VDD,
+ 270825.500000ns, VDD,
+ 270825.600000ns, VSS,
+ 270945.600000ns, VSS,
+ 270945.700000ns, VDD,
+ 271426.000000ns, VDD,
+ 271426.100000ns, VSS,
+ 271546.100000ns, VSS,
+ 271546.200000ns, VDD,
+ 271666.200000ns, VDD,
+ 271666.300000ns, VSS,
+ 272386.800000ns, VSS,
+ 272386.900000ns, VDD,
+ 273347.600000ns, VDD,
+ 273347.700000ns, VSS,
+ 273707.900000ns, VSS,
+ 273708.000000ns, VDD,
+ 274788.800000ns, VDD,
+ 274788.900000ns, VSS,
+ 275629.500000ns, VSS,
+ 275629.600000ns, VDD,
+ 277551.100000ns, VDD,
+ 277551.200000ns, VSS,
+ 278391.800000ns, VSS,
+ 278391.900000ns, VDD,
+ 278872.200000ns, VDD,
+ 278872.300000ns, VSS,
+ 278992.300000ns, VSS,
+ 278992.400000ns, VDD,
+ 279112.400000ns, VDD,
+ 279112.500000ns, VSS,
+ 280193.300000ns, VSS,
+ 280193.400000ns, VDD,
+ 280313.400000ns, VDD,
+ 280313.500000ns, VSS,
+ 280673.700000ns, VSS,
+ 280673.800000ns, VDD,
+ 281154.100000ns, VDD,
+ 281154.200000ns, VSS,
+ 281634.500000ns, VSS,
+ 281634.600000ns, VDD,
+ 282355.100000ns, VDD,
+ 282355.200000ns, VSS,
+ 283075.700000ns, VSS,
+ 283075.800000ns, VDD,
+ 284997.300000ns, VDD,
+ 284997.400000ns, VSS,
+ 285237.500000ns, VSS,
+ 285237.600000ns, VDD,
+ 286918.900000ns, VDD,
+ 286919.000000ns, VSS,
+ 287159.100000ns, VSS,
+ 287159.200000ns, VDD,
+ 287399.300000ns, VDD,
+ 287399.400000ns, VSS,
+ 287759.600000ns, VSS,
+ 287759.700000ns, VDD,
+ 287879.700000ns, VDD,
+ 287879.800000ns, VSS,
+ 287999.800000ns, VSS,
+ 287999.900000ns, VDD,
+ 288840.500000ns, VDD,
+ 288840.600000ns, VSS,
+ 289561.100000ns, VSS,
+ 289561.200000ns, VDD,
+ 290161.600000ns, VDD,
+ 290161.700000ns, VSS,
+ 290762.100000ns, VSS,
+ 290762.200000ns, VDD,
+ 290882.200000ns, VDD,
+ 290882.300000ns, VSS,
+ 291362.600000ns, VSS,
+ 291362.700000ns, VDD,
+ 291722.900000ns, VDD,
+ 291723.000000ns, VSS,
+ 292203.300000ns, VSS,
+ 292203.400000ns, VDD,
+ 293884.700000ns, VDD,
+ 293884.800000ns, VSS,
+ 294004.800000ns, VSS,
+ 294004.900000ns, VDD,
+ 294605.300000ns, VDD,
+ 294605.400000ns, VSS,
+ 295085.700000ns, VSS,
+ 295085.800000ns, VDD,
+ 295446.000000ns, VDD,
+ 295446.100000ns, VSS,
+ 295566.100000ns, VSS,
+ 295566.200000ns, VDD,
+ 296526.900000ns, VDD,
+ 296527.000000ns, VSS,
+ 297007.300000ns, VSS,
+ 297007.400000ns, VDD,
+ 297247.500000ns, VDD,
+ 297247.600000ns, VSS,
+ 297367.600000ns, VSS,
+ 297367.700000ns, VDD,
+ 297607.800000ns, VDD,
+ 297607.900000ns, VSS,
+ 297727.900000ns, VSS,
+ 297728.000000ns, VDD,
+ 298208.300000ns, VDD,
+ 298208.400000ns, VSS,
+ 298568.600000ns, VSS,
+ 298568.700000ns, VDD,
+ 300490.200000ns, VDD,
+ 300490.300000ns, VSS,
+ 301090.700000ns, VSS,
+ 301090.800000ns, VDD,
+ 302652.000000ns, VDD,
+ 302652.100000ns, VSS,
+ 303132.400000ns, VSS,
+ 303132.500000ns, VDD,
+ 303252.500000ns, VDD,
+ 303252.600000ns, VSS,
+ 304213.300000ns, VSS,
+ 304213.400000ns, VDD,
+ 304453.500000ns, VDD,
+ 304453.600000ns, VSS,
+ 304693.700000ns, VSS,
+ 304693.800000ns, VDD,
+ 305654.500000ns, VDD,
+ 305654.600000ns, VSS,
+ 305774.600000ns, VSS,
+ 305774.700000ns, VDD,
+ 305894.700000ns, VDD,
+ 305894.800000ns, VSS,
+ 306735.400000ns, VSS,
+ 306735.500000ns, VDD,
+ 307215.800000ns, VDD,
+ 307215.900000ns, VSS,
+ 308056.500000ns, VSS,
+ 308056.600000ns, VDD,
+ 308536.900000ns, VDD,
+ 308537.000000ns, VSS,
+ 309017.300000ns, VSS,
+ 309017.400000ns, VDD,
+ 309737.900000ns, VDD,
+ 309738.000000ns, VSS,
+ 309858.000000ns, VSS,
+ 309858.100000ns, VDD,
+ 311419.300000ns, VDD,
+ 311419.400000ns, VSS,
+ 312740.400000ns, VSS,
+ 312740.500000ns, VDD,
+ 312980.600000ns, VDD,
+ 312980.700000ns, VSS,
+ 313100.700000ns, VSS,
+ 313100.800000ns, VDD,
+ 315142.400000ns, VDD,
+ 315142.500000ns, VSS,
+ 315863.000000ns, VSS,
+ 315863.100000ns, VDD,
+ 316583.600000ns, VDD,
+ 316583.700000ns, VSS,
+ 316703.700000ns, VSS,
+ 316703.800000ns, VDD,
+ 318265.000000ns, VDD,
+ 318265.100000ns, VSS,
+ 318745.400000ns, VSS,
+ 318745.500000ns, VDD,
+ 319586.100000ns, VDD,
+ 319586.200000ns, VSS,
+ 319706.200000ns, VSS,
+ 319706.300000ns, VDD,
+ 320186.600000ns, VDD,
+ 320186.700000ns, VSS,
+ 321627.800000ns, VSS,
+ 321627.900000ns, VDD,
+ 322588.600000ns, VDD,
+ 322588.700000ns, VSS,
+ 322828.800000ns, VSS,
+ 322828.900000ns, VDD,
+ 323429.300000ns, VDD,
+ 323429.400000ns, VSS,
+ 324390.100000ns, VSS,
+ 324390.200000ns, VDD,
+ 326071.500000ns, VDD,
+ 326071.600000ns, VSS,
+ 326551.900000ns, VSS,
+ 326552.000000ns, VDD,
+ 327032.300000ns, VDD,
+ 327032.400000ns, VSS,
+ 327392.600000ns, VSS,
+ 327392.700000ns, VDD,
+ 327632.800000ns, VDD,
+ 327632.900000ns, VSS,
+ 327873.000000ns, VSS,
+ 327873.100000ns, VDD,
+ 328353.400000ns, VDD,
+ 328353.500000ns, VSS,
+ 328473.500000ns, VSS,
+ 328473.600000ns, VDD,
+ 329074.000000ns, VDD,
+ 329074.100000ns, VSS,
+ 329794.600000ns, VSS,
+ 329794.700000ns, VDD,
+ 331716.200000ns, VDD,
+ 331716.300000ns, VSS,
+ 331836.300000ns, VSS,
+ 331836.400000ns, VDD,
+ 332076.500000ns, VDD,
+ 332076.600000ns, VSS,
+ 332196.600000ns, VSS,
+ 332196.700000ns, VDD,
+ 332316.700000ns, VDD,
+ 332316.800000ns, VSS,
+ 333517.700000ns, VSS,
+ 333517.800000ns, VDD,
+ 334358.400000ns, VDD,
+ 334358.500000ns, VSS,
+ 335199.100000ns, VSS,
+ 335199.200000ns, VDD,
+ 335559.400000ns, VDD,
+ 335559.500000ns, VSS,
+ 335679.500000ns, VSS,
+ 335679.600000ns, VDD,
+ 336280.000000ns, VDD,
+ 336280.100000ns, VSS,
+ 337841.300000ns, VSS,
+ 337841.400000ns, VDD,
+ 338441.800000ns, VDD,
+ 338441.900000ns, VSS,
+ 339642.800000ns, VSS,
+ 339642.900000ns, VDD,
+ 339762.900000ns, VDD,
+ 339763.000000ns, VSS,
+ 340843.800000ns, VSS,
+ 340843.900000ns, VDD,
+ 341324.200000ns, VDD,
+ 341324.300000ns, VSS,
+ 343245.800000ns, VSS,
+ 343245.900000ns, VDD,
+ 344446.800000ns, VDD,
+ 344446.900000ns, VSS,
+ 345407.600000ns, VSS,
+ 345407.700000ns, VDD,
+ 346008.100000ns, VDD,
+ 346008.200000ns, VSS,
+ 347929.700000ns, VSS,
+ 347929.800000ns, VDD,
+ 348650.300000ns, VDD,
+ 348650.400000ns, VSS,
+ 349491.000000ns, VSS,
+ 349491.100000ns, VDD,
+ 350331.700000ns, VDD,
+ 350331.800000ns, VSS,
+ 351532.700000ns, VSS,
+ 351532.800000ns, VDD,
+ 352013.100000ns, VDD,
+ 352013.200000ns, VSS,
+ 352373.400000ns, VSS,
+ 352373.500000ns, VDD,
+ 352853.800000ns, VDD,
+ 352853.900000ns, VSS,
+ 353574.400000ns, VSS,
+ 353574.500000ns, VDD,
+ 354775.400000ns, VDD,
+ 354775.500000ns, VSS,
+ 355736.200000ns, VSS,
+ 355736.300000ns, VDD,
+ 355976.400000ns, VDD,
+ 355976.500000ns, VSS,
+ 356216.600000ns, VSS,
+ 356216.700000ns, VDD,
+ 357057.300000ns, VDD,
+ 357057.400000ns, VSS,
+ 358018.100000ns, VSS,
+ 358018.200000ns, VDD,
+ 358858.800000ns, VDD,
+ 358858.900000ns, VSS,
+ 359339.200000ns, VSS,
+ 359339.300000ns, VDD,
+ 359699.500000ns, VDD,
+ 359699.600000ns, VSS,
+ 359819.600000ns, VSS,
+ 359819.700000ns, VDD,
+ 361501.000000ns, VDD,
+ 361501.100000ns, VSS,
+ 361741.200000ns, VSS,
+ 361741.300000ns, VDD,
+ 362581.900000ns, VDD,
+ 362582.000000ns, VSS,
+ 363662.800000ns, VSS,
+ 363662.900000ns, VDD,
+ 364743.700000ns, VDD,
+ 364743.800000ns, VSS,
+ 365224.100000ns, VSS,
+ 365224.200000ns, VDD,
+ 365584.400000ns, VDD,
+ 365584.500000ns, VSS,
+ 367145.700000ns, VSS,
+ 367145.800000ns, VDD,
+ 367746.200000ns, VDD,
+ 367746.300000ns, VSS,
+ 367986.400000ns, VSS,
+ 367986.500000ns, VDD,
+ 368106.500000ns, VDD,
+ 368106.600000ns, VSS,
+ 368346.700000ns, VSS,
+ 368346.800000ns, VDD,
+ 368466.800000ns, VDD,
+ 368466.900000ns, VSS,
+ 369908.000000ns, VSS,
+ 369908.100000ns, VDD,
+ 370148.200000ns, VDD,
+ 370148.300000ns, VSS,
+ 370388.400000ns, VSS,
+ 370388.500000ns, VDD,
+ 370628.600000ns, VDD,
+ 370628.700000ns, VSS,
+ 374952.200000ns, VSS,
+ 374952.300000ns, VDD,
+ 375192.400000ns, VDD,
+ 375192.500000ns, VSS,
+ 376033.100000ns, VSS,
+ 376033.200000ns, VDD,
+ 376633.600000ns, VDD,
+ 376633.700000ns, VSS,
+ 376993.900000ns, VSS,
+ 376994.000000ns, VDD,
+ 377234.100000ns, VDD,
+ 377234.200000ns, VSS,
+ 378315.000000ns, VSS,
+ 378315.100000ns, VDD,
+ 378795.400000ns, VDD,
+ 378795.500000ns, VSS,
+ 379035.600000ns, VSS,
+ 379035.700000ns, VDD,
+ 379275.800000ns, VDD,
+ 379275.900000ns, VSS,
+ 379996.400000ns, VSS,
+ 379996.500000ns, VDD,
+ 381197.400000ns, VDD,
+ 381197.500000ns, VSS,
+ 381677.800000ns, VSS,
+ 381677.900000ns, VDD,
+ 382398.400000ns, VDD,
+ 382398.500000ns, VSS,
+ 383839.600000ns, VSS,
+ 383839.700000ns, VDD,
+ 384680.300000ns, VDD,
+ 384680.400000ns, VSS,
+ 385040.600000ns, VSS,
+ 385040.700000ns, VDD,
+ 385400.900000ns, VDD,
+ 385401.000000ns, VSS,
+ 386001.400000ns, VSS,
+ 386001.500000ns, VDD,
+ 386121.500000ns, VDD,
+ 386121.600000ns, VSS,
+ 386241.600000ns, VSS,
+ 386241.700000ns, VDD,
+ 387082.300000ns, VDD,
+ 387082.400000ns, VSS,
+ 387322.500000ns, VSS,
+ 387322.600000ns, VDD,
+ 387442.600000ns, VDD,
+ 387442.700000ns, VSS,
+ 388883.800000ns, VSS,
+ 388883.900000ns, VDD,
+ 389364.200000ns, VDD,
+ 389364.300000ns, VSS,
+ 389724.500000ns, VSS,
+ 389724.600000ns, VDD,
+ 391405.900000ns, VDD,
+ 391406.000000ns, VSS,
+ 392006.400000ns, VSS,
+ 392006.500000ns, VDD,
+ 392246.600000ns, VDD,
+ 392246.700000ns, VSS,
+ 392486.800000ns, VSS,
+ 392486.900000ns, VDD,
+ 392967.200000ns, VDD,
+ 392967.300000ns, VSS,
+ 393567.700000ns, VSS,
+ 393567.800000ns, VDD,
+ 394408.400000ns, VDD,
+ 394408.500000ns, VSS,
+ 394888.800000ns, VSS,
+ 394888.900000ns, VDD,
+ 395729.500000ns, VDD,
+ 395729.600000ns, VSS,
+ 396089.800000ns, VSS,
+ 396089.900000ns, VDD,
+ 396810.400000ns, VDD,
+ 396810.500000ns, VSS,
+ 398852.100000ns, VSS,
+ 398852.200000ns, VDD,
+ 400053.100000ns, VDD,
+ 400053.200000ns, VSS,
+ 401374.200000ns, VSS,
+ 401374.300000ns, VDD,
+ 401854.600000ns, VDD,
+ 401854.700000ns, VSS,
+ 402455.100000ns, VSS,
+ 402455.200000ns, VDD,
+ 402935.500000ns, VDD,
+ 402935.600000ns, VSS,
+ 404016.400000ns, VSS,
+ 404016.500000ns, VDD,
+ 404256.600000ns, VDD,
+ 404256.700000ns, VSS,
+ 404496.800000ns, VSS,
+ 404496.900000ns, VDD,
+ 404857.100000ns, VDD,
+ 404857.200000ns, VSS,
+ 406418.400000ns, VSS,
+ 406418.500000ns, VDD,
+ 407379.200000ns, VDD,
+ 407379.300000ns, VSS,
+ 408460.100000ns, VSS,
+ 408460.200000ns, VDD,
+ 408940.500000ns, VDD,
+ 408940.600000ns, VSS,
+ 412063.100000ns, VSS,
+ 412063.200000ns, VDD,
+ 413984.700000ns, VDD,
+ 413984.800000ns, VSS,
+ 414465.100000ns, VSS,
+ 414465.200000ns, VDD,
+ 414585.200000ns, VDD,
+ 414585.300000ns, VSS,
+ 415666.100000ns, VSS,
+ 415666.200000ns, VDD,
+ 415906.300000ns, VDD,
+ 415906.400000ns, VSS,
+ 417227.400000ns, VSS,
+ 417227.500000ns, VDD,
+ 418308.300000ns, VDD,
+ 418308.400000ns, VSS,
+ 418788.700000ns, VSS,
+ 418788.800000ns, VDD,
+ 419509.300000ns, VDD,
+ 419509.400000ns, VSS,
+ 419989.700000ns, VSS,
+ 419989.800000ns, VDD,
+ 420109.800000ns, VDD,
+ 420109.900000ns, VSS,
+ 420710.300000ns, VSS,
+ 420710.400000ns, VDD,
+ 420950.500000ns, VDD,
+ 420950.600000ns, VSS,
+ 421070.600000ns, VSS,
+ 421070.700000ns, VDD,
+ 421190.700000ns, VDD,
+ 421190.800000ns, VSS,
+ 422992.200000ns, VSS,
+ 422992.300000ns, VDD,
+ 423953.000000ns, VDD,
+ 423953.100000ns, VSS,
+ 424193.200000ns, VSS,
+ 424193.300000ns, VDD,
+ 424313.300000ns, VDD,
+ 424313.400000ns, VSS,
+ 425033.900000ns, VSS,
+ 425034.000000ns, VDD,
+ 425514.300000ns, VDD,
+ 425514.400000ns, VSS,
+ 425634.400000ns, VSS,
+ 425634.500000ns, VDD,
+ 426114.800000ns, VDD,
+ 426114.900000ns, VSS,
+ 426355.000000ns, VSS,
+ 426355.100000ns, VDD,
+ 426955.500000ns, VDD,
+ 426955.600000ns, VSS,
+ 427075.600000ns, VSS,
+ 427075.700000ns, VDD,
+ 427435.900000ns, VDD,
+ 427436.000000ns, VSS,
+ 428396.700000ns, VSS,
+ 428396.800000ns, VDD,
+ 429958.000000ns, VDD,
+ 429958.100000ns, VSS,
+ 430198.200000ns, VSS,
+ 430198.300000ns, VDD,
+ 430318.300000ns, VDD,
+ 430318.400000ns, VSS,
+ 430438.400000ns, VSS,
+ 430438.500000ns, VDD,
+ 430918.800000ns, VDD,
+ 430918.900000ns, VSS,
+ 431038.900000ns, VSS,
+ 431039.000000ns, VDD,
+ 431759.500000ns, VDD,
+ 431759.600000ns, VSS,
+ 432600.200000ns, VSS,
+ 432600.300000ns, VDD,
+ 432840.400000ns, VDD,
+ 432840.500000ns, VSS,
+ 433080.600000ns, VSS,
+ 433080.700000ns, VDD,
+ 433320.800000ns, VDD,
+ 433320.900000ns, VSS,
+ 433561.000000ns, VSS,
+ 433561.100000ns, VDD,
+ 434041.400000ns, VDD,
+ 434041.500000ns, VSS,
+ 436683.600000ns, VSS,
+ 436683.700000ns, VDD,
+ 437644.400000ns, VDD,
+ 437644.500000ns, VSS,
+ 438965.500000ns, VSS,
+ 438965.600000ns, VDD,
+ 439445.900000ns, VDD,
+ 439446.000000ns, VSS,
+ 440406.700000ns, VSS,
+ 440406.800000ns, VDD,
+ 440887.100000ns, VDD,
+ 440887.200000ns, VSS,
+ 441127.300000ns, VSS,
+ 441127.400000ns, VDD,
+ 441247.400000ns, VDD,
+ 441247.500000ns, VSS,
+ 441487.600000ns, VSS,
+ 441487.700000ns, VDD,
+ 441607.700000ns, VDD,
+ 441607.800000ns, VSS,
+ 442568.500000ns, VSS,
+ 442568.600000ns, VDD,
+ 442808.700000ns, VDD,
+ 442808.800000ns, VSS,
+ 444970.500000ns, VSS,
+ 444970.600000ns, VDD,
+ 446411.700000ns, VDD,
+ 446411.800000ns, VSS,
+ 446892.100000ns, VSS,
+ 446892.200000ns, VDD,
+ 447492.600000ns, VDD,
+ 447492.700000ns, VSS,
+ 447852.900000ns, VSS,
+ 447853.000000ns, VDD,
+ 448333.300000ns, VDD,
+ 448333.400000ns, VSS,
+ 448573.500000ns, VSS,
+ 448573.600000ns, VDD,
+ 448933.800000ns, VDD,
+ 448933.900000ns, VSS,
+ 449894.600000ns, VSS,
+ 449894.700000ns, VDD,
+ 450134.800000ns, VDD,
+ 450134.900000ns, VSS,
+ 450855.400000ns, VSS,
+ 450855.500000ns, VDD,
+ 450975.500000ns, VDD,
+ 450975.600000ns, VSS,
+ 451335.800000ns, VSS,
+ 451335.900000ns, VDD,
+ 451576.000000ns, VDD,
+ 451576.100000ns, VSS,
+ 452296.600000ns, VSS,
+ 452296.700000ns, VDD,
+ 452777.000000ns, VDD,
+ 452777.100000ns, VSS,
+ 453137.300000ns, VSS,
+ 453137.400000ns, VDD,
+ 453377.500000ns, VDD,
+ 453377.600000ns, VSS,
+ 453978.000000ns, VSS,
+ 453978.100000ns, VDD,
+ 455058.900000ns, VDD,
+ 455059.000000ns, VSS,
+ 455659.400000ns, VSS,
+ 455659.500000ns, VDD,
+ 455899.600000ns, VDD,
+ 455899.700000ns, VSS,
+ 456019.700000ns, VSS,
+ 456019.800000ns, VDD,
+ 456259.900000ns, VDD,
+ 456260.000000ns, VSS,
+ 456740.300000ns, VSS,
+ 456740.400000ns, VDD,
+ 456980.500000ns, VDD,
+ 456980.600000ns, VSS,
+ 457220.700000ns, VSS,
+ 457220.800000ns, VDD,
+ 460463.400000ns, VDD,
+ 460463.500000ns, VSS,
+ 460943.800000ns, VSS,
+ 460943.900000ns, VDD,
+ 463105.600000ns, VDD,
+ 463105.700000ns, VSS,
+ 463586.000000ns, VSS,
+ 463586.100000ns, VDD,
+ 464066.400000ns, VDD,
+ 464066.500000ns, VSS,
+ 464907.100000ns, VSS,
+ 464907.200000ns, VDD,
+ 465627.700000ns, VDD,
+ 465627.800000ns, VSS,
+ 466228.200000ns, VSS,
+ 466228.300000ns, VDD,
+ 466468.400000ns, VDD,
+ 466468.500000ns, VSS,
+ 466948.800000ns, VSS,
+ 466948.900000ns, VDD,
+ 467189.000000ns, VDD,
+ 467189.100000ns, VSS,
+ 467429.200000ns, VSS,
+ 467429.300000ns, VDD,
+ 467789.500000ns, VDD,
+ 467789.600000ns, VSS,
+ 467909.600000ns, VSS,
+ 467909.700000ns, VDD,
+ 468029.700000ns, VDD,
+ 468029.800000ns, VSS,
+ 468750.300000ns, VSS,
+ 468750.400000ns, VDD,
+ 468870.400000ns, VDD,
+ 468870.500000ns, VSS,
+ 470912.100000ns, VSS,
+ 470912.200000ns, VDD,
+ 471632.700000ns, VDD,
+ 471632.800000ns, VSS,
+ 472113.100000ns, VSS,
+ 472113.200000ns, VDD,
+ 472593.500000ns, VDD,
+ 472593.600000ns, VSS,
+ 472713.600000ns, VSS,
+ 472713.700000ns, VDD,
+ 473194.000000ns, VDD,
+ 473194.100000ns, VSS,
+ 473674.400000ns, VSS,
+ 473674.500000ns, VDD,
+ 475115.600000ns, VDD,
+ 475115.700000ns, VSS,
+ 475235.700000ns, VSS,
+ 475235.800000ns, VDD,
+ 475475.900000ns, VDD,
+ 475476.000000ns, VSS,
+ 475596.000000ns, VSS,
+ 475596.100000ns, VDD,
+ 476076.400000ns, VDD,
+ 476076.500000ns, VSS,
+ 476316.600000ns, VSS,
+ 476316.700000ns, VDD,
+ 477037.200000ns, VDD,
+ 477037.300000ns, VSS,
+ 477157.300000ns, VSS,
+ 477157.400000ns, VDD,
+ 477277.400000ns, VDD,
+ 477277.500000ns, VSS,
+ 477757.800000ns, VSS,
+ 477757.900000ns, VDD,
+ 478478.400000ns, VDD,
+ 478478.500000ns, VSS,
+ 478598.500000ns, VSS,
+ 478598.600000ns, VDD,
+ 479919.600000ns, VDD,
+ 479919.700000ns, VSS,
+ 480039.700000ns, VSS,
+ 480039.800000ns, VDD,
+ 480760.300000ns, VDD,
+ 480760.400000ns, VSS,
+ 481480.900000ns, VSS,
+ 481481.000000ns, VDD,
+ 481841.200000ns, VDD,
+ 481841.300000ns, VSS,
+ 481961.300000ns, VSS,
+ 481961.400000ns, VDD,
+ 482561.800000ns, VDD,
+ 482561.900000ns, VSS,
+ 483042.200000ns, VSS,
+ 483042.300000ns, VDD,
+ 484363.300000ns, VDD,
+ 484363.400000ns, VSS,
+ 484963.800000ns, VSS,
+ 484963.900000ns, VDD,
+ 485204.000000ns, VDD,
+ 485204.100000ns, VSS,
+ 485324.100000ns, VSS,
+ 485324.200000ns, VDD,
+ 485804.500000ns, VDD,
+ 485804.600000ns, VSS,
+ 486645.200000ns, VSS,
+ 486645.300000ns, VDD,
+ 486765.300000ns, VDD,
+ 486765.400000ns, VSS,
+ 487726.100000ns, VSS,
+ 487726.200000ns, VDD,
+ 487966.300000ns, VDD,
+ 487966.400000ns, VSS,
+ 488086.400000ns, VSS,
+ 488086.500000ns, VDD,
+ 488446.700000ns, VDD,
+ 488446.800000ns, VSS,
+ 488566.800000ns, VSS,
+ 488566.900000ns, VDD,
+ 488927.100000ns, VDD,
+ 488927.200000ns, VSS,
+ 490008.000000ns, VSS,
+ 490008.100000ns, VDD,
+ 490368.300000ns, VDD,
+ 490368.400000ns, VSS,
+ 490728.600000ns, VSS,
+ 490728.700000ns, VDD,
+ 492049.700000ns, VDD,
+ 492049.800000ns, VSS,
+ 492650.200000ns, VSS,
+ 492650.300000ns, VDD,
+ 493010.500000ns, VDD,
+ 493010.600000ns, VSS,
+ 493611.000000ns, VSS,
+ 493611.100000ns, VDD,
+ 493851.200000ns, VDD,
+ 493851.300000ns, VSS,
+ 494451.700000ns, VSS,
+ 494451.800000ns, VDD,
+ 496133.100000ns, VDD,
+ 496133.200000ns, VSS,
+ 496733.600000ns, VSS,
+ 496733.700000ns, VDD,
+ 496973.800000ns, VDD,
+ 496973.900000ns, VSS,
+ 497093.900000ns, VSS,
+ 497094.000000ns, VDD,
+ 497214.000000ns, VDD,
+ 497214.100000ns, VSS,
+ 497454.200000ns, VSS,
+ 497454.300000ns, VDD,
+ 497574.300000ns, VDD,
+ 497574.400000ns, VSS,
+ 498294.900000ns, VSS,
+ 498295.000000ns, VDD,
+ 499135.600000ns, VDD,
+ 499135.700000ns, VSS,
+ 499736.100000ns, VSS,
+ 499736.200000ns, VDD,
+ 501417.500000ns, VDD,
+ 501417.600000ns, VSS,
+ 502018.000000ns, VSS,
+ 502018.100000ns, VDD,
+ 502978.800000ns, VDD,
+ 502978.900000ns, VSS,
+ 503459.200000ns, VSS,
+ 503459.300000ns, VDD,
+ 503579.300000ns, VDD,
+ 503579.400000ns, VSS,
+ 503819.500000ns, VSS,
+ 503819.600000ns, VDD,
+ 504059.700000ns, VDD,
+ 504059.800000ns, VSS,
+ 505260.700000ns, VSS,
+ 505260.800000ns, VDD,
+ 506101.400000ns, VDD,
+ 506101.500000ns, VSS,
+ 506221.500000ns, VSS,
+ 506221.600000ns, VDD,
+ 506581.800000ns, VDD,
+ 506581.900000ns, VSS,
+ 507062.200000ns, VSS,
+ 507062.300000ns, VDD,
+ 507662.700000ns, VDD,
+ 507662.800000ns, VSS,
+ 507782.800000ns, VSS,
+ 507782.900000ns, VDD,
+ 508143.100000ns, VDD,
+ 508143.200000ns, VSS,
+ 508503.400000ns, VSS,
+ 508503.500000ns, VDD,
+ 508743.600000ns, VDD,
+ 508743.700000ns, VSS,
+ 510184.800000ns, VSS,
+ 510184.900000ns, VDD,
+ 511986.300000ns, VDD,
+ 511986.400000ns, VSS,
+ 512947.100000ns, VSS,
+ 512947.200000ns, VDD,
+ 513547.600000ns, VDD,
+ 513547.700000ns, VSS,
+ 513787.800000ns, VSS,
+ 513787.900000ns, VDD,
+ 513907.900000ns, VDD,
+ 513908.000000ns, VSS,
+ 515349.100000ns, VSS,
+ 515349.200000ns, VDD,
+ 517270.700000ns, VDD,
+ 517270.800000ns, VSS,
+ 517390.800000ns, VSS,
+ 517390.900000ns, VDD,
+ 518111.400000ns, VDD,
+ 518111.500000ns, VSS,
+ 518471.700000ns, VSS,
+ 518471.800000ns, VDD,
+ 518591.800000ns, VDD,
+ 518591.900000ns, VSS,
+ 518711.900000ns, VSS,
+ 518712.000000ns, VDD,
+ 518952.100000ns, VDD,
+ 518952.200000ns, VSS,
+ 519912.900000ns, VSS,
+ 519913.000000ns, VDD,
+ 520033.000000ns, VDD,
+ 520033.100000ns, VSS,
+ 520753.600000ns, VSS,
+ 520753.700000ns, VDD,
+ 522314.900000ns, VDD,
+ 522315.000000ns, VSS,
+ 522435.000000ns, VSS,
+ 522435.100000ns, VDD,
+ 523515.900000ns, VDD,
+ 523516.000000ns, VSS,
+ 523996.300000ns, VSS,
+ 523996.400000ns, VDD,
+ 525077.200000ns, VDD,
+ 525077.300000ns, VSS,
+ 525197.300000ns, VSS,
+ 525197.400000ns, VDD,
+ 525677.700000ns, VDD,
+ 525677.800000ns, VSS,
+ 526998.800000ns, VSS,
+ 526998.900000ns, VDD,
+ 528079.700000ns, VDD,
+ 528079.800000ns, VSS,
+ 528199.800000ns, VSS,
+ 528199.900000ns, VDD,
+ 528800.300000ns, VDD,
+ 528800.400000ns, VSS,
+ 529400.800000ns, VSS,
+ 529400.900000ns, VDD,
+ 530121.400000ns, VDD,
+ 530121.500000ns, VSS,
+ 530601.800000ns, VSS,
+ 530601.900000ns, VDD,
+ 530721.900000ns, VDD,
+ 530722.000000ns, VSS,
+ 531082.200000ns, VSS,
+ 531082.300000ns, VDD,
+ 531562.600000ns, VDD,
+ 531562.700000ns, VSS,
+ 531682.700000ns, VSS,
+ 531682.800000ns, VDD,
+ 532643.500000ns, VDD,
+ 532643.600000ns, VSS,
+ 533123.900000ns, VSS,
+ 533124.000000ns, VDD,
+ 534084.700000ns, VDD,
+ 534084.800000ns, VSS,
+ 534324.900000ns, VSS,
+ 534325.000000ns, VDD,
+ 536967.100000ns, VDD,
+ 536967.200000ns, VSS,
+ 537447.500000ns, VSS,
+ 537447.600000ns, VDD,
+ 538648.500000ns, VDD,
+ 538648.600000ns, VSS,
+ 539128.900000ns, VSS,
+ 539129.000000ns, VDD,
+ 539849.500000ns, VDD,
+ 539849.600000ns, VSS,
+ 539969.600000ns, VSS,
+ 539969.700000ns, VDD,
+ 540690.200000ns, VDD,
+ 540690.300000ns, VSS,
+ 541891.200000ns, VSS,
+ 541891.300000ns, VDD,
+ 543692.700000ns, VDD,
+ 543692.800000ns, VSS,
+ 545854.500000ns, VSS,
+ 545854.600000ns, VDD,
+ 546334.900000ns, VDD,
+ 546335.000000ns, VSS,
+ 546575.100000ns, VSS,
+ 546575.200000ns, VDD,
+ 548376.600000ns, VDD,
+ 548376.700000ns, VSS,
+ 548616.800000ns, VSS,
+ 548616.900000ns, VDD,
+ 548736.900000ns, VDD,
+ 548737.000000ns, VSS,
+ 549817.800000ns, VSS,
+ 549817.900000ns, VDD,
+ 550418.300000ns, VDD,
+ 550418.400000ns, VSS,
+ 551619.300000ns, VSS,
+ 551619.400000ns, VDD,
+ 552099.700000ns, VDD,
+ 552099.800000ns, VSS,
+ 552219.800000ns, VSS,
+ 552219.900000ns, VDD,
+ 553420.800000ns, VDD,
+ 553420.900000ns, VSS,
+ 553661.000000ns, VSS,
+ 553661.100000ns, VDD,
+ 555462.500000ns, VDD,
+ 555462.600000ns, VSS,
+ 555822.800000ns, VSS,
+ 555822.900000ns, VDD,
+ 556663.500000ns, VDD,
+ 556663.600000ns, VSS,
+ 557023.800000ns, VSS,
+ 557023.900000ns, VDD,
+ 557624.300000ns, VDD,
+ 557624.400000ns, VSS,
+ 558104.700000ns, VSS,
+ 558104.800000ns, VDD,
+ 558344.900000ns, VDD,
+ 558345.000000ns, VSS,
+ 558825.300000ns, VSS,
+ 558825.400000ns, VDD,
+ 559065.500000ns, VDD,
+ 559065.600000ns, VSS,
+ 559545.900000ns, VSS,
+ 559546.000000ns, VDD,
+ 560386.600000ns, VDD,
+ 560386.700000ns, VSS,
+ 560506.700000ns, VSS,
+ 560506.800000ns, VDD,
+ 560626.800000ns, VDD,
+ 560626.900000ns, VSS,
+ 560867.000000ns, VSS,
+ 560867.100000ns, VDD,
+ 562548.400000ns, VDD,
+ 562548.500000ns, VSS,
+ 563389.100000ns, VSS,
+ 563389.200000ns, VDD,
+ 565070.500000ns, VDD,
+ 565070.600000ns, VSS,
+ 565190.600000ns, VSS,
+ 565190.700000ns, VDD,
+ 565310.700000ns, VDD,
+ 565310.800000ns, VSS,
+ 566031.300000ns, VSS,
+ 566031.400000ns, VDD,
+ 566511.700000ns, VDD,
+ 566511.800000ns, VSS,
+ 568193.100000ns, VSS,
+ 568193.200000ns, VDD,
+ 569153.900000ns, VDD,
+ 569154.000000ns, VSS,
+ 569274.000000ns, VSS,
+ 569274.100000ns, VDD,
+ 570475.000000ns, VDD,
+ 570475.100000ns, VSS,
+ 570835.300000ns, VSS,
+ 570835.400000ns, VDD,
+ 571075.500000ns, VDD,
+ 571075.600000ns, VSS,
+ 571195.600000ns, VSS,
+ 571195.700000ns, VDD,
+ 571435.800000ns, VDD,
+ 571435.900000ns, VSS,
+ 572877.000000ns, VSS,
+ 572877.100000ns, VDD,
+ 575519.200000ns, VDD,
+ 575519.300000ns, VSS,
+ 575639.300000ns, VSS,
+ 575639.400000ns, VDD,
+ 575759.400000ns, VDD,
+ 575759.500000ns, VSS,
+ 576480.000000ns, VSS,
+ 576480.100000ns, VDD,
+ 576600.100000ns, VDD,
+ 576600.200000ns, VSS,
+ 576960.400000ns, VSS,
+ 576960.500000ns, VDD,
+ 577080.500000ns, VDD,
+ 577080.600000ns, VSS,
+ 577200.600000ns, VSS,
+ 577200.700000ns, VDD,
+ 577681.000000ns, VDD,
+ 577681.100000ns, VSS,
+ 578161.400000ns, VSS,
+ 578161.500000ns, VDD,
+ 578761.900000ns, VDD,
+ 578762.000000ns, VSS,
+ 578882.000000ns, VSS,
+ 578882.100000ns, VDD,
+ 579362.400000ns, VDD,
+ 579362.500000ns, VSS,
+ 580443.300000ns, VSS,
+ 580443.400000ns, VDD,
+ 581043.800000ns, VDD,
+ 581043.900000ns, VSS,
+ 581163.900000ns, VSS,
+ 581164.000000ns, VDD,
+ 581884.500000ns, VDD,
+ 581884.600000ns, VSS,
+ 582364.900000ns, VSS,
+ 582365.000000ns, VDD,
+ 582845.300000ns, VDD,
+ 582845.400000ns, VSS,
+ 583085.500000ns, VSS,
+ 583085.600000ns, VDD,
+ 583686.000000ns, VDD,
+ 583686.100000ns, VSS,
+ 583806.100000ns, VSS,
+ 583806.200000ns, VDD,
+ 583926.200000ns, VDD,
+ 583926.300000ns, VSS,
+ 585247.300000ns, VSS,
+ 585247.400000ns, VDD,
+ 585487.500000ns, VDD,
+ 585487.600000ns, VSS,
+ 585847.800000ns, VSS,
+ 585847.900000ns, VDD,
+ 586088.000000ns, VDD,
+ 586088.100000ns, VSS,
+ 586208.100000ns, VSS,
+ 586208.200000ns, VDD,
+ 586808.600000ns, VDD,
+ 586808.700000ns, VSS,
+ 587409.100000ns, VSS,
+ 587409.200000ns, VDD,
+ 587529.200000ns, VDD,
+ 587529.300000ns, VSS,
+ 587769.400000ns, VSS,
+ 587769.500000ns, VDD,
+ 588249.800000ns, VDD,
+ 588249.900000ns, VSS,
+ 589090.500000ns, VSS,
+ 589090.600000ns, VDD,
+ 589691.000000ns, VDD,
+ 589691.100000ns, VSS,
+ 589931.200000ns, VSS,
+ 589931.300000ns, VDD,
+ 590771.900000ns, VDD,
+ 590772.000000ns, VSS,
+ 591012.100000ns, VSS,
+ 591012.200000ns, VDD,
+ 591132.200000ns, VDD,
+ 591132.300000ns, VSS,
+ 592093.000000ns, VSS,
+ 592093.100000ns, VDD,
+ 592453.300000ns, VDD,
+ 592453.400000ns, VSS,
+ 593294.000000ns, VSS,
+ 593294.100000ns, VDD,
+ 594855.300000ns, VDD,
+ 594855.400000ns, VSS,
+ 595936.200000ns, VSS,
+ 595936.300000ns, VDD,
+ 596656.800000ns, VDD,
+ 596656.900000ns, VSS,
+ 596776.900000ns, VSS,
+ 596777.000000ns, VDD,
+ 597017.100000ns, VDD,
+ 597017.200000ns, VSS,
+ 597257.300000ns, VSS,
+ 597257.400000ns, VDD,
+ 598818.600000ns, VDD,
+ 598818.700000ns, VSS,
+ 599779.400000ns, VSS,
+ 599779.500000ns, VDD,
+ 600500.000000ns, VDD,
+ 600500.100000ns, VSS,
+ 601100.500000ns, VSS,
+ 601100.600000ns, VDD,
+ 602061.300000ns, VDD,
+ 602061.400000ns, VSS,
+ 602301.500000ns, VSS,
+ 602301.600000ns, VDD,
+ 602421.600000ns, VDD,
+ 602421.700000ns, VSS,
+ 603382.400000ns, VSS,
+ 603382.500000ns, VDD,
+ 603502.500000ns, VDD,
+ 603502.600000ns, VSS,
+ 603982.900000ns, VSS,
+ 603983.000000ns, VDD,
+ 605784.400000ns, VDD,
+ 605784.500000ns, VSS,
+ 608066.300000ns, VSS,
+ 608066.400000ns, VDD,
+ 608306.500000ns, VDD,
+ 608306.600000ns, VSS,
+ 609027.100000ns, VSS,
+ 609027.200000ns, VDD,
+ 609267.300000ns, VDD,
+ 609267.400000ns, VSS,
+ 610348.200000ns, VSS,
+ 610348.300000ns, VDD,
+ 610828.600000ns, VDD,
+ 610828.700000ns, VSS,
+ 611549.200000ns, VSS,
+ 611549.300000ns, VDD,
+ 612750.200000ns, VDD,
+ 612750.300000ns, VSS,
+ 613350.700000ns, VSS,
+ 613350.800000ns, VDD,
+ 613951.200000ns, VDD,
+ 613951.300000ns, VSS,
+ 614912.000000ns, VSS,
+ 614912.100000ns, VDD,
+ 615872.800000ns, VDD,
+ 615872.900000ns, VSS,
+ 615992.900000ns, VSS,
+ 615993.000000ns, VDD,
+ 616473.300000ns, VDD,
+ 616473.400000ns, VSS,
+ 617554.200000ns, VSS,
+ 617554.300000ns, VDD,
+ 618034.600000ns, VDD,
+ 618034.700000ns, VSS,
+ 618875.300000ns, VSS,
+ 618875.400000ns, VDD,
+ 621877.800000ns, VDD,
+ 621877.900000ns, VSS,
+ 622118.000000ns, VSS,
+ 622118.100000ns, VDD,
+ 622958.700000ns, VDD,
+ 622958.800000ns, VSS,
+ 624039.600000ns, VSS,
+ 624039.700000ns, VDD,
+ 624159.700000ns, VDD,
+ 624159.800000ns, VSS,
+ 625120.500000ns, VSS,
+ 625120.600000ns, VDD,
+ 626201.400000ns, VDD,
+ 626201.500000ns, VSS,
+ 626922.000000ns, VSS,
+ 626922.100000ns, VDD,
+ 627882.800000ns, VDD,
+ 627882.900000ns, VSS,
+ 628723.500000ns, VSS,
+ 628723.600000ns, VDD,
+ 628963.700000ns, VDD,
+ 628963.800000ns, VSS,
+ 630525.000000ns, VSS,
+ 630525.100000ns, VDD,
+ 630885.300000ns, VDD,
+ 630885.400000ns, VSS,
+ 631125.500000ns, VSS,
+ 631125.600000ns, VDD,
+ 631605.900000ns, VDD,
+ 631606.000000ns, VSS,
+ 631726.000000ns, VSS,
+ 631726.100000ns, VDD,
+ 631846.100000ns, VDD,
+ 631846.200000ns, VSS,
+ 632086.300000ns, VSS,
+ 632086.400000ns, VDD,
+ 632206.400000ns, VDD,
+ 632206.500000ns, VSS,
+ 632686.800000ns, VSS,
+ 632686.900000ns, VDD,
+ 633887.800000ns, VDD,
+ 633887.900000ns, VSS,
+ 634728.500000ns, VSS,
+ 634728.600000ns, VDD,
+ 635449.100000ns, VDD,
+ 635449.200000ns, VSS,
+ 636169.700000ns, VSS,
+ 636169.800000ns, VDD,
+ 636650.100000ns, VDD,
+ 636650.200000ns, VSS,
+ 637010.400000ns, VSS,
+ 637010.500000ns, VDD,
+ 637490.800000ns, VDD,
+ 637490.900000ns, VSS,
+ 637971.200000ns, VSS,
+ 637971.300000ns, VDD,
+ 638451.600000ns, VDD,
+ 638451.700000ns, VSS,
+ 639292.300000ns, VSS,
+ 639292.400000ns, VDD,
+ 639412.400000ns, VDD,
+ 639412.500000ns, VSS,
+ 642895.300000ns, VSS,
+ 642895.400000ns, VDD,
+ 643736.000000ns, VDD,
+ 643736.100000ns, VSS,
+ 643856.100000ns, VSS,
+ 643856.200000ns, VDD,
+ 643976.200000ns, VDD,
+ 643976.300000ns, VSS,
+ 644216.400000ns, VSS,
+ 644216.500000ns, VDD,
+ 644336.500000ns, VDD,
+ 644336.600000ns, VSS,
+ 644816.900000ns, VSS,
+ 644817.000000ns, VDD,
+ 645297.300000ns, VDD,
+ 645297.400000ns, VSS,
+ 646618.400000ns, VSS,
+ 646618.500000ns, VDD,
+ 646978.700000ns, VDD,
+ 646978.800000ns, VSS,
+ 647218.900000ns, VSS,
+ 647219.000000ns, VDD,
+ 649741.000000ns, VDD,
+ 649741.100000ns, VSS,
+ 650341.500000ns, VSS,
+ 650341.600000ns, VDD,
+ 650701.800000ns, VDD,
+ 650701.900000ns, VSS,
+ 651782.700000ns, VSS,
+ 651782.800000ns, VDD,
+ 652623.400000ns, VDD,
+ 652623.500000ns, VSS,
+ 653103.800000ns, VSS,
+ 653103.900000ns, VDD,
+ 653704.300000ns, VDD,
+ 653704.400000ns, VSS,
+ 653944.500000ns, VSS,
+ 653944.600000ns, VDD,
+ 654785.200000ns, VDD,
+ 654785.300000ns, VSS,
+ 654905.300000ns, VSS,
+ 654905.400000ns, VDD,
+ 655025.400000ns, VDD,
+ 655025.500000ns, VSS,
+ 656106.300000ns, VSS,
+ 656106.400000ns, VDD,
+ 657547.500000ns, VDD,
+ 657547.600000ns, VSS,
+ 657787.700000ns, VSS,
+ 657787.800000ns, VDD,
+ 658628.400000ns, VDD,
+ 658628.500000ns, VSS,
+ 659829.400000ns, VSS,
+ 659829.500000ns, VDD,
+ 660189.700000ns, VDD,
+ 660189.800000ns, VSS,
+ 661030.400000ns, VSS,
+ 661030.500000ns, VDD,
+ 661270.600000ns, VDD,
+ 661270.700000ns, VSS,
+ 662231.400000ns, VSS,
+ 662231.500000ns, VDD,
+ 662831.900000ns, VDD,
+ 662832.000000ns, VSS,
+ 663072.100000ns, VSS,
+ 663072.200000ns, VDD,
+ 663552.500000ns, VDD,
+ 663552.600000ns, VSS,
+ 664513.300000ns, VSS,
+ 664513.400000ns, VDD,
+ 664753.500000ns, VDD,
+ 664753.600000ns, VSS,
+ 665594.200000ns, VSS,
+ 665594.300000ns, VDD,
+ 665954.500000ns, VDD,
+ 665954.600000ns, VSS,
+ 666675.100000ns, VSS,
+ 666675.200000ns, VDD,
+ 667035.400000ns, VDD,
+ 667035.500000ns, VSS,
+ 668716.800000ns, VSS,
+ 668716.900000ns, VDD,
+ 669677.600000ns, VDD,
+ 669677.700000ns, VSS,
+ 670398.200000ns, VSS,
+ 670398.300000ns, VDD,
+ 670998.700000ns, VDD,
+ 670998.800000ns, VSS,
+ 671359.000000ns, VSS,
+ 671359.100000ns, VDD,
+ 671479.100000ns, VDD,
+ 671479.200000ns, VSS,
+ 672079.600000ns, VSS,
+ 672079.700000ns, VDD,
+ 673280.600000ns, VDD,
+ 673280.700000ns, VSS,
+ 673520.800000ns, VSS,
+ 673520.900000ns, VDD,
+ 673761.000000ns, VDD,
+ 673761.100000ns, VSS,
+ 674241.400000ns, VSS,
+ 674241.500000ns, VDD,
+ 675562.500000ns, VDD,
+ 675562.600000ns, VSS,
+ 675802.700000ns, VSS,
+ 675802.800000ns, VDD,
+ 675922.800000ns, VDD,
+ 675922.900000ns, VSS,
+ 676283.100000ns, VSS,
+ 676283.200000ns, VDD,
+ 677484.100000ns, VDD,
+ 677484.200000ns, VSS,
+ 678084.600000ns, VSS,
+ 678084.700000ns, VDD,
+ 681807.700000ns, VDD,
+ 681807.800000ns, VSS,
+ 682288.100000ns, VSS,
+ 682288.200000ns, VDD,
+ 683128.800000ns, VDD,
+ 683128.900000ns, VSS,
+ 683609.200000ns, VSS,
+ 683609.300000ns, VDD,
+ 685530.800000ns, VDD,
+ 685530.900000ns, VSS,
+ 685891.100000ns, VSS,
+ 685891.200000ns, VDD,
+ 686131.300000ns, VDD,
+ 686131.400000ns, VSS,
+ 686731.800000ns, VSS,
+ 686731.900000ns, VDD,
+ 687092.100000ns, VDD,
+ 687092.200000ns, VSS,
+ 687212.200000ns, VSS,
+ 687212.300000ns, VDD,
+ 687932.800000ns, VDD,
+ 687932.900000ns, VSS,
+ 688173.000000ns, VSS,
+ 688173.100000ns, VDD,
+ 688293.100000ns, VDD,
+ 688293.200000ns, VSS,
+ 688653.400000ns, VSS,
+ 688653.500000ns, VDD,
+ 689013.700000ns, VDD,
+ 689013.800000ns, VSS,
+ 689374.000000ns, VSS,
+ 689374.100000ns, VDD,
+ 689974.500000ns, VDD,
+ 689974.600000ns, VSS,
+ 690094.600000ns, VSS,
+ 690094.700000ns, VDD,
+ 690575.000000ns, VDD,
+ 690575.100000ns, VSS,
+ 691776.000000ns, VSS,
+ 691776.100000ns, VDD,
+ 692256.400000ns, VDD,
+ 692256.500000ns, VSS,
+ 692736.800000ns, VSS,
+ 692736.900000ns, VDD,
+ 693217.200000ns, VDD,
+ 693217.300000ns, VSS,
+ 693337.300000ns, VSS,
+ 693337.400000ns, VDD,
+ 693457.400000ns, VDD,
+ 693457.500000ns, VSS,
+ 693697.600000ns, VSS,
+ 693697.700000ns, VDD,
+ 693937.800000ns, VDD,
+ 693937.900000ns, VSS,
+ 694178.000000ns, VSS,
+ 694178.100000ns, VDD,
+ 694298.100000ns, VDD,
+ 694298.200000ns, VSS,
+ 694418.200000ns, VSS,
+ 694418.300000ns, VDD,
+ 695258.900000ns, VDD,
+ 695259.000000ns, VSS,
+ 695379.000000ns, VSS,
+ 695379.100000ns, VDD,
+ 696219.700000ns, VDD,
+ 696219.800000ns, VSS,
+ 696700.100000ns, VSS,
+ 696700.200000ns, VDD,
+ 697300.600000ns, VDD,
+ 697300.700000ns, VSS,
+ 697420.700000ns, VSS,
+ 697420.800000ns, VDD,
+ 697540.800000ns, VDD,
+ 697540.900000ns, VSS,
+ 698501.600000ns, VSS,
+ 698501.700000ns, VDD,
+ 698621.700000ns, VDD,
+ 698621.800000ns, VSS,
+ 698982.000000ns, VSS,
+ 698982.100000ns, VDD,
+ 699342.300000ns, VDD,
+ 699342.400000ns, VSS,
+ 699822.700000ns, VSS,
+ 699822.800000ns, VDD,
+ 701504.100000ns, VDD,
+ 701504.200000ns, VSS,
+ 702464.900000ns, VSS,
+ 702465.000000ns, VDD,
+ 703305.600000ns, VDD,
+ 703305.700000ns, VSS,
+ 705467.400000ns, VSS,
+ 705467.500000ns, VDD,
+ 707148.800000ns, VDD,
+ 707148.900000ns, VSS,
+ 709070.400000ns, VSS,
+ 709070.500000ns, VDD,
+ 711112.100000ns, VDD,
+ 711112.200000ns, VSS,
+ 711952.800000ns, VSS,
+ 711952.900000ns, VDD,
+ 713153.800000ns, VDD,
+ 713153.900000ns, VSS,
+ 715435.700000ns, VSS,
+ 715435.800000ns, VDD,
+ 715916.100000ns, VDD,
+ 715916.200000ns, VSS,
+ 716516.600000ns, VSS,
+ 716516.700000ns, VDD,
+ 717957.800000ns, VDD,
+ 717957.900000ns, VSS,
+ 718077.900000ns, VSS,
+ 718078.000000ns, VDD,
+ 718198.000000ns, VDD,
+ 718198.100000ns, VSS,
+ 719879.400000ns, VSS,
+ 719879.500000ns, VDD,
+ 720119.600000ns, VDD,
+ 720119.700000ns, VSS,
+ 720239.700000ns, VSS,
+ 720239.800000ns, VDD,
+ 720359.800000ns, VDD,
+ 720359.900000ns, VSS,
+ 720600.000000ns, VSS,
+ 720600.100000ns, VDD,
+ 721921.100000ns, VDD,
+ 721921.200000ns, VSS,
+ 722401.500000ns, VSS,
+ 722401.600000ns, VDD,
+ 722521.600000ns, VDD,
+ 722521.700000ns, VSS,
+ 722881.900000ns, VSS,
+ 722882.000000ns, VDD,
+ 723362.300000ns, VDD,
+ 723362.400000ns, VSS,
+ 724082.900000ns, VSS,
+ 724083.000000ns, VDD,
+ 725163.800000ns, VDD,
+ 725163.900000ns, VSS,
+ 726725.100000ns, VSS,
+ 726725.200000ns, VDD,
+ 727325.600000ns, VDD,
+ 727325.700000ns, VSS,
+ 727806.000000ns, VSS,
+ 727806.100000ns, VDD,
+ 728046.200000ns, VDD,
+ 728046.300000ns, VSS,
+ 728166.300000ns, VSS,
+ 728166.400000ns, VDD,
+ 729007.000000ns, VDD,
+ 729007.100000ns, VSS,
+ 729967.800000ns, VSS,
+ 729967.900000ns, VDD,
+ 730568.300000ns, VDD,
+ 730568.400000ns, VSS,
+ 730928.600000ns, VSS,
+ 730928.700000ns, VDD,
+ 731048.700000ns, VDD,
+ 731048.800000ns, VSS,
+ 731409.000000ns, VSS,
+ 731409.100000ns, VDD,
+ 732249.700000ns, VDD,
+ 732249.800000ns, VSS,
+ 732489.900000ns, VSS,
+ 732490.000000ns, VDD,
+ 732970.300000ns, VDD,
+ 732970.400000ns, VSS,
+ 733210.500000ns, VSS,
+ 733210.600000ns, VDD,
+ 733330.600000ns, VDD,
+ 733330.700000ns, VSS,
+ 735492.400000ns, VSS,
+ 735492.500000ns, VDD,
+ 735732.600000ns, VDD,
+ 735732.700000ns, VSS,
+ 736573.300000ns, VSS,
+ 736573.400000ns, VDD,
+ 737053.700000ns, VDD,
+ 737053.800000ns, VSS,
+ 737534.100000ns, VSS,
+ 737534.200000ns, VDD,
+ 738615.000000ns, VDD,
+ 738615.100000ns, VSS,
+ 738855.200000ns, VSS,
+ 738855.300000ns, VDD,
+ 739215.500000ns, VDD,
+ 739215.600000ns, VSS,
+ 739455.700000ns, VSS,
+ 739455.800000ns, VDD,
+ 740176.300000ns, VDD,
+ 740176.400000ns, VSS,
+ 741377.300000ns, VSS,
+ 741377.400000ns, VDD,
+ 741617.500000ns, VDD,
+ 741617.600000ns, VSS,
+ 742458.200000ns, VSS,
+ 742458.300000ns, VDD,
+ 743058.700000ns, VDD,
+ 743058.800000ns, VSS,
+ 744620.000000ns, VSS,
+ 744620.100000ns, VDD,
+ 746301.400000ns, VDD,
+ 746301.500000ns, VSS,
+ 747262.200000ns, VSS,
+ 747262.300000ns, VDD,
+ 747622.500000ns, VDD,
+ 747622.600000ns, VSS,
+ 748102.900000ns, VSS,
+ 748103.000000ns, VDD,
+ 748583.300000ns, VDD,
+ 748583.400000ns, VSS,
+ 750504.900000ns, VSS,
+ 750505.000000ns, VDD,
+ 751585.800000ns, VDD,
+ 751585.900000ns, VSS,
+ 752666.700000ns, VSS,
+ 752666.800000ns, VDD,
+ 752786.800000ns, VDD,
+ 752786.900000ns, VSS,
+ 752906.900000ns, VSS,
+ 752907.000000ns, VDD,
+ 753747.600000ns, VDD,
+ 753747.700000ns, VSS,
+ 755308.900000ns, VSS,
+ 755309.000000ns, VDD,
+ 756750.100000ns, VDD,
+ 756750.200000ns, VSS,
+ 757350.600000ns, VSS,
+ 757350.700000ns, VDD,
+ 757470.700000ns, VDD,
+ 757470.800000ns, VSS,
+ 757590.800000ns, VSS,
+ 757590.900000ns, VDD,
+ 758431.500000ns, VDD,
+ 758431.600000ns, VSS,
+ 759992.800000ns, VSS,
+ 759992.900000ns, VDD,
+ 760233.000000ns, VDD,
+ 760233.100000ns, VSS,
+ 760953.600000ns, VSS,
+ 760953.700000ns, VDD,
+ 762394.800000ns, VDD,
+ 762394.900000ns, VSS,
+ 762755.100000ns, VSS,
+ 762755.200000ns, VDD,
+ 762875.200000ns, VDD,
+ 762875.300000ns, VSS,
+ 762995.300000ns, VSS,
+ 762995.400000ns, VDD,
+ 763355.600000ns, VDD,
+ 763355.700000ns, VSS,
+ 763956.100000ns, VSS,
+ 763956.200000ns, VDD,
+ 764436.500000ns, VDD,
+ 764436.600000ns, VSS,
+ 765277.200000ns, VSS,
+ 765277.300000ns, VDD,
+ 765517.400000ns, VDD,
+ 765517.500000ns, VSS,
+ 765877.700000ns, VSS,
+ 765877.800000ns, VDD,
+ 766358.100000ns, VDD,
+ 766358.200000ns, VSS,
+ 767198.800000ns, VSS,
+ 767198.900000ns, VDD,
+ 768279.700000ns, VDD,
+ 768279.800000ns, VSS,
+ 768519.900000ns, VSS,
+ 768520.000000ns, VDD,
+ 768640.000000ns, VDD,
+ 768640.100000ns, VSS,
+ 768760.100000ns, VSS,
+ 768760.200000ns, VDD,
+ 769360.600000ns, VDD,
+ 769360.700000ns, VSS,
+ 769480.700000ns, VSS,
+ 769480.800000ns, VDD,
+ 769600.800000ns, VDD,
+ 769600.900000ns, VSS,
+ 770081.200000ns, VSS,
+ 770081.300000ns, VDD,
+ 770801.800000ns, VDD,
+ 770801.900000ns, VSS,
+ 771042.000000ns, VSS,
+ 771042.100000ns, VDD,
+ 771162.100000ns, VDD,
+ 771162.200000ns, VSS,
+ 771642.500000ns, VSS,
+ 771642.600000ns, VDD,
+ 772122.900000ns, VDD,
+ 772123.000000ns, VSS,
+ 772483.200000ns, VSS,
+ 772483.300000ns, VDD,
+ 774164.600000ns, VDD,
+ 774164.700000ns, VSS,
+ 774524.900000ns, VSS,
+ 774525.000000ns, VDD,
+ 777887.700000ns, VDD,
+ 777887.800000ns, VSS,
+ 778248.000000ns, VSS,
+ 778248.100000ns, VDD,
+ 778608.300000ns, VDD,
+ 778608.400000ns, VSS,
+ 778968.600000ns, VSS,
+ 778968.700000ns, VDD,
+ 779689.200000ns, VDD,
+ 779689.300000ns, VSS,
+ 780650.000000ns, VSS,
+ 780650.100000ns, VDD,
+ 780770.100000ns, VDD,
+ 780770.200000ns, VSS,
+ 781851.000000ns, VSS,
+ 781851.100000ns, VDD,
+ 782571.600000ns, VDD,
+ 782571.700000ns, VSS,
+ 783052.000000ns, VSS,
+ 783052.100000ns, VDD,
+ 783172.100000ns, VDD,
+ 783172.200000ns, VSS,
+ 784132.900000ns, VSS,
+ 784133.000000ns, VDD,
+ 785093.700000ns, VDD,
+ 785093.800000ns, VSS,
+ 785454.000000ns, VSS,
+ 785454.100000ns, VDD,
+ 785934.400000ns, VDD,
+ 785934.500000ns, VSS,
+ 787255.500000ns, VSS,
+ 787255.600000ns, VDD,
+ 788216.300000ns, VDD,
+ 788216.400000ns, VSS,
+ 788696.700000ns, VSS,
+ 788696.800000ns, VDD,
+ 788936.900000ns, VDD,
+ 788937.000000ns, VSS,
+ 789417.300000ns, VSS,
+ 789417.400000ns, VDD,
+ 790618.300000ns, VDD,
+ 790618.400000ns, VSS,
+ 791338.900000ns, VSS,
+ 791339.000000ns, VDD,
+ 791939.400000ns, VDD,
+ 791939.500000ns, VSS,
+ 792539.900000ns, VSS,
+ 792540.000000ns, VDD,
+ 792900.200000ns, VDD,
+ 792900.300000ns, VSS,
+ 793260.500000ns, VSS,
+ 793260.600000ns, VDD,
+ 793500.700000ns, VDD,
+ 793500.800000ns, VSS,
+ 793861.000000ns, VSS,
+ 793861.100000ns, VDD,
+ 794701.700000ns, VDD,
+ 794701.800000ns, VSS,
+ 795182.100000ns, VSS,
+ 795182.200000ns, VDD,
+ 796142.900000ns, VDD,
+ 796143.000000ns, VSS,
+ 796863.500000ns, VSS,
+ 796863.600000ns, VDD,
+ 797944.400000ns, VDD,
+ 797944.500000ns, VSS,
+ 798064.500000ns, VSS,
+ 798064.600000ns, VDD,
+ 798665.000000ns, VDD,
+ 798665.100000ns, VSS,
+ 798785.100000ns, VSS,
+ 798785.200000ns, VDD,
+ 798905.200000ns, VDD,
+ 798905.300000ns, VSS,
+ 799505.700000ns, VSS,
+ 799505.800000ns, VDD,
+ 800106.200000ns, VDD,
+ 800106.300000ns, VSS,
+ 800226.300000ns, VSS,
+ 800226.400000ns, VDD,
+ 800826.800000ns, VDD,
+ 800826.900000ns, VSS,
+ 801787.600000ns, VSS,
+ 801787.700000ns, VDD,
+ 802027.800000ns, VDD,
+ 802027.900000ns, VSS,
+ 802147.900000ns, VSS,
+ 802148.000000ns, VDD,
+ 802268.000000ns, VDD,
+ 802268.100000ns, VSS,
+ 804429.800000ns, VSS,
+ 804429.900000ns, VDD,
+ 805390.600000ns, VDD,
+ 805390.700000ns, VSS,
+ 805991.100000ns, VSS,
+ 805991.200000ns, VDD,
+ 806111.200000ns, VDD,
+ 806111.300000ns, VSS,
+ 806231.300000ns, VSS,
+ 806231.400000ns, VDD,
+ 806471.500000ns, VDD,
+ 806471.600000ns, VSS,
+ 806591.600000ns, VSS,
+ 806591.700000ns, VDD,
+ 807192.100000ns, VDD,
+ 807192.200000ns, VSS,
+ 807312.200000ns, VSS,
+ 807312.300000ns, VDD,
+ 808152.900000ns, VDD,
+ 808153.000000ns, VSS,
+ 808273.000000ns, VSS,
+ 808273.100000ns, VDD,
+ 808393.100000ns, VDD,
+ 808393.200000ns, VSS,
+ 809714.200000ns, VSS,
+ 809714.300000ns, VDD,
+ 810314.700000ns, VDD,
+ 810314.800000ns, VSS,
+ 810675.000000ns, VSS,
+ 810675.100000ns, VDD,
+ 810795.100000ns, VDD,
+ 810795.200000ns, VSS,
+ 811395.600000ns, VSS,
+ 811395.700000ns, VDD,
+ 811515.700000ns, VDD,
+ 811515.800000ns, VSS,
+ 812116.200000ns, VSS,
+ 812116.300000ns, VDD,
+ 812476.500000ns, VDD,
+ 812476.600000ns, VSS,
+ 813677.500000ns, VSS,
+ 813677.600000ns, VDD,
+ 817160.400000ns, VDD,
+ 817160.500000ns, VSS,
+ 817760.900000ns, VSS,
+ 817761.000000ns, VDD,
+ 819562.400000ns, VDD,
+ 819562.500000ns, VSS,
+ 820403.100000ns, VSS,
+ 820403.200000ns, VDD,
+ 820523.200000ns, VDD,
+ 820523.300000ns, VSS,
+ 821123.700000ns, VSS,
+ 821123.800000ns, VDD,
+ 821484.000000ns, VDD,
+ 821484.100000ns, VSS,
+ 821604.100000ns, VSS,
+ 821604.200000ns, VDD,
+ 821724.200000ns, VDD,
+ 821724.300000ns, VSS,
+ 822204.600000ns, VSS,
+ 822204.700000ns, VDD,
+ 822564.900000ns, VDD,
+ 822565.000000ns, VSS,
+ 822685.000000ns, VSS,
+ 822685.100000ns, VDD,
+ 822925.200000ns, VDD,
+ 822925.300000ns, VSS,
+ 823165.400000ns, VSS,
+ 823165.500000ns, VDD,
+ 823645.800000ns, VDD,
+ 823645.900000ns, VSS,
+ 823765.900000ns, VSS,
+ 823766.000000ns, VDD,
+ 825807.600000ns, VDD,
+ 825807.700000ns, VSS,
+ 826288.000000ns, VSS,
+ 826288.100000ns, VDD,
+ 826408.100000ns, VDD,
+ 826408.200000ns, VSS,
+ 826648.300000ns, VSS,
+ 826648.400000ns, VDD,
+ 827248.800000ns, VDD,
+ 827248.900000ns, VSS,
+ 827969.400000ns, VSS,
+ 827969.500000ns, VDD,
+ 829170.400000ns, VDD,
+ 829170.500000ns, VSS,
+ 829770.900000ns, VSS,
+ 829771.000000ns, VDD,
+ 831212.100000ns, VDD,
+ 831212.200000ns, VSS,
+ 832172.900000ns, VSS,
+ 832173.000000ns, VDD,
+ 832293.000000ns, VDD,
+ 832293.100000ns, VSS,
+ 832413.100000ns, VSS,
+ 832413.200000ns, VDD,
+ 832773.400000ns, VDD,
+ 832773.500000ns, VSS,
+ 832893.500000ns, VSS,
+ 832893.600000ns, VDD,
+ 833734.200000ns, VDD,
+ 833734.300000ns, VSS,
+ 835055.300000ns, VSS,
+ 835055.400000ns, VDD,
+ 835415.600000ns, VDD,
+ 835415.700000ns, VSS,
+ 836496.500000ns, VSS,
+ 836496.600000ns, VDD,
+ 837097.000000ns, VDD,
+ 837097.100000ns, VSS,
+ 838298.000000ns, VSS,
+ 838298.100000ns, VDD,
+ 838778.400000ns, VDD,
+ 838778.500000ns, VSS,
+ 841300.500000ns, VSS,
+ 841300.600000ns, VDD,
+ 841420.600000ns, VDD,
+ 841420.700000ns, VSS,
+ 841540.700000ns, VSS,
+ 841540.800000ns, VDD,
+ 842021.100000ns, VDD,
+ 842021.200000ns, VSS,
+ 842261.300000ns, VSS,
+ 842261.400000ns, VDD,
+ 842741.700000ns, VDD,
+ 842741.800000ns, VSS,
+ 843102.000000ns, VSS,
+ 843102.100000ns, VDD,
+ 845143.700000ns, VDD,
+ 845143.800000ns, VSS,
+ 845263.800000ns, VSS,
+ 845263.900000ns, VDD,
+ 845864.300000ns, VDD,
+ 845864.400000ns, VSS,
+ 845984.400000ns, VSS,
+ 845984.500000ns, VDD,
+ 846464.800000ns, VDD,
+ 846464.900000ns, VSS,
+ 846945.200000ns, VSS,
+ 846945.300000ns, VDD,
+ 847785.900000ns, VDD,
+ 847786.000000ns, VSS,
+ 848626.600000ns, VSS,
+ 848626.700000ns, VDD,
+ 849107.000000ns, VDD,
+ 849107.100000ns, VSS,
+ 849587.400000ns, VSS,
+ 849587.500000ns, VDD,
+ 850187.900000ns, VDD,
+ 850188.000000ns, VSS,
+ 851268.800000ns, VSS,
+ 851268.900000ns, VDD,
+ 851869.300000ns, VDD,
+ 851869.400000ns, VSS,
+ 852109.500000ns, VSS,
+ 852109.600000ns, VDD,
+ 852830.100000ns, VDD,
+ 852830.200000ns, VSS,
+ 853070.300000ns, VSS,
+ 853070.400000ns, VDD,
+ 854511.500000ns, VDD,
+ 854511.600000ns, VSS,
+ 854751.700000ns, VSS,
+ 854751.800000ns, VDD,
+ 854871.800000ns, VDD,
+ 854871.900000ns, VSS,
+ 855472.300000ns, VSS,
+ 855472.400000ns, VDD,
+ 858114.500000ns, VDD,
+ 858114.600000ns, VSS,
+ 858234.600000ns, VSS,
+ 858234.700000ns, VDD,
+ 859675.800000ns, VDD,
+ 859675.900000ns, VSS,
+ 860756.700000ns, VSS,
+ 860756.800000ns, VDD,
+ 860876.800000ns, VDD,
+ 860876.900000ns, VSS,
+ 861357.200000ns, VSS,
+ 861357.300000ns, VDD,
+ 862077.800000ns, VDD,
+ 862077.900000ns, VSS,
+ 863278.800000ns, VSS,
+ 863278.900000ns, VDD,
+ 863398.900000ns, VDD,
+ 863399.000000ns, VSS,
+ 863759.200000ns, VSS,
+ 863759.300000ns, VDD,
+ 865440.600000ns, VDD,
+ 865440.700000ns, VSS,
+ 865680.800000ns, VSS,
+ 865680.900000ns, VDD,
+ 866881.800000ns, VDD,
+ 866881.900000ns, VSS,
+ 867362.200000ns, VSS,
+ 867362.300000ns, VDD,
+ 867602.400000ns, VDD,
+ 867602.500000ns, VSS,
+ 868082.800000ns, VSS,
+ 868082.900000ns, VDD,
+ 869163.700000ns, VDD,
+ 869163.800000ns, VSS,
+ 869283.800000ns, VSS,
+ 869283.900000ns, VDD,
+ 869764.200000ns, VDD,
+ 869764.300000ns, VSS,
+ 870124.500000ns, VSS,
+ 870124.600000ns, VDD,
+ 870244.600000ns, VDD,
+ 870244.700000ns, VSS,
+ 870725.000000ns, VSS,
+ 870725.100000ns, VDD,
+ 870845.100000ns, VDD,
+ 870845.200000ns, VSS,
+ 870965.200000ns, VSS,
+ 870965.300000ns, VDD,
+ 871685.800000ns, VDD,
+ 871685.900000ns, VSS,
+ 872046.100000ns, VSS,
+ 872046.200000ns, VDD,
+ 873247.100000ns, VDD,
+ 873247.200000ns, VSS,
+ 873367.200000ns, VSS,
+ 873367.300000ns, VDD,
+ 873967.700000ns, VDD,
+ 873967.800000ns, VSS,
+ 875168.700000ns, VSS,
+ 875168.800000ns, VDD,
+ 876129.500000ns, VDD,
+ 876129.600000ns, VSS,
+ 876249.600000ns, VSS,
+ 876249.700000ns, VDD,
+ 878171.200000ns, VDD,
+ 878171.300000ns, VSS,
+ 878651.600000ns, VSS,
+ 878651.700000ns, VDD,
+ 879372.200000ns, VDD,
+ 879372.300000ns, VSS,
+ 880333.000000ns, VSS,
+ 880333.100000ns, VDD,
+ 881173.700000ns, VDD,
+ 881173.800000ns, VSS,
+ 882374.700000ns, VSS,
+ 882374.800000ns, VDD,
+ 883215.400000ns, VDD,
+ 883215.500000ns, VSS,
+ 883815.900000ns, VSS,
+ 883816.000000ns, VDD,
+ 884296.300000ns, VDD,
+ 884296.400000ns, VSS,
+ 884536.500000ns, VSS,
+ 884536.600000ns, VDD,
+ 884656.600000ns, VDD,
+ 884656.700000ns, VSS,
+ 885617.400000ns, VSS,
+ 885617.500000ns, VDD,
+ 888259.600000ns, VDD,
+ 888259.700000ns, VSS,
+ 888499.800000ns, VSS,
+ 888499.900000ns, VDD,
+ 888980.200000ns, VDD,
+ 888980.300000ns, VSS,
+ 891142.000000ns, VSS,
+ 891142.100000ns, VDD,
+ 891262.100000ns, VDD,
+ 891262.200000ns, VSS,
+ 891382.200000ns, VSS,
+ 891382.300000ns, VDD,
+ 891622.400000ns, VDD,
+ 891622.500000ns, VSS,
+ 892583.200000ns, VSS,
+ 892583.300000ns, VDD,
+ 892703.300000ns, VDD,
+ 892703.400000ns, VSS,
+ 892823.400000ns, VSS,
+ 892823.500000ns, VDD,
+ 893063.600000ns, VDD,
+ 893063.700000ns, VSS,
+ 893183.700000ns, VSS,
+ 893183.800000ns, VDD,
+ 893664.100000ns, VDD,
+ 893664.200000ns, VSS,
+ 893784.200000ns, VSS,
+ 893784.300000ns, VDD,
+ 893904.300000ns, VDD,
+ 893904.400000ns, VSS,
+ 895585.700000ns, VSS,
+ 895585.800000ns, VDD,
+ 896426.400000ns, VDD,
+ 896426.500000ns, VSS,
+ 897387.200000ns, VSS,
+ 897387.300000ns, VDD,
+ 898348.000000ns, VDD,
+ 898348.100000ns, VSS,
+ 898468.100000ns, VSS,
+ 898468.200000ns, VDD,
+ 899068.600000ns, VDD,
+ 899068.700000ns, VSS,
+ 900750.000000ns, VSS,
+ 900750.100000ns, VDD,
+ 901951.000000ns, VDD,
+ 901951.100000ns, VSS,
+ 903031.900000ns, VSS,
+ 903032.000000ns, VDD,
+ 903512.300000ns, VDD,
+ 903512.400000ns, VSS,
+ 904593.200000ns, VSS,
+ 904593.300000ns, VDD,
+ 904833.400000ns, VDD,
+ 904833.500000ns, VSS,
+ 909277.100000ns, VSS,
+ 909277.200000ns, VDD,
+ 909757.500000ns, VDD,
+ 909757.600000ns, VSS,
+ 911318.800000ns, VSS,
+ 911318.900000ns, VDD,
+ 912880.100000ns, VDD,
+ 912880.200000ns, VSS,
+ 913720.800000ns, VSS,
+ 913720.900000ns, VDD,
+ 914921.800000ns, VDD,
+ 914921.900000ns, VSS,
+ 915041.900000ns, VSS,
+ 915042.000000ns, VDD,
+ 915162.000000ns, VDD,
+ 915162.100000ns, VSS,
+ 916122.800000ns, VSS,
+ 916122.900000ns, VDD,
+ 916963.500000ns, VDD,
+ 916963.600000ns, VSS,
+ 917083.600000ns, VSS,
+ 917083.700000ns, VDD,
+ 919125.300000ns, VDD,
+ 919125.400000ns, VSS,
+ 920806.700000ns, VSS,
+ 920806.800000ns, VDD,
+ 921046.900000ns, VDD,
+ 921047.000000ns, VSS,
+ 921287.100000ns, VSS,
+ 921287.200000ns, VDD,
+ 922007.700000ns, VDD,
+ 922007.800000ns, VSS,
+ 922488.100000ns, VSS,
+ 922488.200000ns, VDD,
+ 922968.500000ns, VDD,
+ 922968.600000ns, VSS,
+ 923088.600000ns, VSS,
+ 923088.700000ns, VDD,
+ 923208.700000ns, VDD,
+ 923208.800000ns, VSS,
+ 923448.900000ns, VSS,
+ 923449.000000ns, VDD,
+ 923809.200000ns, VDD,
+ 923809.300000ns, VSS,
+ 924169.500000ns, VSS,
+ 924169.600000ns, VDD,
+ 924649.900000ns, VDD,
+ 924650.000000ns, VSS,
+ 925370.500000ns, VSS,
+ 925370.600000ns, VDD,
+ 925730.800000ns, VDD,
+ 925730.900000ns, VSS,
+ 925850.900000ns, VSS,
+ 925851.000000ns, VDD,
+ 925971.000000ns, VDD,
+ 925971.100000ns, VSS,
+ 926691.600000ns, VSS,
+ 926691.700000ns, VDD,
+ 927412.200000ns, VDD,
+ 927412.300000ns, VSS,
+ 928132.800000ns, VSS,
+ 928132.900000ns, VDD,
+ 928853.400000ns, VDD,
+ 928853.500000ns, VSS,
+ 929574.000000ns, VSS,
+ 929574.100000ns, VDD,
+ 929694.100000ns, VDD,
+ 929694.200000ns, VSS,
+ 930174.500000ns, VSS,
+ 930174.600000ns, VDD,
+ 931015.200000ns, VDD,
+ 931015.300000ns, VSS,
+ 931135.300000ns, VSS,
+ 931135.400000ns, VDD,
+ 931735.800000ns, VDD,
+ 931735.900000ns, VSS,
+ 932696.600000ns, VSS,
+ 932696.700000ns, VDD,
+ 932816.700000ns, VDD,
+ 932816.800000ns, VSS,
+ 933297.100000ns, VSS,
+ 933297.200000ns, VDD,
+ 933417.200000ns, VDD,
+ 933417.300000ns, VSS,
+ 934498.100000ns, VSS,
+ 934498.200000ns, VDD,
+ 934738.300000ns, VDD,
+ 934738.400000ns, VSS,
+ 934858.400000ns, VSS,
+ 934858.500000ns, VDD,
+ 935819.200000ns, VDD,
+ 935819.300000ns, VSS,
+ 936780.000000ns, VSS,
+ 936780.100000ns, VDD,
+ 937380.500000ns, VDD,
+ 937380.600000ns, VSS,
+ 937620.700000ns, VSS,
+ 937620.800000ns, VDD,
+ 937740.800000ns, VDD,
+ 937740.900000ns, VSS,
+ 937860.900000ns, VSS,
+ 937861.000000ns, VDD,
+ 938101.100000ns, VDD,
+ 938101.200000ns, VSS,
+ 938341.300000ns, VSS,
+ 938341.400000ns, VDD,
+ 938941.800000ns, VDD,
+ 938941.900000ns, VSS,
+ 940022.700000ns, VSS,
+ 940022.800000ns, VDD,
+ 940383.000000ns, VDD,
+ 940383.100000ns, VSS,
+ 941584.000000ns, VSS,
+ 941584.100000ns, VDD,
+ 941704.100000ns, VDD,
+ 941704.200000ns, VSS,
+ 942184.500000ns, VSS,
+ 942184.600000ns, VDD,
+ 943145.300000ns, VDD,
+ 943145.400000ns, VSS,
+ 943745.800000ns, VSS,
+ 943745.900000ns, VDD,
+ 944106.100000ns, VDD,
+ 944106.200000ns, VSS,
+ 944586.500000ns, VSS,
+ 944586.600000ns, VDD,
+ 945066.900000ns, VDD,
+ 945067.000000ns, VSS,
+ 945667.400000ns, VSS,
+ 945667.500000ns, VDD,
+ 946147.800000ns, VDD,
+ 946147.900000ns, VSS,
+ 946267.900000ns, VSS,
+ 946268.000000ns, VDD,
+ 946628.200000ns, VDD,
+ 946628.300000ns, VSS,
+ 947949.300000ns, VSS,
+ 947949.400000ns, VDD,
+ 948549.800000ns, VDD,
+ 948549.900000ns, VSS,
+ 949390.500000ns, VSS,
+ 949390.600000ns, VDD,
+ 950231.200000ns, VDD,
+ 950231.300000ns, VSS,
+ 950591.500000ns, VSS,
+ 950591.600000ns, VDD,
+ 951432.200000ns, VDD,
+ 951432.300000ns, VSS,
+ 951552.300000ns, VSS,
+ 951552.400000ns, VDD,
+ 952152.800000ns, VDD,
+ 952152.900000ns, VSS,
+ 952272.900000ns, VSS,
+ 952273.000000ns, VDD,
+ 953233.700000ns, VDD,
+ 953233.800000ns, VSS,
+ 953954.300000ns, VSS,
+ 953954.400000ns, VDD,
+ 954915.100000ns, VDD,
+ 954915.200000ns, VSS,
+ 955996.000000ns, VSS,
+ 955996.100000ns, VDD,
+ 956836.700000ns, VDD,
+ 956836.800000ns, VSS,
+ 956956.800000ns, VSS,
+ 956956.900000ns, VDD,
+ 957076.900000ns, VDD,
+ 957077.000000ns, VSS,
+ 957557.300000ns, VSS,
+ 957557.400000ns, VDD,
+ 957917.600000ns, VDD,
+ 957917.700000ns, VSS,
+ 958157.800000ns, VSS,
+ 958157.900000ns, VDD,
+ 958277.900000ns, VDD,
+ 958278.000000ns, VSS,
+ 958398.000000ns, VSS,
+ 958398.100000ns, VDD,
+ 959238.700000ns, VDD,
+ 959238.800000ns, VSS,
+ 959599.000000ns, VSS,
+ 959599.100000ns, VDD,
+ 961760.800000ns, VDD,
+ 961760.900000ns, VSS,
+ 962721.600000ns, VSS,
+ 962721.700000ns, VDD,
+ 965363.800000ns, VDD,
+ 965363.900000ns, VSS,
+ 965724.100000ns, VSS,
+ 965724.200000ns, VDD,
+ 966204.500000ns, VDD,
+ 966204.600000ns, VSS,
+ 966684.900000ns, VSS,
+ 966685.000000ns, VDD,
+ 966925.100000ns, VDD,
+ 966925.200000ns, VSS,
+ 967045.200000ns, VSS,
+ 967045.300000ns, VDD,
+ 967525.600000ns, VDD,
+ 967525.700000ns, VSS,
+ 968486.400000ns, VSS,
+ 968486.500000ns, VDD,
+ 968966.800000ns, VDD,
+ 968966.900000ns, VSS,
+ 969927.600000ns, VSS,
+ 969927.700000ns, VDD,
+ 970287.900000ns, VDD,
+ 970288.000000ns, VSS,
+ 971128.600000ns, VSS,
+ 971128.700000ns, VDD,
+ 972329.600000ns, VDD,
+ 972329.700000ns, VSS,
+ 972810.000000ns, VSS,
+ 972810.100000ns, VDD,
+ 974131.100000ns, VDD,
+ 974131.200000ns, VSS,
+ 975212.000000ns, VSS,
+ 975212.100000ns, VDD,
+ 975572.300000ns, VDD,
+ 975572.400000ns, VSS,
+ 975812.500000ns, VSS,
+ 975812.600000ns, VDD,
+ 976172.800000ns, VDD,
+ 976172.900000ns, VSS,
+ 976653.200000ns, VSS,
+ 976653.300000ns, VDD,
+ 976773.300000ns, VDD,
+ 976773.400000ns, VSS,
+ 978574.800000ns, VSS,
+ 978574.900000ns, VDD,
+ 978935.100000ns, VDD,
+ 978935.200000ns, VSS,
+ 980736.600000ns, VSS,
+ 980736.700000ns, VDD,
+ 982297.900000ns, VDD,
+ 982298.000000ns, VSS,
+ 983018.500000ns, VSS,
+ 983018.600000ns, VDD,
+ 983138.600000ns, VDD,
+ 983138.700000ns, VSS,
+ 983258.700000ns, VSS,
+ 983258.800000ns, VDD,
+ 983498.900000ns, VDD,
+ 983499.000000ns, VSS,
+ 984940.100000ns, VSS,
+ 984940.200000ns, VDD,
+ 985060.200000ns, VDD,
+ 985060.300000ns, VSS,
+ 985300.400000ns, VSS,
+ 985300.500000ns, VDD,
+ 986261.200000ns, VDD,
+ 986261.300000ns, VSS,
+ 986381.300000ns, VSS,
+ 986381.400000ns, VDD,
+ 987101.900000ns, VDD,
+ 987102.000000ns, VSS,
+ 987462.200000ns, VSS,
+ 987462.300000ns, VDD,
+ 987582.300000ns, VDD,
+ 987582.400000ns, VSS,
+ 987702.400000ns, VSS,
+ 987702.500000ns, VDD,
+ 988182.800000ns, VDD,
+ 988182.900000ns, VSS,
+ 988543.100000ns, VSS,
+ 988543.200000ns, VDD,
+ 989143.600000ns, VDD,
+ 989143.700000ns, VSS,
+ 989864.200000ns, VSS,
+ 989864.300000ns, VDD,
+ 990464.700000ns, VDD,
+ 990464.800000ns, VSS,
+ 990704.900000ns, VSS,
+ 990705.000000ns, VDD,
+ 991185.300000ns, VDD,
+ 991185.400000ns, VSS,
+ 991305.400000ns, VSS,
+ 991305.500000ns, VDD,
+ 992386.300000ns, VDD,
+ 992386.400000ns, VSS,
+ 993106.900000ns, VSS,
+ 993107.000000ns, VDD,
+ 993227.000000ns, VDD,
+ 993227.100000ns, VSS,
+ 993707.400000ns, VSS,
+ 993707.500000ns, VDD,
+ 995148.600000ns, VDD,
+ 995148.700000ns, VSS,
+ 997070.200000ns, VSS,
+ 997070.300000ns, VDD,
+ 997310.400000ns, VDD,
+ 997310.500000ns, VSS,
+ 997670.700000ns, VSS,
+ 997670.800000ns, VDD,
+ 998751.600000ns, VDD,
+ 998751.700000ns, VSS,
+ 999832.500000ns, VSS,
+ 999832.600000ns, VDD,
+ 1001273.700000ns, VDD,
+ 1001273.800000ns, VSS,
+ 1001754.100000ns, VSS,
+ 1001754.200000ns, VDD,
+ 1001994.300000ns, VDD,
+ 1001994.400000ns, VSS,
+ 1002594.800000ns, VSS,
+ 1002594.900000ns, VDD,
+ 1002955.100000ns, VDD,
+ 1002955.200000ns, VSS,
+ 1003435.500000ns, VSS,
+ 1003435.600000ns, VDD,
+ 1005717.400000ns, VDD,
+ 1005717.500000ns, VSS,
+ 1006077.700000ns, VSS,
+ 1006077.800000ns, VDD,
+ 1006438.000000ns, VDD,
+ 1006438.100000ns, VSS,
+ 1006558.100000ns, VSS,
+ 1006558.200000ns, VDD,
+ 1006678.200000ns, VDD,
+ 1006678.300000ns, VSS,
+ 1007639.000000ns, VSS,
+ 1007639.100000ns, VDD,
+ 1007879.200000ns, VDD,
+ 1007879.300000ns, VSS,
+ 1009080.200000ns, VSS,
+ 1009080.300000ns, VDD,
+ 1009560.600000ns, VDD,
+ 1009560.700000ns, VSS,
+ 1009800.800000ns, VSS,
+ 1009800.900000ns, VDD,
+ 1009920.900000ns, VDD,
+ 1009921.000000ns, VSS,
+ 1010161.100000ns, VSS,
+ 1010161.200000ns, VDD,
+ 1011602.300000ns, VDD,
+ 1011602.400000ns, VSS,
+ 1012322.900000ns, VSS,
+ 1012323.000000ns, VDD,
+ 1012803.300000ns, VDD,
+ 1012803.400000ns, VSS,
+ 1014364.600000ns, VSS,
+ 1014364.700000ns, VDD,
+ 1014724.900000ns, VDD,
+ 1014725.000000ns, VSS,
+ 1015685.700000ns, VSS,
+ 1015685.800000ns, VDD,
+ 1016166.100000ns, VDD,
+ 1016166.200000ns, VSS,
+ 1016646.500000ns, VSS,
+ 1016646.600000ns, VDD,
+ 1016766.600000ns, VDD,
+ 1016766.700000ns, VSS,
+ 1017126.900000ns, VSS,
+ 1017127.000000ns, VDD,
+ 1017607.300000ns, VDD,
+ 1017607.400000ns, VSS,
+ 1018448.000000ns, VSS,
+ 1018448.100000ns, VDD,
+ 1019889.200000ns, VDD,
+ 1019889.300000ns, VSS,
+ 1020970.100000ns, VSS,
+ 1020970.200000ns, VDD,
+ 1021570.600000ns, VDD,
+ 1021570.700000ns, VSS,
+ 1021690.700000ns, VSS,
+ 1021690.800000ns, VDD,
+ 1022051.000000ns, VDD,
+ 1022051.100000ns, VSS,
+ 1022171.100000ns, VSS,
+ 1022171.200000ns, VDD,
+ 1024453.000000ns, VDD,
+ 1024453.100000ns, VSS,
+ 1025533.900000ns, VSS,
+ 1025534.000000ns, VDD,
+ 1025654.000000ns, VDD,
+ 1025654.100000ns, VSS,
+ 1026134.400000ns, VSS,
+ 1026134.500000ns, VDD,
+ 1027095.200000ns, VDD,
+ 1027095.300000ns, VSS,
+ 1027335.400000ns, VSS,
+ 1027335.500000ns, VDD,
+ 1027935.900000ns, VDD,
+ 1027936.000000ns, VSS,
+ 1029016.800000ns, VSS,
+ 1029016.900000ns, VDD,
+ 1029257.000000ns, VDD,
+ 1029257.100000ns, VSS,
+ 1029497.200000ns, VSS,
+ 1029497.300000ns, VDD,
+ 1029737.400000ns, VDD,
+ 1029737.500000ns, VSS,
+ 1029857.500000ns, VSS,
+ 1029857.600000ns, VDD,
+ 1030698.200000ns, VDD,
+ 1030698.300000ns, VSS,
+ 1031779.100000ns, VSS,
+ 1031779.200000ns, VDD,
+ 1032139.400000ns, VDD,
+ 1032139.500000ns, VSS,
+ 1033580.600000ns, VSS,
+ 1033580.700000ns, VDD,
+ 1035141.900000ns, VDD,
+ 1035142.000000ns, VSS,
+ 1035862.500000ns, VSS,
+ 1035862.600000ns, VDD,
+ 1036463.000000ns, VDD,
+ 1036463.100000ns, VSS,
+ 1037183.600000ns, VSS,
+ 1037183.700000ns, VDD,
+ 1037664.000000ns, VDD,
+ 1037664.100000ns, VSS,
+ 1038144.400000ns, VSS,
+ 1038144.500000ns, VDD,
+ 1038865.000000ns, VDD,
+ 1038865.100000ns, VSS,
+ 1039225.300000ns, VSS,
+ 1039225.400000ns, VDD,
+ 1039945.900000ns, VDD,
+ 1039946.000000ns, VSS,
+ 1041627.300000ns, VSS,
+ 1041627.400000ns, VDD,
+ 1041747.400000ns, VDD,
+ 1041747.500000ns, VSS,
+ 1041867.500000ns, VSS,
+ 1041867.600000ns, VDD,
+ 1042828.300000ns, VDD,
+ 1042828.400000ns, VSS,
+ 1043068.500000ns, VSS,
+ 1043068.600000ns, VDD,
+ 1043308.700000ns, VDD,
+ 1043308.800000ns, VSS,
+ 1043428.800000ns, VSS,
+ 1043428.900000ns, VDD,
+ 1044269.500000ns, VDD,
+ 1044269.600000ns, VSS,
+ 1044389.600000ns, VSS,
+ 1044389.700000ns, VDD,
+ 1046551.400000ns, VDD,
+ 1046551.500000ns, VSS,
+ 1046791.600000ns, VSS,
+ 1046791.700000ns, VDD,
+ 1047392.100000ns, VDD,
+ 1047392.200000ns, VSS,
+ 1047872.500000ns, VSS,
+ 1047872.600000ns, VDD,
+ 1048352.900000ns, VDD,
+ 1048353.000000ns, VSS,
+ 1048953.400000ns, VSS,
+ 1048953.500000ns, VDD,
+ 1049073.500000ns, VDD,
+ 1049073.600000ns, VSS,
+ 1049193.600000ns, VSS,
+ 1049193.700000ns, VDD,
+ 1049433.800000ns, VDD,
+ 1049433.900000ns, VSS,
+ 1049553.900000ns, VSS,
+ 1049554.000000ns, VDD,
+ 1051355.400000ns, VDD,
+ 1051355.500000ns, VSS,
+ 1052436.300000ns, VSS,
+ 1052436.400000ns, VDD,
+ 1052916.700000ns, VDD,
+ 1052916.800000ns, VSS,
+ 1053156.900000ns, VSS,
+ 1053157.000000ns, VDD,
+ 1053277.000000ns, VDD,
+ 1053277.100000ns, VSS,
+ 1053877.500000ns, VSS,
+ 1053877.600000ns, VDD,
+ 1054357.900000ns, VDD,
+ 1054358.000000ns, VSS,
+ 1056399.600000ns, VSS,
+ 1056399.700000ns, VDD,
+ 1056880.000000ns, VDD,
+ 1056880.100000ns, VSS,
+ 1057840.800000ns, VSS,
+ 1057840.900000ns, VDD,
+ 1058801.600000ns, VDD,
+ 1058801.700000ns, VSS,
+ 1059282.000000ns, VSS,
+ 1059282.100000ns, VDD,
+ 1060963.400000ns, VDD,
+ 1060963.500000ns, VSS,
+ 1061804.100000ns, VSS,
+ 1061804.200000ns, VDD,
+ 1062644.800000ns, VDD,
+ 1062644.900000ns, VSS,
+ 1064686.500000ns, VSS,
+ 1064686.600000ns, VDD,
+ 1065166.900000ns, VDD,
+ 1065167.000000ns, VSS,
+ 1065887.500000ns, VSS,
+ 1065887.600000ns, VDD,
+ 1066127.700000ns, VDD,
+ 1066127.800000ns, VSS,
+ 1067328.700000ns, VSS,
+ 1067328.800000ns, VDD,
+ 1068049.300000ns, VDD,
+ 1068049.400000ns, VSS,
+ 1068649.800000ns, VSS,
+ 1068649.900000ns, VDD,
+ 1069250.300000ns, VDD,
+ 1069250.400000ns, VSS,
+ 1069730.700000ns, VSS,
+ 1069730.800000ns, VDD,
+ 1070451.300000ns, VDD,
+ 1070451.400000ns, VSS,
+ 1071171.900000ns, VSS,
+ 1071172.000000ns, VDD,
+ 1072973.400000ns, VDD,
+ 1072973.500000ns, VSS,
+ 1074054.300000ns, VSS,
+ 1074054.400000ns, VDD,
+ 1074294.500000ns, VDD,
+ 1074294.600000ns, VSS,
+ 1075375.400000ns, VSS,
+ 1075375.500000ns, VDD,
+ 1075615.600000ns, VDD,
+ 1075615.700000ns, VSS,
+ 1077056.800000ns, VSS,
+ 1077056.900000ns, VDD,
+ 1077777.400000ns, VDD,
+ 1077777.500000ns, VSS,
+ 1078377.900000ns, VSS,
+ 1078378.000000ns, VDD,
+ 1079338.700000ns, VDD,
+ 1079338.800000ns, VSS,
+ 1080419.600000ns, VSS,
+ 1080419.700000ns, VDD,
+ 1080539.700000ns, VDD,
+ 1080539.800000ns, VSS,
+ 1081140.200000ns, VSS,
+ 1081140.300000ns, VDD,
+ 1081620.600000ns, VDD,
+ 1081620.700000ns, VSS,
+ 1081980.900000ns, VSS,
+ 1081981.000000ns, VDD,
+ 1082341.200000ns, VDD,
+ 1082341.300000ns, VSS,
+ 1083662.300000ns, VSS,
+ 1083662.400000ns, VDD,
+ 1087985.900000ns, VDD,
+ 1087986.000000ns, VSS,
+ 1088106.000000ns, VSS,
+ 1088106.100000ns, VDD,
+ 1089667.300000ns, VDD,
+ 1089667.400000ns, VSS,
+ 1089787.400000ns, VSS,
+ 1089787.500000ns, VDD,
+ 1090027.600000ns, VDD,
+ 1090027.700000ns, VSS,
+ 1090508.000000ns, VSS,
+ 1090508.100000ns, VDD,
+ 1090988.400000ns, VDD,
+ 1090988.500000ns, VSS,
+ 1092429.600000ns, VSS,
+ 1092429.700000ns, VDD,
+ 1092910.000000ns, VDD,
+ 1092910.100000ns, VSS,
+ 1093030.100000ns, VSS,
+ 1093030.200000ns, VDD,
+ 1093150.200000ns, VDD,
+ 1093150.300000ns, VSS,
+ 1094351.200000ns, VSS,
+ 1094351.300000ns, VDD,
+ 1094831.600000ns, VDD,
+ 1094831.700000ns, VSS,
+ 1096032.600000ns, VSS,
+ 1096032.700000ns, VDD,
+ 1096392.900000ns, VDD,
+ 1096393.000000ns, VSS,
+ 1096753.200000ns, VSS,
+ 1096753.300000ns, VDD,
+ 1098194.400000ns, VDD,
+ 1098194.500000ns, VSS,
+ 1098434.600000ns, VSS,
+ 1098434.700000ns, VDD,
+ 1099155.200000ns, VDD,
+ 1099155.300000ns, VSS,
+ 1099395.400000ns, VSS,
+ 1099395.500000ns, VDD,
+ 1099515.500000ns, VDD,
+ 1099515.600000ns, VSS,
+ 1099635.600000ns, VSS,
+ 1099635.700000ns, VDD,
+ 1100476.300000ns, VDD,
+ 1100476.400000ns, VSS,
+ 1100836.600000ns, VSS,
+ 1100836.700000ns, VDD,
+ 1101196.900000ns, VDD,
+ 1101197.000000ns, VSS,
+ 1101677.300000ns, VSS,
+ 1101677.400000ns, VDD,
+ 1102758.200000ns, VDD,
+ 1102758.300000ns, VSS,
+ 1103478.800000ns, VSS,
+ 1103478.900000ns, VDD,
+ 1103598.900000ns, VDD,
+ 1103599.000000ns, VSS,
+ 1104079.300000ns, VSS,
+ 1104079.400000ns, VDD,
+ 1104799.900000ns, VDD,
+ 1104800.000000ns, VSS,
+ 1105280.300000ns, VSS,
+ 1105280.400000ns, VDD,
+ 1105760.700000ns, VDD,
+ 1105760.800000ns, VSS,
+ 1106241.100000ns, VSS,
+ 1106241.200000ns, VDD,
+ 1106721.500000ns, VDD,
+ 1106721.600000ns, VSS,
+ 1107922.500000ns, VSS,
+ 1107922.600000ns, VDD,
+ 1108282.800000ns, VDD,
+ 1108282.900000ns, VSS,
+ 1108643.100000ns, VSS,
+ 1108643.200000ns, VDD,
+ 1110684.800000ns, VDD,
+ 1110684.900000ns, VSS,
+ 1111765.700000ns, VSS,
+ 1111765.800000ns, VDD,
+ 1112606.400000ns, VDD,
+ 1112606.500000ns, VSS,
+ 1112966.700000ns, VSS,
+ 1112966.800000ns, VDD,
+ 1113086.800000ns, VDD,
+ 1113086.900000ns, VSS,
+ 1113447.100000ns, VSS,
+ 1113447.200000ns, VDD,
+ 1113567.200000ns, VDD,
+ 1113567.300000ns, VSS,
+ 1114167.700000ns, VSS,
+ 1114167.800000ns, VDD,
+ 1114648.100000ns, VDD,
+ 1114648.200000ns, VSS,
+ 1115128.500000ns, VSS,
+ 1115128.600000ns, VDD,
+ 1115969.200000ns, VDD,
+ 1115969.300000ns, VSS,
+ 1116449.600000ns, VSS,
+ 1116449.700000ns, VDD,
+ 1116569.700000ns, VDD,
+ 1116569.800000ns, VSS,
+ 1116689.800000ns, VSS,
+ 1116689.900000ns, VDD,
+ 1116809.900000ns, VDD,
+ 1116810.000000ns, VSS,
+ 1117770.700000ns, VSS,
+ 1117770.800000ns, VDD,
+ 1118010.900000ns, VDD,
+ 1118011.000000ns, VSS,
+ 1118251.100000ns, VSS,
+ 1118251.200000ns, VDD,
+ 1118371.200000ns, VDD,
+ 1118371.300000ns, VSS,
+ 1118851.600000ns, VSS,
+ 1118851.700000ns, VDD,
+ 1119332.000000ns, VDD,
+ 1119332.100000ns, VSS,
+ 1119452.100000ns, VSS,
+ 1119452.200000ns, VDD,
+ 1119572.200000ns, VDD,
+ 1119572.300000ns, VSS,
+ 1119812.400000ns, VSS,
+ 1119812.500000ns, VDD,
+ 1121013.400000ns, VDD,
+ 1121013.500000ns, VSS,
+ 1121373.700000ns, VSS,
+ 1121373.800000ns, VDD,
+ 1121974.200000ns, VDD,
+ 1121974.300000ns, VSS,
+ 1122094.300000ns, VSS,
+ 1122094.400000ns, VDD,
+ 1124136.000000ns, VDD,
+ 1124136.100000ns, VSS,
+ 1124736.500000ns, VSS,
+ 1124736.600000ns, VDD,
+ 1125937.500000ns, VDD,
+ 1125937.600000ns, VSS,
+ 1126297.800000ns, VSS,
+ 1126297.900000ns, VDD,
+ 1128099.300000ns, VDD,
+ 1128099.400000ns, VSS,
+ 1128219.400000ns, VSS,
+ 1128219.500000ns, VDD,
+ 1128579.700000ns, VDD,
+ 1128579.800000ns, VSS,
+ 1130141.000000ns, VSS,
+ 1130141.100000ns, VDD,
+ 1131101.800000ns, VDD,
+ 1131101.900000ns, VSS,
+ 1131221.900000ns, VSS,
+ 1131222.000000ns, VDD,
+ 1131942.500000ns, VDD,
+ 1131942.600000ns, VSS,
+ 1133143.500000ns, VSS,
+ 1133143.600000ns, VDD,
+ 1133383.700000ns, VDD,
+ 1133383.800000ns, VSS,
+ 1133623.900000ns, VSS,
+ 1133624.000000ns, VDD,
+ 1133984.200000ns, VDD,
+ 1133984.300000ns, VSS,
+ 1134464.600000ns, VSS,
+ 1134464.700000ns, VDD,
+ 1134704.800000ns, VDD,
+ 1134704.900000ns, VSS,
+ 1135545.500000ns, VSS,
+ 1135545.600000ns, VDD,
+ 1136386.200000ns, VDD,
+ 1136386.300000ns, VSS,
+ 1136866.600000ns, VSS,
+ 1136866.700000ns, VDD,
+ 1137347.000000ns, VDD,
+ 1137347.100000ns, VSS,
+ 1137827.400000ns, VSS,
+ 1137827.500000ns, VDD,
+ 1138067.600000ns, VDD,
+ 1138067.700000ns, VSS,
+ 1138187.700000ns, VSS,
+ 1138187.800000ns, VDD,
+ 1140349.500000ns, VDD,
+ 1140349.600000ns, VSS,
+ 1140709.800000ns, VSS,
+ 1140709.900000ns, VDD,
+ 1141310.300000ns, VDD,
+ 1141310.400000ns, VSS,
+ 1141670.600000ns, VSS,
+ 1141670.700000ns, VDD,
+ 1142271.100000ns, VDD,
+ 1142271.200000ns, VSS,
+ 1142391.200000ns, VSS,
+ 1142391.300000ns, VDD,
+ 1143712.300000ns, VDD,
+ 1143712.400000ns, VSS,
+ 1143952.500000ns, VSS,
+ 1143952.600000ns, VDD,
+ 1144673.100000ns, VDD,
+ 1144673.200000ns, VSS,
+ 1145513.800000ns, VSS,
+ 1145513.900000ns, VDD,
+ 1147075.100000ns, VDD,
+ 1147075.200000ns, VSS,
+ 1150558.000000ns, VSS,
+ 1150558.100000ns, VDD,
+ 1150678.100000ns, VDD,
+ 1150678.200000ns, VSS,
+ 1150798.200000ns, VSS,
+ 1150798.300000ns, VDD,
+ 1151158.500000ns, VDD,
+ 1151158.600000ns, VSS,
+ 1153800.700000ns, VSS,
+ 1153800.800000ns, VDD,
+ 1154521.300000ns, VDD,
+ 1154521.400000ns, VSS,
+ 1154641.400000ns, VSS,
+ 1154641.500000ns, VDD,
+ 1154761.500000ns, VDD,
+ 1154761.600000ns, VSS,
+ 1155241.900000ns, VSS,
+ 1155242.000000ns, VDD,
+ 1156082.600000ns, VDD,
+ 1156082.700000ns, VSS,
+ 1156563.000000ns, VSS,
+ 1156563.100000ns, VDD,
+ 1157043.400000ns, VDD,
+ 1157043.500000ns, VSS,
+ 1157283.600000ns, VSS,
+ 1157283.700000ns, VDD,
+ 1157523.800000ns, VDD,
+ 1157523.900000ns, VSS,
+ 1159085.100000ns, VSS,
+ 1159085.200000ns, VDD,
+ 1159445.400000ns, VDD,
+ 1159445.500000ns, VSS,
+ 1159685.600000ns, VSS,
+ 1159685.700000ns, VDD,
+ 1161607.200000ns, VDD,
+ 1161607.300000ns, VSS,
+ 1162327.800000ns, VSS,
+ 1162327.900000ns, VDD,
+ 1162568.000000ns, VDD,
+ 1162568.100000ns, VSS,
+ 1162688.100000ns, VSS,
+ 1162688.200000ns, VDD,
+ 1163048.400000ns, VDD,
+ 1163048.500000ns, VSS,
+ 1163168.500000ns, VSS,
+ 1163168.600000ns, VDD,
+ 1164849.900000ns, VDD,
+ 1164850.000000ns, VSS,
+ 1164970.000000ns, VSS,
+ 1164970.100000ns, VDD,
+ 1165690.600000ns, VDD,
+ 1165690.700000ns, VSS,
+ 1166771.500000ns, VSS,
+ 1166771.600000ns, VDD,
+ 1167732.300000ns, VDD,
+ 1167732.400000ns, VSS,
+ 1168212.700000ns, VSS,
+ 1168212.800000ns, VDD,
+ 1168813.200000ns, VDD,
+ 1168813.300000ns, VSS,
+ 1170134.300000ns, VSS,
+ 1170134.400000ns, VDD,
+ 1171095.100000ns, VDD,
+ 1171095.200000ns, VSS,
+ 1171335.300000ns, VSS,
+ 1171335.400000ns, VDD,
+ 1171455.400000ns, VDD,
+ 1171455.500000ns, VSS,
+ 1171575.500000ns, VSS,
+ 1171575.600000ns, VDD,
+ 1173016.700000ns, VDD,
+ 1173016.800000ns, VSS,
+ 1173377.000000ns, VSS,
+ 1173377.100000ns, VDD,
+ 1173737.300000ns, VDD,
+ 1173737.400000ns, VSS,
+ 1174097.600000ns, VSS,
+ 1174097.700000ns, VDD,
+ 1174337.800000ns, VDD,
+ 1174337.900000ns, VSS,
+ 1174457.900000ns, VSS,
+ 1174458.000000ns, VDD,
+ 1174578.000000ns, VDD,
+ 1174578.100000ns, VSS,
+ 1175418.700000ns, VSS,
+ 1175418.800000ns, VDD,
+ 1176019.200000ns, VDD,
+ 1176019.300000ns, VSS,
+ 1176499.600000ns, VSS,
+ 1176499.700000ns, VDD,
+ 1176619.700000ns, VDD,
+ 1176619.800000ns, VSS,
+ 1178661.400000ns, VSS,
+ 1178661.500000ns, VDD,
+ 1178781.500000ns, VDD,
+ 1178781.600000ns, VSS,
+ 1178901.600000ns, VSS,
+ 1178901.700000ns, VDD,
+ 1179382.000000ns, VDD,
+ 1179382.100000ns, VSS,
+ 1179502.100000ns, VSS,
+ 1179502.200000ns, VDD,
+ 1180462.900000ns, VDD,
+ 1180463.000000ns, VSS,
+ 1181303.600000ns, VSS,
+ 1181303.700000ns, VDD,
+ 1181904.100000ns, VDD,
+ 1181904.200000ns, VSS,
+ 1182384.500000ns, VSS,
+ 1182384.600000ns, VDD,
+ 1182744.800000ns, VDD,
+ 1182744.900000ns, VSS,
+ 1183345.300000ns, VSS,
+ 1183345.400000ns, VDD,
+ 1183705.600000ns, VDD,
+ 1183705.700000ns, VSS,
+ 1183945.800000ns, VSS,
+ 1183945.900000ns, VDD,
+ 1184426.200000ns, VDD,
+ 1184426.300000ns, VSS,
+ 1184666.400000ns, VSS,
+ 1184666.500000ns, VDD,
+ 1185146.800000ns, VDD,
+ 1185146.900000ns, VSS,
+ 1185747.300000ns, VSS,
+ 1185747.400000ns, VDD,
+ 1186347.800000ns, VDD,
+ 1186347.900000ns, VSS,
+ 1187308.600000ns, VSS,
+ 1187308.700000ns, VDD,
+ 1187789.000000ns, VDD,
+ 1187789.100000ns, VSS,
+ 1188869.900000ns, VSS,
+ 1188870.000000ns, VDD,
+ 1190551.300000ns, VDD,
+ 1190551.400000ns, VSS,
+ 1190911.600000ns, VSS,
+ 1190911.700000ns, VDD,
+ 1191031.700000ns, VDD,
+ 1191031.800000ns, VSS,
+ 1191271.900000ns, VSS,
+ 1191272.000000ns, VDD,
+ 1191392.000000ns, VDD,
+ 1191392.100000ns, VSS,
+ 1191512.100000ns, VSS,
+ 1191512.200000ns, VDD,
+ 1192352.800000ns, VDD,
+ 1192352.900000ns, VSS,
+ 1192833.200000ns, VSS,
+ 1192833.300000ns, VDD,
+ 1193193.500000ns, VDD,
+ 1193193.600000ns, VSS,
+ 1193914.100000ns, VSS,
+ 1193914.200000ns, VDD,
+ 1194514.600000ns, VDD,
+ 1194514.700000ns, VSS,
+ 1194754.800000ns, VSS,
+ 1194754.900000ns, VDD,
+ 1194995.000000ns, VDD,
+ 1194995.100000ns, VSS,
+ 1195235.200000ns, VSS,
+ 1195235.300000ns, VDD,
+ 1195475.400000ns, VDD,
+ 1195475.500000ns, VSS,
+ 1195715.600000ns, VSS,
+ 1195715.700000ns, VDD,
+ 1196316.100000ns, VDD,
+ 1196316.200000ns, VSS,
+ 1196676.400000ns, VSS,
+ 1196676.500000ns, VDD,
+ 1197156.800000ns, VDD,
+ 1197156.900000ns, VSS,
+ 1197276.900000ns, VSS,
+ 1197277.000000ns, VDD,
+ 1198598.000000ns, VDD,
+ 1198598.100000ns, VSS,
+ 1199198.500000ns, VSS,
+ 1199198.600000ns, VDD,
+ 1201480.400000ns, VDD,
+ 1201480.500000ns, VSS,
+ 1201960.800000ns, VSS,
+ 1201960.900000ns, VDD,
+ 1202080.900000ns, VDD,
+ 1202081.000000ns, VSS,
+ 1202201.000000ns, VSS,
+ 1202201.100000ns, VDD,
+ 1202441.200000ns, VDD,
+ 1202441.300000ns, VSS,
+ 1202561.300000ns, VSS,
+ 1202561.400000ns, VDD,
+ 1203041.700000ns, VDD,
+ 1203041.800000ns, VSS,
+ 1203882.400000ns, VSS,
+ 1203882.500000ns, VDD,
+ 1205083.400000ns, VDD,
+ 1205083.500000ns, VSS,
+ 1205804.000000ns, VSS,
+ 1205804.100000ns, VDD,
+ 1205924.100000ns, VDD,
+ 1205924.200000ns, VSS,
+ 1206044.200000ns, VSS,
+ 1206044.300000ns, VDD,
+ 1206284.400000ns, VDD,
+ 1206284.500000ns, VSS,
+ 1206644.700000ns, VSS,
+ 1206644.800000ns, VDD,
+ 1207365.300000ns, VDD,
+ 1207365.400000ns, VSS,
+ 1207965.800000ns, VSS,
+ 1207965.900000ns, VDD,
+ 1208206.000000ns, VDD,
+ 1208206.100000ns, VSS,
+ 1209046.700000ns, VSS,
+ 1209046.800000ns, VDD,
+ 1210608.000000ns, VDD,
+ 1210608.100000ns, VSS,
+ 1211328.600000ns, VSS,
+ 1211328.700000ns, VDD,
+ 1211568.800000ns, VDD,
+ 1211568.900000ns, VSS,
+ 1212049.200000ns, VSS,
+ 1212049.300000ns, VDD,
+ 1212169.300000ns, VDD,
+ 1212169.400000ns, VSS,
+ 1213850.700000ns, VSS,
+ 1213850.800000ns, VDD,
+ 1214331.100000ns, VDD,
+ 1214331.200000ns, VSS,
+ 1215291.900000ns, VSS,
+ 1215292.000000ns, VDD,
+ 1216012.500000ns, VDD,
+ 1216012.600000ns, VSS,
+ 1216492.900000ns, VSS,
+ 1216493.000000ns, VDD,
+ 1217213.500000ns, VDD,
+ 1217213.600000ns, VSS,
+ 1217573.800000ns, VSS,
+ 1217573.900000ns, VDD,
+ 1218294.400000ns, VDD,
+ 1218294.500000ns, VSS,
+ 1218774.800000ns, VSS,
+ 1218774.900000ns, VDD,
+ 1219255.200000ns, VDD,
+ 1219255.300000ns, VSS,
+ 1220336.100000ns, VSS,
+ 1220336.200000ns, VDD,
+ 1220816.500000ns, VDD,
+ 1220816.600000ns, VSS,
+ 1221056.700000ns, VSS,
+ 1221056.800000ns, VDD,
+ 1221657.200000ns, VDD,
+ 1221657.300000ns, VSS,
+ 1222257.700000ns, VSS,
+ 1222257.800000ns, VDD,
+ 1223698.900000ns, VDD,
+ 1223699.000000ns, VSS,
+ 1224419.500000ns, VSS,
+ 1224419.600000ns, VDD,
+ 1224539.600000ns, VDD,
+ 1224539.700000ns, VSS,
+ 1224899.900000ns, VSS,
+ 1224900.000000ns, VDD,
+ 1226341.100000ns, VDD,
+ 1226341.200000ns, VSS,
+ 1226821.500000ns, VSS,
+ 1226821.600000ns, VDD,
+ 1228142.600000ns, VDD,
+ 1228142.700000ns, VSS,
+ 1228623.000000ns, VSS,
+ 1228623.100000ns, VDD,
+ 1228743.100000ns, VDD,
+ 1228743.200000ns, VSS,
+ 1229223.500000ns, VSS,
+ 1229223.600000ns, VDD,
+ 1229703.900000ns, VDD,
+ 1229704.000000ns, VSS,
+ 1229824.000000ns, VSS,
+ 1229824.100000ns, VDD,
+ 1230424.500000ns, VDD,
+ 1230424.600000ns, VSS,
+ 1232105.900000ns, VSS,
+ 1232106.000000ns, VDD,
+ 1232226.000000ns, VDD,
+ 1232226.100000ns, VSS,
+ 1233186.800000ns, VSS,
+ 1233186.900000ns, VDD,
+ 1233787.300000ns, VDD,
+ 1233787.400000ns, VSS,
+ 1235228.500000ns, VSS,
+ 1235228.600000ns, VDD,
+ 1235949.100000ns, VDD,
+ 1235949.200000ns, VSS,
+ 1236069.200000ns, VSS,
+ 1236069.300000ns, VDD,
+ 1236429.500000ns, VDD,
+ 1236429.600000ns, VSS,
+ 1237030.000000ns, VSS,
+ 1237030.100000ns, VDD,
+ 1237150.100000ns, VDD,
+ 1237150.200000ns, VSS,
+ 1237270.200000ns, VSS,
+ 1237270.300000ns, VDD,
+ 1237750.600000ns, VDD,
+ 1237750.700000ns, VSS,
+ 1237870.700000ns, VSS,
+ 1237870.800000ns, VDD,
+ 1237990.800000ns, VDD,
+ 1237990.900000ns, VSS,
+ 1238110.900000ns, VSS,
+ 1238111.000000ns, VDD,
+ 1239071.700000ns, VDD,
+ 1239071.800000ns, VSS,
+ 1239552.100000ns, VSS,
+ 1239552.200000ns, VDD,
+ 1239912.400000ns, VDD,
+ 1239912.500000ns, VSS,
+ 1240272.700000ns, VSS,
+ 1240272.800000ns, VDD,
+ 1241233.500000ns, VDD,
+ 1241233.600000ns, VSS,
+ 1241473.700000ns, VSS,
+ 1241473.800000ns, VDD,
+ 1241834.000000ns, VDD,
+ 1241834.100000ns, VSS,
+ 1243995.800000ns, VSS,
+ 1243995.900000ns, VDD,
+ 1244236.000000ns, VDD,
+ 1244236.100000ns, VSS,
+ 1245076.700000ns, VSS,
+ 1245076.800000ns, VDD,
+ 1245557.100000ns, VDD,
+ 1245557.200000ns, VSS,
+ 1245797.300000ns, VSS,
+ 1245797.400000ns, VDD,
+ 1246037.500000ns, VDD,
+ 1246037.600000ns, VSS,
+ 1248559.600000ns, VSS,
+ 1248559.700000ns, VDD,
+ 1249160.100000ns, VDD,
+ 1249160.200000ns, VSS,
+ 1251201.800000ns, VSS,
+ 1251201.900000ns, VDD,
+ 1251682.200000ns, VDD,
+ 1251682.300000ns, VSS,
+ 1252162.600000ns, VSS,
+ 1252162.700000ns, VDD,
+ 1252643.000000ns, VDD,
+ 1252643.100000ns, VSS,
+ 1254204.300000ns, VSS,
+ 1254204.400000ns, VDD,
+ 1254924.900000ns, VDD,
+ 1254925.000000ns, VSS,
+ 1256366.100000ns, VSS,
+ 1256366.200000ns, VDD,
+ 1256606.300000ns, VDD,
+ 1256606.400000ns, VSS,
+ 1256846.500000ns, VSS,
+ 1256846.600000ns, VDD,
+ 1258407.800000ns, VDD,
+ 1258407.900000ns, VSS,
+ 1259488.700000ns, VSS,
+ 1259488.800000ns, VDD,
+ 1261170.100000ns, VDD,
+ 1261170.200000ns, VSS,
+ 1261650.500000ns, VSS,
+ 1261650.600000ns, VDD,
+ 1261770.600000ns, VDD,
+ 1261770.700000ns, VSS,
+ 1262130.900000ns, VSS,
+ 1262131.000000ns, VDD,
+ 1262731.400000ns, VDD,
+ 1262731.500000ns, VSS,
+ 1263211.800000ns, VSS,
+ 1263211.900000ns, VDD,
+ 1263812.300000ns, VDD,
+ 1263812.400000ns, VSS,
+ 1264052.500000ns, VSS,
+ 1264052.600000ns, VDD,
+ 1264172.600000ns, VDD,
+ 1264172.700000ns, VSS,
+ 1265133.400000ns, VSS,
+ 1265133.500000ns, VDD,
+ 1265253.500000ns, VDD,
+ 1265253.600000ns, VSS,
+ 1265974.100000ns, VSS,
+ 1265974.200000ns, VDD,
+ 1266334.400000ns, VDD,
+ 1266334.500000ns, VSS,
+ 1266814.800000ns, VSS,
+ 1266814.900000ns, VDD,
+ 1266934.900000ns, VDD,
+ 1266935.000000ns, VSS,
+ 1267175.100000ns, VSS,
+ 1267175.200000ns, VDD,
+ 1267295.200000ns, VDD,
+ 1267295.300000ns, VSS,
+ 1267775.600000ns, VSS,
+ 1267775.700000ns, VDD,
+ 1268015.800000ns, VDD,
+ 1268015.900000ns, VSS,
+ 1268256.000000ns, VSS,
+ 1268256.100000ns, VDD,
+ 1269216.800000ns, VDD,
+ 1269216.900000ns, VSS,
+ 1269336.900000ns, VSS,
+ 1269337.000000ns, VDD,
+ 1269457.000000ns, VDD,
+ 1269457.100000ns, VSS,
+ 1269577.100000ns, VSS,
+ 1269577.200000ns, VDD,
+ 1270297.700000ns, VDD,
+ 1270297.800000ns, VSS,
+ 1270778.100000ns, VSS,
+ 1270778.200000ns, VDD,
+ 1271498.700000ns, VDD,
+ 1271498.800000ns, VSS,
+ 1271618.800000ns, VSS,
+ 1271618.900000ns, VDD,
+ 1271738.900000ns, VDD,
+ 1271739.000000ns, VSS,
+ 1272219.300000ns, VSS,
+ 1272219.400000ns, VDD,
+ 1272459.500000ns, VDD,
+ 1272459.600000ns, VSS,
+ 1273540.400000ns, VSS,
+ 1273540.500000ns, VDD,
+ 1273660.500000ns, VDD,
+ 1273660.600000ns, VSS,
+ 1273780.600000ns, VSS,
+ 1273780.700000ns, VDD,
+ 1275341.900000ns, VDD,
+ 1275342.000000ns, VSS,
+ 1277023.300000ns, VSS,
+ 1277023.400000ns, VDD,
+ 1277503.700000ns, VDD,
+ 1277503.800000ns, VSS,
+ 1278104.200000ns, VSS,
+ 1278104.300000ns, VDD,
+ 1278584.600000ns, VDD,
+ 1278584.700000ns, VSS,
+ 1279905.700000ns, VSS,
+ 1279905.800000ns, VDD,
+ 1280986.600000ns, VDD,
+ 1280986.700000ns, VSS,
+ 1281587.100000ns, VSS,
+ 1281587.200000ns, VDD,
+ 1281947.400000ns, VDD,
+ 1281947.500000ns, VSS,
+ 1283508.700000ns, VSS,
+ 1283508.800000ns, VDD,
+ 1284589.600000ns, VDD,
+ 1284589.700000ns, VSS,
+ 1286271.000000ns, VSS,
+ 1286271.100000ns, VDD,
+ 1287111.700000ns, VDD,
+ 1287111.800000ns, VSS,
+ 1288552.900000ns, VSS,
+ 1288553.000000ns, VDD,
+ 1289033.300000ns, VDD,
+ 1289033.400000ns, VSS,
+ 1289393.600000ns, VSS,
+ 1289393.700000ns, VDD,
+ 1289994.100000ns, VDD,
+ 1289994.200000ns, VSS,
+ 1290834.800000ns, VSS,
+ 1290834.900000ns, VDD,
+ 1291555.400000ns, VDD,
+ 1291555.500000ns, VSS,
+ 1291795.600000ns, VSS,
+ 1291795.700000ns, VDD,
+ 1292276.000000ns, VDD,
+ 1292276.100000ns, VSS,
+ 1293356.900000ns, VSS,
+ 1293357.000000ns, VDD,
+ 1295038.300000ns, VDD,
+ 1295038.400000ns, VSS,
+ 1295518.700000ns, VSS,
+ 1295518.800000ns, VDD,
+ 1295638.800000ns, VDD,
+ 1295638.900000ns, VSS,
+ 1295758.900000ns, VSS,
+ 1295759.000000ns, VDD,
+ 1297320.200000ns, VDD,
+ 1297320.300000ns, VSS,
+ 1298881.500000ns, VSS,
+ 1298881.600000ns, VDD,
+ 1299001.600000ns, VDD,
+ 1299001.700000ns, VSS,
+ 1299722.200000ns, VSS,
+ 1299722.300000ns, VDD,
+ 1300562.900000ns, VDD,
+ 1300563.000000ns, VSS,
+ 1301043.300000ns, VSS,
+ 1301043.400000ns, VDD,
+ 1301523.700000ns, VDD,
+ 1301523.800000ns, VSS,
+ 1302244.300000ns, VSS,
+ 1302244.400000ns, VDD,
+ 1302484.500000ns, VDD,
+ 1302484.600000ns, VSS,
+ 1304886.500000ns, VSS,
+ 1304886.600000ns, VDD,
+ 1305727.200000ns, VDD,
+ 1305727.300000ns, VSS,
+ 1306087.500000ns, VSS,
+ 1306087.600000ns, VDD,
+ 1306928.200000ns, VDD,
+ 1306928.300000ns, VSS,
+ 1308129.200000ns, VSS,
+ 1308129.300000ns, VDD,
+ 1308489.500000ns, VDD,
+ 1308489.600000ns, VSS,
+ 1308969.900000ns, VSS,
+ 1308970.000000ns, VDD,
+ 1310291.000000ns, VDD,
+ 1310291.100000ns, VSS,
+ 1310891.500000ns, VSS,
+ 1310891.600000ns, VDD,
+ 1312933.200000ns, VDD,
+ 1312933.300000ns, VSS,
+ 1313413.600000ns, VSS,
+ 1313413.700000ns, VDD,
+ 1313773.900000ns, VDD,
+ 1313774.000000ns, VSS,
+ 1314614.600000ns, VSS,
+ 1314614.700000ns, VDD,
+ 1315455.300000ns, VDD,
+ 1315455.400000ns, VSS,
+ 1315935.700000ns, VSS,
+ 1315935.800000ns, VDD,
+ 1317256.800000ns, VDD,
+ 1317256.900000ns, VSS,
+ 1318217.600000ns, VSS,
+ 1318217.700000ns, VDD,
+ 1318337.700000ns, VDD,
+ 1318337.800000ns, VSS,
+ 1319058.300000ns, VSS,
+ 1319058.400000ns, VDD,
+ 1319418.600000ns, VDD,
+ 1319418.700000ns, VSS,
+ 1319538.700000ns, VSS,
+ 1319538.800000ns, VDD,
+ 1320019.100000ns, VDD,
+ 1320019.200000ns, VSS,
+ 1320499.500000ns, VSS,
+ 1320499.600000ns, VDD,
+ 1321580.400000ns, VDD,
+ 1321580.500000ns, VSS,
+ 1321820.600000ns, VSS,
+ 1321820.700000ns, VDD,
+ 1322421.100000ns, VDD,
+ 1322421.200000ns, VSS,
+ 1322901.500000ns, VSS,
+ 1322901.600000ns, VDD,
+ 1324462.800000ns, VDD,
+ 1324462.900000ns, VSS,
+ 1326744.700000ns, VSS,
+ 1326744.800000ns, VDD,
+ 1326864.800000ns, VDD,
+ 1326864.900000ns, VSS,
+ 1326984.900000ns, VSS,
+ 1326985.000000ns, VDD,
+ 1327225.100000ns, VDD,
+ 1327225.200000ns, VSS,
+ 1327465.300000ns, VSS,
+ 1327465.400000ns, VDD,
+ 1327585.400000ns, VDD,
+ 1327585.500000ns, VSS,
+ 1327945.700000ns, VSS,
+ 1327945.800000ns, VDD,
+ 1328426.100000ns, VDD,
+ 1328426.200000ns, VSS,
+ 1328546.200000ns, VSS,
+ 1328546.300000ns, VDD,
+ 1328906.500000ns, VDD,
+ 1328906.600000ns, VSS,
+ 1330107.500000ns, VSS,
+ 1330107.600000ns, VDD,
+ 1330467.800000ns, VDD,
+ 1330467.900000ns, VSS,
+ 1330708.000000ns, VSS,
+ 1330708.100000ns, VDD,
+ 1331188.400000ns, VDD,
+ 1331188.500000ns, VSS,
+ 1331308.500000ns, VSS,
+ 1331308.600000ns, VDD,
+ 1332269.300000ns, VDD,
+ 1332269.400000ns, VSS,
+ 1333350.200000ns, VSS,
+ 1333350.300000ns, VDD,
+ 1333710.500000ns, VDD,
+ 1333710.600000ns, VSS,
+ 1335031.600000ns, VSS,
+ 1335031.700000ns, VDD,
+ 1335512.000000ns, VDD,
+ 1335512.100000ns, VSS,
+ 1335752.200000ns, VSS,
+ 1335752.300000ns, VDD,
+ 1336112.500000ns, VDD,
+ 1336112.600000ns, VSS,
+ 1336232.600000ns, VSS,
+ 1336232.700000ns, VDD,
+ 1337313.500000ns, VDD,
+ 1337313.600000ns, VSS,
+ 1337553.700000ns, VSS,
+ 1337553.800000ns, VDD,
+ 1338514.500000ns, VDD,
+ 1338514.600000ns, VSS,
+ 1338994.900000ns, VSS,
+ 1338995.000000ns, VDD,
+ 1339115.000000ns, VDD,
+ 1339115.100000ns, VSS,
+ 1339595.400000ns, VSS,
+ 1339595.500000ns, VDD,
+ 1340075.800000ns, VDD,
+ 1340075.900000ns, VSS,
+ 1340436.100000ns, VSS,
+ 1340436.200000ns, VDD,
+ 1340676.300000ns, VDD,
+ 1340676.400000ns, VSS,
+ 1341156.700000ns, VSS,
+ 1341156.800000ns, VDD,
+ 1341276.800000ns, VDD,
+ 1341276.900000ns, VSS,
+ 1341877.300000ns, VSS,
+ 1341877.400000ns, VDD,
+ 1342718.000000ns, VDD,
+ 1342718.100000ns, VSS,
+ 1343198.400000ns, VSS,
+ 1343198.500000ns, VDD,
+ 1343318.500000ns, VDD,
+ 1343318.600000ns, VSS,
+ 1343558.700000ns, VSS,
+ 1343558.800000ns, VDD,
+ 1345360.200000ns, VDD,
+ 1345360.300000ns, VSS,
+ 1345840.600000ns, VSS,
+ 1345840.700000ns, VDD,
+ 1347041.600000ns, VDD,
+ 1347041.700000ns, VSS,
+ 1347522.000000ns, VSS,
+ 1347522.100000ns, VDD,
+ 1348002.400000ns, VDD,
+ 1348002.500000ns, VSS,
+ 1348122.500000ns, VSS,
+ 1348122.600000ns, VDD,
+ 1348482.800000ns, VDD,
+ 1348482.900000ns, VSS,
+ 1349683.800000ns, VSS,
+ 1349683.900000ns, VDD,
+ 1350284.300000ns, VDD,
+ 1350284.400000ns, VSS,
+ 1351485.300000ns, VSS,
+ 1351485.400000ns, VDD,
+ 1351605.400000ns, VDD,
+ 1351605.500000ns, VSS,
+ 1351965.700000ns, VSS,
+ 1351965.800000ns, VDD,
+ 1352686.300000ns, VDD,
+ 1352686.400000ns, VSS,
+ 1353166.700000ns, VSS,
+ 1353166.800000ns, VDD,
+ 1353406.900000ns, VDD,
+ 1353407.000000ns, VSS,
+ 1353647.100000ns, VSS,
+ 1353647.200000ns, VDD,
+ 1353887.300000ns, VDD,
+ 1353887.400000ns, VSS,
+ 1354367.700000ns, VSS,
+ 1354367.800000ns, VDD,
+ 1355929.000000ns, VDD,
+ 1355929.100000ns, VSS,
+ 1356289.300000ns, VSS,
+ 1356289.400000ns, VDD,
+ 1357250.100000ns, VDD,
+ 1357250.200000ns, VSS,
+ 1357730.500000ns, VSS,
+ 1357730.600000ns, VDD,
+ 1357850.600000ns, VDD,
+ 1357850.700000ns, VSS,
+ 1357970.700000ns, VSS,
+ 1357970.800000ns, VDD,
+ 1359532.000000ns, VDD,
+ 1359532.100000ns, VSS,
+ 1361693.800000ns, VSS,
+ 1361693.900000ns, VDD,
+ 1362534.500000ns, VDD,
+ 1362534.600000ns, VSS,
+ 1363255.100000ns, VSS,
+ 1363255.200000ns, VDD,
+ 1363975.700000ns, VDD,
+ 1363975.800000ns, VSS,
+ 1364696.300000ns, VSS,
+ 1364696.400000ns, VDD,
+ 1365176.700000ns, VDD,
+ 1365176.800000ns, VSS,
+ 1365537.000000ns, VSS,
+ 1365537.100000ns, VDD,
+ 1366497.800000ns, VDD,
+ 1366497.900000ns, VSS,
+ 1366617.900000ns, VSS,
+ 1366618.000000ns, VDD,
+ 1366978.200000ns, VDD,
+ 1366978.300000ns, VSS,
+ 1369380.200000ns, VSS,
+ 1369380.300000ns, VDD,
+ 1369620.400000ns, VDD,
+ 1369620.500000ns, VSS,
+ 1370461.100000ns, VSS,
+ 1370461.200000ns, VDD,
+ 1370581.200000ns, VDD,
+ 1370581.300000ns, VSS,
+ 1371662.100000ns, VSS,
+ 1371662.200000ns, VDD,
+ 1372983.200000ns, VDD,
+ 1372983.300000ns, VSS,
+ 1373463.600000ns, VSS,
+ 1373463.700000ns, VDD,
+ 1373823.900000ns, VDD,
+ 1373824.000000ns, VSS,
+ 1374784.700000ns, VSS,
+ 1374784.800000ns, VDD,
+ 1375505.300000ns, VDD,
+ 1375505.400000ns, VSS,
+ 1375745.500000ns, VSS,
+ 1375745.600000ns, VDD,
+ 1375985.700000ns, VDD,
+ 1375985.800000ns, VSS,
+ 1376105.800000ns, VSS,
+ 1376105.900000ns, VDD,
+ 1377186.700000ns, VDD,
+ 1377186.800000ns, VSS,
+ 1377667.100000ns, VSS,
+ 1377667.200000ns, VDD,
+ 1379108.300000ns, VDD,
+ 1379108.400000ns, VSS,
+ 1379708.800000ns, VSS,
+ 1379708.900000ns, VDD,
+ 1380789.700000ns, VDD,
+ 1380789.800000ns, VSS,
+ 1381029.900000ns, VSS,
+ 1381030.000000ns, VDD,
+ 1381150.000000ns, VDD,
+ 1381150.100000ns, VSS,
+ 1381270.100000ns, VSS,
+ 1381270.200000ns, VDD,
+ 1382351.000000ns, VDD,
+ 1382351.100000ns, VSS,
+ 1383191.700000ns, VSS,
+ 1383191.800000ns, VDD,
+ 1383672.100000ns, VDD,
+ 1383672.200000ns, VSS,
+ 1385713.800000ns, VSS,
+ 1385713.900000ns, VDD,
+ 1386074.100000ns, VDD,
+ 1386074.200000ns, VSS,
+ 1387515.300000ns, VSS,
+ 1387515.400000ns, VDD,
+ 1387875.600000ns, VDD,
+ 1387875.700000ns, VSS,
+ 1388235.900000ns, VSS,
+ 1388236.000000ns, VDD,
+ 1389196.700000ns, VDD,
+ 1389196.800000ns, VSS,
+ 1389677.100000ns, VSS,
+ 1389677.200000ns, VDD,
+ 1390157.500000ns, VDD,
+ 1390157.600000ns, VSS,
+ 1390998.200000ns, VSS,
+ 1390998.300000ns, VDD,
+ 1391959.000000ns, VDD,
+ 1391959.100000ns, VSS,
+ 1392319.300000ns, VSS,
+ 1392319.400000ns, VDD,
+ 1392679.600000ns, VDD,
+ 1392679.700000ns, VSS,
+ 1392919.800000ns, VSS,
+ 1392919.900000ns, VDD,
+ 1393160.000000ns, VDD,
+ 1393160.100000ns, VSS,
+ 1393400.200000ns, VSS,
+ 1393400.300000ns, VDD,
+ 1394721.300000ns, VDD,
+ 1394721.400000ns, VSS,
+ 1395441.900000ns, VSS,
+ 1395442.000000ns, VDD,
+ 1395922.300000ns, VDD,
+ 1395922.400000ns, VSS,
+ 1396162.500000ns, VSS,
+ 1396162.600000ns, VDD,
+ 1396402.700000ns, VDD,
+ 1396402.800000ns, VSS,
+ 1397003.200000ns, VSS,
+ 1397003.300000ns, VDD,
+ 1398324.300000ns, VDD,
+ 1398324.400000ns, VSS,
+ 1398684.600000ns, VSS,
+ 1398684.700000ns, VDD,
+ 1400245.900000ns, VDD,
+ 1400246.000000ns, VSS,
+ 1401086.600000ns, VSS,
+ 1401086.700000ns, VDD,
+ 1401687.100000ns, VDD,
+ 1401687.200000ns, VSS,
+ 1402167.500000ns, VSS,
+ 1402167.600000ns, VDD,
+ 1402407.700000ns, VDD,
+ 1402407.800000ns, VSS,
+ 1402647.900000ns, VSS,
+ 1402648.000000ns, VDD,
+ 1403248.400000ns, VDD,
+ 1403248.500000ns, VSS,
+ 1403848.900000ns, VSS,
+ 1403849.000000ns, VDD,
+ 1404569.500000ns, VDD,
+ 1404569.600000ns, VSS,
+ 1405650.400000ns, VSS,
+ 1405650.500000ns, VDD,
+ 1406491.100000ns, VDD,
+ 1406491.200000ns, VSS,
+ 1406971.500000ns, VSS,
+ 1406971.600000ns, VDD,
+ 1407211.700000ns, VDD,
+ 1407211.800000ns, VSS,
+ 1407451.900000ns, VSS,
+ 1407452.000000ns, VDD,
+ 1407572.000000ns, VDD,
+ 1407572.100000ns, VSS,
+ 1407932.300000ns, VSS,
+ 1407932.400000ns, VDD,
+ 1408412.700000ns, VDD,
+ 1408412.800000ns, VSS,
+ 1411775.500000ns, VSS,
+ 1411775.600000ns, VDD,
+ 1412856.400000ns, VDD,
+ 1412856.500000ns, VSS,
+ 1414778.000000ns, VSS,
+ 1414778.100000ns, VDD,
+ 1415498.600000ns, VDD,
+ 1415498.700000ns, VSS,
+ 1416459.400000ns, VSS,
+ 1416459.500000ns, VDD,
+ 1416579.500000ns, VDD,
+ 1416579.600000ns, VSS,
+ 1417420.200000ns, VSS,
+ 1417420.300000ns, VDD,
+ 1417660.400000ns, VDD,
+ 1417660.500000ns, VSS,
+ 1418140.800000ns, VSS,
+ 1418140.900000ns, VDD,
+ 1418861.400000ns, VDD,
+ 1418861.500000ns, VSS,
+ 1419221.700000ns, VSS,
+ 1419221.800000ns, VDD,
+ 1422464.400000ns, VDD,
+ 1422464.500000ns, VSS,
+ 1422824.700000ns, VSS,
+ 1422824.800000ns, VDD,
+ 1423545.300000ns, VDD,
+ 1423545.400000ns, VSS,
+ 1424025.700000ns, VSS,
+ 1424025.800000ns, VDD,
+ 1425587.000000ns, VDD,
+ 1425587.100000ns, VSS,
+ 1426187.500000ns, VSS,
+ 1426187.600000ns, VDD,
+ 1427028.200000ns, VDD,
+ 1427028.300000ns, VSS,
+ 1427148.300000ns, VSS,
+ 1427148.400000ns, VDD,
+ 1427268.400000ns, VDD,
+ 1427268.500000ns, VSS,
+ 1427628.700000ns, VSS,
+ 1427628.800000ns, VDD,
+ 1427868.900000ns, VDD,
+ 1427869.000000ns, VSS,
+ 1428229.200000ns, VSS,
+ 1428229.300000ns, VDD,
+ 1429190.000000ns, VDD,
+ 1429190.100000ns, VSS,
+ 1430150.800000ns, VSS,
+ 1430150.900000ns, VDD,
+ 1430631.200000ns, VDD,
+ 1430631.300000ns, VSS,
+ 1431111.600000ns, VSS,
+ 1431111.700000ns, VDD,
+ 1432192.500000ns, VDD,
+ 1432192.600000ns, VSS,
+ 1432432.700000ns, VSS,
+ 1432432.800000ns, VDD,
+ 1432672.900000ns, VDD,
+ 1432673.000000ns, VSS,
+ 1432793.000000ns, VSS,
+ 1432793.100000ns, VDD,
+ 1433513.600000ns, VDD,
+ 1433513.700000ns, VSS,
+ 1433633.700000ns, VSS,
+ 1433633.800000ns, VDD,
+ 1435074.900000ns, VDD,
+ 1435075.000000ns, VSS,
+ 1435675.400000ns, VSS,
+ 1435675.500000ns, VDD,
+ 1436275.900000ns, VDD,
+ 1436276.000000ns, VSS,
+ 1436756.300000ns, VSS,
+ 1436756.400000ns, VDD,
+ 1437116.600000ns, VDD,
+ 1437116.700000ns, VSS,
+ 1437236.700000ns, VSS,
+ 1437236.800000ns, VDD,
+ 1437957.300000ns, VDD,
+ 1437957.400000ns, VSS,
+ 1438317.600000ns, VSS,
+ 1438317.700000ns, VDD,
+ 1439518.600000ns, VDD,
+ 1439518.700000ns, VSS,
+ 1440959.800000ns, VSS,
+ 1440959.900000ns, VDD,
+ 1441320.100000ns, VDD,
+ 1441320.200000ns, VSS,
+ 1442280.900000ns, VSS,
+ 1442281.000000ns, VDD,
+ 1442521.100000ns, VDD,
+ 1442521.200000ns, VSS,
+ 1443842.200000ns, VSS,
+ 1443842.300000ns, VDD,
+ 1443962.300000ns, VDD,
+ 1443962.400000ns, VSS,
+ 1444202.500000ns, VSS,
+ 1444202.600000ns, VDD,
+ 1444803.000000ns, VDD,
+ 1444803.100000ns, VSS,
+ 1444923.100000ns, VSS,
+ 1444923.200000ns, VDD,
+ 1445163.300000ns, VDD,
+ 1445163.400000ns, VSS,
+ 1445283.400000ns, VSS,
+ 1445283.500000ns, VDD,
+ 1447205.000000ns, VDD,
+ 1447205.100000ns, VSS,
+ 1450327.600000ns, VSS,
+ 1450327.700000ns, VDD,
+ 1451048.200000ns, VDD,
+ 1451048.300000ns, VSS,
+ 1452129.100000ns, VSS,
+ 1452129.200000ns, VDD,
+ 1453330.100000ns, VDD,
+ 1453330.200000ns, VSS,
+ 1453570.300000ns, VSS,
+ 1453570.400000ns, VDD,
+ 1453690.400000ns, VDD,
+ 1453690.500000ns, VSS,
+ 1454411.000000ns, VSS,
+ 1454411.100000ns, VDD,
+ 1454771.300000ns, VDD,
+ 1454771.400000ns, VSS,
+ 1455251.700000ns, VSS,
+ 1455251.800000ns, VDD,
+ 1455972.300000ns, VDD,
+ 1455972.400000ns, VSS,
+ 1456572.800000ns, VSS,
+ 1456572.900000ns, VDD,
+ 1456933.100000ns, VDD,
+ 1456933.200000ns, VSS,
+ 1457173.300000ns, VSS,
+ 1457173.400000ns, VDD,
+ 1457773.800000ns, VDD,
+ 1457773.900000ns, VSS,
+ 1459695.400000ns, VSS,
+ 1459695.500000ns, VDD,
+ 1460055.700000ns, VDD,
+ 1460055.800000ns, VSS,
+ 1460175.800000ns, VSS,
+ 1460175.900000ns, VDD,
+ 1460896.400000ns, VDD,
+ 1460896.500000ns, VSS,
+ 1462097.400000ns, VSS,
+ 1462097.500000ns, VDD,
+ 1462217.500000ns, VDD,
+ 1462217.600000ns, VSS,
+ 1462337.600000ns, VSS,
+ 1462337.700000ns, VDD,
+ 1462818.000000ns, VDD,
+ 1462818.100000ns, VSS,
+ 1463658.700000ns, VSS,
+ 1463658.800000ns, VDD,
+ 1464139.100000ns, VDD,
+ 1464139.200000ns, VSS,
+ 1464619.500000ns, VSS,
+ 1464619.600000ns, VDD,
+ 1464859.700000ns, VDD,
+ 1464859.800000ns, VSS,
+ 1465700.400000ns, VSS,
+ 1465700.500000ns, VDD,
+ 1466060.700000ns, VDD,
+ 1466060.800000ns, VSS,
+ 1466661.200000ns, VSS,
+ 1466661.300000ns, VDD,
+ 1468342.600000ns, VDD,
+ 1468342.700000ns, VSS,
+ 1468943.100000ns, VSS,
+ 1468943.200000ns, VDD,
+ 1469303.400000ns, VDD,
+ 1469303.500000ns, VSS,
+ 1471225.000000ns, VSS,
+ 1471225.100000ns, VDD,
+ 1471825.500000ns, VDD,
+ 1471825.600000ns, VSS,
+ 1474227.500000ns, VSS,
+ 1474227.600000ns, VDD,
+ 1476269.200000ns, VDD,
+ 1476269.300000ns, VSS,
+ 1476629.500000ns, VSS,
+ 1476629.600000ns, VDD,
+ 1477109.900000ns, VDD,
+ 1477110.000000ns, VSS,
+ 1477470.200000ns, VSS,
+ 1477470.300000ns, VDD,
+ 1477590.300000ns, VDD,
+ 1477590.400000ns, VSS,
+ 1477950.600000ns, VSS,
+ 1477950.700000ns, VDD,
+ 1478310.900000ns, VDD,
+ 1478311.000000ns, VSS,
+ 1478791.300000ns, VSS,
+ 1478791.400000ns, VDD,
+ 1479271.700000ns, VDD,
+ 1479271.800000ns, VSS,
+ 1479391.800000ns, VSS,
+ 1479391.900000ns, VDD,
+ 1479872.200000ns, VDD,
+ 1479872.300000ns, VSS,
+ 1480352.600000ns, VSS,
+ 1480352.700000ns, VDD,
+ 1480953.100000ns, VDD,
+ 1480953.200000ns, VSS,
+ 1481433.500000ns, VSS,
+ 1481433.600000ns, VDD,
+ 1481913.900000ns, VDD,
+ 1481914.000000ns, VSS,
+ 1482274.200000ns, VSS,
+ 1482274.300000ns, VDD,
+ 1482514.400000ns, VDD,
+ 1482514.500000ns, VSS,
+ 1483355.100000ns, VSS,
+ 1483355.200000ns, VDD,
+ 1483835.500000ns, VDD,
+ 1483835.600000ns, VSS,
+ 1485156.600000ns, VSS,
+ 1485156.700000ns, VDD,
+ 1485516.900000ns, VDD,
+ 1485517.000000ns, VSS,
+ 1486117.400000ns, VSS,
+ 1486117.500000ns, VDD,
+ 1486237.500000ns, VDD,
+ 1486237.600000ns, VSS,
+ 1486597.800000ns, VSS,
+ 1486597.900000ns, VDD,
+ 1486958.100000ns, VDD,
+ 1486958.200000ns, VSS,
+ 1487078.200000ns, VSS,
+ 1487078.300000ns, VDD,
+ 1487198.300000ns, VDD,
+ 1487198.400000ns, VSS,
+ 1487678.700000ns, VSS,
+ 1487678.800000ns, VDD,
+ 1488159.100000ns, VDD,
+ 1488159.200000ns, VSS,
+ 1488519.400000ns, VSS,
+ 1488519.500000ns, VDD,
+ 1488999.800000ns, VDD,
+ 1488999.900000ns, VSS,
+ 1489480.200000ns, VSS,
+ 1489480.300000ns, VDD,
+ 1489840.500000ns, VDD,
+ 1489840.600000ns, VSS,
+ 1491762.100000ns, VSS,
+ 1491762.200000ns, VDD,
+ 1492242.500000ns, VDD,
+ 1492242.600000ns, VSS,
+ 1492843.000000ns, VSS,
+ 1492843.100000ns, VDD,
+ 1493323.400000ns, VDD,
+ 1493323.500000ns, VSS,
+ 1494524.400000ns, VSS,
+ 1494524.500000ns, VDD,
+ 1494764.600000ns, VDD,
+ 1494764.700000ns, VSS,
+ 1495124.900000ns, VSS,
+ 1495125.000000ns, VDD,
+ 1495365.100000ns, VDD,
+ 1495365.200000ns, VSS,
+ 1496686.200000ns, VSS,
+ 1496686.300000ns, VDD,
+ 1496806.300000ns, VDD,
+ 1496806.400000ns, VSS,
+ 1497526.900000ns, VSS,
+ 1497527.000000ns, VDD,
+ 1499688.700000ns, VDD,
+ 1499688.800000ns, VSS,
+ 1500769.600000ns, VSS,
+ 1500769.700000ns, VDD,
+ 1501610.300000ns, VDD,
+ 1501610.400000ns, VSS,
+ 1501730.400000ns, VSS,
+ 1501730.500000ns, VDD,
+ 1501850.500000ns, VDD,
+ 1501850.600000ns, VSS,
+ 1502330.900000ns, VSS,
+ 1502331.000000ns, VDD,
+ 1502691.200000ns, VDD,
+ 1502691.300000ns, VSS,
+ 1503291.700000ns, VSS,
+ 1503291.800000ns, VDD,
+ 1503772.100000ns, VDD,
+ 1503772.200000ns, VSS,
+ 1504252.500000ns, VSS,
+ 1504252.600000ns, VDD,
+ 1506654.500000ns, VDD,
+ 1506654.600000ns, VSS,
+ 1507375.100000ns, VSS,
+ 1507375.200000ns, VDD,
+ 1508936.400000ns, VDD,
+ 1508936.500000ns, VSS,
+ 1510137.400000ns, VSS,
+ 1510137.500000ns, VDD,
+ 1510257.500000ns, VDD,
+ 1510257.600000ns, VSS,
+ 1511098.200000ns, VSS,
+ 1511098.300000ns, VDD,
+ 1512659.500000ns, VDD,
+ 1512659.600000ns, VSS,
+ 1512899.700000ns, VSS,
+ 1512899.800000ns, VDD,
+ 1513620.300000ns, VDD,
+ 1513620.400000ns, VSS,
+ 1514100.700000ns, VSS,
+ 1514100.800000ns, VDD,
+ 1514461.000000ns, VDD,
+ 1514461.100000ns, VSS,
+ 1515061.500000ns, VSS,
+ 1515061.600000ns, VDD,
+ 1517343.400000ns, VDD,
+ 1517343.500000ns, VSS,
+ 1519024.800000ns, VSS,
+ 1519024.900000ns, VDD,
+ 1519265.000000ns, VDD,
+ 1519265.100000ns, VSS,
+ 1521426.800000ns, VSS,
+ 1521426.900000ns, VDD,
+ 1521667.000000ns, VDD,
+ 1521667.100000ns, VSS,
+ 1522387.600000ns, VSS,
+ 1522387.700000ns, VDD,
+ 1523708.700000ns, VDD,
+ 1523708.800000ns, VSS,
+ 1524429.300000ns, VSS,
+ 1524429.400000ns, VDD,
+ 1524669.500000ns, VDD,
+ 1524669.600000ns, VSS,
+ 1524909.700000ns, VSS,
+ 1524909.800000ns, VDD,
+ 1525029.800000ns, VDD,
+ 1525029.900000ns, VSS,
+ 1525390.100000ns, VSS,
+ 1525390.200000ns, VDD,
+ 1525510.200000ns, VDD,
+ 1525510.300000ns, VSS,
+ 1526831.300000ns, VSS,
+ 1526831.400000ns, VDD,
+ 1527311.700000ns, VDD,
+ 1527311.800000ns, VSS,
+ 1529353.400000ns, VSS,
+ 1529353.500000ns, VDD,
+ 1529953.900000ns, VDD,
+ 1529954.000000ns, VSS,
+ 1530674.500000ns, VSS,
+ 1530674.600000ns, VDD,
+ 1531395.100000ns, VDD,
+ 1531395.200000ns, VSS,
+ 1531755.400000ns, VSS,
+ 1531755.500000ns, VDD,
+ 1532716.200000ns, VDD,
+ 1532716.300000ns, VSS,
+ 1533196.600000ns, VSS,
+ 1533196.700000ns, VDD,
+ 1533436.800000ns, VDD,
+ 1533436.900000ns, VSS,
+ 1533556.900000ns, VSS,
+ 1533557.000000ns, VDD,
+ 1533677.000000ns, VDD,
+ 1533677.100000ns, VSS,
+ 1534037.300000ns, VSS,
+ 1534037.400000ns, VDD,
+ 1534637.800000ns, VDD,
+ 1534637.900000ns, VSS,
+ 1535238.300000ns, VSS,
+ 1535238.400000ns, VDD,
+ 1535718.700000ns, VDD,
+ 1535718.800000ns, VSS,
+ 1536079.000000ns, VSS,
+ 1536079.100000ns, VDD,
+ 1536559.400000ns, VDD,
+ 1536559.500000ns, VSS,
+ 1538000.600000ns, VSS,
+ 1538000.700000ns, VDD,
+ 1538240.800000ns, VDD,
+ 1538240.900000ns, VSS,
+ 1538360.900000ns, VSS,
+ 1538361.000000ns, VDD,
+ 1538481.000000ns, VDD,
+ 1538481.100000ns, VSS,
+ 1539081.500000ns, VSS,
+ 1539081.600000ns, VDD,
+ 1539321.700000ns, VDD,
+ 1539321.800000ns, VSS,
+ 1540042.300000ns, VSS,
+ 1540042.400000ns, VDD,
+ 1541843.800000ns, VDD,
+ 1541843.900000ns, VSS,
+ 1542804.600000ns, VSS,
+ 1542804.700000ns, VDD,
+ 1544245.800000ns, VDD,
+ 1544245.900000ns, VSS,
+ 1544606.100000ns, VSS,
+ 1544606.200000ns, VDD,
+ 1544726.200000ns, VDD,
+ 1544726.300000ns, VSS,
+ 1545566.900000ns, VSS,
+ 1545567.000000ns, VDD,
+ 1545687.000000ns, VDD,
+ 1545687.100000ns, VSS,
+ 1545807.100000ns, VSS,
+ 1545807.200000ns, VDD,
+ 1546767.900000ns, VDD,
+ 1546768.000000ns, VSS,
+ 1547248.300000ns, VSS,
+ 1547248.400000ns, VDD,
+ 1547728.700000ns, VDD,
+ 1547728.800000ns, VSS,
+ 1548209.100000ns, VSS,
+ 1548209.200000ns, VDD,
+ 1548449.300000ns, VDD,
+ 1548449.400000ns, VSS,
+ 1548569.400000ns, VSS,
+ 1548569.500000ns, VDD,
+ 1549890.500000ns, VDD,
+ 1549890.600000ns, VSS
+)}


.end

