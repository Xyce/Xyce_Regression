**********************************************************************
* Test of core dump from invalid .PRINT line, where the .PRINT
* line does not have a trailing parenthesis, such as V(1), or 
* is mssing the variable, such as V().  These lines would cause
* a core dump, per SON Bug 694.
*
*
*
*
*
*
**********************************************************************
V1 1 0 SIN(0 1 1KHZ)
R1 1 2 1
R2 2 0 1

.TRAN 0 1ms
.PRINT TRAN V(1
.PRINT TRAN V()
.PRINT TRAN V(
.PRINT TRAN I(V1
.PRINT TRAN I()
.PRINT TRAN I(
.PRINT TRAN N(R1
.PRINT TRAN N()
.PRINT TRAN N(
.PRINT TRAN P(R1
.PRINT TRAN P()
.PRINT TRAN P(
.PRINT TRAN W(R1
.PRINT TRAN W()
.PRINT TRAN W(

.END
