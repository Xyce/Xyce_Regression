*Test of BSIM6 output variable feature
*Duplicates BSIM6 gummel_nmos test
.options nonlin abstol=1e-6 reltol=1e-6 
.options device temp=25

*.hdl "bsim6.va"
.include "modelcard_xyce.nmos"

* --- Voltage Sources ---
vdrain drain 0 dc 0
esource source 0 drain 0 -1
vgate gate  0 dc 1.0
vbulk bulk 0 dc 0.0


* --- Transistor ---
M1 drain gate source bulk nmos W=10u L=10u 

* Second transistor for finite differencing
Bdrain drain2 0 V={V(drain)}
Bgate gate2 0  V={V(gate)+((V(gate)==0)?.00000001:(1e-8*abs(v(gate))))}
Bsource source2 0 V={V(source)}
Bbulk bulk2 0 V={V(bulk)}

M2 drain2 gate2 source2 bulk2 nmos W=10u L=10u 

* --- DC Analysis ---
.dc vdrain -0.1 0.1 0.001 vgate 0.0 1.0 0.2
*.probe dc ids=par'-i(vdrain)'
*.probe dc gx=deriv(ids)
*.probe dc gx2=deriv(gx)
*.probe dc gx3=deriv(gx2)
*.probe dc gx4=deriv(gx3)
*.print dc par'ids' par'gx' par'gx2' par'gx3' par 'gx4'
*COMP {N(M1:gm)-{(N(M2:ids)-N(M1:ids))/(V(gate2)-V(gate))}} abstol=1e-9
*COMP {(N(M2:ids)-N(M1:ids))/(V(gate2)-V(gate))} abstol=1e-9
.print dc v(drain) v(gate) N(M1:ids) {(N(M2:ids)-N(M1:ids))/(V(gate2)-V(gate))} N(M1:gm) {N(M1:gm)-{(N(M2:ids)-N(M1:ids))/(V(gate2)-V(gate))}}  N(M1:Vth) N(M1:Vds) N(M1:Vbs) N(M1:Vgs) N(M1:Vdsat)

.end
