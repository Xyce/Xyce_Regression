* AC simulation for xyce
.options device temp=25
.subckt mysub c_x b_x e_x s_x
e_c c_v 0 c_x 0 1
v_c c_v c 0
f_c c_x 0 v_c   -1
e_b b_v 0 b_x 0 1
v_b b_v b 0
f_b b_x 0 v_b   -1
e_e e_v 0 e_x 0 1
v_e e_v e 0
f_e e_x 0 v_e   -1
e_s s_v 0 s_x 0 1
v_s s_v s 0
f_s s_x 0 v_s   -1
q1 c b e s mymodel
.model mymodel npn level=504
+ LEVEL=504.0
+ TREF=25.00
+ DTA=0.000
+ EXMOD=1.000
+ EXPHI=1.000
+ EXAVL=0.000
+ EXSUB=0.000
+ IS=22.0E-18
+ IK=0.1
+ VER=2.5
+ VEF=44.0
+ BF=215.0
+ IBF=2.7E-15
+ MLF=2.000
+ XIBI=0.0
+ IZEB=0.0
+ NZEB=22.0
+ BRI=7.00
+ IBR=1.0E-015
+ VLR=0.2
+ XEXT=0.63
+ WAVL=1.1E-006
+ VAVL=3.0
+ SFH=0.3
+ RE=5.0
+ RBC=23.0
+ RBV=18.0
+ RCC=12.0
+ RCBLX=0.000
+ RCBLI=0.000
+ RCV=150.0
+ SCRCV=1250.0
+ IHC=4.000E-003
+ AXI=0.3
+ CJE=73.0E-015
+ VDE=950.0E-003
+ PE=400.0E-003
+ XCJE=400.0E-003
+ CBEO=0.000
+ CJC=78.0E-015
+ VDC=680.0E-003
+ PC=500.0E-003
+ XP=350.0E-003
+ MC=500.0E-003
+ XCJC=32.0E-003
+ CBCO=0.000
+ MTAU=1.0
+ TAUE=2.0E-012
+ TAUB=4.2E-12
+ TEPI=41.0E-12
+ TAUR=520.0E-012
+ DEG=0.01
+ XREC=0.1
+ AQBO=300.0E-003
+ AE=0.0E-003
+ AB=1.0
+ AEX=620.0E-003
+ AEPI=2.5
+ AC=2.0
+ ACBL=2.0
+ DAIS=0.000
+ DVGBF=50.0E-003
+ DVGBR=45.00E-003
+ VGB=1.17
+ VGC=1.18
+ VGJ=1.15
+ VGZEB=1.15
+ AVGEB=4.73E-4
+ TVGEB=636.0
+ DVGTE=50.0E-003
+ AF=2.000
+ KF=20.0E-012
+ KFN=20.0E-012
+ KAVL=1.000
+ ISS=48.0E-18
+ ICSS=-1.0
+ IKS=250.E-006
+ CJS=315.0E-015
+ VDS=620.0E-003
+ PS=340.0E-003
+ VGS=1.20
+ AS=1.580
+ ASUB=2.0
+ MULT=1.5
.ends
v_c_b c_b 0 2.0
v_b_b b_b 0 0.85 ac 1
v_e_b e_b 0 0
v_s_b s_b 0 0
x_b c_b b_b e_b s_b mysub
.ac dec 1 1e6 1e9
.print ac i(v_c_b)
+ i(v_b_b)
.print ac FILE=b538_6_bl i(v_e_b)
+ i(v_s_b)
.end
