* Test invalid syntaxes for TABLE and POLY forms of
* E and F sources.  This also covers G and H sources,
* since they use the same code blocks for device-line 
* parsing.

B1   1 0 V={2.0*sin(2*pi*TIME) }
R1   1 2 1K
R2   0 2 100

* POLY E-source is missing all expression terms
EPOLY1 3 0 POLY(2) 
R3     3 4 1K
R4     0 4 100

* POLY E-source is missing number after POLY( 
EPOLY2 5 0 POLY( 
R5     5 6 1K
R6     0 6 100

* TABLE E-source is missing = sign after TABLE keyword
ETABLE  7 0 TABLE V(1,0) (0,1) (1,2)
R7      7 8 1K
R8      0 8 100

* POLY F-source is missing all expression terms
FPOLY  9 0 POLY(1)
R9     9 10 1K
R10    0 10 100


.TRAN 0 1
.PRINT TRAN V(1)

.END

