THIS CIRCUIT TESTS THE MOS BSIM3 MODEL AS A CHAIN OF INVERTERS IN SERIES
* This is a chain of 20 1-input CMOS inverters
* The NMOS and PMOS devices have their gates tied 
* together to form a CMOS inverter. VIN1, the input signal, is applied to a 1K
* resistor,RIN, which is connected to the gates of the inverter at node IN.
*
* This version uses the bsim soi version 3.2 model cards from the berkeley
* web site:  http://www-device.eecs.berkeley.edu/~bsimsoi/circuits2.html

.subckt INVERTER IN OUT VDD GND
M2 OUT IN GND GND n1 w=1.8u l=1.2u
M1 OUT IN VDD VDD p1 w=3.6u l=1.2u
.ends

* A small load (R1, C1) is applied to the output node, VOUT. The input signal
* is at 2V for 1.5us and then at 0V for 1.5us. The voltage at VOUT is high 
* when VIN1 is low and vice versa.

.tran 0 1us
.print tran v(vout) v(out20) v(in) v(1)
.print homotopy v(vout) v(out20) v(in) v(1)
.options device vgstconst=3.0 Temp=100.0

************************************
* **** Start Homotopy Setup ****
************************************
.options nonlin maxstep=200 continuation=mos

**********************************
* **** End Homotopy Setup ****
**********************************

VDDdev 	VDD	0	2V 
RIN	IN	1	1K
VIN1  1	0  2V 
R1    VOUT  0  10K  
C2    VOUT  0  0.1p
XINV1 IN OUT2 VDD 0 INVERTER
XINV2 OUT2 OUT3 VDD 0 INVERTER
XINV3 OUT3 OUT4 VDD 0 INVERTER
XINV4 OUT4 OUT5 VDD 0 INVERTER
XINV5 OUT5 OUT6 VDD 0 INVERTER
XINV6 OUT6 OUT7 VDD 0 INVERTER
XINV7 OUT7 OUT8 VDD 0 INVERTER
XINV8 OUT8 OUT9 VDD 0 INVERTER
XINV9 OUT9 OUT10 VDD 0 INVERTER
XINV10 OUT10 OUT11 VDD 0 INVERTER
XINV11 OUT11 OUT12 VDD 0 INVERTER
XINV12 OUT12 OUT13 VDD 0 INVERTER
XINV13 OUT13 OUT14 VDD 0 INVERTER
XINV14 OUT14 OUT15 VDD 0 INVERTER
XINV15 OUT15 OUT16 VDD 0 INVERTER
XINV16 OUT16 OUT17 VDD 0 INVERTER
XINV17 OUT17 OUT18 VDD 0 INVERTER
XINV18 OUT18 OUT19 VDD 0 INVERTER
XINV19 OUT19 OUT20 VDD 0 INVERTER
XINV20 OUT20 VOUT VDD 0 INVERTER

**************************************************************************
.MODEL  N1  NMOS  (LEVEL = 9)
.MODEL  P1  PMOS  (LEVEL = 9)
**************************************************************************

*
.END
