Test of Exponential and Natural Log Functions
********************************************************************************
* Tier No.:     1
* Directory/Circuit Name: ABM_EXPLN/exp_ln.cir
* Description:  Test of the XYCE analog behavioral modeling exponential 
*	and natural log functions
* Input: VS
* Output: V(1), V(2), V(3)
* Analysis:
*	The input voltage, VS, is a piece wise linear source with specified time
*	and voltage pairs.  Two nonlinear dependent voltage sources are used to 
*	define the functions as follows:
*		V(2)=B2=EXP(V(1)) = exponent of input voltage = EXP(V(1)) 
*		V(3)=B3=LN(V(2)) = ln of B2 (EXP function) = V(1)
*	A transient analysis is performed and the output recorded is the node  
*	voltages defined by the input source, V(1),  the exponential, V(2), and 
*	natural log , V(3),  functions. 
*
*	This table is a set of hand calculations for the EXP and LN functions:	
*	 	   X		EXP(X)		LN(EXP(X)) 			
*		 2.500		12.182		2.500	
*		 5.000		148.410		5.000
*		 7.500		1808.00		7.500
*		10.000		2202.60		10.00
*
*********************************************************************************
* This also tests the case of a function that does not contain all the independent
* variables in the definition
.func abc(x,y) {y}
VS  1  0  PWL(0 2.5V 0.5MS 5V 1MS 7.5V 1.5MS 10V 2MS 7.5V)
R1  1  0  {abc(0,1)}
*R1  1  0  1
B2  2  0  V = {EXP(V(1))}
R2  2  0  1
B3  3  0  V = {LN(V(2))}
R3  3  0  1
.TRAN 0.02MS 2.5MS
.PRINT TRAN V(1) V(2) V(3)
.END
