* Transient sensitivity example, SFFM source, analytical derivatives
.param cap=0.1u
.param res=1K

c1 1 0 cap
c2 2 0 cap
R1 1 3 res
R2 1 2 res

Vin 3 0 SFFM(0 1 1MEG 2 250K)

* Transient commands
.tran 0 10us 
.options timeint reltol=1e-6 abstol=1e-6

.print tran v(1) v(2) v(3)

* Sensitivity commands
.print sens 
.SENS objfunc={V(2)} sensdevicename=vin
.options SENSITIVITY direct=1 adjoint=0  forceanalytic=true
.end

