RC ladder circuit 

P1 1 0 port=2
*P2 12 0  port=1  z0=100

C1 2 0 1e-2
Rgs 1 2 0.02

.subckt RCBlock IN OUT GND
R1 IN OUT 20
C1 IN OUT 1p
Cg1 OUT GND 1p
.ends

X1 2 3 0 RCBlock
X2 3 4 0 RCBlock
X3 4 5 0 RCBlock
X4 5 6 0 RCBlock
X5 6 7 0 RCBlock
X6 7 8 0 RCBlock
X7 8 9 0 RCBlock
X8 9 10 0 RCBlock
X9 10 11 0 RCBlock
X10 11 12 0 RCBlock

.AC lin 11 -1e5 1e5

*.AC DEC 10 10  1e5 

.LIN FORMAT=TOUCHSTONE

P2 12 0  port=1  z0=100

.END
