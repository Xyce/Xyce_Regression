*A Simple MOSFET Gain Stage. AC Analysis.

M1 3 2 0 0 nmos w=4u l=1u 
Rsource 1 2 100k
Rload 3 vdd 25k

Vdd1 vdd 0 5 
Vin 1 0 1.44 ac .1 sin(0 1 1e+5 0 0) 

*.ac dec 10 100Hz 1000MegHz 
.ac dec 10 1e7Hz 1000MegHz 
.print ac v(3)

.sens objvars=2 param=m1:w,m1:l
.options sensitivity direct=0 adjoint=1  stdoutput=1  forcedevicefd=1

.print sens 
*format=tecplot

.model nmos nmos level=9

.end

