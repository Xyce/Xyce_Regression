AC test of FORMAT=TECPLOT output format
*
* Trivial resistor circuit, just do a DC sweep and watch the output
*

R1 1 0 10
V1 1 0 DC 0V

.print AC FORMAT=TECPLOT v(1) I(v1)
.ac dec 10 100Hz 1000MegHz

.end
