RAW File Output test for the NSOI MOSFET.
************************************************************
* This test has two purposes:
*   1) Verify that the variable type (e.g., "voltage") and 
*      variable name is correct for the MOSFET. This test
*      just has a gate prime contribution, which is a 
*      voltage contribution.    
*
*   2) Verify that the data is actually correct for all of
*      the time-steps in the .RAW file output 
*
* The "gold" .RAW file output was generated by manually
* comparing that "gold" file with a .PRN file.  It was 
* generated for a limited set of fixed time-steps, so that
* a file comparison could be used to verify the test output's
* .RAW file against that "gold" .RAW file.
*
************************************************************
*
.options device mincap=1uf
.options timeint method=gear
.options nonlin-tran rhstol=1.0e-7

rin in 1 100K
vin   1 0  0V PULSE (0V 4V 1.5us 5ns 5ns 1.5us 3.01us)
cin in 0 1.0p

Rnd   in  nd  1
Rng   in  ng  1
Rns   0   ns  1
Rne   0   ne  1
Rnb   0   nb  1e+8

MN1 nd ng ns ne nb  cmosn L=0.258u W=19.585u

.MODEL cmosn nmos (    LEVEL   = 10
+ soimod = 0
+ rgatemod = 1
+ mobmod = 2  capmod = 2
+ shmod = 1  igmod = 0  paramchk = 0 )

.tran 20ns 3us
.options output initial_interval=0.2us

* .PRINT statement is not actually used for .RAW output.
* It was included in the netslit so that the "gold" .RAW 
* file output could manually verified against a .PRN file
* during test development
.print tran v(1) v(in) N(mn1_gate) v(nb) v(nd) v(ne) 
+ v(ng) v(ns) I(vin)
 
.end

