* AC simulation for xyce
* this is the fgum_ac_npn_full_sh_ac test from the CMC suite
.options device temp=27
.subckt mysub coll_x base_x emit_x subs_x therm_x
e_coll coll_v 0 coll_x 0 1
v_coll coll_v coll 0
f_coll coll_x 0 v_coll   -1
e_base base_v 0 base_x 0 1
v_base base_v base 0
f_base base_x 0 v_base   -1
e_emit emit_v 0 emit_x 0 1
v_emit emit_v emit 0
f_emit emit_x 0 v_emit   -1
e_subs subs_v 0 subs_x 0 1
v_subs subs_v subs 0
f_subs subs_x 0 v_subs   -1
v_therm therm therm_x 0
q1 coll base emit subs therm mymodel
.model mymodel npn level=230
+ mcf= 1 
+ rbi0= 4.444 
+ rbx= 2.568 
+ fgeo= 0.7409 
+ re= 1.511 
+ rcx= 2.483 
+ itss= 0 
+ msf= 1 
+ iscs= 0 
+ msc= 1 
+ cjci0= 3.58e-015 
+ vdci= 0.8201 
+ zci= 0.2857 
+ vptci= 1.79 
+ cjcx0= 6.299e-015 
+ vdcx= 0.8201 
+ zcx= 0.2863 
+ vptcx= 1.977 
+ cjs0= 2.6e-014 
+ vds= 0.9997 
+ zs= 0.4295 
+ vpts= 100 
+ t0= 2.089e-013 
+ dt0h= 8e-014 
+ tbvl= 8.25e-014 
+ tef0= 3.271e-013 
+ thcs= 5.001e-012 
+ ahc= 0.05 
+ rci0= 9.523 
+ vlim= 0.6999 
+ vces= 0.01 
+ vpt= 2 
+ tr= 0 
+ cbepar= 2.609e-014 
+ cbcpar= 1.64512e-014 
+ alqf= 0.166667 
+ alit= 0.333333 
+ flnqs= 0 
+ kf= 0 
+ af= 2 
+ vgb= 0.91 
+ alt0= 0.004 
+ kt0= 6.588e-005 
+ zetaci= 0.58 
+ alvs= 0.001 
+ alces= -0.2286 
+ zetarbi= 0.3002 
+ zetarbx= 0.06011 
+ zetarcx= -0.02768 
+ zetare= -0.9605 
+ vge= 1.17 
+ vgc= 1.17 
+ vgs= 1.17 
+ f1vg= -0.000102377 
+ f2vg= 0.00043215 
+ zetact= 5 
+ zetabet= 4.892 
+ flsh= 1 
+ rth= 1113.4 
+ cth= 6.841e-012 
+ zetarth= 0 
+ tnom= 26.85 
+ zetavgbe= 0.7 
.ends
.global_param coll_voltage=1.5
.global_param base_voltage=1.05
v_coll_coll coll_coll 0 'coll_voltage' ac 1
v_base_coll base_coll 0 'base_voltage'
v_emit_coll emit_coll 0 0
v_subs_coll subs_coll 0 0
i_therm_coll therm_coll 0 0
x_coll coll_coll base_coll emit_coll subs_coll therm_coll mysub
v_coll_base coll_base 0 'coll_voltage'
v_base_base base_base 0 'base_voltage' ac 1
v_emit_base emit_base 0 0
v_subs_base subs_base 0 0
i_therm_base therm_base 0 0
x_base coll_base base_base emit_base subs_base therm_base mysub
.step lin base_voltage 0.75 1.05 0.01
.step coll_voltage list 0.5 1.0 1.5
.ac dec 10 1e+010 2e+010
.print ac 
+ i(v_coll_coll)
+ i(v_base_coll)
+ i(v_emit_coll)
+ i(v_subs_coll)
+ v(therm_coll)
+ i(v_coll_base)
+ i(v_base_base)
+ i(v_emit_base)
+ i(v_subs_base)
+ v(therm_base)
.end
