Local Variation test
*
V1 1 0 1.0

.param random_value=nint(1+10*rand())
.param global_variation=random_value
.param param2=random_value*100+global_variation

r1 1 2 global_variation
r2 2 0 param2

.dc V1 1 1 1
.print dc precision=12 width=21 v(1) v(2) 

.sampling useExpr=true

.options samples numsamples=10 seed=1923635719
+ outputs={v(1)+0.2}
+ sample_type=lhs
+ stdoutput=false

.result {r1:R}
.result {r2:R}

.END

