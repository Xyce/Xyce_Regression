2222 bjt failure test
.MODEL N2222 NPN 
+ LEVEL = 1
+ IS = 2.6E-14  BF = 200      NF = 1.0     VAF = 90.0
+ IKF = 0.14    ISE = 3.4E-15 NE = 1.3     BR = 14
+ NR = 1.0      VAR = 9.0     IKR = 0.1    ISC = 2.0E-14 
+ NC = 4.5      IRB = 0.0004 RBM = 0.002 

V1     node1   0     1.0
E1  coll1 0  node1 0  2
Ib1  0 base1  0.0000
Ve1  emit1 0  0V 
Qtest1  coll1 base1 emit1  N2222

.DC Ib1 0.0 0.0 1.0
.STEP V1 0 1.001 5.0e-3

.PRINT DC V(coll1)  Ic(Qtest1) 

.End

