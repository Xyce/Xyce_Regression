* test the TABLE form of the B source
* The G source in the original netlist is internally converted into this
* B source, so this should be (and is) identical in behavior to the 
* original netlist

*COMP v(node1) OFFSET=.0
*COMP v(node2) OFFSET=3.0

.TRAN 0 1us
.PRINT TRAN V(node1) V(node2)
R1         node2 0  1
B1         node2 0 I={table(v(node1),-1,-3,1,3)}
V1         node1 0 SIN(0V 0.75V 1e6 0 0 0)
