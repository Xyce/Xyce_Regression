Test of expressions on .TRAN line
*******************************************************************************
*
* a few sources of different types
VS1  1  0  SIN(0 1.0 1KHZ 0 0)
VP2  2  0  PULSE( 0 100 0.2ms 0.2ms 0.2ms 1ms 2ms )
VS3  3  0  SIN(0 -1.0 1KHZ 0 0)
VS4  4  0  SIN(-0.5 1.0 1KHZ 0 0.5)
VS5  5  0  SIN(0.5 -1.0 1KHZ 0 0.5)

R1  1  0  100
R2  2  0  100
R3  3  0  100
R4  4  0  100
R5  5  0  100

.param initial_step_value=0.0
.param final_time_value=5ms
.param start_time_value=0.0
.param step_ceiling_value=1.0e-5

.tran {initial_step_value} {final_time_value} {start_time_value} {step_ceiling_value}

.PRINT TRAN V(1) V(2) V(3) V(4) V(5) V(1,0) V(3,0)

.END

