* This .HB analysis was used to generate the Gold standards for the
* ylin-5port-yparam.cir test.  However, it is not run as part of any
* regression test.

* RC ladder circuit

v1 1 0  sin  0 5 1e4
C1 2 0 1e-2
Rgs 1 2 0.02

.subckt RCBlock IN OUT GND
R1 IN OUT 20
C1 IN OUT 1p
Cg1 OUT GND 1p
.ends

X1 2 3 0 RCBlock
X2 3 4 0 RCBlock
X3 4 5 0 RCBlock
X4 5 6 0 RCBlock
X5 6 7 0 RCBlock
X6 7 8 0 RCBlock
X7 8 9 0 RCBlock
X8 9 10 0 RCBlock
X9 10 11 0 RCBlock
X10 11 12 0 RCBlock

.options hbint numfreq=10 tahb=0
.hb 1e4
.print hb v(1) v(2) v(5) v(6) v(7) v(12) i(v1)

.END
