* Transient sensitivity example, pulse source, finite difference version
.param cap=0.1u
.param res=1K
.param v1=0
.param v2=1
.param td=0s
.param tr=10us
.param tf=10us 
.param pw=100us 
.param per=220us

c1 1 0 cap
c2 2 0 cap
R1 1 3 res
R2 1 2 res

Vin 3 0 PULSE({v1} {v2} {td} {tr} {tf} {pw} {per})

* Transient commands
.tran 0 4ms uic
.options timeint reltol=1e-6 abstol=1e-6

.print tran v(1) v(2) v(3)

* Sensitivity commands
.print sens 
.SENS objfunc={V(2)} param=v1,v2,td,tr,tf,pw,per
.options SENSITIVITY direct=1 adjoint=0 forcefd=true
.end

