Netlist to demonstrate TEMP bug
* .global_param foobar={Vt/(1.3806226e-23/1.6021918e-19)}
* .global_param foobaz={TEMP}
B1 2 0 V={Vt/(1.3806226e-23/1.6021918e-19)}
R2 2 0 1

B2 3 0 V={TEMP}
R3 3 0 1

* B3 4 0 V={foobaz}
* R4 4 0 1

* This little circuit here to please xyce_verify and for no other reason
vjunk 5 0 1
rjunk 5 0 1

.OP
*.dc line necessary for xyce_verify to know what to do
.DC vjunk 1 1 1
.step TEMP 27 30 1

*v(5) must be printed because xyce_verify needs a sweep variable
.PRINT DC  v(5) V(2) V(3) {TEMP} {Vt/(1.3806226e-23/1.6021918e-19)}

.END
