*********************************************************
* Test FORMAT=GNUPLOT with .STEP.  This should produce 
* the same .prn files as FORMAT=STD, but with two 
* blank lines before steps 1,2, ... N-1.  Note that
* first step is "step 0".  In this netlist, N is 4.
*
* Also test FORMAT=SPLOT with .STEP. This should
* produce the same files as FORMAT=STD, but
* with one blank line before steps 1,2, ... N-1.
*
* This version uses separate .PRINT lines for the 
* .HB.TD.prn and .HB.FD.prn files.  It will also make 
* a .startup.prn file.
**********************************************************

R1  1 1a 500
R1a 1a 0 500
C1 1 0 1p
D1 2 1 D1N3940
.MODEL D1N3940 D (IS=4e-10 RS=.105 N=1.48 TT=8e-7 CJO=1.95E-11 VJ=.4 M=.38 
+ EG=1.36 XTI=-8 KF=0 AF=1 FC=.9 BV=600 IBV=1e-4)

*            low high td tr  tf  pulsewidth    period
v1 2 0 pulse 1V 2V  0 1e-5 1e-5 {1/1e4/2-1e-5 } {1/1e4}

.print HB_FD FORMAT=GNUPLOT vm(1) vm(1a)
.print HB_TD FORMAT=GNUPLOT vm(1)
.print HB_FD FORMAT=SPLOT FILE=hb-fd-td-step-gnuplot.cir.HB.FD.splot.prn vm(1) vm(1a)
.print HB_TD FORMAT=SPLOT FILE=hb-fd-td-step-gnuplot.cir.HB.TD.splot.prn vm(1)
.hb 1e4
.STEP R1:R 250 750 500
.STEP R1A:R 1000 2000 1000

.options hbint numfreq=10
.options hbint STARTUPPERIODS=5

.end
