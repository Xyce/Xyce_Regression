* Xyce netlist for testing lossless transmission line

.TRAN 0 100ns 0
.PRINT TRAN FORMAT=PROBE V(N15504) V(N15586) V(in_3) V(out_3)

* Lossy transmission lines
R_R1 N15586 0 TC=0,0 R=10
V_V1 N15504 0 PULSE(0 5 0 0.1e-9 0.1e-9 5e-9 25e-9)
O_T1  N15504 0 N15586 0 cable
.MODEL cable LTRA LEN=100 R=0.05 L=1e-8 G=0 C=20e-12

R_R2 out_3 0 R=10 TC=0,0
V_V2  in_3 0 PULSE(0 5 0 0.1e-9 0.1e-9 5e-9 25e-9) 
O_T2  in_3 0 out_3 0 cable

.END

