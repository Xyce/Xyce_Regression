NOISE test of -r output ASCII format with .OP
*
V1  1 0 DC 5.0 AC  1.0   
R1  1 0 100K

* For testing SON Bug 1026, the .OP statement
* precedes the .NOISE statement.
.OP
.NOISE  V(1) V1  DEC  5 100 100K 1
.PRINT NOISE INOISE ONOISE

.END

