CMOS INVERTER, testing sensitivities with .FOUR
*
* The version is nearly the same as bsim3sensFourFD.cir, except that it has 
* additional signals to process.  In an early version of this capability, this 
* extra complexity caused an indexing mistake.
*
.param Vmag=2.0
*
.param lengthN=0.35U
.param lengthP=0.46U

.param dLN={lengthN*1e-10}
.param dLP={lengthP*1e-10}

M1 2 1 0 0 NMOS L={lengthN} W=4.2U AD=4.2P AS=4.2P PD=10U PS=10U
M2 2 1 3 3 PMOS L={lengthP} W=1U  AD=1P   AS=1P   PD=4U  PS=4U
VDD 3 0 {Vmag}
VIN 1 0 SIN {0.5*Vmag} {0.5*Vmag} 20MEG

* FD circuit for M1:L
M1_a 2a 1a 0  0  NMOS L={lengthN+dLN} W=4.2U AD=4.2P AS=4.2P PD=10U PS=10U
M2_a 2a 1a 3a 3a PMOS L={lengthP} W=1U  AD=1P   AS=1P   PD=4U  PS=4U
VDD_a 3a 0 {Vmag}
VIN_a 1a 0 SIN {0.5*Vmag} {0.5*Vmag} 20MEG

* FD circuit for M2:L
M1_b 2b 1b 0  0  NMOS L={lengthN} W=4.2U AD=4.2P AS=4.2P PD=10U PS=10U
M2_b 2b 1b 3b 3b PMOS L={lengthP+dLP} W=1U  AD=1P   AS=1P   PD=4U  PS=4U
VDD_b 3b 0 {Vmag}
VIN_b 1b 0 SIN {0.5*Vmag} {0.5*Vmag} 20MEG

.options timeint reltol=1.0e-7 abstol=1.0e-7

.sens objfunc={V(2)}  param=M1:L,M2:L
.print sens format=tecplot { (V(2a)-V(2))/dLN }  { (V(2b)-V(2))/dLP }  v(1) v(2) v(3)
.options sensitivity direct=1 adjoint=0

.TRAN 1N 100N

.FOUR 20MEG V(2) { (V(2a)-V(2))/dLN } { (V(2b)-V(2))/dLP }
.FOUR 30MEG V(2a) V(2)
.FOUR 40MEG V(2) { (V(2a)-V(2))/dLN } { (V(2b)-V(2))/dLP }

* this is the new feature, in progress:
* Possibly formats:
*
** do every sensitivity:
.FOUR 20MEG sens
.FOUR 40MEG sens

.PRINT TRAN V(2) V(1)

.MODEL NMOS NMOS (                                LEVEL   = 9
+TNOM    = 27             TOX     = 7.9E-9
+XJ      = 1.5E-7         NCH     = 1.7E17         VTH0    = 0.5169662
+K1      = 0.5862027      K2      = 0.0120774      K3      = 16.1323712
+K3B     = 0.8487425      W0      = 2.17449E-6     NLX     = 2.079688E-7
+DVT0W   = 0              DVT1W   = 5.3E6          DVT2W   = -0.032
+DVT0    = 9.7504029      DVT1    = 0.9681505      DVT2    = -0.0235742
+U0      = 438.6895901    UA      = 8.263356E-11   UB      = 2.159824E-18
+UC      = 8.361115E-11   VSAT    = 1.173431E5     A0      = 0.9412879
+AGS     = 0.3886454      B0      = 3.227443E-6    B1      = 4.764379E-6
+KETA    = -5.567324E-3   A1      = 0              A2      = 1
+RDSW    = 923.7832391    PRWG    = -3.089043E-4   PRWB    = -0.094855
+WR      = 1              WINT    = 5.838392E-8    LINT    = 1.759761E-8
+DWG     = -1.288272E-8
+DWB     = 5.449646E-9    VOFF    = -0.1076921     NFACTOR = 0
+CIT     = 0              CDSC    = 8.530932E-4    CDSCD   = 1.554386E-4
+CDSCB   = 1.940792E-4    ETA0    = 0.0298638      ETAB    = -3.113611E-3
+DSUB    = 0.3695329      PCLM    = 1.0357865      PDIBLC1 = 0.0176042
+PDIBLC2 = 4.154589E-3    PDIBLCB = 0.1            DROUT   = 0.5839275
+PSCBE1  = 7.231401E9     PSCBE2  = 5E-10          PVAG    = 0.3898063
+DELTA   = 0.01           MOBMOD  = 1              PRT     = 0
+UTE     = -1.5           KT1     = -0.11          KT1L    = 0
+KT2     = 0.022          UA1     = 4.31E-9        UB1     = -7.61E-18
+UC1     = -5.6E-11       AT      = 3.3E4          WL      = 0
+WLN     = 1              WW      = 0              WWN     = 1
+WWL     = 0              LL      = 0              LLN     = 1
+LW      = 0              LWN     = 1              LWL     = 0
+CAPMOD  = 2              XPART   = 0.4            CGDO    = 3.67E-10
+CGSO    = 3.67E-10       CGBO    = 0              CJ      = 9.366619E-4
+PB      = 0.8472082      MJ      = 0.3782709      CJSW    = 1.705874E-10
+PBSW    = 0.6459681      MJSW    = 0.1595611      PVTH0   = -0.0153794
+PRDSW   = -150.7148427   PK2     = 1.079181E-3    WKETA   = 1.316537E-3
+LKETA   = -2.53398E-3     )
*
.MODEL PMOS PMOS (                                LEVEL   = 9
+TNOM    = 27             TOX     = 7.9E-9
+XJ      = 1.5E-7         NCH     = 1.7E17         VTH0    = -0.5874767
+K1      = 0.6644374      K2      = -0.0114964     K3      = 14.2635744
+K3B     = -3.0055422     W0      = 3.097499E-6    NLX     = 4.063655E-8
+DVT0W   = 0              DVT1W   = 5.3E6          DVT2W   = -0.032
+DVT0    = 1.531602       DVT1    = 0.6223798      DVT2    = -0.15
+U0      = 140.9814676    UA      = 2.073141E-9    UB      = 4.311698E-19
+UC      = -2.47491E-11   VSAT    = 1.907922E5     A0      = 1.1020888
+AGS     = 0.2992066      B0      = 2.685878E-6    B1      = 5E-6
+KETA    = -4.965703E-3   A1      = 0              A2      = 1
+RDSW    = 1.816999E3     PRWG    = -4.79226E-4    PRWB    = -0.0130234
+WR      = 1              WINT    = 6.05421E-8     LINT    = 1.854495E-8
+DWG     = -1.817774E-8
+DWB     = 1.258711E-9    VOFF    = -0.1150203     NFACTOR = 0
+CIT     = 0              CDSC    = 0              CDSCD   = 0
+CDSCB   = 5.062751E-4    ETA0    = 0.087128       ETAB    = -0.108095
+DSUB    = 0.859253       PCLM    = 4.3937251      PDIBLC1 = 2.62547E-3
+PDIBLC2 = 0.0116633      PDIBLCB = 0.016944       DROUT   = 0.0985252
+PSCBE1  = 2.122679E10    PSCBE2  = 9.323911E-9    PVAG    = 10.23015
+DELTA   = 0.01           MOBMOD  = 1              PRT     = 0
+UTE     = -1.5           KT1     = -0.11          KT1L    = 0
+KT2     = 0.022          UA1     = 4.31E-9        UB1     = -7.61E-18
+UC1     = -5.6E-11       AT      = 3.3E4          WL      = 0
+WLN     = 1              WW      = 0              WWN     = 1
+WWL     = 0              LL      = 0              LLN     = 1
+LW      = 0              LWN     = 1              LWL     = 0
+CAPMOD  = 2              XPART   = 0.4            CGDO    = 4.9E-10
+CGSO    = 4.9E-10        CGBO    = 0              CJ      = 8.663825E-4
+PB      = 0.99           MJ      = 0.5738763      CJSW    = 1.877938E-10
+PBSW    = 0.99           MJSW    = 0.2504781      PVTH0   = 0.0159148
+PRDSW   = -282.5443722   PK2     = 5.401242E-4    WKETA   = -1.688757E-3
+LKETA   = -0.018132       )

.END
