Diode test with missing node
VIN 1 0 PULSE ( 5 -1 0.05ms 100ns 100ns 0.1ms 0.2ms )
R1 1 2 2K
D1 3 DMOD
VMON 2 3 0
.MODEL DMOD D (IS=100FA)
.TRAN 0 0.5ms
.PRINT TRAN I(VMON) V(3) {V(3)/I(VMON)}
*
.END
