* Xyce netlist for testing various syntaxes for E-Sources

*controlling voltage
R1 1 0  1 
V1 1 0  SIN(0V 1V 1e3 0 0 0)

* linear form
E2 2 0 1 0 2
r2 2 0 1

* polynomial form
E3 3 0 poly(1) 1 0 0.0 3.0
R3 3 0 1

.tran 10u 1ms
.print tran format=probe V(1) V(2) v(3)

.end

