* Test use of .OPTIONS OUTPUT ADD_STEPNUM_COL=TRUE
*
* See SON Bug 1209 for more details.
**************************************************

V1 1 0 1
R1 1 2 1
R2 2 0 1

* step over two variables
.STEP R1 1 2 1
.STEP R2 3 8 5

.PRINT DC R1:R R2:R V(1) V(2)
.DC V1 1 25 1

.sens objfunc={V(2)} param=R2:R
.print SENS R1:R R2:R
.PRINT SENS FORMAT=NOINDEX FILE=sens-stepnum-col.cir.SENS.noindex.prn R1:R R2:R
.print SENS FORMAT=GNUPLOT FILE=sens-stepnum-col.cir.SENS.gnuplot.prn R1:R R2:R
.PRINT SENS FORMAT=SPLOT FILE=sens-stepnum-col.cir.SENS.splot.prn R1:R R2:R

.OPTIONS OUTPUT ADD_STEPNUM_COL=true
.options SENSITIVITY direct=1 adjoint=0

.end
