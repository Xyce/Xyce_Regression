Testing "sign" functionality

.param res = {sign(3,2) + sign(2,-3) + sign(1000,0)}

I1 1 0 DC -1
R1 1 0 res

.DC I1 -1 -1 -.1
.print DC I(I1) V(1)
.end
