* DC simulation for xyce

.subckt mysub d_x g_x s_x b_x dt_x
e_d d_v 0 d_x 0 1
v_d d_v d 0
f_d d_x 0 v_d   -1
e_g g_v 0 g_x 0 1
v_g g_v g 0
f_g g_x 0 v_g   -1
e_s s_v 0 s_x 0 1
v_s s_v s 0
f_s s_x 0 v_s   -1
e_b b_v 0 b_x 0 1
v_b b_v b 0
f_b b_x 0 v_b   -1
v_dt dt dt_x 0
m1 d g s b dt mymodel
+ W=10.0e-6
+ L=0.1e-6
+ AS=5e-12
+ AD=5e-12
+ PS=21e-6
+ PD=21e-6
.model mymodel nmos level=1031
+ SWJUNASYM=1
+ TR=27.0
+ DTA=0.0
+ SWGEO=1
+ QMC=1.0
+ LVARO=-1.0E-8
+ LVARL=0.0
+ LVARW=0.0
+ LAP=1.0E-8
+ WVARO=1.0E-8
+ WVARL=0.0
+ WVARW=0.0
+ WOT=0.0
+ DLQ=0.0
+ DWQ=0.0
+ VFBO=-1.1
+ VFBL=0.0
+ VFBW=0.0
+ VFBLW=0.0
+ STVFBO=5.0E-4
+ STVFBL=0.0
+ STVFBW=0.0
+ STVFBLW=0.0
+ TOXO=1.5E-9
+ EPSROXO=3.9
+ NSUBO=3.0E+23
+ NSUBW=0.0
+ WSEG=1.5E-10
+ NPCK=1.0E+24
+ NPCKW=0.0
+ WSEGP=9.0E-9
+ LPCK=5.5E-8
+ LPCKW=0.0
+ FOL1=2.0E-2
+ FOL2=5.0E-6
+ FACNEFFACO=0.8
+ FACNEFFACL=0.0
+ FACNEFFACW=0.0
+ FACNEFFACLW=0.0
+ GFACNUDO=0.1
+ GFACNUDL=0.0
+ GFACNUDLEXP=1.0
+ GFACNUDW=0.0
+ GFACNUDLW=0.0
+ VSBNUDO=0.0
+ DVSBNUDO=1.0
+ VNSUBO=0.0
+ NSLPO=0.05
+ DNSUBO=0.0
+ DPHIBO=0.0
+ DPHIBL=0.0
+ DPHIBLEXP=1.0
+ DPHIBW=0.0
+ DPHIBLW=0.0
+ DELVTACO=0.0
+ DELVTACL=0.0
+ DELVTACLEXP=1.0
+ DELVTACW=0.0
+ DELVTACLW=0.0
+ NPO=1.5E+26
+ NPL=1.0E-17
+ CTO=5.0E-15
+ CTL=0.0
+ CTLEXP=1.0
+ CTW=0.0
+ CTLW=0.0
+ TOXOVO=1.5E-9
+ TOXOVDO=2.0E-9
+ LOV=1.0E-8
+ LOVD=0.0
+ NOVO=7.5E+25
+ NOVDO=5.0E+25
+ CFL=1.0E-3
+ CFLEXP=2.0
+ CFW=5.0E-3
+ CFDO=20.0
+ CFBO=0.3
+ PSCEL=4.0E-2
+ PSCELEXP=0.6
+ PSCEW=0.0
+ PSCEBO=0.2
+ PSCEDO=0.1
+ UO=3.5E-2
+ FBET1=-0.3
+ FBET1W=0.15
+ LP1=1.5E-7
+ LP1W=-2.5E-2
+ FBET2=50.0
+ LP2=8.5E-10
+ BETW1=5.0E-2
+ BETW2=-2.0E-2
+ WBET=5.0E-10
+ STBETO=1.75
+ STBETL=-2.0E-2
+ STBETW=-2.0E-3
+ STBETLW=-3.0E-3
+ MUEO=0.6
+ MUEW=-1.2E-2
+ STMUEO=0.5
+ THEMUO=2.75
+ STTHEMUO=-0.1
+ CSO=1.0E-2
+ CSL=0.0
+ CSLEXP=1.0
+ CSW=0.0
+ CSLW=0.0
+ STCSO=-5.0
+ XCORO=0.15
+ XCORL=2.0E-3
+ XCORW=-3.0E-2
+ XCORLW=-3.5E-3
+ STXCORO=1.25
+ FETAO=1.0
+ RSW1=50.0
+ RSW2=5.0E-2
+ STRSO=-2.0
+ RSBO=0.0
+ RSGO=0.0
+ THESATO=1.0E-6
+ THESATL=0.6
+ THESATLEXP=0.75
+ THESATW=-1.0E-2
+ THESATLW=0.0
+ STTHESATO=1.5
+ STTHESATL=-2.5E-2
+ STTHESATW=-2.0E-2
+ STTHESATLW=-5.0E-3
+ THESATBO=0.15
+ THESATGO=0.75
+ AXO=20.0
+ AXL=0.2
+ ALPL=7.0E-3
+ ALPLEXP=0.6
+ ALPW=5.0E-2
+ ALP1L1=2.5E-2
+ ALP1LEXP=0.4
+ ALP1L2=0.1
+ ALP1W=8.5E-3
+ ALP2L1=0.5
+ ALP2LEXP=0.0
+ ALP2L2=0.5
+ ALP2W=-0.2
+ VPO=0.25
+ A1O=1.0
+ A1L=0.0
+ A1W=0.0
+ A2O=10.0
+ STA2O=-0.5
+ A3O=1.0
+ A3L=0.0
+ A3W=0.0
+ A4O=0.0
+ A4L=0.0
+ A4W=0.0
+ GCOO=5.0
+ IGINVLW=50.0
+ IGOVW=10.0
+ IGOVDW=0.0
+ STIGO=1.5
+ GC2O=1.0
+ GC3O=-1.0
+ CHIBO=3.1
+ AGIDLW=50.0
+ AGIDLDW=0.0
+ BGIDLO=35.0
+ BGIDLDO=41.0
+ STBGIDLO=-5.0E-4
+ STBGIDLDO=0.0
+ CGIDLO=0.15
+ CGIDLDO=0.0
+ CGBOVL=0.0
+ CFRW=5.0E-17
+ CFRDW=0.0
+ FNTO=1.0
+ NFALW=8.0E+22
+ NFBLW=3.0E+7
+ NFCLW=0.0
+ EFO=1.0
+ LINTNOI=0.0
+ ALPNOI=2.0
+ WEDGE=5.0E-8
+ WEDGEW=0.0
+ VFBEDGEO=-1.2
+ STVFBEDGEO=1.0E-4
+ STVFBEDGEL=0.0
+ STVFBEDGEW=0.0
+ STVFBEDGELW=0.0
+ DPHIBEDGEO=0.0
+ DPHIBEDGEL=0.0
+ DPHIBEDGELEXP=1.0
+ DPHIBEDGEW=0.0
+ DPHIBEDGELW=0.0
+ NSUBEDGEO=5.0E+23
+ NSUBEDGEL=0.0
+ NSUBEDGEW=0.0
+ NSUBEDGELW=0.0
+ CTEDGEO=0.0
+ CTEDGEL=0.0
+ CTEDGELEXP=1.0
+ FBETEDGE=-0.3
+ LPEDGE=1.5E-7
+ BETEDGEW=0.0
+ STBETEDGEO=1.75
+ STBETEDGEL=-2.0E-2
+ STBETEDGEW=0.0
+ STBETEDGELW=0.0
+ PSCEEDGEL=6.0E-2
+ PSCEEDGELEXP=0.6
+ PSCEEDGEW=-2.0E-3
+ PSCEBEDGEO=0.05
+ PSCEDEDGEO=0.1
+ CFEDGEL=1.0E-3
+ CFEDGELEXP=2.0
+ CFEDGEW=0.0
+ CFDEDGEO=20.0
+ CFBEDGEO=0.3
+ FNTEDGEO=1.0
+ NFAEDGELW=8.0E+22
+ NFBEDGELW=3.0E+7
+ NFCEDGELW=0.0
+ EFEDGEO=1.0
+ KVTHOWEO=0.0
+ KVTHOWEL=0.0
+ KVTHOWEW=0.0
+ KVTHOWELW=0.0
+ KUOWEO=0.0
+ KUOWEL=0.0
+ KUOWEW=0.0
+ KUOWELW=0.0
+ RGO=0.0
+ RINT=0.0
+ RVPOLY=0.0
+ RSHG=0.0
+ DLSIL=0.0
+ RSH=0.0
+ RSHD=0.0
+ RBULKO=0.0
+ RWELLO=0.0
+ RJUNDO=0.0
+ RJUNSO=0.0
+ WLOD=0.0
+ TKUO=0.0
+ LKUO=0.0
+ WKUO=0.0
+ PKUO=0.0
+ LLODKUO=0.0
+ WLODKUO=0.0
+ LKVTHO=0.0
+ WKVTHO=0.0
+ PKVTHO=0.0
+ LLODVTH=0.0
+ WLODVTH=0.0
+ STETAO=0.0
+ LODETAO=1.0
+ SCREF=1.0E-6
+ WEB=0.0
+ WEC=0.0
+ SWJUNEXP=0
+ IMAX=1.0E+3
+ TRJ=27.0
+ FREV=1.0E+3
+ VJUNREF=2.5
+ FJUNQ=0.03
+ CJORBOT=1.0E-3
+ CJORSTI=1.0E-9
+ CJORGAT=5.0E-10
+ VBIRBOT=0.75
+ VBIRSTI=1.0
+ VBIRGAT=0.75
+ PBOT=0.35
+ PSTI=0.35
+ PGAT=0.6
+ PHIGBOT=1.16
+ PHIGSTI=1.16
+ PHIGGAT=1.16
+ IDSATRBOT=5.0E-9
+ IDSATRSTI=1.0E-18
+ IDSATRGAT=1.0E-18
+ CSRHBOT=5.0E+2
+ CSRHSTI=0.0
+ CSRHGAT=1.0E+3
+ XJUNSTI=1.0E-8
+ XJUNGAT=1.0E-9
+ CTATBOT=5.0E+2
+ CTATSTI=0.0
+ CTATGAT=1.0E+3
+ MEFFTATBOT=0.25
+ MEFFTATSTI=0.25
+ MEFFTATGAT=0.25
+ CBBTBOT=1.0E-12
+ CBBTSTI=1.0E-18
+ CBBTGAT=1.0E-18
+ FBBTRBOT=1.0E+9
+ FBBTRSTI=1.0E+9
+ FBBTRGAT=1.0E+9
+ STFBBTBOT=-1.0E-3
+ STFBBTSTI=-1.0E-3
+ STFBBTGAT=-1.0E-2
+ VBRBOT=10.0
+ VBRSTI=10.0
+ VBRGAT=10.0
+ PBRBOT=3.0
+ PBRSTI=4.0
+ PBRGAT=3.0
+ VJUNREFD=2.5
+ FJUNQD=0.03
+ CJORBOTD=1.0E-3
+ CJORSTID=1.0E-9
+ CJORGATD=1.0E-9
+ VBIRBOTD=1.0
+ VBIRSTID=1.0
+ VBIRGATD=1.0
+ PBOTD=0.5
+ PSTID=0.5
+ PGATD=0.5
+ PHIGBOTD=1.16
+ PHIGSTID=1.16
+ PHIGGATD=1.16
+ IDSATRBOTD=1.0E-12
+ IDSATRSTID=1.0E-18
+ IDSATRGATD=1.0E-18
+ CSRHBOTD=1.0E+2
+ CSRHSTID=1.0E-4
+ CSRHGATD=1.0E-4
+ XJUNSTID=1.0E-7
+ XJUNGATD=1.0E-7
+ CTATBOTD=1.0E+2
+ CTATSTID=1.0E-4
+ CTATGATD=1.0E-4
+ MEFFTATBOTD=0.25
+ MEFFTATSTID=0.25
+ MEFFTATGATD=0.25
+ CBBTBOTD=1.0E-12
+ CBBTSTID=1.0E-18
+ CBBTGATD=1.0E-18
+ FBBTRBOTD=1.0E+9
+ FBBTRSTID=1.0E+9
+ FBBTRGATD=1.0E+9
+ STFBBTBOTD=-1.0E-3
+ STFBBTSTID=-1.0E-3
+ STFBBTGATD=-1.0E-3
+ VBRBOTD=10.0
+ VBRSTID=10.0
+ VBRGATD=10.0
+ PBRBOTD=4.0
+ PBRSTID=4.0
+ PBRGATD=4.0
+ RTHO=1.1E+4
+ RTHW1=990.5
+ RTHW2=14.4
+ RTHLW=15.0
+ CTHO=1.0E-7
+ CTHW1=1.0E-8
+ CTHW2=1.5
+ CTHLW=4.0
+ STRTHO=1.3
+ SWIGATE=1
+ SWIMPACT=1
+ SWGIDL=1
+ SWJUNCAP=3
+ SWEDGE=0
.ends
v_d d 0 -0.01
v_g g 0 1.0
v_s s 0 0
v_b b 0 -1.0
i_dt dt 0 0
x1 d g s b dt mysub
.step temp list 27 100
.dc v_d 0 1.2 0.01 list v_g 0.15 0.25 0.5 0.75 1.0
.print dc V(d) v(g) TEMP
+ v(dt)
.end
