Basic diode circuit testing simple parameter use in model statement

.param IS0=100FA

D1 1 0 DMOD1
V1 1 0 DC 5V

.model DMOD1 D (IS={IS0} RS=2K)
.dc V1 0 5 1
.print DC v(1) I(v1)
.end
