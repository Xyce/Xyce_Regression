Testing to make sure that "int" take integer part of real argument

.param res = {int(3.14159265)}

I1 1 0 DC -1
R1 1 0 res

.DC I1 -1 -1 -.1
.print DC I(I1) V(1)
.end
