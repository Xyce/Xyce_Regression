Test various forms of inline comments.  See README file for more details.
;inline comment followed by a non-comment line
v1 11 0 0
v2 20 0 0
r1 30 5 1k ; inline comment on a line that is not continued.
v3 5 0 0
MNORMA 11 20 30 30 MOSNORM 
;inline comment followed by continuation line
+ L=1E-4 W=1000

.dc v1 1 2 1
.print dc v(11) i(v1) i(v3)
;inline comment followed by a blank line and another inline commnt 

;another inline comment after whitespace
.MODEL MOSNORM NMOS (
+      LEVEL = 1
+        VTO = 128
+         KP = .00002
+      GAMMA = 0
+        PHI = .6
+     LAMBDA = 0
+         RD = 0.16
+         RS = 0.001
+        CBD = 10pF
+        CBS = 10pF
+         IS = 1E-14
+         PB = .8
+       CGSO = 5pF ;controls trigger pulse width at 50V & firing
+       CGDO = 10pF; la de da
+       CGBO = 10pF
+        RSH = 0.001
+         CJ = 10pF
; next continution line starts with white space
 +         MJ = .5
+       CJSW = 0.1pF
+       MJSW = .33
+         JS = 0
+ )
