Basic dual diode circuit for baseline calculation

*Tests use of subcircuit parameters  used in .model statements, when the
* parameter on the call line is also an expression.
*THIS TEST FAILS WITH RELEASE 1.1 OF XYCE, but passes with the (newer) version 
* of Xyce that's at the head of the repository when I wrote the test!  

.param IS0=100FA
V1 1 0 DC 5V
R1 1 2 2K
Vmon1 2 3 0V
XD1 3 0 DMODsub IS0={IS0}
Vmon2 2 4 0V
XD2 4 0 DMODsub IS0={2*IS0}

.subckt DMODsub 1 2 IS0=1A
.model DMOD1 D (IS={IS0})
D1 1 2 DMOD1
.ends

.dc V1 0 5 1
.print DC v(1) I(v1) I(vmon1) I(vmon2)
.end
