Testing .MEASURE lines that are mismatched with the Analysis Types
*********************************************************************
* This tests the error messages that should occur if a TRAN, NOISE or
* DC mode measure is requested for a netlist that is doing a
* .AC analysis. 
* 
* See SON Bug 889 for more details.
*
*
*********************************************************************

* Trivial high-pass filter (V-C-R) circuit
R1 b 0 2
C1 a b 1u
V1 a 0 DC 0V AC 1

.print AC v(b) 

.ac dec 5 100Hz 10e6

* Test what happens when a TRAN, NOISE or DC measure is requested for a .AC netlist
.MEASURE DC dcmax max v(b)
.MEASURE TRAN tranmax max v(b)
.MEASURE NOISE noisemax max v(b)

.END

