****************************************************
* Test allowed data formats (RI, MA and DB) in
* Touchstone2 output using a 2-Port S-Parameter
* analysis.  Also test the PRECISION and
* FILE/FILENAME qualifiers.  This test uses lower
* case for ri, ma and db.
*
* This netlist also tests that:
*
*  1) FORMAT=STD defaults to FORMAT=TOUCHSTONE2
*
*  2) The parameters DELIMITER=<val>, FREQDIGIT=<val>
*     and SPARDIGIT=<val>are all ignored
*
*  3) the .PRINT AC line should produce no output
*
****************************************************

* RC ladder circuit
* Note that all ports (P devices) must use a common
* Reference Node, which is 0 here.
P1 1  0  port=1  z0=50
P2 12 0  port=2  z0=50

C1 2 0 1e-2
Rgs 1 2 0.02

.subckt RCBlock IN OUT GND
R1 IN OUT 20
C1 IN OUT 1p
Cg1 OUT GND 1p
.ends

X1 2 3 0 RCBlock
X2 3 4 0 RCBlock
X3 4 5 0 RCBlock
X4 5 6 0 RCBlock
X5 6 7 0 RCBlock
X6 7 8 0 RCBlock
X7 8 9 0 RCBlock
X8 9 10 0 RCBlock
X9 10 11 0 RCBlock
X10 11 12 0 RCBlock

.AC DEC 10 10  1e5

* the .PRINT AC line should produce no output
.PRINT AC V(1)

* The first line requests FORMAT=STD.  That should default to TOUCHSTONE2 format.
* That first line also tests that the DELIMITER, SPARDIGIT and FREQDIGIT parameters
* are all ignored on a .LIN line.
.LIN FORMAT=STD FILE=sparams-ts2-dataFormat.cir.ri.s2p dataformat=ri PRECISION=6
+ DELIMITER=COMMA SPARDIGIT=8 FREQDIGIT=8
.LIN FORMAT=TOUCHSTONE2 FILENAME=sparams-ts2-dataFormat.cir.ma.s2p DATAFORMAT=ma PRECISION=6
.LIN FORMAT=TOUCHSTONE2 FILE=sparams-ts2-dataFormat.cir.db.s2p DATAFORMAT=db PRECISION=6

.END
