embedded sampling version of a CMOS inverter
*
* This "circuit" exists to provide a meaningful .PRINT line to xyce_verify.pl.
*
* It isn't supposed to be run, and will exit with error.
*

*COMP {v(1)}_mean       OFFSET=1.0 RELTOL=0.1
*COMP {v(1)}_meanPlus   OFFSET=1.0 RELTOL=0.1
*COMP {v(1)}_meanMinus  OFFSET=1.0 RELTOL=0.1
*COMP {v(1)}_stddev     OFFSET=1.0 RELTOL=0.1
*COMP {v(1)}_variance   OFFSET=1.0 RELTOL=0.1

.PRINT TRAN {v(1)}_mean {v(1)}_meanPlus {v(1)}_meanMinus {v(1)}_stddev {v(1)}_variance

.tran 1ns 1.5e-6

