simple RC to test HB with .STEP output
.hb 1e5
.print hb FORMAT=CSV v(1) v(2) i(v1)
.step r1 0.5k 1.5k 0.5k

.options hbint numfreq=5 saveicdata=1
.options linsol-hb prec_type=block_jacobi

v1 1 0 sin 0 1V 1e5 0 0
r1 1 2 1k
c1 2 0 2u
.end
