** NMOSFET: Benchmarking Implementation of BSIM4.6.0 by Mohan V. Dunga 12/13/2006.

** Circuit Description **
m1 2 1 0 0 p1 L=0.09u W=10.0u rgeoMod=1
vgs 1 0 -1.2 
vds 2 0 -1.2 

.dc vds 0 -1.18 -0.02 vgs 0 -1.2 -0.2

.options device Temp=100.0

.print dc v(2) v(1) i(vds)
*COMP i(vds) abstol=1e-5

.include modelcard.pmos
.end
