RAW File Output test for the N-Type JFET.
************************************************************
* This test has two purposes:
*   1) Verify that the variable type (e.g., "voltage") and 
*      variable name is correct for the JFET. This test
*      just has a non-zero source conductivity.  So, sourceprime 
*      properly shows up as an internal voltage node.  It 
*      does not test for a non-zero drain conductivity, which 
*      would also contribute an internal variable to the 
*      solution vector for the J device.
*
*   2) Verify that the data is actually correct for all of
*      the time-steps in the .RAW file output 
*
* The "gold" .RAW file output was generated by manually
* comparing that "gold" file with a .PRN file.  It was 
* generated for a limited set of fixed time-steps, so that
* a file comparison could be used to verify the test output's
* .RAW file against that "gold" .RAW file.
*
************************************************************
*
*Drain curves
Vds 1 0 5V
Vgs 2 0 pulse (0 1 1ns 1ns 1ns 1us 2us)
.options timeint method=gear newbpstepping=0
.options output initial_interval=0.5us
.tran 1ns 10us
*
Vidmon 1 1a 0
Vigmon 2 2a 0
Vismon 0 3 0

*
Jtest 1a 2a 3 SA2109 
*
.MODEL SA2109 NJF
+ LEVEL=2
+ BETA= 0.0003790
+ VTO = -3.760
+ PB = 0.650
+ LAMBDA = 0.01240
+ DELTA = 0.370;
+ THETA = 0.01120;
+ RD = 0.0
+ RS = 104.5
+ FC = 0.5
+ IS = 1.393E-10
+ AF = 1.0
+ KF = 0.05
+ CGS= 1uf
+ CGD= 1uf
*

* .PRINT statement is not actually used for .RAW output.
* It was included in the netlist so that the "gold" .RAW 
* file output could manually verified against a .PRN file
* during test development
.print tran v(1) v(1a) v(2) v(2a) v(3) N(jtest_sourceprime)
+ I(VDS) I(VGS) I(VIDMON) I(VIGMON) I(VISMON) 
 
.end

