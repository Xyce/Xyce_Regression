RAW File Output test for the BJT.
************************************************************
* This test has two purposes:
*   1) Verify that the variable type (e.g., "voltage") and 
*      variable name is correct for the BJT.  This test
*      just has a non-zero base resistance.  So, baseprime 
*      properly shows up as an internal voltage node.  It 
*      does not test for a non-zero emitter or collector 
*      resistance, which would also contribute internal 
*      variables to the solution vector for the Q device.
*
*   2) Verify that the data is actually correct for all of
*      the time-steps in the .RAW file output 
*
* The "gold" .RAW file output was generated by manually
* comparing that "gold" file with a .PRN file.  It was 
* generated for a limited set of fixed time-steps, so that
* a file comparison could be used to verify the test output's
* .RAW file against that "gold" .RAW file.
*
************************************************************
*
vie 0 1 0
vic 0 3 5
vib 0 2 pulse(0 1 1ns 1ns 1ns 1us) 
q1 3 2 1 qjunk 

.model qjunk npn
+bf=130 br=1 is=3e-14
+tf=1e-8 vjs=0.68 ne=1.6 nc=2.0 rb=450
+cje=1uf cjc=1uf cjs=1uf ikf=0.002 ikr=0.002 vaf=50 var=50
+nf=1.0 ise=0 nr=1 isc=0 irb=0 rbm=450 re=0 rc=0 vje=0.75 
+mje=0.33 xtf=0 vtf=100 itf=0 ptf=0 vjc=0.75 mjs=0 xtb=0 
+eg=1.11 xti=3 kf=0 af=1 fc=0.5 tnom=27

.options timeint method=8
.options nonlin-tran rhstol=1.0e-7
.options output initial_interval=1us
.tran 1ns 20us

* .PRINT statement is not actually used for .RAW output.
* It was included in the netslit so that the "gold" .RAW 
* file output could manually verified against a .PRN file
* during test development
.print tran v(1) v(2) v(3) n(q1_baseprime)
+ I(vib) I(vic) I(vie) 
 
.end

