* Verilog-A vbic_3T_et_cf test circuit
*.verilog "vbic_3T_et_cf.vla"

vbe bx 0  0
vcb cx bx 0
vib bx b  0
vic cx c  0
rxth dt 0 1e12
q1 c  b  0  dt vbicmodel

.model vbicmodel npn
+ level=11
+ RCX=10 RCI=10 RBX=1 RBI=10 RE=1 RBP=10 RS=10
+ IBEN=1.0e-13 RTH=100

.dc vbe 0.5 1.0 0.02
.print dc v(bx) i(vib) i(vic)
.end
