Regression test for simple normal distribution sampling

c1 1 0 1uF IC=1
R1 1 2 1K
v1 2 0 0V
*.print tran format=tecplot v(1)
.print tran v(1)
.tran 0 5ms
.options timeint reltol=1e-6 abstol=1e-6

.SAMPLING NORMAL R1 3K 1K 10

.end

