* Verilog-A vbic_3T_et_cf test circuit
* This test simulates two identical VBIC devices in parallel using the "M=2"
* instance parameter

vbe bx 0  0
vcb cx bx 0
vib bx b  0
vic cx c  0

*simulated two in parallel, but separate self-heating nodes
q1 c  b  0 vbicmodel M=2

.model vbicmodel NPN
+ level=11
+ RCX=10 RCI=10 RBX=1 RBI=10 RE=1 RBP=10 RS=10
+ IBEN=1.0e-13 RTH=100

.dc vbe 0.5 1.0 0.02
.print dc v(bx) i(vib) i(vic)
.end
