Lead current test for 2D PDE device
*
* Also tests the three allowed forms (in .print) for lead currents
* for this type of device
*
VPOS  1 0 DC 5V
*VBB   6 0 DC -2V
BBB   6 0 V={-V(T1)}
RE    1 2 2K
RB    3 4 190K

YPDE BJT 5 3 7 PDEBJT meshfile=internal.msh 
+ node = {name = collector, base, emitter}
+ sgplotlevel=0 tecplotlevel=0
+ l=2.0e-3  w=1.0e-3
+ nx=30     ny=15
+ mobmodel=carr
* The old intrinsic calculation was used to generate gold standard.
* It is inaccurate, however. 
+ useOldNi=true


* Zero volt sources acting as an ammeter to measure the
* base, collector, and emmitter currents, respectively
VMONB 6 4 0
VMONC 0 5 0
VMONE 2 7 0 

VBB T1 0 2V
RBB T1 0 1.0

.MODEL PDEBJT   ZOD  level=2

*.DC VPOS 0.0 2.0 1.0 VBB 0.0 -0.5 -0.5 

************************************
* **** Start Homotopy Setup ****
************************************
.options nonlin nlstrategy=0 searchmethod=2
+ maxstep=30 maxsearchstep=1 in_forcing=0 AZ_Tol=1.0e-6 memory=0
+ continuation=1

.options loca stepper=0 predictor=0 stepcontrol=0
+ conparam=VPOS,VBB
+ initialvalue=0.0,0.0 minvalue=0.0,0.0 maxvalue=2.0,2.0
+ initialstepsize=0.2,0.2 minstepsize=1.0e-4,1.0e-4 maxstepsize=0.2,0.2
+ aggressiveness=1.0,1.0
+ maxsteps=5000 maxnliters=200
**********************************
* **** End Homotopy Setup ****
**********************************

.options LINSOL type=klu
*.options NONLIN maxstep=70 maxsearchstep=1 searchmethod=2 
*+in_forcing=0 nlstrategy=0 debuglevel=-1

.options TIMEINT reltol=1.0e-3 abstol=1.0e-6 doubledcop=drift_diffusion
.options DEVICE numjac=0 debuglevel=0

.DC VMONC 0.0 0.0 1.0
.PRINT DC V(5) V(1) V(6) {I(VMONC)-I1(Y%PDE%BJT)} {I(VMONB)-I2(YPDE BJT)} {I(VMONE)-I3(BJT)}

.END

