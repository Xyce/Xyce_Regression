sqrt.sp SPICE FILE
.model nenh nmos
+ level = 2
+   vto = 0.779   kp = 3.52e-05   gamma = 1.04
+   phi = 0.6
+
+   cgso = 5.2e-10   cgdo = 5.2e-10
+   rsh = 25   cj = 0.00042
+   mj = 0.5   cjsw = 9e-12   mjsw = 0.33
+   tox = 5e-08   nsub = 1e+16
+   nss = 0   nfs = 1.306e+11   tpg = 1
+   xj = 3.85e-08   ld = 1e-07   uo = 400
+   ucrit = 999000   uexp = 0.001001
+   vmax = 32585.3   neff = 0.01001
+
+   delta = 1.33
.model penh pmos
+ level = 2
+   vto = -0.988   kp = 1.206e-05   gamma = 0.619
+   phi = 0.6
+
+   cgso = 4e-10   cgdo = 4e-10
+   rsh = 95   cj = 0.00025
+   mj = 0.5   cjsw = 4.5e-12   mjsw = 0.33
+   tox = 5e-08   nsub = 8.158e+14
+   nss = 0   nfs = 5.55e+09   tpg = -1
+   xj = 1.46e-07   ld = 2.52e-07   uo = 150
+   ucrit = 54941   uexp = 0.17
+   vmax = 100000   neff = 0.01001
+
+   delta = 1.129
.subckt cell 1 2 3 4 5
+ 6 7 8 9 10 11
+ 12 13 14 15 16 17
+ 18 19 20 21 22 23
+ 24 25 26 27 28 29
+ 30 31 32 33 34 35
md1 36 27 10 26 nenh l=3e-06 w=1.8e-05 
+ as=1.44e-10 ad=1.64571e-10 ps=7.8e-05 pd=6e-05 
+ nrs=0.444444 nrd=0.507936 
md2 36 28 10 35 penh l=3e-06 w=2.55e-05 
+ as=1.5075e-10 ad=9.675e-11 ps=9e-05 pd=5.7e-05 
+ nrs=0.231834 nrd=0.148789 
md3 26 38 37 26 nenh l=3e-06 w=2.85e-05 
+ as=1.1025e-10 ad=3.62499e-11 ps=6.9e-05 pd=1.66666e-05 
+ nrs=0.135734 nrd=0.044629 
md4 35 38 37 35 penh l=3e-06 w=2.25e-05 
+ as=1.6875e-10 ad=4.91666e-11 ps=6e-05 pd=2.13889e-05 
+ nrs=0.333333 nrd=0.0971192 
md5 26 31 36 26 nenh l=3e-06 w=1.35e-05 
+ as=1.23428e-10 ad=1.7171e-11 ps=4.5e-05 pd=7.89473e-06 
+ nrs=0.677248 nrd=0.0942169 
md6 26 36 39 26 nenh l=3e-06 w=1.8e-05 
+ as=8.19641e-11 ad=2.28947e-11 ps=3.98571e-05 pd=1.05263e-05 
+ nrs=0.252975 nrd=0.0706626 
md7 40 22 26 26 nenh l=3e-06 w=9e-06 
+ as=1.14474e-11 ad=4.725e-11 ps=5.26315e-06 pd=1.8e-05 
+ nrs=0.141325 nrd=0.583333 
md8 41 19 26 26 nenh l=3e-06 w=2.85e-05 
+ as=3.62499e-11 ad=1.12371e-10 ps=1.66666e-05 pd=4.88571e-05 
+ nrs=0.044629 nrd=0.138346 
md9 6 42 26 26 nenh l=3e-06 w=2.25e-05 
+ as=2.86184e-11 ad=6.40085e-11 ps=1.31579e-05 pd=3.10345e-05 
+ nrs=0.0565301 nrd=0.126437 
md10 26 8 43 26 nenh l=3e-06 w=2.7e-05 
+ as=1.06875e-10 ad=3.05263e-11 ps=4.8e-05 pd=1.40351e-05 
+ nrs=0.11875 nrd=0.0529971 
md11 26 4 3 26 nenh l=3e-06 w=3e-05 
+ as=1.31351e-10 ad=3.81578e-11 ps=7.62162e-05 pd=1.75438e-05 
+ nrs=0.145946 nrd=0.0423976 
md12 44 3 26 26 nenh l=3e-06 w=2.7e-05 
+ as=3.4342e-11 ad=8.33822e-11 ps=1.57895e-05 pd=3.49411e-05 
+ nrs=0.0471085 nrd=0.114379 
md13 26 13 45 26 nenh l=3e-06 w=3.15e-05 
+ as=4.725e-11 ad=4.00657e-11 ps=3.45e-05 pd=1.84211e-05 
+ nrs=0.047619 nrd=0.0403787 
md14 13 5 26 26 nenh l=3e-06 w=2.4e-05 
+ as=3.05263e-11 ad=9.9e-11 ps=1.40351e-05 pd=5.4e-05 
+ nrs=0.0529971 nrd=0.171875 
md15 39 29 42 26 nenh l=3e-06 w=2.4e-05 
+ as=9.9e-11 ad=1.09286e-10 ps=5.4e-05 pd=5.31428e-05 
+ nrs=0.171875 nrd=0.189732 
md16 39 30 42 35 penh l=3e-06 w=1.5e-05 
+ as=9.9e-11 ad=4.67307e-11 ps=4.5e-05 pd=2.1923e-05 
+ nrs=0.44 nrd=0.207692 
md17 35 36 39 35 penh l=3e-06 w=2.4e-05 
+ as=7.4769e-11 ad=5.24444e-11 ps=3.50769e-05 pd=2.28148e-05 
+ nrs=0.129807 nrd=0.0910493 
md18 16 38 17 26 nenh l=3e-06 w=2.1e-05 
+ as=1.53e-10 ad=1.4175e-10 ps=8.4e-05 pd=6.9e-05 
+ nrs=0.346939 nrd=0.321428 
md19 3 7 38 26 nenh l=3e-06 w=2.55e-05 
+ as=1.17068e-10 ad=1.11649e-10 ps=3.70909e-05 pd=6.47837e-05 
+ nrs=0.180035 nrd=0.171701 
md20 38 9 44 26 nenh l=3e-06 w=2.4e-05 
+ as=7.41176e-11 ad=1.10182e-10 ps=3.10588e-05 pd=3.49091e-05 
+ nrs=0.128676 nrd=0.191288 
md21 3 9 38 35 penh l=3e-06 w=1.95e-05 
+ as=7.60499e-11 ad=1.56e-10 ps=2.73e-05 pd=6.93333e-05 
+ nrs=0.2 nrd=0.410256 
md22 38 7 44 35 penh l=3e-06 w=2.55e-05 
+ as=9.83569e-11 ad=9.94498e-11 ps=4.80857e-05 pd=3.57e-05 
+ nrs=0.15126 nrd=0.152941 
md23 35 38 15 35 penh l=3e-06 w=1.05e-05 
+ as=6.3e-11 ad=2.29444e-11 ps=4.2e-05 pd=9.98148e-06 
+ nrs=0.571428 nrd=0.208113 
md24 40 22 35 35 penh l=3e-06 w=9e-06 
+ as=1.96667e-11 ad=3.65294e-11 ps=8.55554e-06 pd=1.8e-05 
+ nrs=0.242798 nrd=0.45098 
md25 41 19 35 35 penh l=3e-06 w=2.7e-05 
+ as=5.89999e-11 ad=9.98999e-11 ps=2.56666e-05 pd=3.96e-05 
+ nrs=0.0809326 nrd=0.137037 
md26 6 42 35 35 penh l=3e-06 w=1.65e-05 
+ as=3.60555e-11 ad=3.84051e-11 ps=1.56852e-05 pd=2.27586e-05 
+ nrs=0.132435 nrd=0.141066 
md27 35 8 43 35 penh l=3e-06 w=3e-05 
+ as=7.07142e-11 ad=6.55555e-11 ps=3.77142e-05 pd=2.85185e-05 
+ nrs=0.0785713 nrd=0.0728395 
md28 35 4 3 35 penh l=3e-06 w=2.1e-05 
+ as=1.68e-10 ad=4.58889e-11 ps=7.46666e-05 pd=1.9963e-05 
+ nrs=0.380952 nrd=0.104056 
md29 44 3 35 35 penh l=3e-06 w=2.7e-05 
+ as=5.89999e-11 ad=1.04143e-10 ps=2.56666e-05 pd=5.09142e-05 
+ nrs=0.0809326 nrd=0.142857 
md30 35 13 46 35 penh l=3e-06 w=2.7e-05 
+ as=4.5439e-11 ad=5.89999e-11 ps=3.29268e-05 pd=2.56666e-05 
+ nrs=0.0623305 nrd=0.0809326 
md31 13 5 35 35 penh l=3e-06 w=2.85e-05 
+ as=6.22777e-11 ad=1.1475e-10 ps=2.70926e-05 pd=6.6e-05 
+ nrs=0.076673 nrd=0.141274 
md32 22 37 34 26 nenh l=3e-06 w=2.7e-05 
+ as=1.85143e-10 ad=6.36428e-11 ps=7.13571e-05 pd=3.54857e-05 
+ nrs=0.253968 nrd=0.0873015 
md33 23 38 22 26 nenh l=3e-06 w=2.55e-05 
+ as=6.01071e-11 ad=5.43552e-11 ps=3.35142e-05 pd=3.08684e-05 
+ nrs=0.0924368 nrd=0.0835912 
md34 22 38 34 35 penh l=3e-06 w=1.8e-05 
+ as=7.16086e-11 ad=8.1e-11 ps=2.66086e-05 pd=2.81739e-05 
+ nrs=0.221014 nrd=0.25 
md35 23 37 22 35 penh l=3e-06 w=1.65e-05 
+ as=7.425e-11 ad=4.51323e-11 ps=2.5826e-05 pd=2.42647e-05 
+ nrs=0.272727 nrd=0.165775 
md36 34 38 40 26 nenh l=3e-06 w=1.5e-05 
+ as=7.875e-11 ad=1.02857e-10 ps=3e-05 pd=3.96428e-05 
+ nrs=0.35 nrd=0.457142 
md37 34 37 40 35 penh l=3e-06 w=1.65e-05 
+ as=6.69705e-11 ad=6.56412e-11 ps=3.3e-05 pd=2.43913e-05 
+ nrs=0.245989 nrd=0.241107 
md38 18 27 19 26 nenh l=3e-06 w=2.25e-05 
+ as=1.845e-10 ad=1.215e-10 ps=6.9e-05 pd=6e-05 
+ nrs=0.364444 nrd=0.24 
md39 19 28 18 35 penh l=3e-06 w=2.4e-05 
+ as=1.3275e-10 ad=1.17e-10 ps=6.3e-05 pd=5.7e-05 
+ nrs=0.230469 nrd=0.203125 
md40 4 29 41 26 nenh l=3e-06 w=2.4e-05 
+ as=9.46285e-11 ad=1.1475e-10 ps=4.11428e-05 pd=6.6e-05 
+ nrs=0.164286 nrd=0.199219 
md41 4 30 41 35 penh l=3e-06 w=1.8e-05 
+ as=6.65999e-11 ad=9.9e-11 ps=2.64e-05 pd=5.1e-05 
+ nrs=0.205555 nrd=0.305555 
md42 5 12 6 26 nenh l=3e-06 w=2.1e-05 
+ as=5.97413e-11 ad=4.63235e-11 ps=2.89655e-05 pd=2.71765e-05 
+ nrs=0.135468 nrd=0.105042 
md43 5 2 6 35 penh l=3e-06 w=2.7e-05 
+ as=6.28448e-11 ad=8.95908e-11 ps=3.72413e-05 pd=3.6e-05 
+ nrs=0.0862068 nrd=0.122896 
md44 43 11 5 26 nenh l=3e-06 w=3e-05 
+ as=6.61764e-11 ad=1.06875e-10 ps=3.88235e-05 pd=4.8e-05 
+ nrs=0.0735292 nrd=0.11875 
md45 43 1 5 35 penh l=3e-06 w=2.25e-05 
+ as=7.46589e-11 ad=5.30356e-11 ps=3e-05 pd=2.82857e-05 
+ nrs=0.147474 nrd=0.104762 
md46 45 14 23 26 nenh l=3e-06 w=3.15e-05 
+ as=6.71447e-11 ad=4.725e-11 ps=3.81315e-05 pd=3.45e-05 
+ nrs=0.0676692 nrd=0.047619 
md47 46 14 23 35 penh l=3e-06 w=3.45e-05 
+ as=9.43676e-11 ad=5.80609e-11 ps=5.07352e-05 pd=4.20731e-05 
+ nrs=0.0792838 nrd=0.0487804 
c1 21 26 8e-18
c2 24 26 4e-18
c3 26 33 1e-17
c4 26 32 9e-18
c5 7 26 4e-18
c6 9 26 1.4e-17
c7 13 26 2.10751e-14
c8 26 28 2.4e-17
c9 23 26 1.50012e-15
c10 8 26 7e-18
c11 44 26 1.52525e-15
c12 14 26 1.5e-17
c13 26 31 2.5e-17
c14 3 26 1.19855e-14
c15 43 26 2.16525e-15
c16 11 26 5e-18
c17 5 26 3.45852e-14
c18 12 26 4e-18
c19 6 26 3.18512e-15
c20 4 26 1.25801e-14
c21 26 30 1.2e-17
c22 26 29 1.2e-17
c23 18 26 4.26012e-15
c24 26 34 4.16525e-15
c25 26 27 2.3e-17
c26 41 26 1.62025e-15
c27 19 26 1.67401e-14
c28 40 26 1.47512e-15
c29 22 26 7.01512e-15
c30 15 26 4.335e-15
c31 16 26 6.53e-15
c32 26 38 4.04802e-14
c33 17 26 9.80125e-16
c34 39 26 8.7025e-16
c35 42 26 9.86012e-15
c36 36 26 1.25852e-14
c37 25 26 3.3e-17
c38 26 37 2.55751e-14
c39 10 26 1.14525e-15
.ends cell
.subckt boost 1 2 3 4 5
+ 6 7 8 9 10 11
+ 12 13 14 15 16 17
+ 18
md48 5 10 19 9 nenh l=3e-06 w=2.25e-05 
+ as=6.27692e-11 ad=1.74687e-10 ps=4.44615e-05 pd=6.06666e-05 
+ nrs=0.0965308 nrd=0.459401 
md49 20 4 5 9 nenh l=3e-06 w=3.45e-05 
+ as=3.09062e-10 ad=5.39062e-11 ps=0.000107333 pd=3.88125e-05 
+ nrs=0.259662 nrd=0.0452898 
md50 21 6 5 18 penh l=3e-06 w=3.9e-05 
+ as=5.83536e-10 ad=5.85e-11 ps=0.0002184 pd=4.2e-05 
+ nrs=0.383653 nrd=0.0384615 
md51 22 10 5 18 penh l=3e-06 w=2.1e-05 
+ as=3.14212e-10 ad=5.16922e-11 ps=0.0001176 pd=3.01538e-05 
+ nrs=0.712499 nrd=0.117216 
md52 19 6 9 9 nenh l=3e-06 w=3.3e-05 
+ as=7.31417e-11 ad=8.12307e-11 ps=2.7582e-05 pd=5.75384e-05 
+ nrs=0.0671641 nrd=0.074592 
md53 9 6 23 9 nenh l=3e-06 w=3e-05 
+ as=1.26e-10 ad=6.64924e-11 ps=7.2e-05 pd=2.50746e-05 
+ nrs=0.14 nrd=0.0738804 
md54 9 23 20 9 nenh l=3e-06 w=3.75e-05 
+ as=5.85937e-11 ad=8.31155e-11 ps=4.21874e-05 pd=3.13433e-05 
+ nrs=0.0416666 nrd=0.0591044 
md55 18 4 21 18 penh l=3e-06 w=3.9e-05 
+ as=5.85e-11 ad=5.85e-11 ps=4.2e-05 pd=3.19091e-05 
+ nrs=0.0384615 nrd=0.0384615 
md56 18 23 22 18 penh l=3e-06 w=3.75e-05 
+ as=9.23076e-11 ad=5.625e-11 ps=5.38461e-05 pd=3.06818e-05 
+ nrs=0.0656409 nrd=0.04 
md57 18 6 23 18 penh l=3e-06 w=2.25e-05 
+ as=1.6875e-10 ad=3.375e-11 ps=6e-05 pd=1.84091e-05 
+ nrs=0.333333 nrd=0.0666666 
c40 5 9 8.69499e-15
c41 9 13 2e-18
c42 9 14 2e-18
c43 9 11 2e-18
c44 9 15 3e-18
c45 3 9 5e-18
c46 9 17 3e-18
c47 20 9 1.60063e-16
c48 23 9 2.60751e-14
c49 4 9 1.3e-17
c50 9 10 1.4e-17
c51 21 9 1.4e-16
c52 6 9 3.8e-17
.ends boost
xcell#2 3 4 5 6 7
+ 8 7 8 9 10 4
+ 3 9 5 11 12 13
+ 14 15 14 16 17 18
+ 4 3 0 19 20 21
+ 22 23 24 10 25 1 cell
xcell#3 3 4 37 38 39
+ 40 41 40 39 8 4
+ 3 41 38 11 42 12
+ 16 43 14 25 18 44
+ 4 3 0 19 20 21
+ 22 23 24 10 45 1 cell
xcell#4 3 4 57 58 59
+ 60 61 60 59 40 4
+ 3 61 58 11 11 42
+ 25 62 14 45 44 63
+ 4 3 0 19 20 21
+ 22 23 24 10 64 1 cell
xboost#0 64 45 60 14 76
+ 11 4 3 0 63 19
+ 20 21 22 23 24 10
+ 1
+ boost
xcell#5 4 3 82 83 84
+ 85 84 85 86 60 3
+ 4 86 82 87 88 0
+ 45 89 76 64 76 90
+ 4 3 0 19 20 21
+ 22 23 24 10 91 1 cell
xcell#6 4 3 103 104 105
+ 106 105 106 107 85 3
+ 4 107 103 87 108 88
+ 64 109 76 91 90 110
+ 4 3 0 19 20 21
+ 22 23 24 10 111 1 cell
xcell#7 4 3 123 124 125
+ 126 127 126 125 106 3
+ 4 127 124 87 128 108
+ 91 129 76 111 110 130
+ 4 3 0 19 20 21
+ 22 23 24 10 131 1 cell
xcell#8 4 3 143 144 145
+ 146 147 146 145 126 3
+ 4 147 144 87 87 128
+ 111 148 76 131 130 149
+ 4 3 0 19 20 21
+ 22 23 24 10 150 1 cell
xboost#1 150 131 146 76 162
+ 87 4 3 0 149 19
+ 20 21 22 23 24 10
+ 1
+ boost
xcell#9 3 4 168 169 170
+ 171 170 171 172 146 4
+ 3 172 168 173 174 0
+ 131 175 162 150 162 176
+ 4 3 0 19 20 21
+ 22 23 24 10 177 1 cell
xcell#10 3 4 189 190 191
+ 192 191 192 193 171 4
+ 3 193 189 173 194 174
+ 150 195 162 177 176 196
+ 4 3 0 19 20 21
+ 22 23 24 10 197 1 cell
xcell#11 3 4 209 210 211
+ 212 213 212 211 192 4
+ 3 213 210 173 214 194
+ 177 215 162 197 196 216
+ 4 3 0 19 20 21
+ 22 23 24 10 217 1 cell
xcell#12 3 4 229 230 231
+ 232 233 232 231 212 4
+ 3 233 230 173 173 214
+ 197 234 162 217 216 235
+ 4 3 0 19 20 21
+ 22 23 24 10 236 1 cell
xboost#2 236 217 232 162 248
+ 173 4 3 0 235 19
+ 20 21 22 23 24 10
+ 1
+ boost
xcell#13 4 3 254 255 256
+ 257 256 257 258 232 3
+ 4 258 254 259 260 0
+ 217 261 248 236 248 262
+ 4 3 0 19 20 21
+ 22 23 24 10 263 1 cell
xcell#14 4 3 275 276 277
+ 278 277 278 279 257 3
+ 4 279 275 259 280 260
+ 236 281 248 263 262 282
+ 4 3 0 19 20 21
+ 22 23 24 10 283 1 cell
xcell#15 4 3 295 296 297
+ 298 299 298 297 278 3
+ 4 299 296 259 300 280
+ 263 301 248 283 282 302
+ 4 3 0 19 20 21
+ 22 23 24 10 303 1 cell
xcell#16 4 3 315 316 317
+ 318 319 318 317 298 3
+ 4 319 316 259 259 300
+ 283 320 248 303 302 321
+ 4 3 0 19 20 21
+ 22 23 24 10 322 1 cell
xboost#3 322 303 318 248 334
+ 259 4 3 0 321 19
+ 20 21 22 23 24 10
+ 1
+ boost
xcell#17 3 4 340 341 342
+ 343 342 343 344 318 4
+ 3 344 340 345 346 0
+ 303 347 334 322 334 348
+ 4 3 0 19 20 21
+ 22 23 24 10 349 1 cell
xcell#18 3 4 361 362 363
+ 364 363 364 365 343 4
+ 3 365 361 345 366 346
+ 322 367 334 349 348 368
+ 4 3 0 19 20 21
+ 22 23 24 10 369 1 cell
xcell#19 3 4 381 382 383
+ 384 385 384 383 364 4
+ 3 385 382 345 386 366
+ 349 387 334 369 368 388
+ 4 3 0 19 20 21
+ 22 23 24 10 389 1 cell
xcell#20 3 4 401 402 403
+ 404 405 404 403 384 4
+ 3 405 402 345 345 386
+ 369 406 334 389 388 407
+ 4 3 0 19 20 21
+ 22 23 24 10 408 1 cell
xboost#4 408 389 404 334 420
+ 345 4 3 0 407 19
+ 20 21 22 23 24 10
+ 1
+ boost
xcell#21 4 3 426 427 428
+ 429 428 429 430 404 3
+ 4 430 426 431 432 0
+ 389 433 420 408 420 434
+ 4 3 0 19 20 21
+ 22 23 24 10 435 1 cell
xcell#22 4 3 447 448 449
+ 450 449 450 451 429 3
+ 4 451 447 431 452 432
+ 408 453 420 435 434 454
+ 4 3 0 19 20 21
+ 22 23 24 10 455 1 cell
xcell#23 4 3 467 468 469
+ 470 471 470 469 450 3
+ 4 471 468 431 472 452
+ 435 473 420 455 454 474
+ 4 3 0 19 20 21
+ 22 23 24 10 475 1 cell
xcell#24 4 3 487 488 489
+ 490 491 490 489 470 3
+ 4 491 488 431 431 472
+ 455 492 420 475 474 493
+ 4 3 0 19 20 21
+ 22 23 24 10 494 1 cell
md58 0 507 506 0 nenh l=3e-06 w=2.85e-05 
+ as=1.1025e-10 ad=1.19893e-11 ps=6.9e-05 pd=4.52124e-06 
+ nrs=0.135734 nrd=0.0147607 
md59 0 4 3 0 nenh l=3e-06 w=3.45e-05 
+ as=2.2275e-10 ad=1.45134e-11 ps=8.4e-05 pd=5.47308e-06 
+ nrs=0.187145 nrd=0.0121936 
md60 4 508 0 0 nenh l=3e-06 w=3.45e-05 
+ as=1.45134e-11 ad=3.3075e-10 ps=5.47308e-06 pd=0.000108 
+ nrs=0.0121936 nrd=0.277883 
md61 509 14 0 0 nenh l=3e-06 w=9e-06 
+ as=3.78611e-12 ad=4.725e-11 ps=1.42776e-06 pd=1.8e-05 
+ nrs=0.0467421 nrd=0.583333 
md62 0 511 510 0 nenh l=3e-06 w=3.15e-05 
+ as=1.50609e-10 ad=1.32514e-11 ps=7.48125e-05 pd=4.99716e-06 
+ nrs=0.151786 nrd=0.0133549 
md63 13 506 0 0 nenh l=3e-06 w=2.1e-05 
+ as=8.83426e-12 ad=6.3e-11 ps=3.33144e-06 pd=4.8e-05 
+ nrs=0.0200323 nrd=0.142857 
md64 0 23 43 0 nenh l=3e-06 w=2.25e-05 
+ as=8.325e-11 ad=9.46529e-12 ps=5.1e-05 pd=3.5694e-06 
+ nrs=0.164444 nrd=0.0186968 
md65 0 23 62 0 nenh l=3e-06 w=2.25e-05 
+ as=8.325e-11 ad=9.46529e-12 ps=5.1e-05 pd=3.5694e-06 
+ nrs=0.164444 nrd=0.0186968 
md66 0 23 89 0 nenh l=3e-06 w=2.25e-05 
+ as=8.325e-11 ad=9.46529e-12 ps=5.1e-05 pd=3.5694e-06 
+ nrs=0.164444 nrd=0.0186968 
md67 0 23 109 0 nenh l=3e-06 w=2.25e-05 
+ as=8.325e-11 ad=9.46529e-12 ps=5.1e-05 pd=3.5694e-06 
+ nrs=0.164444 nrd=0.0186968 
md68 0 23 215 0 nenh l=3e-06 w=2.25e-05 
+ as=8.325e-11 ad=9.46529e-12 ps=5.1e-05 pd=3.5694e-06 
+ nrs=0.164444 nrd=0.0186968 
md69 0 23 234 0 nenh l=3e-06 w=2.25e-05 
+ as=8.325e-11 ad=9.46529e-12 ps=5.1e-05 pd=3.5694e-06 
+ nrs=0.164444 nrd=0.0186968 
md70 0 23 261 0 nenh l=3e-06 w=2.25e-05 
+ as=8.325e-11 ad=9.46529e-12 ps=5.1e-05 pd=3.5694e-06 
+ nrs=0.164444 nrd=0.0186968 
md71 0 23 281 0 nenh l=3e-06 w=2.25e-05 
+ as=8.325e-11 ad=9.46529e-12 ps=5.1e-05 pd=3.5694e-06 
+ nrs=0.164444 nrd=0.0186968 
md72 0 23 387 0 nenh l=3e-06 w=2.25e-05 
+ as=8.325e-11 ad=9.46529e-12 ps=5.1e-05 pd=3.5694e-06 
+ nrs=0.164444 nrd=0.0186968 
md73 0 23 406 0 nenh l=3e-06 w=2.25e-05 
+ as=8.325e-11 ad=9.46529e-12 ps=5.1e-05 pd=3.5694e-06 
+ nrs=0.164444 nrd=0.0186968 
md74 0 23 433 0 nenh l=3e-06 w=2.25e-05 
+ as=8.325e-11 ad=9.46529e-12 ps=5.1e-05 pd=3.5694e-06 
+ nrs=0.164444 nrd=0.0186968 
md75 0 23 453 0 nenh l=3e-06 w=2.25e-05 
+ as=8.325e-11 ad=9.46529e-12 ps=5.1e-05 pd=3.5694e-06 
+ nrs=0.164444 nrd=0.0186968 
md76 512 431 0 0 nenh l=3e-06 w=3.3e-05 
+ as=1.38824e-11 ad=8.12307e-11 ps=5.23512e-06 pd=5.75384e-05 
+ nrs=0.0127479 nrd=0.074592 
md77 0 431 513 0 nenh l=3e-06 w=3e-05 
+ as=1.2375e-10 ad=1.26204e-11 ps=7.2e-05 pd=4.7592e-06 
+ nrs=0.1375 nrd=0.0140226 
md78 0 513 514 0 nenh l=3e-06 w=3.75e-05 
+ as=5.85937e-11 ad=1.57755e-11 ps=4.21874e-05 pd=5.94901e-06 
+ nrs=0.0416666 nrd=0.0112181 
md79 1 507 506 1 penh l=3e-06 w=3.3e-05 
+ as=1.1925e-10 ad=8.39845e-12 ps=7.2e-05 pd=4.58097e-06 
+ nrs=0.109504 nrd=0.00771207 
md80 1 4 3 1 penh l=3e-06 w=3.45e-05 
+ as=2.6775e-10 ad=8.7802e-12 ps=8.7e-05 pd=4.78919e-06 
+ nrs=0.224953 nrd=0.00737677 
md81 4 508 1 1 penh l=3e-06 w=3.45e-05 
+ as=8.7802e-12 ad=2.5875e-10 ps=4.78919e-06 pd=8.4e-05 
+ nrs=0.00737677 nrd=0.217391 
md82 509 14 1 1 penh l=3e-06 w=9e-06 
+ as=2.29049e-12 ad=3.65294e-11 ps=1.24936e-06 pd=1.8e-05 
+ nrs=0.0282776 nrd=0.45098 
md83 1 511 510 1 penh l=3e-06 w=2.1e-05 
+ as=1.20167e-10 ad=5.34447e-12 ps=4.2e-05 pd=2.91516e-06 
+ nrs=0.272486 nrd=0.012119 
md84 511 24 1 1 penh l=3e-06 w=2.25e-05 
+ as=5.72622e-12 ad=1.0125e-10 ps=3.12339e-06 pd=4.78125e-05 
+ nrs=0.011311 nrd=0.2 
md85 1 506 17 1 penh l=3e-06 w=3.45e-05 
+ as=1.36985e-10 ad=8.7802e-12 ps=5.88529e-05 pd=4.78919e-06 
+ nrs=0.115089 nrd=0.00737677 
md86 11 506 1 1 penh l=3e-06 w=1.5e-05 
+ as=3.81748e-12 ad=9.9e-11 ps=2.08226e-06 pd=5.4e-05 
+ nrs=0.0169666 nrd=0.44 
md87 1 24 15 1 penh l=3e-06 w=2.55e-05 
+ as=7.65e-11 ad=6.48971e-12 ps=5.7e-05 pd=3.53984e-06 
+ nrs=0.117647 nrd=0.00998032 
md88 1 24 129 1 penh l=3e-06 w=2.55e-05 
+ as=7.65e-11 ad=6.48971e-12 ps=5.7e-05 pd=3.53984e-06 
+ nrs=0.117647 nrd=0.00998032 
md89 1 24 148 1 penh l=3e-06 w=2.55e-05 
+ as=7.65e-11 ad=6.48971e-12 ps=5.7e-05 pd=3.53984e-06 
+ nrs=0.117647 nrd=0.00998032 
md90 1 24 175 1 penh l=3e-06 w=2.55e-05 
+ as=7.65e-11 ad=6.48971e-12 ps=5.7e-05 pd=3.53984e-06 
+ nrs=0.117647 nrd=0.00998032 
md91 1 24 195 1 penh l=3e-06 w=2.55e-05 
+ as=7.65e-11 ad=6.48971e-12 ps=5.7e-05 pd=3.53984e-06 
+ nrs=0.117647 nrd=0.00998032 
md92 1 24 301 1 penh l=3e-06 w=2.55e-05 
+ as=7.65e-11 ad=6.48971e-12 ps=5.7e-05 pd=3.53984e-06 
+ nrs=0.117647 nrd=0.00998032 
md93 1 24 320 1 penh l=3e-06 w=2.55e-05 
+ as=7.65e-11 ad=6.48971e-12 ps=5.7e-05 pd=3.53984e-06 
+ nrs=0.117647 nrd=0.00998032 
md94 1 24 347 1 penh l=3e-06 w=2.55e-05 
+ as=7.65e-11 ad=6.48971e-12 ps=5.7e-05 pd=3.53984e-06 
+ nrs=0.117647 nrd=0.00998032 
md95 1 24 367 1 penh l=3e-06 w=2.55e-05 
+ as=7.65e-11 ad=6.48971e-12 ps=5.7e-05 pd=3.53984e-06 
+ nrs=0.117647 nrd=0.00998032 
md96 1 24 473 1 penh l=3e-06 w=2.55e-05 
+ as=7.65e-11 ad=6.48971e-12 ps=5.7e-05 pd=3.53984e-06 
+ nrs=0.117647 nrd=0.00998032 
md97 1 24 492 1 penh l=3e-06 w=2.55e-05 
+ as=7.65e-11 ad=6.48971e-12 ps=5.7e-05 pd=3.53984e-06 
+ nrs=0.117647 nrd=0.00998032 
md98 1 420 515 1 penh l=3e-06 w=3.9e-05 
+ as=5.85e-11 ad=9.92543e-12 ps=4.2e-05 pd=5.41388e-06 
+ nrs=0.0384615 nrd=0.0065256 
md99 1 513 516 1 penh l=3e-06 w=3.75e-05 
+ as=9.23076e-11 ad=9.54369e-12 ps=5.38461e-05 pd=5.20565e-06 
+ nrs=0.0656409 nrd=0.00678661 
md100 1 431 513 1 penh l=3e-06 w=2.25e-05 
+ as=1.6875e-10 ad=5.72622e-12 ps=6e-05 pd=3.12339e-06 
+ nrs=0.333333 nrd=0.011311 
md101 14 507 16 0 nenh l=3e-06 w=2.7e-05 
+ as=2.08286e-10 ad=6.36428e-11 ps=6.75e-05 pd=3.54857e-05 
+ nrs=0.285714 nrd=0.0873015 
md102 17 506 14 0 nenh l=3e-06 w=2.55e-05 
+ as=6.01071e-11 ad=1.3275e-10 ps=3.35142e-05 pd=6.6e-05 
+ nrs=0.0924368 nrd=0.204152 
md103 14 506 16 1 penh l=3e-06 w=1.8e-05 
+ as=7.16086e-11 ad=8.1e-11 ps=2.66086e-05 pd=2.81739e-05 
+ nrs=0.221014 nrd=0.25 
md104 17 507 14 1 penh l=3e-06 w=1.65e-05 
+ as=7.425e-11 ad=6.55146e-11 ps=2.5826e-05 pd=2.8147e-05 
+ nrs=0.272727 nrd=0.240642 
md105 16 506 509 0 nenh l=3e-06 w=1.5e-05 
+ as=7.875e-11 ad=1.15714e-10 ps=3e-05 pd=3.75e-05 
+ nrs=0.35 nrd=0.514285 
md106 16 507 509 1 penh l=3e-06 w=1.65e-05 
+ as=6.69705e-11 ad=6.56412e-11 ps=3.3e-05 pd=2.43913e-05 
+ nrs=0.245989 nrd=0.241107 
md107 510 21 508 0 nenh l=3e-06 w=1.65e-05 
+ as=1.2375e-10 ad=7.88906e-11 ps=4.8e-05 pd=3.91875e-05 
+ nrs=0.454545 nrd=0.289773 
md108 510 22 508 1 penh l=3e-06 w=1.95e-05 
+ as=1.4625e-10 ad=1.11583e-10 ps=5.4e-05 pd=3.9e-05 
+ nrs=0.384615 nrd=0.293447 
md109 10 19 511 0 nenh l=3e-06 w=1.8e-05 
+ as=1.35e-10 ad=1.20938e-10 ps=7.5e-05 pd=4.2e-05 
+ nrs=0.416667 nrd=0.373264 
md110 10 20 511 1 penh l=3e-06 w=2.55e-05 
+ as=1.1475e-10 ad=7.65e-11 ps=5.41875e-05 pd=5.7e-05 
+ nrs=0.176471 nrd=0.117647 
md111 10 493 512 0 nenh l=3e-06 w=2.25e-05 
+ as=6.27692e-11 ad=1.31015e-10 ps=4.44615e-05 pd=4.54999e-05 
+ nrs=0.0965308 nrd=0.344551 
md112 514 420 10 0 nenh l=3e-06 w=3.45e-05 
+ as=2.31797e-10 ad=5.39062e-11 ps=8.04999e-05 pd=3.88125e-05 
+ nrs=0.194746 nrd=0.0452898 
md113 515 431 10 1 penh l=3e-06 w=3.9e-05 
+ as=4.95787e-10 ad=5.85e-11 ps=0.00020085 pd=4.2e-05 
+ nrs=0.325961 nrd=0.0384615 
md114 516 493 10 1 penh l=3e-06 w=2.1e-05 
+ as=2.66962e-10 ad=5.16922e-11 ps=0.00010815 pd=3.01538e-05 
+ nrs=0.605356 nrd=0.117216 
c53 0 21 1.8e-17
c54 0 22 1.7e-17
c55 0 19 2.4e-17
c56 0 23 1.5e-17
c57 0 24 2.4e-17
c58 0 20 2.2e-17
c59 3 0 7.76725e-15
c60 490 0 2e-18
c61 4 0 1.3059e-14
c62 514 0 1.60063e-16
c63 513 0 2.5805e-14
c64 420 0 1.3e-17
c65 0 493 1.4e-17
c66 515 0 1.4e-16
c67 0 10 7.00959e-14
c68 431 0 3.8e-17
c69 492 0 5.5e-17
c70 473 0 5.5e-17
c71 367 0 5.5e-17
c72 347 0 5.5e-17
c73 320 0 5.5e-17
c74 301 0 5.5e-17
c75 195 0 5.5e-17
c76 175 0 5.5e-17
c77 148 0 5.5e-17
c78 129 0 5.5e-17
c79 15 0 5.5e-17
c80 11 0 6.30063e-16
c81 17 0 2.60025e-15
c82 0 16 3.0455e-15
c83 0 511 1.1e-14
c84 0 510 3.56525e-15
c85 508 0 7.38499e-15
c86 0 509 1.47512e-15
c87 0 14 2.20151e-14
c88 0 506 3.94101e-14
c89 0 507 2.6e-17
c90 6 0 1e-15
c91 37 0 1e-15
c92 57 0 1e-15
c93 83 0 1e-15
c94 104 0 1e-15
c95 123 0 1e-15
c96 143 0 1e-15
c97 169 0 1e-15
c98 190 0 1e-15
c99 209 0 1e-15
c100 229 0 1e-15
c101 255 0 1e-15
c102 276 0 1e-15
c103 295 0 1e-15
c104 315 0 1e-15
c105 341 0 1e-15
c106 362 0 1e-15
c107 381 0 1e-15
c108 401 0 1e-15
c109 427 0 1e-15
c110 448 0 1e-15
c111 467 0 1e-15
c112 487 0 1e-15
VNResetQ1H 19 0 pwl (0 0 1.4e-07 0 1.41e-07 5 2.2e-07 5 
+ 2.21e-07 0 3.4e-07 0 3.41e-07 5 4.2e-07 5 
+ 4.21e-07 0 5.4e-07 0 5.41e-07 5 6.2e-07 5 
+ 6.21e-07 0 7.4e-07 0 7.41e-07 5 8.2e-07 5 
+ 8.21e-07 0 9e-07 0 )
VNResetQ1L 20 0 pwl (0 5 1.4e-07 5 1.41e-07 0 2.2e-07 0 
+ 2.21e-07 5 3.4e-07 5 3.41e-07 0 4.2e-07 0 
+ 4.21e-07 5 5.4e-07 5 5.41e-07 0 6.2e-07 0 
+ 6.21e-07 5 7.4e-07 5 7.41e-07 0 8.2e-07 0 
+ 8.21e-07 5 9e-07 5 )
VPhi2H 21 0 pwl (0 5 1.2e-07 5 1.21e-07 0 2.4e-07 0 
+ 2.41e-07 5 3.2e-07 5 3.21e-07 0 4.4e-07 0 
+ 4.41e-07 5 5.2e-07 5 5.21e-07 0 6.4e-07 0 
+ 6.41e-07 5 7.2e-07 5 7.21e-07 0 8.4e-07 0 
+ 8.41e-07 5 9e-07 5 )
VPhi2L 22 0 pwl (0 0 1.2e-07 0 1.21e-07 5 2.4e-07 5 
+ 2.41e-07 0 3.2e-07 0 3.21e-07 5 4.4e-07 5 
+ 4.41e-07 0 5.2e-07 0 5.21e-07 5 6.4e-07 5 
+ 6.41e-07 0 7.2e-07 0 7.21e-07 5 8.4e-07 5 
+ 8.41e-07 0 9e-07 0 )
VResetQ1H 23 0 pwl (0 5 6e-08 5 6.1e-08 0 9e-07 0 
+ 9.01e-07 5 )
VResetQ1L 24 0 pwl (0 0 6e-08 0 6.1e-08 5 8.06e-06 5 
+ 8.061e-06 0 )
VInput0 14 0 pwl (0 0 6e-08 0 6.1e-08 5 8e-08 5 
+ 8.1e-08 0 1.4e-07 0 1.41e-07 5 1.6e-07 5 
+ 1.61e-07 0 2.2e-07 0 2.21e-07 5 2.4e-07 5 
+ 2.41e-07 0 3e-07 0 3.01e-07 5 3.2e-07 5 
+ 3.21e-07 0 3.8e-07 0 3.81e-07 5 4e-07 5 
+ 4.01e-07 0 4.6e-07 0 4.61e-07 5 4.8e-07 5 
+ 4.81e-07 0 5.4e-07 0 5.41e-07 5 5.6e-07 5 
+ 5.61e-07 0 6.2e-07 0 6.21e-07 5 6.4e-07 5 
+ 6.41e-07 0 7e-07 0 7.01e-07 5 7.2e-07 5 
+ 7.21e-07 0 7.8e-07 0 7.81e-07 5 8e-07 5 
+ 8.01e-07 0 8.6e-07 0 8.61e-07 5 8.8e-07 5 
+ 8.81e-07 0 9.4e-07 0 )
VInput1 507 0 pwl (0 0 8e-08 0 1.6e-07 0 2.4e-07 0 
+ 3.2e-07 0 4e-07 0 4.8e-07 0 5.6e-07 0 
+ 6.4e-07 0 7.2e-07 0 8e-07 0 8.8e-07 0 
+ 9.6e-07 0 )
VVDD 1 0 5
.print TRAN v(19) v(20) v(21) v(22) v(23) v(24) 
+v(14) v(507) v(10) 
*.options limpts=50000 itl5=50000
.TRAN 1e-10 9e-07
.end
