
* test for subcircuit instance parameters, when they refer to each other.
*
* this test also tests precedence rules for subcircuit parameters.   
* The resistor Rinside uses the parameter 'par3'.  It is defined in 3 places.  
* The one with highest priority is on the Xtest line.
*
* This version applies a .step sweep to one of the independent Xtest parameters 
* (par1), to test if the updated value will propagate properly all the way 
* thru to the device Rinside.
*
* This is slightly different than test2, in that the Xtest params don't include a par3.  
* So, the correct par3 is the one on the subckt simple line, but it needs to use the
* par1 and par2 values from the Xtest line.
*
.subckt simple in out 
Rinside in out 88.0
.ends

V1 1 0 1.0
R1 1 2 1.0
Xtest 2 0  simple 

*.step fred list 2.0 3.0 4.0

.dc v1 1.0 1.0 1.0
.print dc v(*) i(*)  {Xtest:Rinside:R}

