A test of the measure duty functionality
*******************************************************************************
*
* a few sources of different types
VS1  1  0  SIN(0 1.0 100HZ 0 0)
VP   2  0  PULSE( 0 100 0ms 1ms 1ms 10ms 20ms )
VS3  3  0  SIN(-0.5 1.0 100HZ 0 0.5)
VS4  4  0  SIN(0.5 -1.0 100HZ 0 0.5)

R1  1  0  100
R2  2  0  100
R3  3  0  100
R4  4  0  100

.TRAN 0  0.1
.PRINT TRAN FORMAT=NOINDEX V(1) V(2) V(3) V(4) V(1,0)

.measure tran dutyAll DUTY V(1) ON=0.75 OFF=0.25
.measure tran duty10All DUTY V(1,0) ON=0.75 OFF=0.25
.measure tran dutyTop Duty V(2) ON=75 OFF=25

* add TO-FROM modifiers
.measure tran sineHalfInterval duty V(1) on=0.75 off=0.25 from=0 to=0.005

* mix in TDs before and after FROM value.
.measure tran sineTDbetween duty V(1) ON=0.75 OFF=0.25 FROM=0 TO=0.025 TD=0.02
.measure tran sineTDbefore duty V(1) ON=0.75 OFF=0.25 FROM=0.02 TO=0.025 TD=0.01

* these tests should return -1 and -100
.measure tran returnNegOne duty V(1) ON=0.75 OFF=0.25 FROM=0.2e-3 TO=0.25e-3 TD=0.5e-3
.measure tran returnNeg100 duty V(1) ON=0.75 OFF=0.25 FROM=0.2e-3 TO=0.25e-3 TD=0.5e-3 default_val=-100

*this test should return 0
.measure tran dutyZero DUTY V(1) ON=2.0 OFF=1.5

* add tests for rise/fall/cross.  V3 and VS4 have a DC offset
* and are damped sinusoids
.measure tran dutyv3fall2 duty v(3) fall=2
.measure tran dutyv4rise1 duty v(4) rise=1
.measure tran dutyv3cross2 duty v(3) cross=2 ON=-0.5 OFF=-1

* test LAST for rise/fall/cross
.measure tran duty3falllast duty v(3) fall=last ON=-0.75 OFF=-1.0
.measure tran duty4riselast duty v(4) rise=last ON=1.0 OFF=0.75
.measure tran duty3crosslast duty v(3) cross=last ON=-0.75 OFF=-1.0
.measure tran duty4crosslast duty v(4) cross=last ON=1.0 OFF=0.75

* test RFC_LEVEL keyword
.measure tran duty1Rise1RFClevel25 duty V(1) RFC_LEVEL=0.25 RISE=1 ON=0.75 OFF=0.5
.measure tran duty1Fall1RFClevel75 duty V(1) RFC_LEVEL=0.75 FALL=1 ON=0.50 OFF=0.25
.measure tran duty1Cross1RFClevel25 duty V(1) RFC_LEVEL=0.25 CROSS=1 ON=0.75 OFF=0.5

*test Failed measures for rise/fall/cross
.measure tran duty3fallfail duty v(3) fall=250
.measure tran duty4risefail duty v(4) rise=250
.measure tran dutyv3crossfail duty v(3) cross=250

.END

