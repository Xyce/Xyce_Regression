Test Circuit for Mutually Coupled, Nonlinear Inductors

VS 1 0 SIN(0 169.7 60HZ)
R1 1 2 1K
R2 3 0 1K
L1 2 0 200
L2 3 0 100
K1 L1 L2 1 nlcore

.model nlcore core level=2 gap=0

.step nlcore:gap 0.25 0.75 0.25
.TRAN 100US 25MS

* Xyce option needed when default is changed to 1 (Backward Euler).
* Also serves as useful test of non-default method.
*.OPTIONS TIMEINT METHOD=2

* Note. The two voltage signals are offset by 0.2 to avoid crossing
* the zero axis.  Axis crossings cause problems for xyce_verify.
.PRINT TRAN I(VS) {V(2)+0.2} {V(3)+0.2} I(L1) I(L2)

*COMP V(2) reltol=0.02
*COMP V(3) reltol=0.02
.END

