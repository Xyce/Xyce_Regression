* simple subcircuit test for issue 24, reference circuit

* sampling 
.sampling useExpr=true
.options SAMPLES numsamples=10
+ outputs={v(2)}
+ sample_type=lhs
+ stdoutput=true
+ seed=1923635719

rtest 0 2 1.0
xtest 1 2 test
v1 0 1 1.0

.subckt test in out
.param fixed_value=aunif(1000,400)
.param other_fixed_value=aunif(1000,400)
r1 in 11 fixed_value
r2 11 out other_fixed_value
.ends

.dc v1 1 1 1
.print dc v(1) v(2) v(xtest:11)

