***************************************************************
* Output both the direct and adjoint sensitivities for
* the case of two objective functions and two parameters.
* This file has both a .PRINT AC and a .PRINT SENS line.
*
* Netlist tests that AC sensitivity output in an unsupported
* format (RAW, PROBE, TOUCHSTONE and TOUCHSTONE2) defaults
* to STD format (.prn file with an Index column)
*
* See SON Bug 1170 for more details.
***************************************************************

* Trivial high-pass filter

R2 c 0 1
R1 b c 1
C1 a b 1u
V1 a 0 DC 0V AC 1

.SENS OBJVARS=b,C PARAM=R1:R,c1:c
.options sensitivity direct=1 adjoint=1 stdoutput=1
.print AC vr(b) vi(b) vp(b) vm(b) R1:R C1:C

.PRINT SENS FILE=ac-sens-formats-default-to-prn.cir.raw FORMAT=RAW
+ vr(b) vi(b) vp(b) vm(b) R1:R R2:R C1:C
.PRINT SENS FILE=ac-sens-formats-default-to-prn.cir.probe FORMAT=PROBE
+ vr(b) vi(b) vp(b) vm(b) R1:R R2:R C1:C
.PRINT SENS FILE=ac-sens-formats-default-to-prn.cir.ts1 FORMAT=TOUCHSTONE
+ vr(b) vi(b) vp(b) vm(b) R1:R R2:R C1:C
.PRINT SENS FILE=ac-sens-formats-default-to-prn.cir.ts2 FORMAT=TOUCHSTONE2
+ vr(b) vi(b) vp(b) vm(b) R1:R R2:R C1:C

.ac dec 5 100Hz 1e6

.end
