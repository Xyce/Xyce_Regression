********************************************************
* Test Embedded Sampling output for .DC for FORMAT =
* STD, CSV and NOINDEX. This covers projection_pce=true
* with one output variable.
*
* See SON Bug 1201 for more details.
********************************************************

*Regression test for simple normal distribution sampling

R2 1 0 3K
R1 1 2 2K
v1 2 0 10V

.dc v1 10 10 1

.print dc v(1)
.PRINT ES

.EMBEDDEDSAMPLING
+ param=R1,R2
+ type=normal,normal
+ means=3K,2K
+ std_deviations=0.1K,0.2K

.options EMBEDDEDSAMPLES numsamples=50
+ projection_pce=true
+ order=3
+ outputs={v(1)}
+ sample_type=lhs
+ stdoutput=true

.PRINT ES PRECISION=6
.PRINT ES PRECISION=6 FORMAT=CSV FILE=es-proj-pce-dc-prn.cir.ES.csv
.PRINT ES PRECISION=6 FORMAT=NOINDEX FILE=es-proj-pce-dc-prn.cir.ES.noindex.prn

.END
