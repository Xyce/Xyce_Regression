* Test syntax for function specified with .param keyword.
* Xyce functions were originally implemented with 
* the .func keyword, but some simulators specify 
* functions as a special type of .param.

* This test exercises multiple function params on the same line, 
* with a conventional parameter in the middle of the list.
* The old .func specification only allowed a single function per line.
* In this case the functions are NOT comma-separated, and the 
* functions have multiple arguments.

.param a=1.0
.param ftest(x,y)={2*x+y}  b=12.0  ftest2(x,y)={3*x+y}

v1 1 0 1.0
r1 1 2 {ftest(2.0,a)*b}
r2 2 0 {ftest2(2.0,a)*b}

.dc v1 1 1 1
.print dc v(1) v(2) {r1:r} {r2:r}

