Test

R1 1 nodename 1k
V1 1 0 1

B1 nodename 0 I={V(nodename)/10}

.DC V1 1 1 1
.PRINT DC V(1) V(nodename)

.END
