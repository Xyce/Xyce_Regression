sram.sp SPICE FILE
.model nenh nmos
+ level = 2
+   vto = 0.59073   kp = 6.12449e-05   gamma = 0.420929
+   phi = 0.7
+
+   cgso = 2.42e-10   cgdo = 2.42e-10
+   rsh = 85   cj = 0.000839
+   mj = 0.796   cjsw = 2.07e-10   mjsw = 0.284
+   tox = 1.75e-08   nsub = 1.50672e+17
+   nss = 3e+10   nfs = 2556.07   tpg = 1
+   xj = 1.73914e-09   ld = 4e-08   uo = 578.411
+   ucrit = 324603   uexp = 0.242015
+   vmax = 128159   neff = 1.22049
+
+   delta = 3.02002
.model penh pmos
+ level = 2
+   vto = -0.59379   kp = 2.35643e-05   gamma = 0.81466
+   phi = 1
+
+   cgso = 2.42e-10   cgdo = 2.42e-10
+   rsh = 154   cj = 0.00054
+   mj = 0.3426   cjsw = 2.15e-10   mjsw = 0.2315
+   tox = 1.75e-08   nsub = 3.36196e+15
+   nss = 3e+10   nfs = 1e+11   tpg = -1
+   xj = 7.41512e-09   ld = 4e-08   uo = 641.842
+   ucrit = 6408.27   uexp = 0.0998923
+   vmax = 132350   neff = 21.4017
+
+   delta = 6.35195
m0 3 5 4 1 penh l=8e-07 w=1e-05 
+ as=1.086e-11 ad=9.39e-12 ps=1.413e-05 pd=1.239e-05 
+ nrs=0.11 nrd=0.09 
m1 4 5 3 1 penh l=8e-07 w=1.08e-05 
+ as=1.015e-11 ad=1.173e-11 ps=1.338e-05 pd=1.526e-05 
+ nrs=0.09 nrd=0.1 
m2 3 5 4 1 penh l=8e-07 w=1e-05 
+ as=1.086e-11 ad=9.39e-12 ps=1.413e-05 pd=1.239e-05 
+ nrs=0.11 nrd=0.09 
m3 4 5 3 1 penh l=8e-07 w=1.1e-05 
+ as=1.033e-11 ad=1.195e-11 ps=1.363e-05 pd=1.554e-05 
+ nrs=0.09 nrd=0.1 
m4 3 5 4 1 penh l=8e-07 w=1e-05 
+ as=1.086e-11 ad=9.39e-12 ps=1.413e-05 pd=1.239e-05 
+ nrs=0.11 nrd=0.09 
m5 3 6 4 0 nenh l=8e-07 w=1e-05 
+ as=7.44e-12 ad=2.334e-11 ps=1.147e-05 pd=1.729e-05 
+ nrs=0.07 nrd=0.23 
m6 4 6 3 0 nenh l=8e-07 w=1.12e-05 
+ as=2.614e-11 ad=8.33e-12 ps=1.936e-05 pd=1.285e-05 
+ nrs=0.21 nrd=0.07 
m7 6 5 0 0 nenh l=8e-07 w=2.2e-06 
+ as=4.04e-12 ad=2.059e-11 ps=5.33e-06 pd=9.94e-06 
+ nrs=0.83 nrd=4.25 
m8 3 6 4 0 nenh l=8e-07 w=1e-05 
+ as=7.44e-12 ad=2.334e-11 ps=1.147e-05 pd=1.729e-05 
+ nrs=0.07 nrd=0.23 
m9 1 5 6 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.889e-11 ps=1.845e-05 pd=2.323e-05 
+ nrs=0.23 nrd=0.3 
m10 4 6 3 0 nenh l=8e-07 w=1.12e-05 
+ as=2.614e-11 ad=8.33e-12 ps=1.936e-05 pd=1.285e-05 
+ nrs=0.21 nrd=0.07 
m11 7 8 6 1 penh l=8e-07 w=2.2e-06 
+ as=7.48e-12 ad=5.19e-12 ps=1.12e-05 pd=6.39e-06 
+ nrs=1.55 nrd=1.07 
m12 9 8 6 1 penh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=5.19e-12 ps=4.4e-06 pd=6.39e-06 
+ nrs=0.5 nrd=1.07 
m13 9 4 6 0 nenh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=4.04e-12 ps=4.4e-06 pd=5.33e-06 
+ nrs=0.5 nrd=0.83 
m14 7 4 6 0 nenh l=8e-07 w=2.2e-06 
+ as=7.48e-12 ad=4.04e-12 ps=1.12e-05 pd=5.33e-06 
+ nrs=1.55 nrd=0.83 
m15 5 9 1 1 penh l=8e-07 w=8e-06 
+ as=1.76e-11 ad=1.465e-11 ps=2.04e-05 pd=1.845e-05 
+ nrs=0.28 nrd=0.23 
m16 3 6 4 0 nenh l=8e-07 w=1e-05 
+ as=7.44e-12 ad=2.334e-11 ps=1.147e-05 pd=1.729e-05 
+ nrs=0.07 nrd=0.23 
m17 0 5 3 0 nenh l=8e-07 w=1.14e-05 
+ as=1.067e-10 ad=8.48e-12 ps=5.151e-05 pd=1.308e-05 
+ nrs=0.82 nrd=0.07 
m18 10 11 9 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=2.42e-12 ps=6.3e-06 pd=4.4e-06 
+ nrs=1 nrd=0.5 
m19 4 13 12 1 penh l=8e-07 w=1e-05 
+ as=9.39e-12 ad=1.112e-11 ps=1.239e-05 pd=1.419e-05 
+ nrs=0.09 nrd=0.11 
m20 12 13 0 0 nenh l=8e-07 w=1.14e-05 
+ as=8.48e-12 ad=1.067e-10 ps=1.308e-05 pd=5.151e-05 
+ nrs=0.07 nrd=0.82 
m21 12 13 4 1 penh l=8e-07 w=1.1e-05 
+ as=1.223e-11 ad=1.033e-11 ps=1.56e-05 pd=1.363e-05 
+ nrs=0.1 nrd=0.09 
m22 4 13 12 1 penh l=8e-07 w=1e-05 
+ as=9.39e-12 ad=1.112e-11 ps=1.239e-05 pd=1.419e-05 
+ nrs=0.09 nrd=0.11 
m23 12 13 4 1 penh l=8e-07 w=1.06e-05 
+ as=1.178e-11 ad=9.96e-12 ps=1.504e-05 pd=1.313e-05 
+ nrs=0.1 nrd=0.09 
m24 4 13 12 1 penh l=8e-07 w=1e-05 
+ as=9.39e-12 ad=1.112e-11 ps=1.239e-05 pd=1.419e-05 
+ nrs=0.09 nrd=0.11 
m25 4 14 12 0 nenh l=8e-07 w=1e-05 
+ as=2.334e-11 ad=7.44e-12 ps=1.729e-05 pd=1.147e-05 
+ nrs=0.23 nrd=0.07 
m26 1 15 13 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.76e-11 ps=1.845e-05 pd=2.04e-05 
+ nrs=0.23 nrd=0.28 
m27 12 14 4 0 nenh l=8e-07 w=1.12e-05 
+ as=8.33e-12 ad=2.614e-11 ps=1.285e-05 pd=1.936e-05 
+ nrs=0.07 nrd=0.21 
m28 4 14 12 0 nenh l=8e-07 w=1e-05 
+ as=2.334e-11 ad=7.44e-12 ps=1.729e-05 pd=1.147e-05 
+ nrs=0.23 nrd=0.07 
m29 14 13 1 1 penh l=8e-07 w=8e-06 
+ as=1.848e-11 ad=1.465e-11 ps=2.323e-05 pd=1.845e-05 
+ nrs=0.29 nrd=0.23 
m30 15 11 16 1 penh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=4.84e-12 ps=4.4e-06 pd=6.3e-06 
+ nrs=0.5 nrd=1 
m31 10 17 9 0 nenh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=2.42e-12 ps=8.8e-06 pd=4.4e-06 
+ nrs=1 nrd=0.5 
m32 0 9 5 0 nenh l=8e-07 w=9e-06 
+ as=8.424e-11 ad=1.248e-11 ps=4.066e-05 pd=1.64e-05 
+ nrs=1.04 nrd=0.15 
m33 16 18 0 0 nenh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=2.059e-11 ps=8.8e-06 pd=9.94e-06 
+ nrs=1 nrd=4.25 
m34 1 18 16 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.76e-11 ps=1.845e-05 pd=2.29e-05 
+ nrs=0.23 nrd=0.28 
m35 18 7 0 0 nenh l=8e-07 w=8e-06 
+ as=1.508e-11 ad=7.488e-11 ps=2.4e-05 pd=3.615e-05 
+ nrs=0.24 nrd=1.17 
m36 18 7 1 1 penh l=8e-07 w=8e-06 
+ as=1.76e-11 ad=1.465e-11 ps=2.04e-05 pd=1.845e-05 
+ nrs=0.28 nrd=0.23 
m37 15 17 16 0 nenh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=4.84e-12 ps=4.4e-06 pd=8.8e-06 
+ nrs=0.5 nrd=1 
m38 19 20 0 0 nenh l=8e-07 w=8e-06 
+ as=1.772e-11 ad=7.488e-11 ps=2.4e-05 pd=3.615e-05 
+ nrs=0.28 nrd=1.17 
m39 1 20 19 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.76e-11 ps=1.845e-05 pd=2.04e-05 
+ nrs=0.23 nrd=0.28 
m40 14 8 20 1 penh l=8e-07 w=2.2e-06 
+ as=5.08e-12 ad=7.48e-12 ps=6.39e-06 pd=1.12e-05 
+ nrs=1.05 nrd=1.55 
m41 14 8 15 1 penh l=8e-07 w=2.2e-06 
+ as=5.08e-12 ad=2.42e-12 ps=6.39e-06 pd=4.4e-06 
+ nrs=1.05 nrd=0.5 
m42 14 4 15 0 nenh l=8e-07 w=2.2e-06 
+ as=3.68e-12 ad=2.42e-12 ps=5.2e-06 pd=4.4e-06 
+ nrs=0.76 nrd=0.5 
m43 14 4 20 0 nenh l=8e-07 w=2.2e-06 
+ as=3.68e-12 ad=1.408e-11 ps=5.2e-06 pd=1.72e-05 
+ nrs=0.76 nrd=2.91 
m44 12 14 4 0 nenh l=8e-07 w=1.12e-05 
+ as=8.33e-12 ad=2.614e-11 ps=1.285e-05 pd=1.936e-05 
+ nrs=0.07 nrd=0.21 
m45 4 14 12 0 nenh l=8e-07 w=1e-05 
+ as=2.334e-11 ad=7.44e-12 ps=1.729e-05 pd=1.147e-05 
+ nrs=0.23 nrd=0.07 
m46 0 13 14 0 nenh l=8e-07 w=2.2e-06 
+ as=2.059e-11 ad=3.68e-12 ps=9.94e-06 pd=5.2e-06 
+ nrs=4.25 nrd=0.76 
m47 0 15 13 0 nenh l=8e-07 w=9e-06 
+ as=8.424e-11 ad=1.224e-11 ps=4.066e-05 pd=1.64e-05 
+ nrs=1.04 nrd=0.15 
m48 21 19 1 1 penh l=8e-07 w=8e-06 
+ as=1.76e-11 ad=1.465e-11 ps=2.04e-05 pd=1.845e-05 
+ nrs=0.28 nrd=0.23 
m49 0 19 21 0 nenh l=8e-07 w=2.2e-06 
+ as=2.059e-11 ad=4.84e-12 ps=9.94e-06 pd=8.8e-06 
+ nrs=4.25 nrd=1 
m50 22 23 4 1 penh l=8e-07 w=1e-05 
+ as=1.086e-11 ad=9.39e-12 ps=1.413e-05 pd=1.239e-05 
+ nrs=0.11 nrd=0.09 
m51 4 23 22 1 penh l=8e-07 w=1.08e-05 
+ as=1.015e-11 ad=1.173e-11 ps=1.338e-05 pd=1.526e-05 
+ nrs=0.09 nrd=0.1 
m52 22 23 4 1 penh l=8e-07 w=1e-05 
+ as=1.086e-11 ad=9.39e-12 ps=1.413e-05 pd=1.239e-05 
+ nrs=0.11 nrd=0.09 
m53 4 23 22 1 penh l=8e-07 w=1.1e-05 
+ as=1.033e-11 ad=1.195e-11 ps=1.363e-05 pd=1.554e-05 
+ nrs=0.09 nrd=0.1 
m54 22 23 4 1 penh l=8e-07 w=1e-05 
+ as=1.086e-11 ad=9.39e-12 ps=1.413e-05 pd=1.239e-05 
+ nrs=0.11 nrd=0.09 
m55 22 24 4 0 nenh l=8e-07 w=1e-05 
+ as=7.44e-12 ad=2.334e-11 ps=1.147e-05 pd=1.729e-05 
+ nrs=0.07 nrd=0.23 
m56 4 24 22 0 nenh l=8e-07 w=1.12e-05 
+ as=2.614e-11 ad=8.33e-12 ps=1.936e-05 pd=1.285e-05 
+ nrs=0.21 nrd=0.07 
m57 24 23 0 0 nenh l=8e-07 w=2.2e-06 
+ as=4.04e-12 ad=2.059e-11 ps=5.33e-06 pd=9.94e-06 
+ nrs=0.83 nrd=4.25 
m58 22 24 4 0 nenh l=8e-07 w=1e-05 
+ as=7.44e-12 ad=2.334e-11 ps=1.147e-05 pd=1.729e-05 
+ nrs=0.07 nrd=0.23 
m59 1 23 24 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.889e-11 ps=1.845e-05 pd=2.323e-05 
+ nrs=0.23 nrd=0.3 
m60 4 24 22 0 nenh l=8e-07 w=1.12e-05 
+ as=2.614e-11 ad=8.33e-12 ps=1.936e-05 pd=1.285e-05 
+ nrs=0.21 nrd=0.07 
m61 25 8 24 1 penh l=8e-07 w=2.2e-06 
+ as=7.48e-12 ad=5.19e-12 ps=1.12e-05 pd=6.39e-06 
+ nrs=1.55 nrd=1.07 
m62 26 8 24 1 penh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=5.19e-12 ps=4.4e-06 pd=6.39e-06 
+ nrs=0.5 nrd=1.07 
m63 26 4 24 0 nenh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=4.04e-12 ps=4.4e-06 pd=5.33e-06 
+ nrs=0.5 nrd=0.83 
m64 25 4 24 0 nenh l=8e-07 w=2.2e-06 
+ as=7.48e-12 ad=4.04e-12 ps=1.12e-05 pd=5.33e-06 
+ nrs=1.55 nrd=0.83 
m65 23 26 1 1 penh l=8e-07 w=8e-06 
+ as=1.76e-11 ad=1.465e-11 ps=2.04e-05 pd=1.845e-05 
+ nrs=0.28 nrd=0.23 
m66 22 24 4 0 nenh l=8e-07 w=1e-05 
+ as=7.44e-12 ad=2.334e-11 ps=1.147e-05 pd=1.729e-05 
+ nrs=0.07 nrd=0.23 
m67 0 23 22 0 nenh l=8e-07 w=1.14e-05 
+ as=1.067e-10 ad=8.48e-12 ps=5.151e-05 pd=1.308e-05 
+ nrs=0.82 nrd=0.07 
m68 27 11 26 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=2.42e-12 ps=6.3e-06 pd=4.4e-06 
+ nrs=1 nrd=0.5 
m69 4 29 28 1 penh l=8e-07 w=1e-05 
+ as=9.39e-12 ad=1.112e-11 ps=1.239e-05 pd=1.419e-05 
+ nrs=0.09 nrd=0.11 
m70 28 29 0 0 nenh l=8e-07 w=1.14e-05 
+ as=8.48e-12 ad=1.067e-10 ps=1.308e-05 pd=5.151e-05 
+ nrs=0.07 nrd=0.82 
m71 28 29 4 1 penh l=8e-07 w=1.1e-05 
+ as=1.223e-11 ad=1.033e-11 ps=1.56e-05 pd=1.363e-05 
+ nrs=0.1 nrd=0.09 
m72 4 29 28 1 penh l=8e-07 w=1e-05 
+ as=9.39e-12 ad=1.112e-11 ps=1.239e-05 pd=1.419e-05 
+ nrs=0.09 nrd=0.11 
m73 28 29 4 1 penh l=8e-07 w=1.06e-05 
+ as=1.178e-11 ad=9.96e-12 ps=1.504e-05 pd=1.313e-05 
+ nrs=0.1 nrd=0.09 
m74 4 29 28 1 penh l=8e-07 w=1e-05 
+ as=9.39e-12 ad=1.112e-11 ps=1.239e-05 pd=1.419e-05 
+ nrs=0.09 nrd=0.11 
m75 4 30 28 0 nenh l=8e-07 w=1e-05 
+ as=2.334e-11 ad=7.44e-12 ps=1.729e-05 pd=1.147e-05 
+ nrs=0.23 nrd=0.07 
m76 1 31 29 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.76e-11 ps=1.845e-05 pd=2.04e-05 
+ nrs=0.23 nrd=0.28 
m77 28 30 4 0 nenh l=8e-07 w=1.12e-05 
+ as=8.33e-12 ad=2.614e-11 ps=1.285e-05 pd=1.936e-05 
+ nrs=0.07 nrd=0.21 
m78 4 30 28 0 nenh l=8e-07 w=1e-05 
+ as=2.334e-11 ad=7.44e-12 ps=1.729e-05 pd=1.147e-05 
+ nrs=0.23 nrd=0.07 
m79 30 29 1 1 penh l=8e-07 w=8e-06 
+ as=1.848e-11 ad=1.465e-11 ps=2.323e-05 pd=1.845e-05 
+ nrs=0.29 nrd=0.23 
m80 31 11 32 1 penh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=4.84e-12 ps=4.4e-06 pd=6.3e-06 
+ nrs=0.5 nrd=1 
m81 27 17 26 0 nenh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=2.42e-12 ps=8.8e-06 pd=4.4e-06 
+ nrs=1 nrd=0.5 
m82 0 26 23 0 nenh l=8e-07 w=9e-06 
+ as=8.424e-11 ad=1.248e-11 ps=4.066e-05 pd=1.64e-05 
+ nrs=1.04 nrd=0.15 
m83 32 33 0 0 nenh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=2.059e-11 ps=8.8e-06 pd=9.94e-06 
+ nrs=1 nrd=4.25 
m84 1 33 32 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.76e-11 ps=1.845e-05 pd=2.29e-05 
+ nrs=0.23 nrd=0.28 
m85 33 25 0 0 nenh l=8e-07 w=8e-06 
+ as=1.508e-11 ad=7.488e-11 ps=2.4e-05 pd=3.615e-05 
+ nrs=0.24 nrd=1.17 
m86 33 25 1 1 penh l=8e-07 w=8e-06 
+ as=1.76e-11 ad=1.465e-11 ps=2.04e-05 pd=1.845e-05 
+ nrs=0.28 nrd=0.23 
m87 31 17 32 0 nenh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=4.84e-12 ps=4.4e-06 pd=8.8e-06 
+ nrs=0.5 nrd=1 
m88 34 35 0 0 nenh l=8e-07 w=8e-06 
+ as=1.772e-11 ad=7.488e-11 ps=2.4e-05 pd=3.615e-05 
+ nrs=0.28 nrd=1.17 
m89 1 35 34 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.76e-11 ps=1.845e-05 pd=2.04e-05 
+ nrs=0.23 nrd=0.28 
m90 30 8 35 1 penh l=8e-07 w=2.2e-06 
+ as=5.08e-12 ad=7.48e-12 ps=6.39e-06 pd=1.12e-05 
+ nrs=1.05 nrd=1.55 
m91 30 8 31 1 penh l=8e-07 w=2.2e-06 
+ as=5.08e-12 ad=2.42e-12 ps=6.39e-06 pd=4.4e-06 
+ nrs=1.05 nrd=0.5 
m92 30 4 31 0 nenh l=8e-07 w=2.2e-06 
+ as=3.68e-12 ad=2.42e-12 ps=5.2e-06 pd=4.4e-06 
+ nrs=0.76 nrd=0.5 
m93 30 4 35 0 nenh l=8e-07 w=2.2e-06 
+ as=3.68e-12 ad=1.408e-11 ps=5.2e-06 pd=1.72e-05 
+ nrs=0.76 nrd=2.91 
m94 28 30 4 0 nenh l=8e-07 w=1.12e-05 
+ as=8.33e-12 ad=2.614e-11 ps=1.285e-05 pd=1.936e-05 
+ nrs=0.07 nrd=0.21 
m95 4 30 28 0 nenh l=8e-07 w=1e-05 
+ as=2.334e-11 ad=7.44e-12 ps=1.729e-05 pd=1.147e-05 
+ nrs=0.23 nrd=0.07 
m96 0 29 30 0 nenh l=8e-07 w=2.2e-06 
+ as=2.059e-11 ad=3.68e-12 ps=9.94e-06 pd=5.2e-06 
+ nrs=4.25 nrd=0.76 
m97 0 31 29 0 nenh l=8e-07 w=9e-06 
+ as=8.424e-11 ad=1.224e-11 ps=4.066e-05 pd=1.64e-05 
+ nrs=1.04 nrd=0.15 
m98 10 34 1 1 penh l=8e-07 w=8e-06 
+ as=1.76e-11 ad=1.465e-11 ps=2.29e-05 pd=1.845e-05 
+ nrs=0.28 nrd=0.23 
m99 0 34 10 0 nenh l=8e-07 w=2.2e-06 
+ as=2.059e-11 ad=4.84e-12 ps=9.94e-06 pd=8.8e-06 
+ nrs=4.25 nrd=1 
m100 36 37 4 1 penh l=8e-07 w=1e-05 
+ as=1.086e-11 ad=9.39e-12 ps=1.413e-05 pd=1.239e-05 
+ nrs=0.11 nrd=0.09 
m101 4 37 36 1 penh l=8e-07 w=1.08e-05 
+ as=1.015e-11 ad=1.173e-11 ps=1.338e-05 pd=1.526e-05 
+ nrs=0.09 nrd=0.1 
m102 36 37 4 1 penh l=8e-07 w=1e-05 
+ as=1.086e-11 ad=9.39e-12 ps=1.413e-05 pd=1.239e-05 
+ nrs=0.11 nrd=0.09 
m103 4 37 36 1 penh l=8e-07 w=1.1e-05 
+ as=1.033e-11 ad=1.195e-11 ps=1.363e-05 pd=1.554e-05 
+ nrs=0.09 nrd=0.1 
m104 36 37 4 1 penh l=8e-07 w=1e-05 
+ as=1.086e-11 ad=9.39e-12 ps=1.413e-05 pd=1.239e-05 
+ nrs=0.11 nrd=0.09 
m105 36 38 4 0 nenh l=8e-07 w=1e-05 
+ as=7.44e-12 ad=2.334e-11 ps=1.147e-05 pd=1.729e-05 
+ nrs=0.07 nrd=0.23 
m106 4 38 36 0 nenh l=8e-07 w=1.12e-05 
+ as=2.614e-11 ad=8.33e-12 ps=1.936e-05 pd=1.285e-05 
+ nrs=0.21 nrd=0.07 
m107 38 37 0 0 nenh l=8e-07 w=2.2e-06 
+ as=4.04e-12 ad=2.059e-11 ps=5.33e-06 pd=9.94e-06 
+ nrs=0.83 nrd=4.25 
m108 36 38 4 0 nenh l=8e-07 w=1e-05 
+ as=7.44e-12 ad=2.334e-11 ps=1.147e-05 pd=1.729e-05 
+ nrs=0.07 nrd=0.23 
m109 1 37 38 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.889e-11 ps=1.845e-05 pd=2.323e-05 
+ nrs=0.23 nrd=0.3 
m110 4 38 36 0 nenh l=8e-07 w=1.12e-05 
+ as=2.614e-11 ad=8.33e-12 ps=1.936e-05 pd=1.285e-05 
+ nrs=0.21 nrd=0.07 
m111 39 8 38 1 penh l=8e-07 w=2.2e-06 
+ as=7.48e-12 ad=5.19e-12 ps=1.12e-05 pd=6.39e-06 
+ nrs=1.55 nrd=1.07 
m112 40 8 38 1 penh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=5.19e-12 ps=4.4e-06 pd=6.39e-06 
+ nrs=0.5 nrd=1.07 
m113 40 4 38 0 nenh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=4.04e-12 ps=4.4e-06 pd=5.33e-06 
+ nrs=0.5 nrd=0.83 
m114 39 4 38 0 nenh l=8e-07 w=2.2e-06 
+ as=7.48e-12 ad=4.04e-12 ps=1.12e-05 pd=5.33e-06 
+ nrs=1.55 nrd=0.83 
m115 37 40 1 1 penh l=8e-07 w=8e-06 
+ as=1.76e-11 ad=1.465e-11 ps=2.04e-05 pd=1.845e-05 
+ nrs=0.28 nrd=0.23 
m116 36 38 4 0 nenh l=8e-07 w=1e-05 
+ as=7.44e-12 ad=2.334e-11 ps=1.147e-05 pd=1.729e-05 
+ nrs=0.07 nrd=0.23 
m117 0 37 36 0 nenh l=8e-07 w=1.14e-05 
+ as=1.067e-10 ad=8.48e-12 ps=5.151e-05 pd=1.308e-05 
+ nrs=0.82 nrd=0.07 
m118 41 11 40 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=2.42e-12 ps=6.3e-06 pd=4.4e-06 
+ nrs=1 nrd=0.5 
m119 4 43 42 1 penh l=8e-07 w=1e-05 
+ as=9.39e-12 ad=1.112e-11 ps=1.239e-05 pd=1.419e-05 
+ nrs=0.09 nrd=0.11 
m120 42 43 0 0 nenh l=8e-07 w=1.14e-05 
+ as=8.48e-12 ad=1.067e-10 ps=1.308e-05 pd=5.151e-05 
+ nrs=0.07 nrd=0.82 
m121 42 43 4 1 penh l=8e-07 w=1.1e-05 
+ as=1.223e-11 ad=1.033e-11 ps=1.56e-05 pd=1.363e-05 
+ nrs=0.1 nrd=0.09 
m122 4 43 42 1 penh l=8e-07 w=1e-05 
+ as=9.39e-12 ad=1.112e-11 ps=1.239e-05 pd=1.419e-05 
+ nrs=0.09 nrd=0.11 
m123 42 43 4 1 penh l=8e-07 w=1.06e-05 
+ as=1.178e-11 ad=9.96e-12 ps=1.504e-05 pd=1.313e-05 
+ nrs=0.1 nrd=0.09 
m124 4 43 42 1 penh l=8e-07 w=1e-05 
+ as=9.39e-12 ad=1.112e-11 ps=1.239e-05 pd=1.419e-05 
+ nrs=0.09 nrd=0.11 
m125 4 44 42 0 nenh l=8e-07 w=1e-05 
+ as=2.334e-11 ad=7.44e-12 ps=1.729e-05 pd=1.147e-05 
+ nrs=0.23 nrd=0.07 
m126 1 45 43 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.76e-11 ps=1.845e-05 pd=2.04e-05 
+ nrs=0.23 nrd=0.28 
m127 42 44 4 0 nenh l=8e-07 w=1.12e-05 
+ as=8.33e-12 ad=2.614e-11 ps=1.285e-05 pd=1.936e-05 
+ nrs=0.07 nrd=0.21 
m128 4 44 42 0 nenh l=8e-07 w=1e-05 
+ as=2.334e-11 ad=7.44e-12 ps=1.729e-05 pd=1.147e-05 
+ nrs=0.23 nrd=0.07 
m129 44 43 1 1 penh l=8e-07 w=8e-06 
+ as=1.848e-11 ad=1.465e-11 ps=2.323e-05 pd=1.845e-05 
+ nrs=0.29 nrd=0.23 
m130 45 11 46 1 penh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=4.84e-12 ps=4.4e-06 pd=6.3e-06 
+ nrs=0.5 nrd=1 
m131 41 17 40 0 nenh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=2.42e-12 ps=8.8e-06 pd=4.4e-06 
+ nrs=1 nrd=0.5 
m132 0 40 37 0 nenh l=8e-07 w=9e-06 
+ as=8.424e-11 ad=1.248e-11 ps=4.066e-05 pd=1.64e-05 
+ nrs=1.04 nrd=0.15 
m133 46 47 0 0 nenh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=2.059e-11 ps=8.8e-06 pd=9.94e-06 
+ nrs=1 nrd=4.25 
m134 1 47 46 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.76e-11 ps=1.845e-05 pd=2.29e-05 
+ nrs=0.23 nrd=0.28 
m135 47 39 0 0 nenh l=8e-07 w=8e-06 
+ as=1.508e-11 ad=7.488e-11 ps=2.4e-05 pd=3.615e-05 
+ nrs=0.24 nrd=1.17 
m136 47 39 1 1 penh l=8e-07 w=8e-06 
+ as=1.76e-11 ad=1.465e-11 ps=2.04e-05 pd=1.845e-05 
+ nrs=0.28 nrd=0.23 
m137 45 17 46 0 nenh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=4.84e-12 ps=4.4e-06 pd=8.8e-06 
+ nrs=0.5 nrd=1 
m138 48 49 0 0 nenh l=8e-07 w=8e-06 
+ as=1.772e-11 ad=7.488e-11 ps=2.4e-05 pd=3.615e-05 
+ nrs=0.28 nrd=1.17 
m139 1 49 48 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.76e-11 ps=1.845e-05 pd=2.04e-05 
+ nrs=0.23 nrd=0.28 
m140 44 8 49 1 penh l=8e-07 w=2.2e-06 
+ as=5.08e-12 ad=7.48e-12 ps=6.39e-06 pd=1.12e-05 
+ nrs=1.05 nrd=1.55 
m141 44 8 45 1 penh l=8e-07 w=2.2e-06 
+ as=5.08e-12 ad=2.42e-12 ps=6.39e-06 pd=4.4e-06 
+ nrs=1.05 nrd=0.5 
m142 44 4 45 0 nenh l=8e-07 w=2.2e-06 
+ as=3.68e-12 ad=2.42e-12 ps=5.2e-06 pd=4.4e-06 
+ nrs=0.76 nrd=0.5 
m143 44 4 49 0 nenh l=8e-07 w=2.2e-06 
+ as=3.68e-12 ad=1.408e-11 ps=5.2e-06 pd=1.72e-05 
+ nrs=0.76 nrd=2.91 
m144 42 44 4 0 nenh l=8e-07 w=1.12e-05 
+ as=8.33e-12 ad=2.614e-11 ps=1.285e-05 pd=1.936e-05 
+ nrs=0.07 nrd=0.21 
m145 4 44 42 0 nenh l=8e-07 w=1e-05 
+ as=2.334e-11 ad=7.44e-12 ps=1.729e-05 pd=1.147e-05 
+ nrs=0.23 nrd=0.07 
m146 0 43 44 0 nenh l=8e-07 w=2.2e-06 
+ as=2.059e-11 ad=3.68e-12 ps=9.94e-06 pd=5.2e-06 
+ nrs=4.25 nrd=0.76 
m147 0 45 43 0 nenh l=8e-07 w=9e-06 
+ as=8.424e-11 ad=1.224e-11 ps=4.066e-05 pd=1.64e-05 
+ nrs=1.04 nrd=0.15 
m148 27 48 1 1 penh l=8e-07 w=8e-06 
+ as=1.76e-11 ad=1.465e-11 ps=2.29e-05 pd=1.845e-05 
+ nrs=0.28 nrd=0.23 
m149 0 48 27 0 nenh l=8e-07 w=2.2e-06 
+ as=2.059e-11 ad=4.84e-12 ps=9.94e-06 pd=8.8e-06 
+ nrs=4.25 nrd=1 
m150 50 51 4 1 penh l=8e-07 w=1e-05 
+ as=1.086e-11 ad=9.39e-12 ps=1.413e-05 pd=1.239e-05 
+ nrs=0.11 nrd=0.09 
m151 4 51 50 1 penh l=8e-07 w=1.08e-05 
+ as=1.015e-11 ad=1.173e-11 ps=1.338e-05 pd=1.526e-05 
+ nrs=0.09 nrd=0.1 
m152 50 51 4 1 penh l=8e-07 w=1e-05 
+ as=1.086e-11 ad=9.39e-12 ps=1.413e-05 pd=1.239e-05 
+ nrs=0.11 nrd=0.09 
m153 4 51 50 1 penh l=8e-07 w=1.1e-05 
+ as=1.033e-11 ad=1.195e-11 ps=1.363e-05 pd=1.554e-05 
+ nrs=0.09 nrd=0.1 
m154 50 51 4 1 penh l=8e-07 w=1e-05 
+ as=1.086e-11 ad=9.39e-12 ps=1.413e-05 pd=1.239e-05 
+ nrs=0.11 nrd=0.09 
m155 50 52 4 0 nenh l=8e-07 w=1e-05 
+ as=7.44e-12 ad=2.334e-11 ps=1.147e-05 pd=1.729e-05 
+ nrs=0.07 nrd=0.23 
m156 4 52 50 0 nenh l=8e-07 w=1.12e-05 
+ as=2.614e-11 ad=8.33e-12 ps=1.936e-05 pd=1.285e-05 
+ nrs=0.21 nrd=0.07 
m157 52 51 0 0 nenh l=8e-07 w=2.2e-06 
+ as=4.04e-12 ad=2.059e-11 ps=5.33e-06 pd=9.94e-06 
+ nrs=0.83 nrd=4.25 
m158 50 52 4 0 nenh l=8e-07 w=1e-05 
+ as=7.44e-12 ad=2.334e-11 ps=1.147e-05 pd=1.729e-05 
+ nrs=0.07 nrd=0.23 
m159 1 51 52 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.889e-11 ps=1.845e-05 pd=2.323e-05 
+ nrs=0.23 nrd=0.3 
m160 4 52 50 0 nenh l=8e-07 w=1.12e-05 
+ as=2.614e-11 ad=8.33e-12 ps=1.936e-05 pd=1.285e-05 
+ nrs=0.21 nrd=0.07 
m161 53 8 52 1 penh l=8e-07 w=2.2e-06 
+ as=7.48e-12 ad=5.19e-12 ps=1.12e-05 pd=6.39e-06 
+ nrs=1.55 nrd=1.07 
m162 54 8 52 1 penh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=5.19e-12 ps=4.4e-06 pd=6.39e-06 
+ nrs=0.5 nrd=1.07 
m163 54 4 52 0 nenh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=4.04e-12 ps=4.4e-06 pd=5.33e-06 
+ nrs=0.5 nrd=0.83 
m164 53 4 52 0 nenh l=8e-07 w=2.2e-06 
+ as=7.48e-12 ad=4.04e-12 ps=1.12e-05 pd=5.33e-06 
+ nrs=1.55 nrd=0.83 
m165 51 54 1 1 penh l=8e-07 w=8e-06 
+ as=1.76e-11 ad=1.465e-11 ps=2.04e-05 pd=1.845e-05 
+ nrs=0.28 nrd=0.23 
m166 50 52 4 0 nenh l=8e-07 w=1e-05 
+ as=7.44e-12 ad=2.334e-11 ps=1.147e-05 pd=1.729e-05 
+ nrs=0.07 nrd=0.23 
m167 0 51 50 0 nenh l=8e-07 w=1.14e-05 
+ as=1.067e-10 ad=8.48e-12 ps=5.151e-05 pd=1.308e-05 
+ nrs=0.82 nrd=0.07 
m168 55 11 54 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=2.42e-12 ps=7.52e-06 pd=4.4e-06 
+ nrs=1 nrd=0.5 
m169 4 57 56 1 penh l=8e-07 w=1e-05 
+ as=9.39e-12 ad=1.112e-11 ps=1.239e-05 pd=1.419e-05 
+ nrs=0.09 nrd=0.11 
m170 56 57 0 0 nenh l=8e-07 w=1.14e-05 
+ as=8.48e-12 ad=1.067e-10 ps=1.308e-05 pd=5.151e-05 
+ nrs=0.07 nrd=0.82 
m171 56 57 4 1 penh l=8e-07 w=1.1e-05 
+ as=1.223e-11 ad=1.033e-11 ps=1.56e-05 pd=1.363e-05 
+ nrs=0.1 nrd=0.09 
m172 4 57 56 1 penh l=8e-07 w=1e-05 
+ as=9.39e-12 ad=1.112e-11 ps=1.239e-05 pd=1.419e-05 
+ nrs=0.09 nrd=0.11 
m173 56 57 4 1 penh l=8e-07 w=1.06e-05 
+ as=1.178e-11 ad=9.96e-12 ps=1.504e-05 pd=1.313e-05 
+ nrs=0.1 nrd=0.09 
m174 4 57 56 1 penh l=8e-07 w=1e-05 
+ as=9.39e-12 ad=1.112e-11 ps=1.239e-05 pd=1.419e-05 
+ nrs=0.09 nrd=0.11 
m175 4 58 56 0 nenh l=8e-07 w=1e-05 
+ as=2.334e-11 ad=7.44e-12 ps=1.729e-05 pd=1.147e-05 
+ nrs=0.23 nrd=0.07 
m176 1 59 57 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.76e-11 ps=1.845e-05 pd=2.04e-05 
+ nrs=0.23 nrd=0.28 
m177 56 58 4 0 nenh l=8e-07 w=1.12e-05 
+ as=8.33e-12 ad=2.614e-11 ps=1.285e-05 pd=1.936e-05 
+ nrs=0.07 nrd=0.21 
m178 4 58 56 0 nenh l=8e-07 w=1e-05 
+ as=2.334e-11 ad=7.44e-12 ps=1.729e-05 pd=1.147e-05 
+ nrs=0.23 nrd=0.07 
m179 58 57 1 1 penh l=8e-07 w=8e-06 
+ as=1.848e-11 ad=1.465e-11 ps=2.323e-05 pd=1.845e-05 
+ nrs=0.29 nrd=0.23 
m180 59 11 60 1 penh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=4.84e-12 ps=4.4e-06 pd=6.3e-06 
+ nrs=0.5 nrd=1 
m181 55 17 54 0 nenh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=2.42e-12 ps=7.52e-06 pd=4.4e-06 
+ nrs=1 nrd=0.5 
m182 0 54 51 0 nenh l=8e-07 w=9e-06 
+ as=8.424e-11 ad=1.248e-11 ps=4.066e-05 pd=1.64e-05 
+ nrs=1.04 nrd=0.15 
m183 60 61 0 0 nenh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=2.059e-11 ps=8.8e-06 pd=9.94e-06 
+ nrs=1 nrd=4.25 
m184 1 61 60 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.76e-11 ps=1.845e-05 pd=2.29e-05 
+ nrs=0.23 nrd=0.28 
m185 61 53 0 0 nenh l=8e-07 w=8e-06 
+ as=1.508e-11 ad=7.488e-11 ps=2.4e-05 pd=3.615e-05 
+ nrs=0.24 nrd=1.17 
m186 61 53 1 1 penh l=8e-07 w=8e-06 
+ as=1.76e-11 ad=1.465e-11 ps=2.04e-05 pd=1.845e-05 
+ nrs=0.28 nrd=0.23 
m187 59 17 60 0 nenh l=8e-07 w=2.2e-06 
+ as=2.42e-12 ad=4.84e-12 ps=4.4e-06 pd=8.8e-06 
+ nrs=0.5 nrd=1 
m188 62 63 0 0 nenh l=8e-07 w=8e-06 
+ as=1.772e-11 ad=7.488e-11 ps=2.4e-05 pd=3.615e-05 
+ nrs=0.28 nrd=1.17 
m189 1 63 62 1 penh l=8e-07 w=8e-06 
+ as=1.465e-11 ad=1.76e-11 ps=1.845e-05 pd=2.04e-05 
+ nrs=0.23 nrd=0.28 
m190 58 8 63 1 penh l=8e-07 w=2.2e-06 
+ as=5.08e-12 ad=7.48e-12 ps=6.39e-06 pd=1.12e-05 
+ nrs=1.05 nrd=1.55 
m191 58 8 59 1 penh l=8e-07 w=2.2e-06 
+ as=5.08e-12 ad=2.42e-12 ps=6.39e-06 pd=4.4e-06 
+ nrs=1.05 nrd=0.5 
m192 58 4 59 0 nenh l=8e-07 w=2.2e-06 
+ as=3.68e-12 ad=2.42e-12 ps=5.2e-06 pd=4.4e-06 
+ nrs=0.76 nrd=0.5 
m193 58 4 63 0 nenh l=8e-07 w=2.2e-06 
+ as=3.68e-12 ad=1.408e-11 ps=5.2e-06 pd=1.72e-05 
+ nrs=0.76 nrd=2.91 
m194 56 58 4 0 nenh l=8e-07 w=1.12e-05 
+ as=8.33e-12 ad=2.614e-11 ps=1.285e-05 pd=1.936e-05 
+ nrs=0.07 nrd=0.21 
m195 4 58 56 0 nenh l=8e-07 w=1e-05 
+ as=2.334e-11 ad=7.44e-12 ps=1.729e-05 pd=1.147e-05 
+ nrs=0.23 nrd=0.07 
m196 0 57 58 0 nenh l=8e-07 w=2.2e-06 
+ as=2.059e-11 ad=3.68e-12 ps=9.94e-06 pd=5.2e-06 
+ nrs=4.25 nrd=0.76 
m197 0 59 57 0 nenh l=8e-07 w=9e-06 
+ as=8.424e-11 ad=1.224e-11 ps=4.066e-05 pd=1.64e-05 
+ nrs=1.04 nrd=0.15 
m198 41 62 1 1 penh l=8e-07 w=8e-06 
+ as=1.76e-11 ad=1.465e-11 ps=2.29e-05 pd=1.845e-05 
+ nrs=0.28 nrd=0.23 
m199 0 62 41 0 nenh l=8e-07 w=2.2e-06 
+ as=2.059e-11 ad=4.84e-12 ps=9.94e-06 pd=8.8e-06 
+ nrs=4.25 nrd=1 
m200 64 65 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m201 65 64 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m202 66 67 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m203 67 66 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m204 64 65 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m205 68 3 64 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m206 65 64 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m207 66 67 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m208 69 3 65 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m209 70 3 66 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m210 67 66 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m211 71 3 67 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m212 72 12 68 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m213 72 73 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m214 73 12 69 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m215 74 12 70 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m216 0 72 73 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m217 74 75 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m218 75 12 71 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m219 0 74 75 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m220 1 73 72 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m221 1 72 73 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m222 1 75 74 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m223 1 74 75 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m224 76 77 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m225 77 76 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m226 78 79 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m227 79 78 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m228 76 77 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m229 68 22 76 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m230 77 76 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m231 78 79 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m232 69 22 77 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m233 70 22 78 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m234 79 78 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m235 71 22 79 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m236 80 28 68 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m237 80 81 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m238 81 28 69 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m239 82 28 70 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m240 0 80 81 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m241 82 83 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m242 83 28 71 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m243 0 82 83 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m244 1 81 80 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m245 1 80 81 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m246 1 83 82 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m247 1 82 83 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m248 84 85 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m249 85 84 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m250 86 87 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m251 87 86 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m252 84 85 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m253 68 36 84 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m254 85 84 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m255 86 87 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m256 69 36 85 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m257 70 36 86 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m258 87 86 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m259 71 36 87 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m260 88 42 68 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m261 88 89 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m262 89 42 69 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m263 90 42 70 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m264 0 88 89 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m265 90 91 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m266 91 42 71 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m267 0 90 91 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m268 1 89 88 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m269 1 88 89 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m270 1 91 90 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m271 1 90 91 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m272 92 93 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m273 93 92 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m274 94 95 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m275 95 94 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m276 92 93 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m277 68 50 92 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m278 93 92 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m279 94 95 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m280 69 50 93 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m281 70 50 94 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m282 95 94 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m283 71 50 95 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m284 96 56 68 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m285 96 97 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m286 97 56 69 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m287 98 56 70 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m288 0 96 97 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m289 98 99 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m290 99 56 71 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m291 0 98 99 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m292 1 97 96 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m293 1 96 97 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m294 1 99 98 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m295 1 98 99 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m296 100 101 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m297 101 100 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m298 102 103 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m299 103 102 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m300 100 101 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m301 104 3 100 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m302 101 100 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m303 102 103 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m304 105 3 101 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m305 106 3 102 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m306 103 102 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m307 107 3 103 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m308 108 12 104 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m309 108 109 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m310 109 12 105 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m311 110 12 106 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m312 0 108 109 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m313 110 111 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m314 111 12 107 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m315 0 110 111 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m316 1 109 108 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m317 1 108 109 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m318 1 111 110 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m319 1 110 111 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m320 112 113 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m321 113 112 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m322 114 115 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m323 115 114 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m324 112 113 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m325 104 22 112 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m326 113 112 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m327 114 115 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m328 105 22 113 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m329 106 22 114 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m330 115 114 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m331 107 22 115 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m332 116 28 104 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m333 116 117 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m334 117 28 105 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m335 118 28 106 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m336 0 116 117 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m337 118 119 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m338 119 28 107 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m339 0 118 119 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m340 1 117 116 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m341 1 116 117 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m342 1 119 118 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m343 1 118 119 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m344 120 121 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m345 121 120 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m346 122 123 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m347 123 122 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m348 120 121 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m349 104 36 120 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m350 121 120 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m351 122 123 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m352 105 36 121 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m353 106 36 122 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m354 123 122 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m355 107 36 123 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m356 124 42 104 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m357 124 125 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m358 125 42 105 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m359 126 42 106 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m360 0 124 125 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m361 126 127 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m362 127 42 107 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m363 0 126 127 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m364 1 125 124 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m365 1 124 125 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m366 1 127 126 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m367 1 126 127 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m368 128 129 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m369 129 128 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m370 130 131 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m371 131 130 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m372 128 129 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m373 104 50 128 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m374 129 128 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m375 130 131 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m376 105 50 129 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m377 106 50 130 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m378 131 130 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m379 107 50 131 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m380 132 56 104 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m381 132 133 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m382 133 56 105 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m383 134 56 106 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m384 0 132 133 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m385 134 135 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m386 135 56 107 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m387 0 134 135 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m388 1 133 132 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m389 1 132 133 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m390 1 135 134 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m391 1 134 135 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m392 136 137 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m393 137 136 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m394 138 139 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m395 139 138 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m396 136 137 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m397 140 3 136 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m398 137 136 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m399 138 139 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m400 141 3 137 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m401 142 3 138 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m402 139 138 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m403 143 3 139 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m404 144 12 140 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m405 144 145 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m406 145 12 141 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m407 146 12 142 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m408 0 144 145 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m409 146 147 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m410 147 12 143 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m411 0 146 147 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m412 1 145 144 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m413 1 144 145 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m414 1 147 146 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m415 1 146 147 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m416 148 149 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m417 149 148 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m418 150 151 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m419 151 150 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m420 148 149 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m421 140 22 148 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m422 149 148 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m423 150 151 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m424 141 22 149 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m425 142 22 150 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m426 151 150 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m427 143 22 151 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m428 152 28 140 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m429 152 153 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m430 153 28 141 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m431 154 28 142 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m432 0 152 153 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m433 154 155 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m434 155 28 143 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m435 0 154 155 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m436 1 153 152 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m437 1 152 153 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m438 1 155 154 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m439 1 154 155 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m440 156 157 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m441 157 156 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m442 158 159 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m443 159 158 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m444 156 157 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m445 140 36 156 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m446 157 156 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m447 158 159 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m448 141 36 157 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m449 142 36 158 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m450 159 158 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m451 143 36 159 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m452 160 42 140 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m453 160 161 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m454 161 42 141 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m455 162 42 142 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m456 0 160 161 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m457 162 163 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m458 163 42 143 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m459 0 162 163 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m460 1 161 160 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m461 1 160 161 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m462 1 163 162 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m463 1 162 163 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m464 164 165 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m465 165 164 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m466 166 167 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m467 167 166 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m468 164 165 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m469 140 50 164 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m470 165 164 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m471 166 167 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m472 141 50 165 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m473 142 50 166 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m474 167 166 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m475 143 50 167 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m476 168 56 140 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m477 168 169 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m478 169 56 141 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m479 170 56 142 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m480 0 168 169 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m481 170 171 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m482 171 56 143 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m483 0 170 171 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m484 1 169 168 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m485 1 168 169 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m486 1 171 170 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m487 1 170 171 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m488 172 173 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m489 173 172 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m490 174 175 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m491 175 174 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m492 172 173 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m493 176 3 172 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m494 173 172 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m495 174 175 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m496 177 3 173 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m497 178 3 174 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m498 175 174 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m499 179 3 175 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m500 180 12 176 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m501 180 181 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m502 181 12 177 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m503 182 12 178 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m504 0 180 181 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m505 182 183 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m506 183 12 179 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m507 0 182 183 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m508 1 181 180 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m509 1 180 181 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m510 1 183 182 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m511 1 182 183 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m512 184 185 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m513 185 184 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m514 186 187 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m515 187 186 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m516 184 185 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m517 176 22 184 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m518 185 184 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m519 186 187 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m520 177 22 185 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m521 178 22 186 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m522 187 186 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m523 179 22 187 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m524 188 28 176 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m525 188 189 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m526 189 28 177 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m527 190 28 178 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m528 0 188 189 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m529 190 191 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m530 191 28 179 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m531 0 190 191 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m532 1 189 188 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m533 1 188 189 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m534 1 191 190 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m535 1 190 191 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m536 192 193 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m537 193 192 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m538 194 195 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m539 195 194 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m540 192 193 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m541 176 36 192 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m542 193 192 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m543 194 195 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m544 177 36 193 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m545 178 36 194 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m546 195 194 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m547 179 36 195 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m548 196 42 176 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m549 196 197 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m550 197 42 177 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m551 198 42 178 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m552 0 196 197 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m553 198 199 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m554 199 42 179 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m555 0 198 199 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m556 1 197 196 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m557 1 196 197 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m558 1 199 198 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m559 1 198 199 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m560 200 201 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m561 201 200 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m562 202 203 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m563 203 202 1 1 penh l=8e-07 w=2.2e-06 
+ as=4.84e-12 ad=3.03e-12 ps=8.8e-06 pd=5.5e-06 
+ nrs=1 nrd=0.63 
m564 200 201 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m565 176 50 200 0 nenh l=8e-07 w=3.2e-06 
+ as=4.39e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m566 201 200 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m567 202 203 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m568 177 50 201 0 nenh l=8e-07 w=3.2e-06 
+ as=4.33e-12 ad=3.39e-12 ps=5.75e-06 pd=6.78e-06 
+ nrs=0.42 nrd=0.33 
m569 178 50 202 0 nenh l=8e-07 w=3.2e-06 
+ as=4.45e-12 ad=3.39e-12 ps=5.78e-06 pd=6.78e-06 
+ nrs=0.43 nrd=0.33 
m570 203 202 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m571 179 50 203 0 nenh l=8e-07 w=3.2e-06 
+ as=4.47e-12 ad=3.39e-12 ps=6.1e-06 pd=6.78e-06 
+ nrs=0.44 nrd=0.33 
m572 204 56 176 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.39e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.43 
m573 204 205 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m574 205 56 177 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.33e-12 ps=6.78e-06 pd=5.75e-06 
+ nrs=0.33 nrd=0.42 
m575 206 56 178 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.45e-12 ps=6.78e-06 pd=5.78e-06 
+ nrs=0.33 nrd=0.43 
m576 0 204 205 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m577 206 207 0 0 nenh l=8e-07 w=6.8e-06 
+ as=7.21e-12 ad=9.44e-12 ps=1.442e-05 pd=1.28e-05 
+ nrs=0.16 nrd=0.2 
m578 207 56 179 0 nenh l=8e-07 w=3.2e-06 
+ as=3.39e-12 ad=4.47e-12 ps=6.78e-06 pd=6.1e-06 
+ nrs=0.33 nrd=0.44 
m579 0 206 207 0 nenh l=8e-07 w=6.8e-06 
+ as=9.44e-12 ad=7.21e-12 ps=1.28e-05 pd=1.442e-05 
+ nrs=0.2 nrd=0.16 
m580 1 205 204 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m581 1 204 205 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m582 1 207 206 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m583 1 206 207 1 penh l=8e-07 w=2.2e-06 
+ as=3.03e-12 ad=4.84e-12 ps=5.5e-06 pd=8.8e-06 
+ nrs=0.63 nrd=1 
m584 68 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.63e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.26 nrd=0.44 
m585 69 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.73e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.27 nrd=0.44 
m586 70 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.84e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.27 nrd=0.44 
m587 71 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.56e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.26 nrd=0.44 
m588 1 208 68 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.63e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.26 
m589 1 208 69 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.73e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.27 
m590 1 208 70 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.84e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.27 
m591 1 208 71 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.56e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.26 
m592 104 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.63e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.26 nrd=0.44 
m593 105 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.73e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.27 nrd=0.44 
m594 106 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.84e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.27 nrd=0.44 
m595 107 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.56e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.26 nrd=0.44 
m596 1 208 104 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.63e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.26 
m597 1 208 105 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.73e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.27 
m598 1 208 106 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.84e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.27 
m599 1 208 107 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.56e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.26 
m600 140 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.63e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.26 nrd=0.44 
m601 141 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.73e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.27 nrd=0.44 
m602 142 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.84e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.27 nrd=0.44 
m603 143 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.56e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.26 nrd=0.44 
m604 1 208 140 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.63e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.26 
m605 1 208 141 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.73e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.27 
m606 1 208 142 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.84e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.27 
m607 1 208 143 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.56e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.26 
m608 176 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.63e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.26 nrd=0.44 
m609 177 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.73e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.27 nrd=0.44 
m610 178 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.84e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.27 nrd=0.44 
m611 179 208 1 1 penh l=8e-07 w=4.2e-06 
+ as=4.56e-12 ad=7.69e-12 ps=6.81e-06 pd=9.68e-06 
+ nrs=0.26 nrd=0.44 
m612 1 208 176 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.63e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.26 
m613 1 208 177 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.73e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.27 
m614 1 208 178 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.84e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.27 
m615 1 208 179 1 penh l=8e-07 w=4.2e-06 
+ as=7.69e-12 ad=4.56e-12 ps=9.68e-06 pd=6.81e-06 
+ nrs=0.44 nrd=0.26 
m616 1 210 209 1 penh l=8e-07 w=6.8e-06 
+ as=1.245e-11 ad=1.128e-11 ps=1.568e-05 pd=1.8e-05 
+ nrs=0.27 nrd=0.24 
m617 210 209 1 1 penh l=8e-07 w=6.8e-06 
+ as=1.172e-11 ad=1.245e-11 ps=1.84e-05 pd=1.568e-05 
+ nrs=0.25 nrd=0.27 
m618 1 212 211 1 penh l=8e-07 w=6.8e-06 
+ as=1.245e-11 ad=1.128e-11 ps=1.568e-05 pd=1.8e-05 
+ nrs=0.27 nrd=0.24 
m619 212 211 1 1 penh l=8e-07 w=6.8e-06 
+ as=1.128e-11 ad=1.245e-11 ps=1.8e-05 pd=1.568e-05 
+ nrs=0.24 nrd=0.27 
m620 213 68 209 0 nenh l=8e-07 w=2.4e-06 
+ as=3.6e-12 ad=5.28e-12 ps=5.04e-06 pd=9.2e-06 
+ nrs=0.62 nrd=0.92 
m621 210 69 213 0 nenh l=8e-07 w=2.4e-06 
+ as=5.24e-12 ad=3.6e-12 ps=9.2e-06 pd=5.04e-06 
+ nrs=0.91 nrd=0.62 
m622 214 70 211 0 nenh l=8e-07 w=2.4e-06 
+ as=3.6e-12 ad=5.28e-12 ps=5.04e-06 pd=9.2e-06 
+ nrs=0.62 nrd=0.92 
m623 212 71 214 0 nenh l=8e-07 w=2.4e-06 
+ as=5.28e-12 ad=3.6e-12 ps=9.2e-06 pd=5.04e-06 
+ nrs=0.92 nrd=0.62 
m624 0 1 213 0 nenh l=1.2e-06 w=3.2e-06 
+ as=2.995e-11 ad=4.8e-12 ps=1.446e-05 pd=6.72e-06 
+ nrs=2.92 nrd=0.47 
m625 0 1 214 0 nenh l=1.2e-06 w=3.2e-06 
+ as=2.995e-11 ad=4.8e-12 ps=1.446e-05 pd=6.72e-06 
+ nrs=2.92 nrd=0.47 
m626 215 216 0 0 nenh l=8e-07 w=4.4e-06 
+ as=9.68e-12 ad=4.118e-11 ps=1.32e-05 pd=1.988e-05 
+ nrs=0.5 nrd=2.13 
m627 217 218 0 0 nenh l=8e-07 w=4.4e-06 
+ as=9.68e-12 ad=4.118e-11 ps=1.32e-05 pd=1.988e-05 
+ nrs=0.5 nrd=2.13 
m628 1 216 215 1 penh l=8e-07 w=9.4e-06 
+ as=1.721e-11 ad=1.368e-11 ps=2.168e-05 pd=1.72e-05 
+ nrs=0.19 nrd=0.15 
m629 1 218 217 1 penh l=8e-07 w=9.4e-06 
+ as=1.721e-11 ad=1.336e-11 ps=2.168e-05 pd=1.72e-05 
+ nrs=0.19 nrd=0.15 
m630 219 216 220 1 penh l=8e-07 w=3.8e-06 
+ as=4.46e-12 ad=6.44e-12 ps=6.17e-06 pd=1.2e-05 
+ nrs=0.31 nrd=0.45 
m631 221 215 219 1 penh l=8e-07 w=5e-06 
+ as=7.64e-12 ad=5.87e-12 ps=1.44e-05 pd=8.12e-06 
+ nrs=0.31 nrd=0.23 
m632 219 218 222 1 penh l=8e-07 w=4.2e-06 
+ as=4.93e-12 ad=1.428e-11 ps=6.82e-06 pd=1.52e-05 
+ nrs=0.28 nrd=0.81 
m633 223 217 219 1 penh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=4.7e-12 ps=1.24e-05 pd=6.49e-06 
+ nrs=0.55 nrd=0.29 
m634 68 220 0 0 nenh l=8e-07 w=1.34e-05 
+ as=1.84e-11 ad=1.2542e-10 ps=2.556e-05 pd=6.054e-05 
+ nrs=0.1 nrd=0.7 
m635 0 221 69 0 nenh l=8e-07 w=1.38e-05 
+ as=1.2917e-10 ad=1.869e-11 ps=6.235e-05 pd=2.48e-05 
+ nrs=0.68 nrd=0.1 
m636 0 222 70 0 nenh l=8e-07 w=1.38e-05 
+ as=1.2917e-10 ad=1.919e-11 ps=6.235e-05 pd=2.494e-05 
+ nrs=0.68 nrd=0.1 
m637 221 215 0 0 nenh l=8e-07 w=5.6e-06 
+ as=9.23e-12 ad=5.242e-11 ps=1.269e-05 pd=2.53e-05 
+ nrs=0.29 nrd=1.67 
m638 219 216 221 0 nenh l=8e-07 w=3.4e-06 
+ as=4.758e-11 ad=5.61e-12 ps=2.305e-05 pd=7.71e-06 
+ nrs=4.12 nrd=0.48 
m639 220 216 0 0 nenh l=8e-07 w=3.2e-06 
+ as=3.52e-12 ad=2.995e-11 ps=5.4e-06 pd=1.446e-05 
+ nrs=0.34 nrd=2.92 
m640 219 215 220 0 nenh l=8e-07 w=3.2e-06 
+ as=4.478e-11 ad=3.52e-12 ps=2.17e-05 pd=5.4e-06 
+ nrs=4.37 nrd=0.34 
m641 222 218 0 0 nenh l=8e-07 w=5.6e-06 
+ as=8.64e-12 ad=5.242e-11 ps=1.244e-05 pd=2.53e-05 
+ nrs=0.28 nrd=1.67 
m642 0 223 71 0 nenh l=8e-07 w=1.34e-05 
+ as=1.2542e-10 ad=1.871e-11 ps=6.054e-05 pd=2.556e-05 
+ nrs=0.7 nrd=0.1 
m643 219 217 222 0 nenh l=8e-07 w=3.4e-06 
+ as=4.758e-11 ad=5.24e-12 ps=2.305e-05 pd=7.56e-06 
+ nrs=4.12 nrd=0.45 
m644 223 218 219 0 nenh l=8e-07 w=3.2e-06 
+ as=3.52e-12 ad=4.478e-11 ps=5.4e-06 pd=2.17e-05 
+ nrs=0.34 nrd=4.37 
m645 0 217 223 0 nenh l=8e-07 w=3.2e-06 
+ as=2.995e-11 ad=3.52e-12 ps=1.446e-05 pd=5.4e-06 
+ nrs=2.92 nrd=0.34 
m646 224 216 225 0 nenh l=8e-07 w=5.2e-06 
+ as=4.9e-11 ad=7.84e-12 ps=2.31e-05 pd=1.48e-05 
+ nrs=1.81 nrd=0.29 
m647 226 215 224 0 nenh l=8e-07 w=4.2e-06 
+ as=6.84e-12 ad=3.958e-11 ps=1.28e-05 pd=1.865e-05 
+ nrs=0.39 nrd=2.24 
m648 224 218 227 0 nenh l=8e-07 w=4.2e-06 
+ as=3.958e-11 ad=6.84e-12 ps=1.865e-05 pd=1.28e-05 
+ nrs=2.24 nrd=0.39 
m649 228 217 224 0 nenh l=8e-07 w=5.2e-06 
+ as=7.84e-12 ad=4.9e-11 ps=1.48e-05 pd=2.31e-05 
+ nrs=0.29 nrd=1.81 
m650 224 215 225 1 penh l=8e-07 w=3e-06 
+ as=3.3e-12 ad=5.54e-12 ps=5.2e-06 pd=8.12e-06 
+ nrs=0.37 nrd=0.62 
m651 226 216 224 1 penh l=8e-07 w=3e-06 
+ as=2.94e-12 ad=3.3e-12 ps=4.24e-06 pd=5.2e-06 
+ nrs=0.33 nrd=0.37 
m652 1 215 226 1 penh l=8e-07 w=5.2e-06 
+ as=9.52e-12 ad=5.1e-12 ps=1.199e-05 pd=7.36e-06 
+ nrs=0.35 nrd=0.19 
m653 224 217 227 1 penh l=8e-07 w=3e-06 
+ as=3.3e-12 ad=2.94e-12 ps=5.2e-06 pd=4.24e-06 
+ nrs=0.37 nrd=0.33 
m654 228 218 224 1 penh l=8e-07 w=3e-06 
+ as=5.27e-12 ad=3.3e-12 ps=7.78e-06 pd=5.2e-06 
+ nrs=0.59 nrd=0.37 
m655 1 218 227 1 penh l=8e-07 w=5.2e-06 
+ as=9.52e-12 ad=5.1e-12 ps=1.199e-05 pd=7.36e-06 
+ nrs=0.35 nrd=0.19 
m656 1 216 225 1 penh l=8e-07 w=3.8e-06 
+ as=6.96e-12 ad=7.02e-12 ps=8.76e-06 pd=1.028e-05 
+ nrs=0.48 nrd=0.49 
m657 1 217 228 1 penh l=8e-07 w=4.4e-06 
+ as=8.06e-12 ad=7.73e-12 ps=1.015e-05 pd=1.142e-05 
+ nrs=0.42 nrd=0.4 
m658 68 225 1 1 penh l=8e-07 w=6.4e-06 
+ as=7.06e-12 ad=1.172e-11 ps=1.038e-05 pd=1.476e-05 
+ nrs=0.17 nrd=0.29 
m659 1 226 69 1 penh l=8e-07 w=6.4e-06 
+ as=1.172e-11 ad=7.21e-12 ps=1.476e-05 pd=1.038e-05 
+ nrs=0.29 nrd=0.18 
m660 1 227 70 1 penh l=8e-07 w=6.4e-06 
+ as=1.172e-11 ad=7.37e-12 ps=1.476e-05 pd=1.038e-05 
+ nrs=0.29 nrd=0.18 
m661 1 228 71 1 penh l=8e-07 w=6.4e-06 
+ as=1.172e-11 ad=6.95e-12 ps=1.476e-05 pd=1.038e-05 
+ nrs=0.29 nrd=0.17 
m662 1 230 229 1 penh l=8e-07 w=6.8e-06 
+ as=1.245e-11 ad=1.128e-11 ps=1.568e-05 pd=1.8e-05 
+ nrs=0.27 nrd=0.24 
m663 230 229 1 1 penh l=8e-07 w=6.8e-06 
+ as=1.172e-11 ad=1.245e-11 ps=1.84e-05 pd=1.568e-05 
+ nrs=0.25 nrd=0.27 
m664 1 232 231 1 penh l=8e-07 w=6.8e-06 
+ as=1.245e-11 ad=1.128e-11 ps=1.568e-05 pd=1.8e-05 
+ nrs=0.27 nrd=0.24 
m665 232 231 1 1 penh l=8e-07 w=6.8e-06 
+ as=1.128e-11 ad=1.245e-11 ps=1.8e-05 pd=1.568e-05 
+ nrs=0.24 nrd=0.27 
m666 233 104 229 0 nenh l=8e-07 w=2.4e-06 
+ as=3.6e-12 ad=5.28e-12 ps=5.04e-06 pd=9.2e-06 
+ nrs=0.62 nrd=0.92 
m667 230 105 233 0 nenh l=8e-07 w=2.4e-06 
+ as=5.24e-12 ad=3.6e-12 ps=9.2e-06 pd=5.04e-06 
+ nrs=0.91 nrd=0.62 
m668 234 106 231 0 nenh l=8e-07 w=2.4e-06 
+ as=3.6e-12 ad=5.28e-12 ps=5.04e-06 pd=9.2e-06 
+ nrs=0.62 nrd=0.92 
m669 232 107 234 0 nenh l=8e-07 w=2.4e-06 
+ as=5.28e-12 ad=3.6e-12 ps=9.2e-06 pd=5.04e-06 
+ nrs=0.92 nrd=0.62 
m670 0 1 233 0 nenh l=1.2e-06 w=3.2e-06 
+ as=2.995e-11 ad=4.8e-12 ps=1.446e-05 pd=6.72e-06 
+ nrs=2.92 nrd=0.47 
m671 0 1 234 0 nenh l=1.2e-06 w=3.2e-06 
+ as=2.995e-11 ad=4.8e-12 ps=1.446e-05 pd=6.72e-06 
+ nrs=2.92 nrd=0.47 
m672 235 236 0 0 nenh l=8e-07 w=4.4e-06 
+ as=9.68e-12 ad=4.118e-11 ps=1.32e-05 pd=1.988e-05 
+ nrs=0.5 nrd=2.13 
m673 237 238 0 0 nenh l=8e-07 w=4.4e-06 
+ as=9.68e-12 ad=4.118e-11 ps=1.32e-05 pd=1.988e-05 
+ nrs=0.5 nrd=2.13 
m674 1 236 235 1 penh l=8e-07 w=9.4e-06 
+ as=1.721e-11 ad=1.368e-11 ps=2.168e-05 pd=1.72e-05 
+ nrs=0.19 nrd=0.15 
m675 1 238 237 1 penh l=8e-07 w=9.4e-06 
+ as=1.721e-11 ad=1.336e-11 ps=2.168e-05 pd=1.72e-05 
+ nrs=0.19 nrd=0.15 
m676 219 236 239 1 penh l=8e-07 w=3.8e-06 
+ as=4.46e-12 ad=6.44e-12 ps=6.17e-06 pd=1.2e-05 
+ nrs=0.31 nrd=0.45 
m677 240 235 219 1 penh l=8e-07 w=5e-06 
+ as=7.64e-12 ad=5.87e-12 ps=1.44e-05 pd=8.12e-06 
+ nrs=0.31 nrd=0.23 
m678 219 238 241 1 penh l=8e-07 w=4.2e-06 
+ as=4.93e-12 ad=1.428e-11 ps=6.82e-06 pd=1.52e-05 
+ nrs=0.28 nrd=0.81 
m679 242 237 219 1 penh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=4.7e-12 ps=1.24e-05 pd=6.49e-06 
+ nrs=0.55 nrd=0.29 
m680 104 239 0 0 nenh l=8e-07 w=1.34e-05 
+ as=1.84e-11 ad=1.2542e-10 ps=2.556e-05 pd=6.054e-05 
+ nrs=0.1 nrd=0.7 
m681 0 240 105 0 nenh l=8e-07 w=1.38e-05 
+ as=1.2917e-10 ad=1.869e-11 ps=6.235e-05 pd=2.48e-05 
+ nrs=0.68 nrd=0.1 
m682 0 241 106 0 nenh l=8e-07 w=1.38e-05 
+ as=1.2917e-10 ad=1.919e-11 ps=6.235e-05 pd=2.494e-05 
+ nrs=0.68 nrd=0.1 
m683 240 235 0 0 nenh l=8e-07 w=5.6e-06 
+ as=9.23e-12 ad=5.242e-11 ps=1.269e-05 pd=2.53e-05 
+ nrs=0.29 nrd=1.67 
m684 219 236 240 0 nenh l=8e-07 w=3.4e-06 
+ as=4.758e-11 ad=5.61e-12 ps=2.305e-05 pd=7.71e-06 
+ nrs=4.12 nrd=0.48 
m685 239 236 0 0 nenh l=8e-07 w=3.2e-06 
+ as=3.52e-12 ad=2.995e-11 ps=5.4e-06 pd=1.446e-05 
+ nrs=0.34 nrd=2.92 
m686 219 235 239 0 nenh l=8e-07 w=3.2e-06 
+ as=4.478e-11 ad=3.52e-12 ps=2.17e-05 pd=5.4e-06 
+ nrs=4.37 nrd=0.34 
m687 241 238 0 0 nenh l=8e-07 w=5.6e-06 
+ as=8.64e-12 ad=5.242e-11 ps=1.244e-05 pd=2.53e-05 
+ nrs=0.28 nrd=1.67 
m688 0 242 107 0 nenh l=8e-07 w=1.34e-05 
+ as=1.2542e-10 ad=1.871e-11 ps=6.054e-05 pd=2.556e-05 
+ nrs=0.7 nrd=0.1 
m689 219 237 241 0 nenh l=8e-07 w=3.4e-06 
+ as=4.758e-11 ad=5.24e-12 ps=2.305e-05 pd=7.56e-06 
+ nrs=4.12 nrd=0.45 
m690 242 238 219 0 nenh l=8e-07 w=3.2e-06 
+ as=3.52e-12 ad=4.478e-11 ps=5.4e-06 pd=2.17e-05 
+ nrs=0.34 nrd=4.37 
m691 0 237 242 0 nenh l=8e-07 w=3.2e-06 
+ as=2.995e-11 ad=3.52e-12 ps=1.446e-05 pd=5.4e-06 
+ nrs=2.92 nrd=0.34 
m692 224 236 243 0 nenh l=8e-07 w=5.2e-06 
+ as=4.9e-11 ad=7.84e-12 ps=2.31e-05 pd=1.48e-05 
+ nrs=1.81 nrd=0.29 
m693 244 235 224 0 nenh l=8e-07 w=4.2e-06 
+ as=6.84e-12 ad=3.958e-11 ps=1.28e-05 pd=1.865e-05 
+ nrs=0.39 nrd=2.24 
m694 224 238 245 0 nenh l=8e-07 w=4.2e-06 
+ as=3.958e-11 ad=6.84e-12 ps=1.865e-05 pd=1.28e-05 
+ nrs=2.24 nrd=0.39 
m695 246 237 224 0 nenh l=8e-07 w=5.2e-06 
+ as=7.84e-12 ad=4.9e-11 ps=1.48e-05 pd=2.31e-05 
+ nrs=0.29 nrd=1.81 
m696 224 235 243 1 penh l=8e-07 w=3e-06 
+ as=3.3e-12 ad=5.54e-12 ps=5.2e-06 pd=8.12e-06 
+ nrs=0.37 nrd=0.62 
m697 244 236 224 1 penh l=8e-07 w=3e-06 
+ as=2.94e-12 ad=3.3e-12 ps=4.24e-06 pd=5.2e-06 
+ nrs=0.33 nrd=0.37 
m698 1 235 244 1 penh l=8e-07 w=5.2e-06 
+ as=9.52e-12 ad=5.1e-12 ps=1.199e-05 pd=7.36e-06 
+ nrs=0.35 nrd=0.19 
m699 224 237 245 1 penh l=8e-07 w=3e-06 
+ as=3.3e-12 ad=2.94e-12 ps=5.2e-06 pd=4.24e-06 
+ nrs=0.37 nrd=0.33 
m700 246 238 224 1 penh l=8e-07 w=3e-06 
+ as=5.27e-12 ad=3.3e-12 ps=7.78e-06 pd=5.2e-06 
+ nrs=0.59 nrd=0.37 
m701 1 238 245 1 penh l=8e-07 w=5.2e-06 
+ as=9.52e-12 ad=5.1e-12 ps=1.199e-05 pd=7.36e-06 
+ nrs=0.35 nrd=0.19 
m702 1 236 243 1 penh l=8e-07 w=3.8e-06 
+ as=6.96e-12 ad=7.02e-12 ps=8.76e-06 pd=1.028e-05 
+ nrs=0.48 nrd=0.49 
m703 1 237 246 1 penh l=8e-07 w=4.4e-06 
+ as=8.06e-12 ad=7.73e-12 ps=1.015e-05 pd=1.142e-05 
+ nrs=0.42 nrd=0.4 
m704 104 243 1 1 penh l=8e-07 w=6.4e-06 
+ as=7.06e-12 ad=1.172e-11 ps=1.038e-05 pd=1.476e-05 
+ nrs=0.17 nrd=0.29 
m705 1 244 105 1 penh l=8e-07 w=6.4e-06 
+ as=1.172e-11 ad=7.21e-12 ps=1.476e-05 pd=1.038e-05 
+ nrs=0.29 nrd=0.18 
m706 1 245 106 1 penh l=8e-07 w=6.4e-06 
+ as=1.172e-11 ad=7.37e-12 ps=1.476e-05 pd=1.038e-05 
+ nrs=0.29 nrd=0.18 
m707 1 246 107 1 penh l=8e-07 w=6.4e-06 
+ as=1.172e-11 ad=6.95e-12 ps=1.476e-05 pd=1.038e-05 
+ nrs=0.29 nrd=0.17 
m708 1 248 247 1 penh l=8e-07 w=6.8e-06 
+ as=1.245e-11 ad=1.128e-11 ps=1.568e-05 pd=1.8e-05 
+ nrs=0.27 nrd=0.24 
m709 248 247 1 1 penh l=8e-07 w=6.8e-06 
+ as=1.172e-11 ad=1.245e-11 ps=1.84e-05 pd=1.568e-05 
+ nrs=0.25 nrd=0.27 
m710 1 250 249 1 penh l=8e-07 w=6.8e-06 
+ as=1.245e-11 ad=1.128e-11 ps=1.568e-05 pd=1.8e-05 
+ nrs=0.27 nrd=0.24 
m711 250 249 1 1 penh l=8e-07 w=6.8e-06 
+ as=1.128e-11 ad=1.245e-11 ps=1.8e-05 pd=1.568e-05 
+ nrs=0.24 nrd=0.27 
m712 251 140 247 0 nenh l=8e-07 w=2.4e-06 
+ as=3.6e-12 ad=5.28e-12 ps=5.04e-06 pd=9.2e-06 
+ nrs=0.62 nrd=0.92 
m713 248 141 251 0 nenh l=8e-07 w=2.4e-06 
+ as=5.24e-12 ad=3.6e-12 ps=9.2e-06 pd=5.04e-06 
+ nrs=0.91 nrd=0.62 
m714 252 142 249 0 nenh l=8e-07 w=2.4e-06 
+ as=3.6e-12 ad=5.28e-12 ps=5.04e-06 pd=9.2e-06 
+ nrs=0.62 nrd=0.92 
m715 250 143 252 0 nenh l=8e-07 w=2.4e-06 
+ as=5.28e-12 ad=3.6e-12 ps=9.2e-06 pd=5.04e-06 
+ nrs=0.92 nrd=0.62 
m716 0 1 251 0 nenh l=1.2e-06 w=3.2e-06 
+ as=2.995e-11 ad=4.8e-12 ps=1.446e-05 pd=6.72e-06 
+ nrs=2.92 nrd=0.47 
m717 0 1 252 0 nenh l=1.2e-06 w=3.2e-06 
+ as=2.995e-11 ad=4.8e-12 ps=1.446e-05 pd=6.72e-06 
+ nrs=2.92 nrd=0.47 
m718 253 254 0 0 nenh l=8e-07 w=4.4e-06 
+ as=9.68e-12 ad=4.118e-11 ps=1.32e-05 pd=1.988e-05 
+ nrs=0.5 nrd=2.13 
m719 255 256 0 0 nenh l=8e-07 w=4.4e-06 
+ as=9.68e-12 ad=4.118e-11 ps=1.32e-05 pd=1.988e-05 
+ nrs=0.5 nrd=2.13 
m720 1 254 253 1 penh l=8e-07 w=9.4e-06 
+ as=1.721e-11 ad=1.368e-11 ps=2.168e-05 pd=1.72e-05 
+ nrs=0.19 nrd=0.15 
m721 1 256 255 1 penh l=8e-07 w=9.4e-06 
+ as=1.721e-11 ad=1.336e-11 ps=2.168e-05 pd=1.72e-05 
+ nrs=0.19 nrd=0.15 
m722 219 254 257 1 penh l=8e-07 w=3.8e-06 
+ as=4.46e-12 ad=6.44e-12 ps=6.17e-06 pd=1.2e-05 
+ nrs=0.31 nrd=0.45 
m723 258 253 219 1 penh l=8e-07 w=5e-06 
+ as=7.64e-12 ad=5.87e-12 ps=1.44e-05 pd=8.12e-06 
+ nrs=0.31 nrd=0.23 
m724 219 256 259 1 penh l=8e-07 w=4.2e-06 
+ as=4.93e-12 ad=1.428e-11 ps=6.82e-06 pd=1.52e-05 
+ nrs=0.28 nrd=0.81 
m725 260 255 219 1 penh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=4.7e-12 ps=1.24e-05 pd=6.49e-06 
+ nrs=0.55 nrd=0.29 
m726 140 257 0 0 nenh l=8e-07 w=1.34e-05 
+ as=1.84e-11 ad=1.2542e-10 ps=2.556e-05 pd=6.054e-05 
+ nrs=0.1 nrd=0.7 
m727 0 258 141 0 nenh l=8e-07 w=1.38e-05 
+ as=1.2917e-10 ad=1.869e-11 ps=6.235e-05 pd=2.48e-05 
+ nrs=0.68 nrd=0.1 
m728 0 259 142 0 nenh l=8e-07 w=1.38e-05 
+ as=1.2917e-10 ad=1.919e-11 ps=6.235e-05 pd=2.494e-05 
+ nrs=0.68 nrd=0.1 
m729 258 253 0 0 nenh l=8e-07 w=5.6e-06 
+ as=9.23e-12 ad=5.242e-11 ps=1.269e-05 pd=2.53e-05 
+ nrs=0.29 nrd=1.67 
m730 219 254 258 0 nenh l=8e-07 w=3.4e-06 
+ as=4.758e-11 ad=5.61e-12 ps=2.305e-05 pd=7.71e-06 
+ nrs=4.12 nrd=0.48 
m731 257 254 0 0 nenh l=8e-07 w=3.2e-06 
+ as=3.52e-12 ad=2.995e-11 ps=5.4e-06 pd=1.446e-05 
+ nrs=0.34 nrd=2.92 
m732 219 253 257 0 nenh l=8e-07 w=3.2e-06 
+ as=4.478e-11 ad=3.52e-12 ps=2.17e-05 pd=5.4e-06 
+ nrs=4.37 nrd=0.34 
m733 259 256 0 0 nenh l=8e-07 w=5.6e-06 
+ as=8.64e-12 ad=5.242e-11 ps=1.244e-05 pd=2.53e-05 
+ nrs=0.28 nrd=1.67 
m734 0 260 143 0 nenh l=8e-07 w=1.34e-05 
+ as=1.2542e-10 ad=1.871e-11 ps=6.054e-05 pd=2.556e-05 
+ nrs=0.7 nrd=0.1 
m735 219 255 259 0 nenh l=8e-07 w=3.4e-06 
+ as=4.758e-11 ad=5.24e-12 ps=2.305e-05 pd=7.56e-06 
+ nrs=4.12 nrd=0.45 
m736 260 256 219 0 nenh l=8e-07 w=3.2e-06 
+ as=3.52e-12 ad=4.478e-11 ps=5.4e-06 pd=2.17e-05 
+ nrs=0.34 nrd=4.37 
m737 0 255 260 0 nenh l=8e-07 w=3.2e-06 
+ as=2.995e-11 ad=3.52e-12 ps=1.446e-05 pd=5.4e-06 
+ nrs=2.92 nrd=0.34 
m738 224 254 261 0 nenh l=8e-07 w=5.2e-06 
+ as=4.9e-11 ad=7.84e-12 ps=2.31e-05 pd=1.48e-05 
+ nrs=1.81 nrd=0.29 
m739 262 253 224 0 nenh l=8e-07 w=4.2e-06 
+ as=6.84e-12 ad=3.958e-11 ps=1.28e-05 pd=1.865e-05 
+ nrs=0.39 nrd=2.24 
m740 224 256 263 0 nenh l=8e-07 w=4.2e-06 
+ as=3.958e-11 ad=6.84e-12 ps=1.865e-05 pd=1.28e-05 
+ nrs=2.24 nrd=0.39 
m741 264 255 224 0 nenh l=8e-07 w=5.2e-06 
+ as=7.84e-12 ad=4.9e-11 ps=1.48e-05 pd=2.31e-05 
+ nrs=0.29 nrd=1.81 
m742 224 253 261 1 penh l=8e-07 w=3e-06 
+ as=3.3e-12 ad=5.54e-12 ps=5.2e-06 pd=8.12e-06 
+ nrs=0.37 nrd=0.62 
m743 262 254 224 1 penh l=8e-07 w=3e-06 
+ as=2.94e-12 ad=3.3e-12 ps=4.24e-06 pd=5.2e-06 
+ nrs=0.33 nrd=0.37 
m744 1 253 262 1 penh l=8e-07 w=5.2e-06 
+ as=9.52e-12 ad=5.1e-12 ps=1.199e-05 pd=7.36e-06 
+ nrs=0.35 nrd=0.19 
m745 224 255 263 1 penh l=8e-07 w=3e-06 
+ as=3.3e-12 ad=2.94e-12 ps=5.2e-06 pd=4.24e-06 
+ nrs=0.37 nrd=0.33 
m746 264 256 224 1 penh l=8e-07 w=3e-06 
+ as=5.27e-12 ad=3.3e-12 ps=7.78e-06 pd=5.2e-06 
+ nrs=0.59 nrd=0.37 
m747 1 256 263 1 penh l=8e-07 w=5.2e-06 
+ as=9.52e-12 ad=5.1e-12 ps=1.199e-05 pd=7.36e-06 
+ nrs=0.35 nrd=0.19 
m748 1 254 261 1 penh l=8e-07 w=3.8e-06 
+ as=6.96e-12 ad=7.02e-12 ps=8.76e-06 pd=1.028e-05 
+ nrs=0.48 nrd=0.49 
m749 1 255 264 1 penh l=8e-07 w=4.4e-06 
+ as=8.06e-12 ad=7.73e-12 ps=1.015e-05 pd=1.142e-05 
+ nrs=0.42 nrd=0.4 
m750 140 261 1 1 penh l=8e-07 w=6.4e-06 
+ as=7.06e-12 ad=1.172e-11 ps=1.038e-05 pd=1.476e-05 
+ nrs=0.17 nrd=0.29 
m751 1 262 141 1 penh l=8e-07 w=6.4e-06 
+ as=1.172e-11 ad=7.21e-12 ps=1.476e-05 pd=1.038e-05 
+ nrs=0.29 nrd=0.18 
m752 1 263 142 1 penh l=8e-07 w=6.4e-06 
+ as=1.172e-11 ad=7.37e-12 ps=1.476e-05 pd=1.038e-05 
+ nrs=0.29 nrd=0.18 
m753 1 264 143 1 penh l=8e-07 w=6.4e-06 
+ as=1.172e-11 ad=6.95e-12 ps=1.476e-05 pd=1.038e-05 
+ nrs=0.29 nrd=0.17 
m754 1 266 265 1 penh l=8e-07 w=6.8e-06 
+ as=1.245e-11 ad=1.128e-11 ps=1.568e-05 pd=1.8e-05 
+ nrs=0.27 nrd=0.24 
m755 266 265 1 1 penh l=8e-07 w=6.8e-06 
+ as=1.172e-11 ad=1.245e-11 ps=1.84e-05 pd=1.568e-05 
+ nrs=0.25 nrd=0.27 
m756 1 268 267 1 penh l=8e-07 w=6.8e-06 
+ as=1.245e-11 ad=1.128e-11 ps=1.568e-05 pd=1.8e-05 
+ nrs=0.27 nrd=0.24 
m757 268 267 1 1 penh l=8e-07 w=6.8e-06 
+ as=1.128e-11 ad=1.245e-11 ps=1.8e-05 pd=1.568e-05 
+ nrs=0.24 nrd=0.27 
m758 269 176 265 0 nenh l=8e-07 w=2.4e-06 
+ as=3.6e-12 ad=5.28e-12 ps=5.04e-06 pd=9.2e-06 
+ nrs=0.62 nrd=0.92 
m759 266 177 269 0 nenh l=8e-07 w=2.4e-06 
+ as=5.24e-12 ad=3.6e-12 ps=9.2e-06 pd=5.04e-06 
+ nrs=0.91 nrd=0.62 
m760 270 178 267 0 nenh l=8e-07 w=2.4e-06 
+ as=3.6e-12 ad=5.28e-12 ps=5.04e-06 pd=9.2e-06 
+ nrs=0.62 nrd=0.92 
m761 268 179 270 0 nenh l=8e-07 w=2.4e-06 
+ as=5.28e-12 ad=3.6e-12 ps=9.2e-06 pd=5.04e-06 
+ nrs=0.92 nrd=0.62 
m762 0 1 269 0 nenh l=1.2e-06 w=3.2e-06 
+ as=2.995e-11 ad=4.8e-12 ps=1.446e-05 pd=6.72e-06 
+ nrs=2.92 nrd=0.47 
m763 0 1 270 0 nenh l=1.2e-06 w=3.2e-06 
+ as=2.995e-11 ad=4.8e-12 ps=1.446e-05 pd=6.72e-06 
+ nrs=2.92 nrd=0.47 
m764 271 272 0 0 nenh l=8e-07 w=4.4e-06 
+ as=9.68e-12 ad=4.118e-11 ps=1.32e-05 pd=1.988e-05 
+ nrs=0.5 nrd=2.13 
m765 273 274 0 0 nenh l=8e-07 w=4.4e-06 
+ as=9.68e-12 ad=4.118e-11 ps=1.32e-05 pd=1.988e-05 
+ nrs=0.5 nrd=2.13 
m766 1 272 271 1 penh l=8e-07 w=9.4e-06 
+ as=1.721e-11 ad=1.368e-11 ps=2.168e-05 pd=1.72e-05 
+ nrs=0.19 nrd=0.15 
m767 1 274 273 1 penh l=8e-07 w=9.4e-06 
+ as=1.721e-11 ad=1.336e-11 ps=2.168e-05 pd=1.72e-05 
+ nrs=0.19 nrd=0.15 
m768 219 272 275 1 penh l=8e-07 w=3.8e-06 
+ as=4.46e-12 ad=6.44e-12 ps=6.17e-06 pd=1.2e-05 
+ nrs=0.31 nrd=0.45 
m769 276 271 219 1 penh l=8e-07 w=5e-06 
+ as=7.64e-12 ad=5.87e-12 ps=1.44e-05 pd=8.12e-06 
+ nrs=0.31 nrd=0.23 
m770 219 274 277 1 penh l=8e-07 w=4.2e-06 
+ as=4.93e-12 ad=1.428e-11 ps=6.82e-06 pd=1.52e-05 
+ nrs=0.28 nrd=0.81 
m771 278 273 219 1 penh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=4.7e-12 ps=1.24e-05 pd=6.49e-06 
+ nrs=0.55 nrd=0.29 
m772 176 275 0 0 nenh l=8e-07 w=1.34e-05 
+ as=1.84e-11 ad=1.2542e-10 ps=2.556e-05 pd=6.054e-05 
+ nrs=0.1 nrd=0.7 
m773 0 276 177 0 nenh l=8e-07 w=1.38e-05 
+ as=1.2917e-10 ad=1.869e-11 ps=6.235e-05 pd=2.48e-05 
+ nrs=0.68 nrd=0.1 
m774 0 277 178 0 nenh l=8e-07 w=1.38e-05 
+ as=1.2917e-10 ad=1.919e-11 ps=6.235e-05 pd=2.494e-05 
+ nrs=0.68 nrd=0.1 
m775 276 271 0 0 nenh l=8e-07 w=5.6e-06 
+ as=9.23e-12 ad=5.242e-11 ps=1.269e-05 pd=2.53e-05 
+ nrs=0.29 nrd=1.67 
m776 219 272 276 0 nenh l=8e-07 w=3.4e-06 
+ as=4.758e-11 ad=5.61e-12 ps=2.305e-05 pd=7.71e-06 
+ nrs=4.12 nrd=0.48 
m777 275 272 0 0 nenh l=8e-07 w=3.2e-06 
+ as=3.52e-12 ad=2.995e-11 ps=5.4e-06 pd=1.446e-05 
+ nrs=0.34 nrd=2.92 
m778 219 271 275 0 nenh l=8e-07 w=3.2e-06 
+ as=4.478e-11 ad=3.52e-12 ps=2.17e-05 pd=5.4e-06 
+ nrs=4.37 nrd=0.34 
m779 277 274 0 0 nenh l=8e-07 w=5.6e-06 
+ as=8.64e-12 ad=5.242e-11 ps=1.244e-05 pd=2.53e-05 
+ nrs=0.28 nrd=1.67 
m780 0 278 179 0 nenh l=8e-07 w=1.34e-05 
+ as=1.2542e-10 ad=1.871e-11 ps=6.054e-05 pd=2.556e-05 
+ nrs=0.7 nrd=0.1 
m781 219 273 277 0 nenh l=8e-07 w=3.4e-06 
+ as=4.758e-11 ad=5.24e-12 ps=2.305e-05 pd=7.56e-06 
+ nrs=4.12 nrd=0.45 
m782 278 274 219 0 nenh l=8e-07 w=3.2e-06 
+ as=3.52e-12 ad=4.478e-11 ps=5.4e-06 pd=2.17e-05 
+ nrs=0.34 nrd=4.37 
m783 0 273 278 0 nenh l=8e-07 w=3.2e-06 
+ as=2.995e-11 ad=3.52e-12 ps=1.446e-05 pd=5.4e-06 
+ nrs=2.92 nrd=0.34 
m784 224 272 279 0 nenh l=8e-07 w=5.2e-06 
+ as=4.9e-11 ad=7.84e-12 ps=2.31e-05 pd=1.48e-05 
+ nrs=1.81 nrd=0.29 
m785 280 271 224 0 nenh l=8e-07 w=4.2e-06 
+ as=6.84e-12 ad=3.958e-11 ps=1.28e-05 pd=1.865e-05 
+ nrs=0.39 nrd=2.24 
m786 224 274 281 0 nenh l=8e-07 w=4.2e-06 
+ as=3.958e-11 ad=6.84e-12 ps=1.865e-05 pd=1.28e-05 
+ nrs=2.24 nrd=0.39 
m787 282 273 224 0 nenh l=8e-07 w=5.2e-06 
+ as=7.84e-12 ad=4.9e-11 ps=1.48e-05 pd=2.31e-05 
+ nrs=0.29 nrd=1.81 
m788 224 271 279 1 penh l=8e-07 w=3e-06 
+ as=3.3e-12 ad=5.54e-12 ps=5.2e-06 pd=8.12e-06 
+ nrs=0.37 nrd=0.62 
m789 280 272 224 1 penh l=8e-07 w=3e-06 
+ as=2.94e-12 ad=3.3e-12 ps=4.24e-06 pd=5.2e-06 
+ nrs=0.33 nrd=0.37 
m790 1 271 280 1 penh l=8e-07 w=5.2e-06 
+ as=9.52e-12 ad=5.1e-12 ps=1.199e-05 pd=7.36e-06 
+ nrs=0.35 nrd=0.19 
m791 224 273 281 1 penh l=8e-07 w=3e-06 
+ as=3.3e-12 ad=2.94e-12 ps=5.2e-06 pd=4.24e-06 
+ nrs=0.37 nrd=0.33 
m792 282 274 224 1 penh l=8e-07 w=3e-06 
+ as=5.27e-12 ad=3.3e-12 ps=7.78e-06 pd=5.2e-06 
+ nrs=0.59 nrd=0.37 
m793 1 274 281 1 penh l=8e-07 w=5.2e-06 
+ as=9.52e-12 ad=5.1e-12 ps=1.199e-05 pd=7.36e-06 
+ nrs=0.35 nrd=0.19 
m794 1 272 279 1 penh l=8e-07 w=3.8e-06 
+ as=6.96e-12 ad=7.02e-12 ps=8.76e-06 pd=1.028e-05 
+ nrs=0.48 nrd=0.49 
m795 1 273 282 1 penh l=8e-07 w=4.4e-06 
+ as=8.06e-12 ad=7.73e-12 ps=1.015e-05 pd=1.142e-05 
+ nrs=0.42 nrd=0.4 
m796 176 279 1 1 penh l=8e-07 w=6.4e-06 
+ as=7.06e-12 ad=1.172e-11 ps=1.038e-05 pd=1.476e-05 
+ nrs=0.17 nrd=0.29 
m797 1 280 177 1 penh l=8e-07 w=6.4e-06 
+ as=1.172e-11 ad=7.21e-12 ps=1.476e-05 pd=1.038e-05 
+ nrs=0.29 nrd=0.18 
m798 1 281 178 1 penh l=8e-07 w=6.4e-06 
+ as=1.172e-11 ad=7.37e-12 ps=1.476e-05 pd=1.038e-05 
+ nrs=0.29 nrd=0.18 
m799 1 282 179 1 penh l=8e-07 w=6.4e-06 
+ as=1.172e-11 ad=6.95e-12 ps=1.476e-05 pd=1.038e-05 
+ nrs=0.29 nrd=0.17 
m800 283 285 284 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.59 nrd=0.67 
m801 283 285 286 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.59 nrd=1 
m802 0 287 283 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=5.22e-12 ps=1.807e-05 pd=7.62e-06 
+ nrs=2.34 nrd=0.33 
m803 288 285 289 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.59 nrd=0.67 
m804 283 208 286 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.6 nrd=1 
m805 288 285 290 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.59 nrd=1 
m806 0 291 288 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=5.22e-12 ps=1.807e-05 pd=7.62e-06 
+ nrs=2.34 nrd=0.33 
m807 283 208 284 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.6 nrd=0.67 
m808 1 287 283 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=5.28e-12 ps=9.22e-06 pd=7.62e-06 
+ nrs=0.46 nrd=0.33 
m809 288 208 290 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.6 nrd=1 
m810 288 208 289 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.6 nrd=0.67 
m811 1 291 288 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=5.28e-12 ps=9.22e-06 pd=7.62e-06 
+ nrs=0.46 nrd=0.33 
m812 1 284 287 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=8.8e-12 ps=9.22e-06 pd=1.24e-05 
+ nrs=0.46 nrd=0.55 
m813 292 286 1 1 penh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=7.32e-12 ps=1.24e-05 pd=9.22e-06 
+ nrs=0.55 nrd=0.46 
m814 1 289 291 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=8.8e-12 ps=9.22e-06 pd=1.24e-05 
+ nrs=0.46 nrd=0.55 
m815 293 290 1 1 penh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=7.32e-12 ps=1.24e-05 pd=9.22e-06 
+ nrs=0.55 nrd=0.46 
m816 0 284 287 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=6.64e-12 ps=1.807e-05 pd=1.24e-05 
+ nrs=2.34 nrd=0.42 
m817 292 286 0 0 nenh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=3.744e-11 ps=1.24e-05 pd=1.807e-05 
+ nrs=0.55 nrd=2.34 
m818 0 289 291 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=6.64e-12 ps=1.807e-05 pd=1.24e-05 
+ nrs=2.34 nrd=0.42 
m819 293 290 0 0 nenh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=3.744e-11 ps=1.24e-05 pd=1.807e-05 
+ nrs=0.55 nrd=2.34 
m820 284 295 294 0 nenh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=4.84e-12 ps=5.87e-06 pd=7.52e-06 
+ nrs=0.67 nrd=1 
m821 296 297 284 0 nenh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m822 0 209 296 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=4.28e-12 ps=1.807e-05 pd=8e-06 
+ nrs=2.34 nrd=0.27 
m823 216 292 0 0 nenh l=8e-07 w=4e-06 
+ as=4.28e-12 ad=3.744e-11 ps=8e-06 pd=1.807e-05 
+ nrs=0.27 nrd=2.34 
m824 289 295 216 0 nenh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=2.36e-12 ps=5.87e-06 pd=4.4e-06 
+ nrs=0.67 nrd=0.49 
m825 298 297 289 0 nenh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m826 0 211 298 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=4.28e-12 ps=1.807e-05 pd=8e-06 
+ nrs=2.34 nrd=0.27 
m827 218 293 0 0 nenh l=8e-07 w=4e-06 
+ as=4.28e-12 ad=3.744e-11 ps=8e-06 pd=1.807e-05 
+ nrs=0.27 nrd=2.34 
m828 284 299 294 1 penh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=4.84e-12 ps=5.87e-06 pd=7.52e-06 
+ nrs=0.67 nrd=1 
m829 296 300 284 1 penh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m830 1 209 296 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=4.28e-12 ps=9.22e-06 pd=8e-06 
+ nrs=0.46 nrd=0.27 
m831 216 292 1 1 penh l=8e-07 w=4e-06 
+ as=4.28e-12 ad=7.32e-12 ps=8e-06 pd=9.22e-06 
+ nrs=0.27 nrd=0.46 
m832 289 299 216 1 penh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=2.36e-12 ps=5.87e-06 pd=4.4e-06 
+ nrs=0.67 nrd=0.49 
m833 298 300 289 1 penh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m834 1 211 298 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=4.28e-12 ps=9.22e-06 pd=8e-06 
+ nrs=0.46 nrd=0.27 
m835 218 293 1 1 penh l=8e-07 w=4e-06 
+ as=4.28e-12 ad=7.32e-12 ps=8e-06 pd=9.22e-06 
+ nrs=0.27 nrd=0.46 
m836 301 285 302 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.59 nrd=0.67 
m837 301 285 303 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.59 nrd=1 
m838 0 304 301 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=5.22e-12 ps=1.807e-05 pd=7.62e-06 
+ nrs=2.34 nrd=0.33 
m839 305 285 306 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.59 nrd=0.67 
m840 301 208 303 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.6 nrd=1 
m841 305 285 307 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.59 nrd=1 
m842 0 308 305 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=5.22e-12 ps=1.807e-05 pd=7.62e-06 
+ nrs=2.34 nrd=0.33 
m843 301 208 302 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.6 nrd=0.67 
m844 1 304 301 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=5.28e-12 ps=9.22e-06 pd=7.62e-06 
+ nrs=0.46 nrd=0.33 
m845 305 208 307 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.6 nrd=1 
m846 305 208 306 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.6 nrd=0.67 
m847 1 308 305 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=5.28e-12 ps=9.22e-06 pd=7.62e-06 
+ nrs=0.46 nrd=0.33 
m848 1 302 304 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=8.8e-12 ps=9.22e-06 pd=1.24e-05 
+ nrs=0.46 nrd=0.55 
m849 309 303 1 1 penh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=7.32e-12 ps=1.24e-05 pd=9.22e-06 
+ nrs=0.55 nrd=0.46 
m850 1 306 308 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=8.8e-12 ps=9.22e-06 pd=1.24e-05 
+ nrs=0.46 nrd=0.55 
m851 310 307 1 1 penh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=7.32e-12 ps=1.24e-05 pd=9.22e-06 
+ nrs=0.55 nrd=0.46 
m852 0 302 304 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=6.64e-12 ps=1.807e-05 pd=1.24e-05 
+ nrs=2.34 nrd=0.42 
m853 309 303 0 0 nenh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=3.744e-11 ps=1.24e-05 pd=1.807e-05 
+ nrs=0.55 nrd=2.34 
m854 0 306 308 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=6.64e-12 ps=1.807e-05 pd=1.24e-05 
+ nrs=2.34 nrd=0.42 
m855 310 307 0 0 nenh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=3.744e-11 ps=1.24e-05 pd=1.807e-05 
+ nrs=0.55 nrd=2.34 
m856 302 295 218 0 nenh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=2.36e-12 ps=5.87e-06 pd=4.4e-06 
+ nrs=0.67 nrd=0.49 
m857 311 297 302 0 nenh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m858 0 229 311 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=4.28e-12 ps=1.807e-05 pd=8e-06 
+ nrs=2.34 nrd=0.27 
m859 236 309 0 0 nenh l=8e-07 w=4e-06 
+ as=4.28e-12 ad=3.744e-11 ps=8e-06 pd=1.807e-05 
+ nrs=0.27 nrd=2.34 
m860 306 295 236 0 nenh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=2.36e-12 ps=5.87e-06 pd=4.4e-06 
+ nrs=0.67 nrd=0.49 
m861 312 297 306 0 nenh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m862 0 231 312 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=4.28e-12 ps=1.807e-05 pd=8e-06 
+ nrs=2.34 nrd=0.27 
m863 238 310 0 0 nenh l=8e-07 w=4e-06 
+ as=4.28e-12 ad=3.744e-11 ps=8e-06 pd=1.807e-05 
+ nrs=0.27 nrd=2.34 
m864 302 299 218 1 penh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=2.36e-12 ps=5.87e-06 pd=4.4e-06 
+ nrs=0.67 nrd=0.49 
m865 311 300 302 1 penh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m866 1 229 311 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=4.28e-12 ps=9.22e-06 pd=8e-06 
+ nrs=0.46 nrd=0.27 
m867 236 309 1 1 penh l=8e-07 w=4e-06 
+ as=4.28e-12 ad=7.32e-12 ps=8e-06 pd=9.22e-06 
+ nrs=0.27 nrd=0.46 
m868 306 299 236 1 penh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=2.36e-12 ps=5.87e-06 pd=4.4e-06 
+ nrs=0.67 nrd=0.49 
m869 312 300 306 1 penh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m870 1 231 312 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=4.28e-12 ps=9.22e-06 pd=8e-06 
+ nrs=0.46 nrd=0.27 
m871 238 310 1 1 penh l=8e-07 w=4e-06 
+ as=4.28e-12 ad=7.32e-12 ps=8e-06 pd=9.22e-06 
+ nrs=0.27 nrd=0.46 
m872 313 285 314 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.59 nrd=0.67 
m873 313 285 315 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.59 nrd=1 
m874 0 316 313 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=5.22e-12 ps=1.807e-05 pd=7.62e-06 
+ nrs=2.34 nrd=0.33 
m875 317 285 318 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.59 nrd=0.67 
m876 313 208 315 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.6 nrd=1 
m877 317 285 319 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.59 nrd=1 
m878 0 320 317 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=5.22e-12 ps=1.807e-05 pd=7.62e-06 
+ nrs=2.34 nrd=0.33 
m879 313 208 314 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.6 nrd=0.67 
m880 1 316 313 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=5.28e-12 ps=9.22e-06 pd=7.62e-06 
+ nrs=0.46 nrd=0.33 
m881 317 208 319 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.6 nrd=1 
m882 317 208 318 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.6 nrd=0.67 
m883 1 320 317 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=5.28e-12 ps=9.22e-06 pd=7.62e-06 
+ nrs=0.46 nrd=0.33 
m884 1 314 316 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=8.8e-12 ps=9.22e-06 pd=1.24e-05 
+ nrs=0.46 nrd=0.55 
m885 321 315 1 1 penh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=7.32e-12 ps=1.24e-05 pd=9.22e-06 
+ nrs=0.55 nrd=0.46 
m886 1 318 320 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=8.8e-12 ps=9.22e-06 pd=1.24e-05 
+ nrs=0.46 nrd=0.55 
m887 322 319 1 1 penh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=7.32e-12 ps=1.24e-05 pd=9.22e-06 
+ nrs=0.55 nrd=0.46 
m888 0 314 316 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=6.64e-12 ps=1.807e-05 pd=1.24e-05 
+ nrs=2.34 nrd=0.42 
m889 321 315 0 0 nenh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=3.744e-11 ps=1.24e-05 pd=1.807e-05 
+ nrs=0.55 nrd=2.34 
m890 0 318 320 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=6.64e-12 ps=1.807e-05 pd=1.24e-05 
+ nrs=2.34 nrd=0.42 
m891 322 319 0 0 nenh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=3.744e-11 ps=1.24e-05 pd=1.807e-05 
+ nrs=0.55 nrd=2.34 
m892 314 295 238 0 nenh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=2.36e-12 ps=5.87e-06 pd=4.4e-06 
+ nrs=0.67 nrd=0.49 
m893 323 297 314 0 nenh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m894 0 247 323 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=4.28e-12 ps=1.807e-05 pd=8e-06 
+ nrs=2.34 nrd=0.27 
m895 254 321 0 0 nenh l=8e-07 w=4e-06 
+ as=4.28e-12 ad=3.744e-11 ps=8e-06 pd=1.807e-05 
+ nrs=0.27 nrd=2.34 
m896 318 295 254 0 nenh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=2.36e-12 ps=5.87e-06 pd=4.4e-06 
+ nrs=0.67 nrd=0.49 
m897 324 297 318 0 nenh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m898 0 249 324 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=4.28e-12 ps=1.807e-05 pd=8e-06 
+ nrs=2.34 nrd=0.27 
m899 256 322 0 0 nenh l=8e-07 w=4e-06 
+ as=4.28e-12 ad=3.744e-11 ps=8e-06 pd=1.807e-05 
+ nrs=0.27 nrd=2.34 
m900 314 299 238 1 penh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=2.36e-12 ps=5.87e-06 pd=4.4e-06 
+ nrs=0.67 nrd=0.49 
m901 323 300 314 1 penh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m902 1 247 323 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=4.28e-12 ps=9.22e-06 pd=8e-06 
+ nrs=0.46 nrd=0.27 
m903 254 321 1 1 penh l=8e-07 w=4e-06 
+ as=4.28e-12 ad=7.32e-12 ps=8e-06 pd=9.22e-06 
+ nrs=0.27 nrd=0.46 
m904 318 299 254 1 penh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=2.36e-12 ps=5.87e-06 pd=4.4e-06 
+ nrs=0.67 nrd=0.49 
m905 324 300 318 1 penh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m906 1 249 324 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=4.28e-12 ps=9.22e-06 pd=8e-06 
+ nrs=0.46 nrd=0.27 
m907 256 322 1 1 penh l=8e-07 w=4e-06 
+ as=4.28e-12 ad=7.32e-12 ps=8e-06 pd=9.22e-06 
+ nrs=0.27 nrd=0.46 
m908 325 285 326 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.59 nrd=0.67 
m909 325 285 327 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.59 nrd=1 
m910 0 328 325 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=5.22e-12 ps=1.807e-05 pd=7.62e-06 
+ nrs=2.34 nrd=0.33 
m911 329 285 330 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.59 nrd=0.67 
m912 325 208 327 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.6 nrd=1 
m913 329 285 331 0 nenh l=8e-07 w=2.2e-06 
+ as=2.87e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.59 nrd=1 
m914 0 332 329 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=5.22e-12 ps=1.807e-05 pd=7.62e-06 
+ nrs=2.34 nrd=0.33 
m915 325 208 326 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.6 nrd=0.67 
m916 1 328 325 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=5.28e-12 ps=9.22e-06 pd=7.62e-06 
+ nrs=0.46 nrd=0.33 
m917 329 208 331 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=4.84e-12 ps=4.19e-06 pd=8.8e-06 
+ nrs=0.6 nrd=1 
m918 329 208 330 1 penh l=8e-07 w=2.2e-06 
+ as=2.9e-12 ad=3.23e-12 ps=4.19e-06 pd=5.87e-06 
+ nrs=0.6 nrd=0.67 
m919 1 332 329 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=5.28e-12 ps=9.22e-06 pd=7.62e-06 
+ nrs=0.46 nrd=0.33 
m920 1 326 328 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=8.8e-12 ps=9.22e-06 pd=1.24e-05 
+ nrs=0.46 nrd=0.55 
m921 333 327 1 1 penh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=7.32e-12 ps=1.24e-05 pd=9.22e-06 
+ nrs=0.55 nrd=0.46 
m922 1 330 332 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=8.8e-12 ps=9.22e-06 pd=1.24e-05 
+ nrs=0.46 nrd=0.55 
m923 334 331 1 1 penh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=7.32e-12 ps=1.24e-05 pd=9.22e-06 
+ nrs=0.55 nrd=0.46 
m924 0 326 328 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=6.64e-12 ps=1.807e-05 pd=1.24e-05 
+ nrs=2.34 nrd=0.42 
m925 333 327 0 0 nenh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=3.744e-11 ps=1.24e-05 pd=1.807e-05 
+ nrs=0.55 nrd=2.34 
m926 0 330 332 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=6.64e-12 ps=1.807e-05 pd=1.24e-05 
+ nrs=2.34 nrd=0.42 
m927 334 331 0 0 nenh l=8e-07 w=4e-06 
+ as=8.8e-12 ad=3.744e-11 ps=1.24e-05 pd=1.807e-05 
+ nrs=0.55 nrd=2.34 
m928 326 295 256 0 nenh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=2.36e-12 ps=5.87e-06 pd=4.4e-06 
+ nrs=0.67 nrd=0.49 
m929 335 297 326 0 nenh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m930 0 265 335 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=4.28e-12 ps=1.807e-05 pd=8e-06 
+ nrs=2.34 nrd=0.27 
m931 272 333 0 0 nenh l=8e-07 w=4e-06 
+ as=4.28e-12 ad=3.744e-11 ps=8e-06 pd=1.807e-05 
+ nrs=0.27 nrd=2.34 
m932 330 295 272 0 nenh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=2.36e-12 ps=5.87e-06 pd=4.4e-06 
+ nrs=0.67 nrd=0.49 
m933 336 297 330 0 nenh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m934 0 267 336 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=4.28e-12 ps=1.807e-05 pd=8e-06 
+ nrs=2.34 nrd=0.27 
m935 274 334 0 0 nenh l=8e-07 w=4e-06 
+ as=6.64e-12 ad=3.744e-11 ps=1.24e-05 pd=1.807e-05 
+ nrs=0.42 nrd=2.34 
m936 326 299 256 1 penh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=2.36e-12 ps=5.87e-06 pd=4.4e-06 
+ nrs=0.67 nrd=0.49 
m937 335 300 326 1 penh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m938 1 265 335 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=4.28e-12 ps=9.22e-06 pd=8e-06 
+ nrs=0.46 nrd=0.27 
m939 272 333 1 1 penh l=8e-07 w=4e-06 
+ as=4.28e-12 ad=7.32e-12 ps=8e-06 pd=9.22e-06 
+ nrs=0.27 nrd=0.46 
m940 330 299 272 1 penh l=8e-07 w=2.2e-06 
+ as=3.23e-12 ad=2.36e-12 ps=5.87e-06 pd=4.4e-06 
+ nrs=0.67 nrd=0.49 
m941 336 300 330 1 penh l=8e-07 w=2.2e-06 
+ as=2.36e-12 ad=3.23e-12 ps=4.4e-06 pd=5.87e-06 
+ nrs=0.49 nrd=0.67 
m942 1 267 336 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=4.28e-12 ps=9.22e-06 pd=8e-06 
+ nrs=0.46 nrd=0.27 
m943 274 334 1 1 penh l=8e-07 w=4e-06 
+ as=6.64e-12 ad=7.32e-12 ps=1.24e-05 pd=9.22e-06 
+ nrs=0.42 nrd=0.46 
m944 0 21 337 0 nenh l=8e-07 w=1.2e-05 
+ as=1.1232e-10 ad=2.64e-11 ps=5.422e-05 pd=2.84e-05 
+ nrs=0.78 nrd=0.18 
m945 337 21 0 0 nenh l=8e-07 w=1.2e-05 
+ as=2.64e-11 ad=1.1232e-10 ps=2.84e-05 pd=5.422e-05 
+ nrs=0.18 nrd=0.78 
m946 0 337 338 0 nenh l=8e-07 w=1.2e-05 
+ as=1.1232e-10 ad=1.54e-11 ps=5.422e-05 pd=1.657e-05 
+ nrs=0.78 nrd=0.11 
m947 338 337 0 0 nenh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=1.1232e-10 ps=1.657e-05 pd=5.422e-05 
+ nrs=0.11 nrd=0.78 
m948 0 337 338 0 nenh l=8e-07 w=1.2e-05 
+ as=1.1232e-10 ad=1.54e-11 ps=5.422e-05 pd=1.657e-05 
+ nrs=0.78 nrd=0.11 
m949 338 337 0 0 nenh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=1.1232e-10 ps=1.657e-05 pd=5.422e-05 
+ nrs=0.11 nrd=0.78 
m950 0 337 338 0 nenh l=8e-07 w=1.2e-05 
+ as=1.1232e-10 ad=1.54e-11 ps=5.422e-05 pd=1.657e-05 
+ nrs=0.78 nrd=0.11 
m951 338 337 0 0 nenh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=1.1232e-10 ps=1.657e-05 pd=5.422e-05 
+ nrs=0.11 nrd=0.78 
m952 0 337 338 0 nenh l=8e-07 w=1.2e-05 
+ as=1.1232e-10 ad=1.54e-11 ps=5.422e-05 pd=1.657e-05 
+ nrs=0.78 nrd=0.11 
m953 338 337 0 0 nenh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=1.1232e-10 ps=1.657e-05 pd=5.422e-05 
+ nrs=0.11 nrd=0.78 
m954 0 337 338 0 nenh l=8e-07 w=1.2e-05 
+ as=1.1232e-10 ad=1.54e-11 ps=5.422e-05 pd=1.657e-05 
+ nrs=0.78 nrd=0.11 
m955 338 337 0 0 nenh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=1.1232e-10 ps=1.657e-05 pd=5.422e-05 
+ nrs=0.11 nrd=0.78 
m956 0 337 338 0 nenh l=8e-07 w=1.2e-05 
+ as=1.1232e-10 ad=1.54e-11 ps=5.422e-05 pd=1.657e-05 
+ nrs=0.78 nrd=0.11 
m957 338 337 0 0 nenh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=1.1232e-10 ps=1.657e-05 pd=5.422e-05 
+ nrs=0.11 nrd=0.78 
m958 1 21 337 1 penh l=8e-07 w=1.2e-05 
+ as=2.197e-11 ad=2.64e-11 ps=2.767e-05 pd=2.84e-05 
+ nrs=0.15 nrd=0.18 
m959 337 21 1 1 penh l=8e-07 w=1.2e-05 
+ as=2.64e-11 ad=2.197e-11 ps=2.84e-05 pd=2.767e-05 
+ nrs=0.18 nrd=0.15 
m960 1 337 338 1 penh l=8e-07 w=1.2e-05 
+ as=2.197e-11 ad=1.54e-11 ps=2.767e-05 pd=1.657e-05 
+ nrs=0.15 nrd=0.11 
m961 338 337 1 1 penh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=2.197e-11 ps=1.657e-05 pd=2.767e-05 
+ nrs=0.11 nrd=0.15 
m962 1 337 338 1 penh l=8e-07 w=1.2e-05 
+ as=2.197e-11 ad=1.54e-11 ps=2.767e-05 pd=1.657e-05 
+ nrs=0.15 nrd=0.11 
m963 338 337 1 1 penh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=2.197e-11 ps=1.657e-05 pd=2.767e-05 
+ nrs=0.11 nrd=0.15 
m964 1 337 338 1 penh l=8e-07 w=1.2e-05 
+ as=2.197e-11 ad=1.54e-11 ps=2.767e-05 pd=1.657e-05 
+ nrs=0.15 nrd=0.11 
m965 338 337 1 1 penh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=2.197e-11 ps=1.657e-05 pd=2.767e-05 
+ nrs=0.11 nrd=0.15 
m966 1 337 338 1 penh l=8e-07 w=1.2e-05 
+ as=2.197e-11 ad=1.54e-11 ps=2.767e-05 pd=1.657e-05 
+ nrs=0.15 nrd=0.11 
m967 338 337 1 1 penh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=2.197e-11 ps=1.657e-05 pd=2.767e-05 
+ nrs=0.11 nrd=0.15 
m968 1 337 338 1 penh l=8e-07 w=1.2e-05 
+ as=2.197e-11 ad=1.54e-11 ps=2.767e-05 pd=1.657e-05 
+ nrs=0.15 nrd=0.11 
m969 338 337 1 1 penh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=2.197e-11 ps=1.657e-05 pd=2.767e-05 
+ nrs=0.11 nrd=0.15 
m970 1 337 338 1 penh l=8e-07 w=1.2e-05 
+ as=2.197e-11 ad=1.54e-11 ps=2.767e-05 pd=1.657e-05 
+ nrs=0.15 nrd=0.11 
m971 338 337 1 1 penh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=2.197e-11 ps=1.657e-05 pd=2.767e-05 
+ nrs=0.11 nrd=0.15 
m972 0 339 55 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=8.8e-12 ps=1.807e-05 pd=1.368e-05 
+ nrs=2.34 nrd=0.55 
m973 339 340 0 0 nenh l=1.6e-06 w=4e-06 
+ as=8.8e-12 ad=3.744e-11 ps=1.24e-05 pd=1.807e-05 
+ nrs=0.55 nrd=2.34 
m974 1 339 55 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=8.8e-12 ps=9.22e-06 pd=1.368e-05 
+ nrs=0.46 nrd=0.55 
m975 339 340 1 1 penh l=1.6e-06 w=4e-06 
+ as=8.8e-12 ad=7.32e-12 ps=1.24e-05 pd=9.22e-06 
+ nrs=0.55 nrd=0.46 
m976 0 274 341 0 nenh l=8e-07 w=1.2e-05 
+ as=1.1232e-10 ad=2.64e-11 ps=5.422e-05 pd=2.84e-05 
+ nrs=0.78 nrd=0.18 
m977 341 274 0 0 nenh l=8e-07 w=1.2e-05 
+ as=2.64e-11 ad=1.1232e-10 ps=2.84e-05 pd=5.422e-05 
+ nrs=0.18 nrd=0.78 
m978 0 341 342 0 nenh l=8e-07 w=1.2e-05 
+ as=1.1232e-10 ad=1.54e-11 ps=5.422e-05 pd=1.657e-05 
+ nrs=0.78 nrd=0.11 
m979 342 341 0 0 nenh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=1.1232e-10 ps=1.657e-05 pd=5.422e-05 
+ nrs=0.11 nrd=0.78 
m980 0 341 342 0 nenh l=8e-07 w=1.2e-05 
+ as=1.1232e-10 ad=1.54e-11 ps=5.422e-05 pd=1.657e-05 
+ nrs=0.78 nrd=0.11 
m981 342 341 0 0 nenh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=1.1232e-10 ps=1.657e-05 pd=5.422e-05 
+ nrs=0.11 nrd=0.78 
m982 0 341 342 0 nenh l=8e-07 w=1.2e-05 
+ as=1.1232e-10 ad=1.54e-11 ps=5.422e-05 pd=1.657e-05 
+ nrs=0.78 nrd=0.11 
m983 342 341 0 0 nenh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=1.1232e-10 ps=1.657e-05 pd=5.422e-05 
+ nrs=0.11 nrd=0.78 
m984 0 341 342 0 nenh l=8e-07 w=1.2e-05 
+ as=1.1232e-10 ad=1.54e-11 ps=5.422e-05 pd=1.657e-05 
+ nrs=0.78 nrd=0.11 
m985 342 341 0 0 nenh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=1.1232e-10 ps=1.657e-05 pd=5.422e-05 
+ nrs=0.11 nrd=0.78 
m986 0 341 342 0 nenh l=8e-07 w=1.2e-05 
+ as=1.1232e-10 ad=1.54e-11 ps=5.422e-05 pd=1.657e-05 
+ nrs=0.78 nrd=0.11 
m987 342 341 0 0 nenh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=1.1232e-10 ps=1.657e-05 pd=5.422e-05 
+ nrs=0.11 nrd=0.78 
m988 0 341 342 0 nenh l=8e-07 w=1.2e-05 
+ as=1.1232e-10 ad=1.54e-11 ps=5.422e-05 pd=1.657e-05 
+ nrs=0.78 nrd=0.11 
m989 342 341 0 0 nenh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=1.1232e-10 ps=1.657e-05 pd=5.422e-05 
+ nrs=0.11 nrd=0.78 
m990 1 274 341 1 penh l=8e-07 w=1.2e-05 
+ as=2.197e-11 ad=2.64e-11 ps=2.767e-05 pd=2.84e-05 
+ nrs=0.15 nrd=0.18 
m991 341 274 1 1 penh l=8e-07 w=1.2e-05 
+ as=2.64e-11 ad=2.197e-11 ps=2.84e-05 pd=2.767e-05 
+ nrs=0.18 nrd=0.15 
m992 1 341 342 1 penh l=8e-07 w=1.2e-05 
+ as=2.197e-11 ad=1.54e-11 ps=2.767e-05 pd=1.657e-05 
+ nrs=0.15 nrd=0.11 
m993 342 341 1 1 penh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=2.197e-11 ps=1.657e-05 pd=2.767e-05 
+ nrs=0.11 nrd=0.15 
m994 1 341 342 1 penh l=8e-07 w=1.2e-05 
+ as=2.197e-11 ad=1.54e-11 ps=2.767e-05 pd=1.657e-05 
+ nrs=0.15 nrd=0.11 
m995 342 341 1 1 penh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=2.197e-11 ps=1.657e-05 pd=2.767e-05 
+ nrs=0.11 nrd=0.15 
m996 1 341 342 1 penh l=8e-07 w=1.2e-05 
+ as=2.197e-11 ad=1.54e-11 ps=2.767e-05 pd=1.657e-05 
+ nrs=0.15 nrd=0.11 
m997 342 341 1 1 penh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=2.197e-11 ps=1.657e-05 pd=2.767e-05 
+ nrs=0.11 nrd=0.15 
m998 1 341 342 1 penh l=8e-07 w=1.2e-05 
+ as=2.197e-11 ad=1.54e-11 ps=2.767e-05 pd=1.657e-05 
+ nrs=0.15 nrd=0.11 
m999 342 341 1 1 penh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=2.197e-11 ps=1.657e-05 pd=2.767e-05 
+ nrs=0.11 nrd=0.15 
m1000 1 341 342 1 penh l=8e-07 w=1.2e-05 
+ as=2.197e-11 ad=1.54e-11 ps=2.767e-05 pd=1.657e-05 
+ nrs=0.15 nrd=0.11 
m1001 342 341 1 1 penh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=2.197e-11 ps=1.657e-05 pd=2.767e-05 
+ nrs=0.11 nrd=0.15 
m1002 1 341 342 1 penh l=8e-07 w=1.2e-05 
+ as=2.197e-11 ad=1.54e-11 ps=2.767e-05 pd=1.657e-05 
+ nrs=0.15 nrd=0.11 
m1003 342 341 1 1 penh l=8e-07 w=1.2e-05 
+ as=1.54e-11 ad=2.197e-11 ps=1.657e-05 pd=2.767e-05 
+ nrs=0.11 nrd=0.15 
m1004 0 343 294 0 nenh l=8e-07 w=4e-06 
+ as=3.744e-11 ad=8.8e-12 ps=1.807e-05 pd=1.368e-05 
+ nrs=2.34 nrd=0.55 
m1005 343 344 0 0 nenh l=1.6e-06 w=4e-06 
+ as=8.8e-12 ad=3.744e-11 ps=1.24e-05 pd=1.807e-05 
+ nrs=0.55 nrd=2.34 
m1006 1 343 294 1 penh l=8e-07 w=4e-06 
+ as=7.32e-12 ad=8.8e-12 ps=9.22e-06 pd=1.368e-05 
+ nrs=0.46 nrd=0.55 
m1007 343 344 1 1 penh l=1.6e-06 w=4e-06 
+ as=8.8e-12 ad=7.32e-12 ps=1.24e-05 pd=9.22e-06 
+ nrs=0.55 nrd=0.46 
c0 344 0 6.57e-13
c1 285 0 9.11e-13
c2 208 0 9.73e-13
c3 295 0 8.91e-13
c4 297 0 8.2e-13
c5 299 0 7.51e-13
c6 342 0 5.25e-13
c7 300 0 7.51e-13
c8 219 0 8.13e-13
c9 224 0 8.38e-13
c10 340 0 6.57e-13
c11 17 0 1.369e-12
c12 21 0 6.66e-13
c13 338 0 5.25e-13
c14 1 0 3.379e-12
c15 11 0 1.336e-12
c16 8 0 1.435e-12
c21 294 0 5.95e-13
c22 1 0 7.851e-12
c23 0 0 6.046e-12
c24 1 1 1.83e-13
c25 0 1 3.487e-12
c26 0 4 2.549e-12
c27 0 55 7.77e-13
VQ1H 285 0 pwl (0 0 2.6e-08 0 2.9e-08 3 4.9e-08 3 
+ 5.2e-08 0 7.8e-08 0 8.1e-08 3 1.01e-07 3 
+ 1.04e-07 0 1.3e-07 0 1.33e-07 3 1.53e-07 3 
+ 1.56e-07 0 1.82e-07 0 1.85e-07 3 2.05e-07 3 
+ 2.08e-07 0 2.34e-07 0 2.37e-07 3 2.57e-07 3 
+ 2.6e-07 0 2.86e-07 0 2.89e-07 3 3.09e-07 3 
+ 3.12e-07 0 3.38e-07 0 3.41e-07 3 3.61e-07 3 
+ 3.64e-07 0 3.9e-07 0 3.93e-07 3 4.13e-07 3 
+ 4.16e-07 0 4.42e-07 0 4.45e-07 3 4.65e-07 3 
+ 4.68e-07 0 4.94e-07 0 4.97e-07 3 5.17e-07 3 
+ 5.2e-07 0 5.46e-07 0 5.49e-07 3 5.69e-07 3 
+ 5.72e-07 0 5.98e-07 0 6.01e-07 3 6.21e-07 3 
+ 6.24e-07 0 6.5e-07 0 6.53e-07 3 6.73e-07 3 
+ 6.76e-07 0 7.02e-07 0 7.05e-07 3 7.25e-07 3 
+ 7.28e-07 0 7.54e-07 0 7.57e-07 3 7.77e-07 3 
+ 7.8e-07 0 8.06e-07 0 8.09e-07 3 8.29e-07 3 
+ 8.32e-07 0 8.58e-07 0 8.61e-07 3 8.81e-07 3 
+ 8.84e-07 0 9.1e-07 0 9.13e-07 3 9.33e-07 3 
+ 9.36e-07 0 9.62e-07 0 9.65e-07 3 9.85e-07 3 
+ 9.88e-07 0 1.014e-06 0 1.017e-06 3 1.037e-06 3 
+ 1.04e-06 0 1.066e-06 0 1.069e-06 3 1.089e-06 3 
+ 1.092e-06 0 1.118e-06 0 1.121e-06 3 1.141e-06 3 
+ 1.144e-06 0 1.17e-06 0 1.173e-06 3 1.193e-06 3 
+ 1.196e-06 0 1.222e-06 0 1.225e-06 3 1.245e-06 3 
+ 1.248e-06 0 1.274e-06 0 1.277e-06 3 1.297e-06 3 
+ 1.3e-06 0 1.326e-06 0 1.329e-06 3 1.349e-06 3 
+ 1.352e-06 0 1.378e-06 0 1.381e-06 3 1.401e-06 3 
+ 1.404e-06 0 1.43e-06 0 1.433e-06 3 1.453e-06 3 
+ 1.456e-06 0 1.482e-06 0 1.485e-06 3 1.505e-06 3 
+ 1.508e-06 0 1.534e-06 0 1.537e-06 3 1.557e-06 3 
+ 1.56e-06 0 1.586e-06 0 1.589e-06 3 1.609e-06 3 
+ 1.612e-06 0 1.638e-06 0 1.641e-06 3 1.661e-06 3 
+ 1.664e-06 0 1.69e-06 0 1.693e-06 3 1.713e-06 3 
+ 1.716e-06 0 1.742e-06 0 1.745e-06 3 1.765e-06 3 
+ 1.768e-06 0 1.794e-06 0 1.797e-06 3 1.817e-06 3 
+ 1.82e-06 0 1.846e-06 0 1.849e-06 3 1.869e-06 3 
+ 1.872e-06 0 1.898e-06 0 1.901e-06 3 1.921e-06 3 
+ 1.924e-06 0 1.95e-06 0 1.953e-06 3 1.973e-06 3 
+ 1.976e-06 0 2.002e-06 0 2.005e-06 3 2.025e-06 3 
+ 2.028e-06 0 2.054e-06 0 2.057e-06 3 2.077e-06 3 
+ 2.08e-06 0 2.106e-06 0 2.109e-06 3 2.129e-06 3 
+ 2.132e-06 0 2.158e-06 0 2.161e-06 3 2.181e-06 3 
+ 2.184e-06 0 2.21e-06 0 2.213e-06 3 2.233e-06 3 
+ 2.236e-06 0 2.262e-06 0 2.265e-06 3 2.285e-06 3 
+ 2.288e-06 0 2.314e-06 0 2.317e-06 3 2.337e-06 3 
+ 2.34e-06 0 2.366e-06 0 2.369e-06 3 2.389e-06 3 
+ 2.392e-06 0 2.418e-06 0 2.421e-06 3 2.441e-06 3 
+ 2.444e-06 0 2.47e-06 0 2.473e-06 3 2.493e-06 3 
+ 2.496e-06 0 2.522e-06 0 2.525e-06 3 2.545e-06 3 
+ 2.548e-06 0 2.574e-06 0 2.577e-06 3 2.597e-06 3 
+ 2.6e-06 0 2.626e-06 0 2.629e-06 3 2.649e-06 3 
+ 2.652e-06 0 2.678e-06 0 2.681e-06 3 2.701e-06 3 
+ 2.704e-06 0 2.73e-06 0 2.733e-06 3 2.753e-06 3 
+ 2.756e-06 0 2.782e-06 0 2.785e-06 3 2.805e-06 3 
+ 2.808e-06 0 2.834e-06 0 2.837e-06 3 2.857e-06 3 
+ 2.86e-06 0 2.886e-06 0 2.889e-06 3 2.909e-06 3 
+ 2.912e-06 0 2.938e-06 0 2.941e-06 3 2.961e-06 3 
+ 2.964e-06 0 2.99e-06 0 2.993e-06 3 3.013e-06 3 
+ 3.016e-06 0 3.042e-06 0 3.045e-06 3 3.065e-06 3 
+ 3.068e-06 0 3.094e-06 0 3.097e-06 3 3.117e-06 3 
+ 3.12e-06 0 3.146e-06 0 3.149e-06 3 3.169e-06 3 
+ 3.172e-06 0 3.198e-06 0 3.201e-06 3 3.221e-06 3 
+ 3.224e-06 0 3.25e-06 0 3.253e-06 3 3.273e-06 3 
+ 3.276e-06 0 3.302e-06 0 3.305e-06 3 3.325e-06 3 
+ 3.328e-06 0 3.354e-06 0 3.357e-06 3 3.377e-06 3 
+ 3.38e-06 0 3.406e-06 0 3.409e-06 3 3.429e-06 3 
+ 3.432e-06 0 3.458e-06 0 3.461e-06 3 3.481e-06 3 
+ 3.484e-06 0 3.51e-06 0 3.513e-06 3 3.533e-06 3 
+ 3.536e-06 0 3.562e-06 0 3.565e-06 3 3.585e-06 3 
+ 3.588e-06 0 3.614e-06 0 3.617e-06 3 3.637e-06 3 
+ 3.64e-06 0 3.666e-06 0 3.669e-06 3 3.689e-06 3 
+ 3.692e-06 0 3.718e-06 0 3.721e-06 3 3.741e-06 3 
+ 3.744e-06 0 3.77e-06 0 3.773e-06 3 3.793e-06 3 
+ 3.796e-06 0 3.822e-06 0 3.825e-06 3 3.845e-06 3 
+ 3.848e-06 0 3.874e-06 0 3.877e-06 3 3.897e-06 3 
+ 3.9e-06 0 3.926e-06 0 3.929e-06 3 3.949e-06 3 
+ 3.952e-06 0 3.978e-06 0 3.981e-06 3 4.001e-06 3 
+ 4.004e-06 0 4.03e-06 0 4.033e-06 3 4.053e-06 3 
+ 4.056e-06 0 4.082e-06 0 4.085e-06 3 4.105e-06 3 
+ 4.108e-06 0 4.134e-06 0 4.137e-06 3 4.157e-06 3 
+ 4.16e-06 0 4.186e-06 0 4.189e-06 3 4.209e-06 3 
+ 4.212e-06 0 4.238e-06 0 4.241e-06 3 4.261e-06 3 
+ 4.264e-06 0 4.29e-06 0 4.293e-06 3 4.313e-06 3 
+ 4.316e-06 0 4.342e-06 0 4.345e-06 3 4.365e-06 3 
+ 4.368e-06 0 4.394e-06 0 4.397e-06 3 4.417e-06 3 
+ 4.42e-06 0 4.446e-06 0 4.449e-06 3 4.469e-06 3 
+ 4.472e-06 0 4.498e-06 0 4.501e-06 3 4.521e-06 3 
+ 4.524e-06 0 4.55e-06 0 4.553e-06 3 4.573e-06 3 
+ 4.576e-06 0 4.602e-06 0 4.605e-06 3 4.625e-06 3 
+ 4.628e-06 0 4.654e-06 0 4.657e-06 3 4.677e-06 3 
+ 4.68e-06 0 4.706e-06 0 4.709e-06 3 4.729e-06 3 
+ 4.732e-06 0 4.758e-06 0 4.761e-06 3 4.781e-06 3 
+ 4.784e-06 0 4.81e-06 0 4.813e-06 3 4.833e-06 3 
+ 4.836e-06 0 4.862e-06 0 4.865e-06 3 4.885e-06 3 
+ 4.888e-06 0 4.914e-06 0 4.917e-06 3 4.937e-06 3 
+ 4.94e-06 0 4.966e-06 0 4.969e-06 3 4.989e-06 3 
+ 4.992e-06 0 5.018e-06 0 5.021e-06 3 5.041e-06 3 
+ 5.044e-06 0 5.07e-06 0 5.073e-06 3 5.093e-06 3 
+ 5.096e-06 0 5.122e-06 0 5.125e-06 3 5.145e-06 3 
+ 5.148e-06 0 5.174e-06 0 5.177e-06 3 5.197e-06 3 
+ 5.2e-06 0 5.226e-06 0 5.229e-06 3 5.249e-06 3 
+ 5.252e-06 0 5.278e-06 0 5.281e-06 3 5.301e-06 3 
+ 5.304e-06 0 5.33e-06 0 5.333e-06 3 5.353e-06 3 
+ 5.356e-06 0 5.382e-06 0 5.385e-06 3 5.405e-06 3 
+ 5.408e-06 0 5.434e-06 0 5.437e-06 3 5.457e-06 3 
+ 5.46e-06 0 5.486e-06 0 5.489e-06 3 5.509e-06 3 
+ 5.512e-06 0 5.538e-06 0 5.541e-06 3 5.561e-06 3 
+ 5.564e-06 0 5.59e-06 0 5.593e-06 3 5.613e-06 3 
+ 5.616e-06 0 5.642e-06 0 5.645e-06 3 5.665e-06 3 
+ 5.668e-06 0 5.694e-06 0 5.697e-06 3 5.717e-06 3 
+ 5.72e-06 0 5.746e-06 0 5.749e-06 3 5.769e-06 3 
+ 5.772e-06 0 5.798e-06 0 5.801e-06 3 5.821e-06 3 
+ 5.824e-06 0 5.85e-06 0 5.853e-06 3 5.873e-06 3 
+ 5.876e-06 0 5.902e-06 0 5.905e-06 3 5.925e-06 3 
+ 5.928e-06 0 5.954e-06 0 5.957e-06 3 5.977e-06 3 
+ 5.98e-06 0 6.006e-06 0 6.009e-06 3 6.029e-06 3 
+ 6.032e-06 0 6.058e-06 0 6.061e-06 3 6.081e-06 3 
+ 6.084e-06 0 6.11e-06 0 6.113e-06 3 6.133e-06 3 
+ 6.136e-06 0 6.162e-06 0 6.165e-06 3 6.185e-06 3 
+ 6.188e-06 0 6.214e-06 0 6.217e-06 3 6.237e-06 3 
+ 6.24e-06 0 6.266e-06 0 6.269e-06 3 6.289e-06 3 
+ 6.292e-06 0 6.318e-06 0 6.321e-06 3 6.341e-06 3 
+ 6.344e-06 0 6.37e-06 0 6.373e-06 3 6.393e-06 3 
+ 6.396e-06 0 6.422e-06 0 6.425e-06 3 6.445e-06 3 
+ 6.448e-06 0 6.474e-06 0 6.477e-06 3 6.497e-06 3 
+ 6.5e-06 0 )
VQ1L 208 0 pwl (0 3 2.6e-08 3 2.9e-08 0 4.9e-08 0 
+ 5.2e-08 3 7.8e-08 3 8.1e-08 0 1.01e-07 0 
+ 1.04e-07 3 1.3e-07 3 1.33e-07 0 1.53e-07 0 
+ 1.56e-07 3 1.82e-07 3 1.85e-07 0 2.05e-07 0 
+ 2.08e-07 3 2.34e-07 3 2.37e-07 0 2.57e-07 0 
+ 2.6e-07 3 2.86e-07 3 2.89e-07 0 3.09e-07 0 
+ 3.12e-07 3 3.38e-07 3 3.41e-07 0 3.61e-07 0 
+ 3.64e-07 3 3.9e-07 3 3.93e-07 0 4.13e-07 0 
+ 4.16e-07 3 4.42e-07 3 4.45e-07 0 4.65e-07 0 
+ 4.68e-07 3 4.94e-07 3 4.97e-07 0 5.17e-07 0 
+ 5.2e-07 3 5.46e-07 3 5.49e-07 0 5.69e-07 0 
+ 5.72e-07 3 5.98e-07 3 6.01e-07 0 6.21e-07 0 
+ 6.24e-07 3 6.5e-07 3 6.53e-07 0 6.73e-07 0 
+ 6.76e-07 3 7.02e-07 3 7.05e-07 0 7.25e-07 0 
+ 7.28e-07 3 7.54e-07 3 7.57e-07 0 7.77e-07 0 
+ 7.8e-07 3 8.06e-07 3 8.09e-07 0 8.29e-07 0 
+ 8.32e-07 3 8.58e-07 3 8.61e-07 0 8.81e-07 0 
+ 8.84e-07 3 9.1e-07 3 9.13e-07 0 9.33e-07 0 
+ 9.36e-07 3 9.62e-07 3 9.65e-07 0 9.85e-07 0 
+ 9.88e-07 3 1.014e-06 3 1.017e-06 0 1.037e-06 0 
+ 1.04e-06 3 1.066e-06 3 1.069e-06 0 1.089e-06 0 
+ 1.092e-06 3 1.118e-06 3 1.121e-06 0 1.141e-06 0 
+ 1.144e-06 3 1.17e-06 3 1.173e-06 0 1.193e-06 0 
+ 1.196e-06 3 1.222e-06 3 1.225e-06 0 1.245e-06 0 
+ 1.248e-06 3 1.274e-06 3 1.277e-06 0 1.297e-06 0 
+ 1.3e-06 3 1.326e-06 3 1.329e-06 0 1.349e-06 0 
+ 1.352e-06 3 1.378e-06 3 1.381e-06 0 1.401e-06 0 
+ 1.404e-06 3 1.43e-06 3 1.433e-06 0 1.453e-06 0 
+ 1.456e-06 3 1.482e-06 3 1.485e-06 0 1.505e-06 0 
+ 1.508e-06 3 1.534e-06 3 1.537e-06 0 1.557e-06 0 
+ 1.56e-06 3 1.586e-06 3 1.589e-06 0 1.609e-06 0 
+ 1.612e-06 3 1.638e-06 3 1.641e-06 0 1.661e-06 0 
+ 1.664e-06 3 1.69e-06 3 1.693e-06 0 1.713e-06 0 
+ 1.716e-06 3 1.742e-06 3 1.745e-06 0 1.765e-06 0 
+ 1.768e-06 3 1.794e-06 3 1.797e-06 0 1.817e-06 0 
+ 1.82e-06 3 1.846e-06 3 1.849e-06 0 1.869e-06 0 
+ 1.872e-06 3 1.898e-06 3 1.901e-06 0 1.921e-06 0 
+ 1.924e-06 3 1.95e-06 3 1.953e-06 0 1.973e-06 0 
+ 1.976e-06 3 2.002e-06 3 2.005e-06 0 2.025e-06 0 
+ 2.028e-06 3 2.054e-06 3 2.057e-06 0 2.077e-06 0 
+ 2.08e-06 3 2.106e-06 3 2.109e-06 0 2.129e-06 0 
+ 2.132e-06 3 2.158e-06 3 2.161e-06 0 2.181e-06 0 
+ 2.184e-06 3 2.21e-06 3 2.213e-06 0 2.233e-06 0 
+ 2.236e-06 3 2.262e-06 3 2.265e-06 0 2.285e-06 0 
+ 2.288e-06 3 2.314e-06 3 2.317e-06 0 2.337e-06 0 
+ 2.34e-06 3 2.366e-06 3 2.369e-06 0 2.389e-06 0 
+ 2.392e-06 3 2.418e-06 3 2.421e-06 0 2.441e-06 0 
+ 2.444e-06 3 2.47e-06 3 2.473e-06 0 2.493e-06 0 
+ 2.496e-06 3 2.522e-06 3 2.525e-06 0 2.545e-06 0 
+ 2.548e-06 3 2.574e-06 3 2.577e-06 0 2.597e-06 0 
+ 2.6e-06 3 2.626e-06 3 2.629e-06 0 2.649e-06 0 
+ 2.652e-06 3 2.678e-06 3 2.681e-06 0 2.701e-06 0 
+ 2.704e-06 3 2.73e-06 3 2.733e-06 0 2.753e-06 0 
+ 2.756e-06 3 2.782e-06 3 2.785e-06 0 2.805e-06 0 
+ 2.808e-06 3 2.834e-06 3 2.837e-06 0 2.857e-06 0 
+ 2.86e-06 3 2.886e-06 3 2.889e-06 0 2.909e-06 0 
+ 2.912e-06 3 2.938e-06 3 2.941e-06 0 2.961e-06 0 
+ 2.964e-06 3 2.99e-06 3 2.993e-06 0 3.013e-06 0 
+ 3.016e-06 3 3.042e-06 3 3.045e-06 0 3.065e-06 0 
+ 3.068e-06 3 3.094e-06 3 3.097e-06 0 3.117e-06 0 
+ 3.12e-06 3 3.146e-06 3 3.149e-06 0 3.169e-06 0 
+ 3.172e-06 3 3.198e-06 3 3.201e-06 0 3.221e-06 0 
+ 3.224e-06 3 3.25e-06 3 3.253e-06 0 3.273e-06 0 
+ 3.276e-06 3 3.302e-06 3 3.305e-06 0 3.325e-06 0 
+ 3.328e-06 3 3.354e-06 3 3.357e-06 0 3.377e-06 0 
+ 3.38e-06 3 3.406e-06 3 3.409e-06 0 3.429e-06 0 
+ 3.432e-06 3 3.458e-06 3 3.461e-06 0 3.481e-06 0 
+ 3.484e-06 3 3.51e-06 3 3.513e-06 0 3.533e-06 0 
+ 3.536e-06 3 3.562e-06 3 3.565e-06 0 3.585e-06 0 
+ 3.588e-06 3 3.614e-06 3 3.617e-06 0 3.637e-06 0 
+ 3.64e-06 3 3.666e-06 3 3.669e-06 0 3.689e-06 0 
+ 3.692e-06 3 3.718e-06 3 3.721e-06 0 3.741e-06 0 
+ 3.744e-06 3 3.77e-06 3 3.773e-06 0 3.793e-06 0 
+ 3.796e-06 3 3.822e-06 3 3.825e-06 0 3.845e-06 0 
+ 3.848e-06 3 3.874e-06 3 3.877e-06 0 3.897e-06 0 
+ 3.9e-06 3 3.926e-06 3 3.929e-06 0 3.949e-06 0 
+ 3.952e-06 3 3.978e-06 3 3.981e-06 0 4.001e-06 0 
+ 4.004e-06 3 4.03e-06 3 4.033e-06 0 4.053e-06 0 
+ 4.056e-06 3 4.082e-06 3 4.085e-06 0 4.105e-06 0 
+ 4.108e-06 3 4.134e-06 3 4.137e-06 0 4.157e-06 0 
+ 4.16e-06 3 4.186e-06 3 4.189e-06 0 4.209e-06 0 
+ 4.212e-06 3 4.238e-06 3 4.241e-06 0 4.261e-06 0 
+ 4.264e-06 3 4.29e-06 3 4.293e-06 0 4.313e-06 0 
+ 4.316e-06 3 4.342e-06 3 4.345e-06 0 4.365e-06 0 
+ 4.368e-06 3 4.394e-06 3 4.397e-06 0 4.417e-06 0 
+ 4.42e-06 3 4.446e-06 3 4.449e-06 0 4.469e-06 0 
+ 4.472e-06 3 4.498e-06 3 4.501e-06 0 4.521e-06 0 
+ 4.524e-06 3 4.55e-06 3 4.553e-06 0 4.573e-06 0 
+ 4.576e-06 3 4.602e-06 3 4.605e-06 0 4.625e-06 0 
+ 4.628e-06 3 4.654e-06 3 4.657e-06 0 4.677e-06 0 
+ 4.68e-06 3 4.706e-06 3 4.709e-06 0 4.729e-06 0 
+ 4.732e-06 3 4.758e-06 3 4.761e-06 0 4.781e-06 0 
+ 4.784e-06 3 4.81e-06 3 4.813e-06 0 4.833e-06 0 
+ 4.836e-06 3 4.862e-06 3 4.865e-06 0 4.885e-06 0 
+ 4.888e-06 3 4.914e-06 3 4.917e-06 0 4.937e-06 0 
+ 4.94e-06 3 4.966e-06 3 4.969e-06 0 4.989e-06 0 
+ 4.992e-06 3 5.018e-06 3 5.021e-06 0 5.041e-06 0 
+ 5.044e-06 3 5.07e-06 3 5.073e-06 0 5.093e-06 0 
+ 5.096e-06 3 5.122e-06 3 5.125e-06 0 5.145e-06 0 
+ 5.148e-06 3 5.174e-06 3 5.177e-06 0 5.197e-06 0 
+ 5.2e-06 3 5.226e-06 3 5.229e-06 0 5.249e-06 0 
+ 5.252e-06 3 5.278e-06 3 5.281e-06 0 5.301e-06 0 
+ 5.304e-06 3 5.33e-06 3 5.333e-06 0 5.353e-06 0 
+ 5.356e-06 3 5.382e-06 3 5.385e-06 0 5.405e-06 0 
+ 5.408e-06 3 5.434e-06 3 5.437e-06 0 5.457e-06 0 
+ 5.46e-06 3 5.486e-06 3 5.489e-06 0 5.509e-06 0 
+ 5.512e-06 3 5.538e-06 3 5.541e-06 0 5.561e-06 0 
+ 5.564e-06 3 5.59e-06 3 5.593e-06 0 5.613e-06 0 
+ 5.616e-06 3 5.642e-06 3 5.645e-06 0 5.665e-06 0 
+ 5.668e-06 3 5.694e-06 3 5.697e-06 0 5.717e-06 0 
+ 5.72e-06 3 5.746e-06 3 5.749e-06 0 5.769e-06 0 
+ 5.772e-06 3 5.798e-06 3 5.801e-06 0 5.821e-06 0 
+ 5.824e-06 3 5.85e-06 3 5.853e-06 0 5.873e-06 0 
+ 5.876e-06 3 5.902e-06 3 5.905e-06 0 5.925e-06 0 
+ 5.928e-06 3 5.954e-06 3 5.957e-06 0 5.977e-06 0 
+ 5.98e-06 3 6.006e-06 3 6.009e-06 0 6.029e-06 0 
+ 6.032e-06 3 6.058e-06 3 6.061e-06 0 6.081e-06 0 
+ 6.084e-06 3 6.11e-06 3 6.113e-06 0 6.133e-06 0 
+ 6.136e-06 3 6.162e-06 3 6.165e-06 0 6.185e-06 0 
+ 6.188e-06 3 6.214e-06 3 6.217e-06 0 6.237e-06 0 
+ 6.24e-06 3 6.266e-06 3 6.269e-06 0 6.289e-06 0 
+ 6.292e-06 3 6.318e-06 3 6.321e-06 0 6.341e-06 0 
+ 6.344e-06 3 6.37e-06 3 6.373e-06 0 6.393e-06 0 
+ 6.396e-06 3 6.422e-06 3 6.425e-06 0 6.445e-06 0 
+ 6.448e-06 3 6.474e-06 3 6.477e-06 0 6.497e-06 0 
+ 6.5e-06 3 )
VQ2H 4 0 pwl (0 0 5.2e-08 0 5.5e-08 3 7.5e-08 3 
+ 7.8e-08 0 1.04e-07 0 1.07e-07 3 1.27e-07 3 
+ 1.3e-07 0 1.56e-07 0 1.59e-07 3 1.79e-07 3 
+ 1.82e-07 0 2.08e-07 0 2.11e-07 3 2.31e-07 3 
+ 2.34e-07 0 2.6e-07 0 2.63e-07 3 2.83e-07 3 
+ 2.86e-07 0 3.12e-07 0 3.15e-07 3 3.35e-07 3 
+ 3.38e-07 0 3.64e-07 0 3.67e-07 3 3.87e-07 3 
+ 3.9e-07 0 4.16e-07 0 4.19e-07 3 4.39e-07 3 
+ 4.42e-07 0 4.68e-07 0 4.71e-07 3 4.91e-07 3 
+ 4.94e-07 0 5.2e-07 0 5.23e-07 3 5.43e-07 3 
+ 5.46e-07 0 5.72e-07 0 5.75e-07 3 5.95e-07 3 
+ 5.98e-07 0 6.24e-07 0 6.27e-07 3 6.47e-07 3 
+ 6.5e-07 0 6.76e-07 0 6.79e-07 3 6.99e-07 3 
+ 7.02e-07 0 7.28e-07 0 7.31e-07 3 7.51e-07 3 
+ 7.54e-07 0 7.8e-07 0 7.83e-07 3 8.03e-07 3 
+ 8.06e-07 0 8.32e-07 0 8.35e-07 3 8.55e-07 3 
+ 8.58e-07 0 8.84e-07 0 8.87e-07 3 9.07e-07 3 
+ 9.1e-07 0 9.36e-07 0 9.39e-07 3 9.59e-07 3 
+ 9.62e-07 0 9.88e-07 0 9.91e-07 3 1.011e-06 3 
+ 1.014e-06 0 1.04e-06 0 1.043e-06 3 1.063e-06 3 
+ 1.066e-06 0 1.092e-06 0 1.095e-06 3 1.115e-06 3 
+ 1.118e-06 0 1.144e-06 0 1.147e-06 3 1.167e-06 3 
+ 1.17e-06 0 1.196e-06 0 1.199e-06 3 1.219e-06 3 
+ 1.222e-06 0 1.248e-06 0 1.251e-06 3 1.271e-06 3 
+ 1.274e-06 0 1.3e-06 0 1.303e-06 3 1.323e-06 3 
+ 1.326e-06 0 1.352e-06 0 1.355e-06 3 1.375e-06 3 
+ 1.378e-06 0 1.404e-06 0 1.407e-06 3 1.427e-06 3 
+ 1.43e-06 0 1.456e-06 0 1.459e-06 3 1.479e-06 3 
+ 1.482e-06 0 1.508e-06 0 1.511e-06 3 1.531e-06 3 
+ 1.534e-06 0 1.56e-06 0 1.563e-06 3 1.583e-06 3 
+ 1.586e-06 0 1.612e-06 0 1.615e-06 3 1.635e-06 3 
+ 1.638e-06 0 1.664e-06 0 1.667e-06 3 1.687e-06 3 
+ 1.69e-06 0 1.716e-06 0 1.719e-06 3 1.739e-06 3 
+ 1.742e-06 0 1.768e-06 0 1.771e-06 3 1.791e-06 3 
+ 1.794e-06 0 1.82e-06 0 1.823e-06 3 1.843e-06 3 
+ 1.846e-06 0 1.872e-06 0 1.875e-06 3 1.895e-06 3 
+ 1.898e-06 0 1.924e-06 0 1.927e-06 3 1.947e-06 3 
+ 1.95e-06 0 1.976e-06 0 1.979e-06 3 1.999e-06 3 
+ 2.002e-06 0 2.028e-06 0 2.031e-06 3 2.051e-06 3 
+ 2.054e-06 0 2.08e-06 0 2.083e-06 3 2.103e-06 3 
+ 2.106e-06 0 2.132e-06 0 2.135e-06 3 2.155e-06 3 
+ 2.158e-06 0 2.184e-06 0 2.187e-06 3 2.207e-06 3 
+ 2.21e-06 0 2.236e-06 0 2.239e-06 3 2.259e-06 3 
+ 2.262e-06 0 2.288e-06 0 2.291e-06 3 2.311e-06 3 
+ 2.314e-06 0 2.34e-06 0 2.343e-06 3 2.363e-06 3 
+ 2.366e-06 0 2.392e-06 0 2.395e-06 3 2.415e-06 3 
+ 2.418e-06 0 2.444e-06 0 2.447e-06 3 2.467e-06 3 
+ 2.47e-06 0 2.496e-06 0 2.499e-06 3 2.519e-06 3 
+ 2.522e-06 0 2.548e-06 0 2.551e-06 3 2.571e-06 3 
+ 2.574e-06 0 2.6e-06 0 2.603e-06 3 2.623e-06 3 
+ 2.626e-06 0 2.652e-06 0 2.655e-06 3 2.675e-06 3 
+ 2.678e-06 0 2.704e-06 0 2.707e-06 3 2.727e-06 3 
+ 2.73e-06 0 2.756e-06 0 2.759e-06 3 2.779e-06 3 
+ 2.782e-06 0 2.808e-06 0 2.811e-06 3 2.831e-06 3 
+ 2.834e-06 0 2.86e-06 0 2.863e-06 3 2.883e-06 3 
+ 2.886e-06 0 2.912e-06 0 2.915e-06 3 2.935e-06 3 
+ 2.938e-06 0 2.964e-06 0 2.967e-06 3 2.987e-06 3 
+ 2.99e-06 0 3.016e-06 0 3.019e-06 3 3.039e-06 3 
+ 3.042e-06 0 3.068e-06 0 3.071e-06 3 3.091e-06 3 
+ 3.094e-06 0 3.12e-06 0 3.123e-06 3 3.143e-06 3 
+ 3.146e-06 0 3.172e-06 0 3.175e-06 3 3.195e-06 3 
+ 3.198e-06 0 3.224e-06 0 3.227e-06 3 3.247e-06 3 
+ 3.25e-06 0 3.276e-06 0 3.279e-06 3 3.299e-06 3 
+ 3.302e-06 0 3.328e-06 0 3.331e-06 3 3.351e-06 3 
+ 3.354e-06 0 3.38e-06 0 3.383e-06 3 3.403e-06 3 
+ 3.406e-06 0 3.432e-06 0 3.435e-06 3 3.455e-06 3 
+ 3.458e-06 0 3.484e-06 0 3.487e-06 3 3.507e-06 3 
+ 3.51e-06 0 3.536e-06 0 3.539e-06 3 3.559e-06 3 
+ 3.562e-06 0 3.588e-06 0 3.591e-06 3 3.611e-06 3 
+ 3.614e-06 0 3.64e-06 0 3.643e-06 3 3.663e-06 3 
+ 3.666e-06 0 3.692e-06 0 3.695e-06 3 3.715e-06 3 
+ 3.718e-06 0 3.744e-06 0 3.747e-06 3 3.767e-06 3 
+ 3.77e-06 0 3.796e-06 0 3.799e-06 3 3.819e-06 3 
+ 3.822e-06 0 3.848e-06 0 3.851e-06 3 3.871e-06 3 
+ 3.874e-06 0 3.9e-06 0 3.903e-06 3 3.923e-06 3 
+ 3.926e-06 0 3.952e-06 0 3.955e-06 3 3.975e-06 3 
+ 3.978e-06 0 4.004e-06 0 4.007e-06 3 4.027e-06 3 
+ 4.03e-06 0 4.056e-06 0 4.059e-06 3 4.079e-06 3 
+ 4.082e-06 0 4.108e-06 0 4.111e-06 3 4.131e-06 3 
+ 4.134e-06 0 4.16e-06 0 4.163e-06 3 4.183e-06 3 
+ 4.186e-06 0 4.212e-06 0 4.215e-06 3 4.235e-06 3 
+ 4.238e-06 0 4.264e-06 0 4.267e-06 3 4.287e-06 3 
+ 4.29e-06 0 4.316e-06 0 4.319e-06 3 4.339e-06 3 
+ 4.342e-06 0 4.368e-06 0 4.371e-06 3 4.391e-06 3 
+ 4.394e-06 0 4.42e-06 0 4.423e-06 3 4.443e-06 3 
+ 4.446e-06 0 4.472e-06 0 4.475e-06 3 4.495e-06 3 
+ 4.498e-06 0 4.524e-06 0 4.527e-06 3 4.547e-06 3 
+ 4.55e-06 0 4.576e-06 0 4.579e-06 3 4.599e-06 3 
+ 4.602e-06 0 4.628e-06 0 4.631e-06 3 4.651e-06 3 
+ 4.654e-06 0 4.68e-06 0 4.683e-06 3 4.703e-06 3 
+ 4.706e-06 0 4.732e-06 0 4.735e-06 3 4.755e-06 3 
+ 4.758e-06 0 4.784e-06 0 4.787e-06 3 4.807e-06 3 
+ 4.81e-06 0 4.836e-06 0 4.839e-06 3 4.859e-06 3 
+ 4.862e-06 0 4.888e-06 0 4.891e-06 3 4.911e-06 3 
+ 4.914e-06 0 4.94e-06 0 4.943e-06 3 4.963e-06 3 
+ 4.966e-06 0 4.992e-06 0 4.995e-06 3 5.015e-06 3 
+ 5.018e-06 0 5.044e-06 0 5.047e-06 3 5.067e-06 3 
+ 5.07e-06 0 5.096e-06 0 5.099e-06 3 5.119e-06 3 
+ 5.122e-06 0 5.148e-06 0 5.151e-06 3 5.171e-06 3 
+ 5.174e-06 0 5.2e-06 0 5.203e-06 3 5.223e-06 3 
+ 5.226e-06 0 5.252e-06 0 5.255e-06 3 5.275e-06 3 
+ 5.278e-06 0 5.304e-06 0 5.307e-06 3 5.327e-06 3 
+ 5.33e-06 0 5.356e-06 0 5.359e-06 3 5.379e-06 3 
+ 5.382e-06 0 5.408e-06 0 5.411e-06 3 5.431e-06 3 
+ 5.434e-06 0 5.46e-06 0 5.463e-06 3 5.483e-06 3 
+ 5.486e-06 0 5.512e-06 0 5.515e-06 3 5.535e-06 3 
+ 5.538e-06 0 5.564e-06 0 5.567e-06 3 5.587e-06 3 
+ 5.59e-06 0 5.616e-06 0 5.619e-06 3 5.639e-06 3 
+ 5.642e-06 0 5.668e-06 0 5.671e-06 3 5.691e-06 3 
+ 5.694e-06 0 5.72e-06 0 5.723e-06 3 5.743e-06 3 
+ 5.746e-06 0 5.772e-06 0 5.775e-06 3 5.795e-06 3 
+ 5.798e-06 0 5.824e-06 0 5.827e-06 3 5.847e-06 3 
+ 5.85e-06 0 5.876e-06 0 5.879e-06 3 5.899e-06 3 
+ 5.902e-06 0 5.928e-06 0 5.931e-06 3 5.951e-06 3 
+ 5.954e-06 0 5.98e-06 0 5.983e-06 3 6.003e-06 3 
+ 6.006e-06 0 6.032e-06 0 6.035e-06 3 6.055e-06 3 
+ 6.058e-06 0 6.084e-06 0 6.087e-06 3 6.107e-06 3 
+ 6.11e-06 0 6.136e-06 0 6.139e-06 3 6.159e-06 3 
+ 6.162e-06 0 6.188e-06 0 6.191e-06 3 6.211e-06 3 
+ 6.214e-06 0 6.24e-06 0 6.243e-06 3 6.263e-06 3 
+ 6.266e-06 0 6.292e-06 0 6.295e-06 3 6.315e-06 3 
+ 6.318e-06 0 6.344e-06 0 6.347e-06 3 6.367e-06 3 
+ 6.37e-06 0 6.396e-06 0 6.399e-06 3 6.419e-06 3 
+ 6.422e-06 0 6.448e-06 0 6.451e-06 3 6.471e-06 3 
+ 6.474e-06 0 6.5e-06 0 )
VQ2L 8 0 pwl (0 3 5.2e-08 3 5.5e-08 0 7.5e-08 0 
+ 7.8e-08 3 1.04e-07 3 1.07e-07 0 1.27e-07 0 
+ 1.3e-07 3 1.56e-07 3 1.59e-07 0 1.79e-07 0 
+ 1.82e-07 3 2.08e-07 3 2.11e-07 0 2.31e-07 0 
+ 2.34e-07 3 2.6e-07 3 2.63e-07 0 2.83e-07 0 
+ 2.86e-07 3 3.12e-07 3 3.15e-07 0 3.35e-07 0 
+ 3.38e-07 3 3.64e-07 3 3.67e-07 0 3.87e-07 0 
+ 3.9e-07 3 4.16e-07 3 4.19e-07 0 4.39e-07 0 
+ 4.42e-07 3 4.68e-07 3 4.71e-07 0 4.91e-07 0 
+ 4.94e-07 3 5.2e-07 3 5.23e-07 0 5.43e-07 0 
+ 5.46e-07 3 5.72e-07 3 5.75e-07 0 5.95e-07 0 
+ 5.98e-07 3 6.24e-07 3 6.27e-07 0 6.47e-07 0 
+ 6.5e-07 3 6.76e-07 3 6.79e-07 0 6.99e-07 0 
+ 7.02e-07 3 7.28e-07 3 7.31e-07 0 7.51e-07 0 
+ 7.54e-07 3 7.8e-07 3 7.83e-07 0 8.03e-07 0 
+ 8.06e-07 3 8.32e-07 3 8.35e-07 0 8.55e-07 0 
+ 8.58e-07 3 8.84e-07 3 8.87e-07 0 9.07e-07 0 
+ 9.1e-07 3 9.36e-07 3 9.39e-07 0 9.59e-07 0 
+ 9.62e-07 3 9.88e-07 3 9.91e-07 0 1.011e-06 0 
+ 1.014e-06 3 1.04e-06 3 1.043e-06 0 1.063e-06 0 
+ 1.066e-06 3 1.092e-06 3 1.095e-06 0 1.115e-06 0 
+ 1.118e-06 3 1.144e-06 3 1.147e-06 0 1.167e-06 0 
+ 1.17e-06 3 1.196e-06 3 1.199e-06 0 1.219e-06 0 
+ 1.222e-06 3 1.248e-06 3 1.251e-06 0 1.271e-06 0 
+ 1.274e-06 3 1.3e-06 3 1.303e-06 0 1.323e-06 0 
+ 1.326e-06 3 1.352e-06 3 1.355e-06 0 1.375e-06 0 
+ 1.378e-06 3 1.404e-06 3 1.407e-06 0 1.427e-06 0 
+ 1.43e-06 3 1.456e-06 3 1.459e-06 0 1.479e-06 0 
+ 1.482e-06 3 1.508e-06 3 1.511e-06 0 1.531e-06 0 
+ 1.534e-06 3 1.56e-06 3 1.563e-06 0 1.583e-06 0 
+ 1.586e-06 3 1.612e-06 3 1.615e-06 0 1.635e-06 0 
+ 1.638e-06 3 1.664e-06 3 1.667e-06 0 1.687e-06 0 
+ 1.69e-06 3 1.716e-06 3 1.719e-06 0 1.739e-06 0 
+ 1.742e-06 3 1.768e-06 3 1.771e-06 0 1.791e-06 0 
+ 1.794e-06 3 1.82e-06 3 1.823e-06 0 1.843e-06 0 
+ 1.846e-06 3 1.872e-06 3 1.875e-06 0 1.895e-06 0 
+ 1.898e-06 3 1.924e-06 3 1.927e-06 0 1.947e-06 0 
+ 1.95e-06 3 1.976e-06 3 1.979e-06 0 1.999e-06 0 
+ 2.002e-06 3 2.028e-06 3 2.031e-06 0 2.051e-06 0 
+ 2.054e-06 3 2.08e-06 3 2.083e-06 0 2.103e-06 0 
+ 2.106e-06 3 2.132e-06 3 2.135e-06 0 2.155e-06 0 
+ 2.158e-06 3 2.184e-06 3 2.187e-06 0 2.207e-06 0 
+ 2.21e-06 3 2.236e-06 3 2.239e-06 0 2.259e-06 0 
+ 2.262e-06 3 2.288e-06 3 2.291e-06 0 2.311e-06 0 
+ 2.314e-06 3 2.34e-06 3 2.343e-06 0 2.363e-06 0 
+ 2.366e-06 3 2.392e-06 3 2.395e-06 0 2.415e-06 0 
+ 2.418e-06 3 2.444e-06 3 2.447e-06 0 2.467e-06 0 
+ 2.47e-06 3 2.496e-06 3 2.499e-06 0 2.519e-06 0 
+ 2.522e-06 3 2.548e-06 3 2.551e-06 0 2.571e-06 0 
+ 2.574e-06 3 2.6e-06 3 2.603e-06 0 2.623e-06 0 
+ 2.626e-06 3 2.652e-06 3 2.655e-06 0 2.675e-06 0 
+ 2.678e-06 3 2.704e-06 3 2.707e-06 0 2.727e-06 0 
+ 2.73e-06 3 2.756e-06 3 2.759e-06 0 2.779e-06 0 
+ 2.782e-06 3 2.808e-06 3 2.811e-06 0 2.831e-06 0 
+ 2.834e-06 3 2.86e-06 3 2.863e-06 0 2.883e-06 0 
+ 2.886e-06 3 2.912e-06 3 2.915e-06 0 2.935e-06 0 
+ 2.938e-06 3 2.964e-06 3 2.967e-06 0 2.987e-06 0 
+ 2.99e-06 3 3.016e-06 3 3.019e-06 0 3.039e-06 0 
+ 3.042e-06 3 3.068e-06 3 3.071e-06 0 3.091e-06 0 
+ 3.094e-06 3 3.12e-06 3 3.123e-06 0 3.143e-06 0 
+ 3.146e-06 3 3.172e-06 3 3.175e-06 0 3.195e-06 0 
+ 3.198e-06 3 3.224e-06 3 3.227e-06 0 3.247e-06 0 
+ 3.25e-06 3 3.276e-06 3 3.279e-06 0 3.299e-06 0 
+ 3.302e-06 3 3.328e-06 3 3.331e-06 0 3.351e-06 0 
+ 3.354e-06 3 3.38e-06 3 3.383e-06 0 3.403e-06 0 
+ 3.406e-06 3 3.432e-06 3 3.435e-06 0 3.455e-06 0 
+ 3.458e-06 3 3.484e-06 3 3.487e-06 0 3.507e-06 0 
+ 3.51e-06 3 3.536e-06 3 3.539e-06 0 3.559e-06 0 
+ 3.562e-06 3 3.588e-06 3 3.591e-06 0 3.611e-06 0 
+ 3.614e-06 3 3.64e-06 3 3.643e-06 0 3.663e-06 0 
+ 3.666e-06 3 3.692e-06 3 3.695e-06 0 3.715e-06 0 
+ 3.718e-06 3 3.744e-06 3 3.747e-06 0 3.767e-06 0 
+ 3.77e-06 3 3.796e-06 3 3.799e-06 0 3.819e-06 0 
+ 3.822e-06 3 3.848e-06 3 3.851e-06 0 3.871e-06 0 
+ 3.874e-06 3 3.9e-06 3 3.903e-06 0 3.923e-06 0 
+ 3.926e-06 3 3.952e-06 3 3.955e-06 0 3.975e-06 0 
+ 3.978e-06 3 4.004e-06 3 4.007e-06 0 4.027e-06 0 
+ 4.03e-06 3 4.056e-06 3 4.059e-06 0 4.079e-06 0 
+ 4.082e-06 3 4.108e-06 3 4.111e-06 0 4.131e-06 0 
+ 4.134e-06 3 4.16e-06 3 4.163e-06 0 4.183e-06 0 
+ 4.186e-06 3 4.212e-06 3 4.215e-06 0 4.235e-06 0 
+ 4.238e-06 3 4.264e-06 3 4.267e-06 0 4.287e-06 0 
+ 4.29e-06 3 4.316e-06 3 4.319e-06 0 4.339e-06 0 
+ 4.342e-06 3 4.368e-06 3 4.371e-06 0 4.391e-06 0 
+ 4.394e-06 3 4.42e-06 3 4.423e-06 0 4.443e-06 0 
+ 4.446e-06 3 4.472e-06 3 4.475e-06 0 4.495e-06 0 
+ 4.498e-06 3 4.524e-06 3 4.527e-06 0 4.547e-06 0 
+ 4.55e-06 3 4.576e-06 3 4.579e-06 0 4.599e-06 0 
+ 4.602e-06 3 4.628e-06 3 4.631e-06 0 4.651e-06 0 
+ 4.654e-06 3 4.68e-06 3 4.683e-06 0 4.703e-06 0 
+ 4.706e-06 3 4.732e-06 3 4.735e-06 0 4.755e-06 0 
+ 4.758e-06 3 4.784e-06 3 4.787e-06 0 4.807e-06 0 
+ 4.81e-06 3 4.836e-06 3 4.839e-06 0 4.859e-06 0 
+ 4.862e-06 3 4.888e-06 3 4.891e-06 0 4.911e-06 0 
+ 4.914e-06 3 4.94e-06 3 4.943e-06 0 4.963e-06 0 
+ 4.966e-06 3 4.992e-06 3 4.995e-06 0 5.015e-06 0 
+ 5.018e-06 3 5.044e-06 3 5.047e-06 0 5.067e-06 0 
+ 5.07e-06 3 5.096e-06 3 5.099e-06 0 5.119e-06 0 
+ 5.122e-06 3 5.148e-06 3 5.151e-06 0 5.171e-06 0 
+ 5.174e-06 3 5.2e-06 3 5.203e-06 0 5.223e-06 0 
+ 5.226e-06 3 5.252e-06 3 5.255e-06 0 5.275e-06 0 
+ 5.278e-06 3 5.304e-06 3 5.307e-06 0 5.327e-06 0 
+ 5.33e-06 3 5.356e-06 3 5.359e-06 0 5.379e-06 0 
+ 5.382e-06 3 5.408e-06 3 5.411e-06 0 5.431e-06 0 
+ 5.434e-06 3 5.46e-06 3 5.463e-06 0 5.483e-06 0 
+ 5.486e-06 3 5.512e-06 3 5.515e-06 0 5.535e-06 0 
+ 5.538e-06 3 5.564e-06 3 5.567e-06 0 5.587e-06 0 
+ 5.59e-06 3 5.616e-06 3 5.619e-06 0 5.639e-06 0 
+ 5.642e-06 3 5.668e-06 3 5.671e-06 0 5.691e-06 0 
+ 5.694e-06 3 5.72e-06 3 5.723e-06 0 5.743e-06 0 
+ 5.746e-06 3 5.772e-06 3 5.775e-06 0 5.795e-06 0 
+ 5.798e-06 3 5.824e-06 3 5.827e-06 0 5.847e-06 0 
+ 5.85e-06 3 5.876e-06 3 5.879e-06 0 5.899e-06 0 
+ 5.902e-06 3 5.928e-06 3 5.931e-06 0 5.951e-06 0 
+ 5.954e-06 3 5.98e-06 3 5.983e-06 0 6.003e-06 0 
+ 6.006e-06 3 6.032e-06 3 6.035e-06 0 6.055e-06 0 
+ 6.058e-06 3 6.084e-06 3 6.087e-06 0 6.107e-06 0 
+ 6.11e-06 3 6.136e-06 3 6.139e-06 0 6.159e-06 0 
+ 6.162e-06 3 6.188e-06 3 6.191e-06 0 6.211e-06 0 
+ 6.214e-06 3 6.24e-06 3 6.243e-06 0 6.263e-06 0 
+ 6.266e-06 3 6.292e-06 3 6.295e-06 0 6.315e-06 0 
+ 6.318e-06 3 6.344e-06 3 6.347e-06 0 6.367e-06 0 
+ 6.37e-06 3 6.396e-06 3 6.399e-06 0 6.419e-06 0 
+ 6.422e-06 3 6.448e-06 3 6.451e-06 0 6.471e-06 0 
+ 6.474e-06 3 6.5e-06 3 )
VWriteH 219 0 pwl (0 0 4.68e-07 0 4.71e-07 3 4.91e-07 3 
+ 4.94e-07 0 5.72e-07 0 5.75e-07 3 5.95e-07 3 
+ 5.98e-07 0 6.76e-07 0 6.79e-07 3 6.99e-07 3 
+ 7.02e-07 0 7.8e-07 0 7.83e-07 3 8.03e-07 3 
+ 8.06e-07 0 8.84e-07 0 8.87e-07 3 9.07e-07 3 
+ 9.1e-07 0 9.88e-07 0 9.91e-07 3 1.011e-06 3 
+ 1.014e-06 0 1.092e-06 0 1.095e-06 3 1.115e-06 3 
+ 1.118e-06 0 1.196e-06 0 1.199e-06 3 1.219e-06 3 
+ 1.222e-06 0 6.5e-06 0 )
VWriteL 224 0 pwl (0 3 4.68e-07 3 4.71e-07 0 4.91e-07 0 
+ 4.94e-07 3 5.72e-07 3 5.75e-07 0 5.95e-07 0 
+ 5.98e-07 3 6.76e-07 3 6.79e-07 0 6.99e-07 0 
+ 7.02e-07 3 7.8e-07 3 7.83e-07 0 8.03e-07 0 
+ 8.06e-07 3 8.84e-07 3 8.87e-07 0 9.07e-07 0 
+ 9.1e-07 3 9.88e-07 3 9.91e-07 0 1.011e-06 0 
+ 1.014e-06 3 1.092e-06 3 1.095e-06 0 1.115e-06 0 
+ 1.118e-06 3 1.196e-06 3 1.199e-06 0 1.219e-06 0 
+ 1.222e-06 3 6.5e-06 3 )
VALoadH 17 0 pwl (0 0 2.6e-08 0 2.9e-08 3 4.9e-08 3 
+ 5.2e-08 0 7.8e-08 0 8.1e-08 3 1.01e-07 3 
+ 1.04e-07 0 1.3e-07 0 1.33e-07 3 1.53e-07 3 
+ 1.56e-07 0 1.82e-07 0 1.85e-07 3 2.05e-07 3 
+ 2.08e-07 0 2.34e-07 0 2.37e-07 3 2.57e-07 3 
+ 2.6e-07 0 2.86e-07 0 2.89e-07 3 3.09e-07 3 
+ 3.12e-07 0 3.38e-07 0 3.41e-07 3 3.61e-07 3 
+ 3.64e-07 0 3.9e-07 0 3.93e-07 3 4.13e-07 3 
+ 4.16e-07 0 4.94e-07 0 4.97e-07 3 5.17e-07 3 
+ 5.2e-07 0 5.98e-07 0 6.01e-07 3 6.21e-07 3 
+ 6.24e-07 0 7.02e-07 0 7.05e-07 3 7.25e-07 3 
+ 7.28e-07 0 8.06e-07 0 8.09e-07 3 8.29e-07 3 
+ 8.32e-07 0 9.1e-07 0 9.13e-07 3 9.33e-07 3 
+ 9.36e-07 0 1.014e-06 0 1.017e-06 3 1.037e-06 3 
+ 1.04e-06 0 1.118e-06 0 1.121e-06 3 1.141e-06 3 
+ 1.144e-06 0 1.222e-06 0 1.225e-06 3 1.245e-06 3 
+ 1.248e-06 0 1.274e-06 0 1.277e-06 3 1.297e-06 3 
+ 1.3e-06 0 1.742e-06 0 1.745e-06 3 1.765e-06 3 
+ 1.768e-06 0 2.21e-06 0 2.213e-06 3 2.233e-06 3 
+ 2.236e-06 0 2.678e-06 0 2.681e-06 3 2.701e-06 3 
+ 2.704e-06 0 3.146e-06 0 3.149e-06 3 3.169e-06 3 
+ 3.172e-06 0 3.614e-06 0 3.617e-06 3 3.637e-06 3 
+ 3.64e-06 0 4.082e-06 0 4.085e-06 3 4.105e-06 3 
+ 4.108e-06 0 4.55e-06 0 4.553e-06 3 4.573e-06 3 
+ 4.576e-06 0 6.5e-06 0 )
VALoadL 11 0 pwl (0 3 2.6e-08 3 2.9e-08 0 4.9e-08 0 
+ 5.2e-08 3 7.8e-08 3 8.1e-08 0 1.01e-07 0 
+ 1.04e-07 3 1.3e-07 3 1.33e-07 0 1.53e-07 0 
+ 1.56e-07 3 1.82e-07 3 1.85e-07 0 2.05e-07 0 
+ 2.08e-07 3 2.34e-07 3 2.37e-07 0 2.57e-07 0 
+ 2.6e-07 3 2.86e-07 3 2.89e-07 0 3.09e-07 0 
+ 3.12e-07 3 3.38e-07 3 3.41e-07 0 3.61e-07 0 
+ 3.64e-07 3 3.9e-07 3 3.93e-07 0 4.13e-07 0 
+ 4.16e-07 3 4.94e-07 3 4.97e-07 0 5.17e-07 0 
+ 5.2e-07 3 5.98e-07 3 6.01e-07 0 6.21e-07 0 
+ 6.24e-07 3 7.02e-07 3 7.05e-07 0 7.25e-07 0 
+ 7.28e-07 3 8.06e-07 3 8.09e-07 0 8.29e-07 0 
+ 8.32e-07 3 9.1e-07 3 9.13e-07 0 9.33e-07 0 
+ 9.36e-07 3 1.014e-06 3 1.017e-06 0 1.037e-06 0 
+ 1.04e-06 3 1.118e-06 3 1.121e-06 0 1.141e-06 0 
+ 1.144e-06 3 1.222e-06 3 1.225e-06 0 1.245e-06 0 
+ 1.248e-06 3 1.274e-06 3 1.277e-06 0 1.297e-06 0 
+ 1.3e-06 3 1.742e-06 3 1.745e-06 0 1.765e-06 0 
+ 1.768e-06 3 2.21e-06 3 2.213e-06 0 2.233e-06 0 
+ 2.236e-06 3 2.678e-06 3 2.681e-06 0 2.701e-06 0 
+ 2.704e-06 3 3.146e-06 3 3.149e-06 0 3.169e-06 0 
+ 3.172e-06 3 3.614e-06 3 3.617e-06 0 3.637e-06 0 
+ 3.64e-06 3 4.082e-06 3 4.085e-06 0 4.105e-06 0 
+ 4.108e-06 3 4.55e-06 3 4.553e-06 0 4.573e-06 0 
+ 4.576e-06 3 6.5e-06 3 )
VDLoadH 295 0 pwl (0 0 5.2e-08 0 5.5e-08 3 7.5e-08 3 
+ 7.8e-08 0 1.04e-07 0 1.07e-07 3 1.27e-07 3 
+ 1.3e-07 0 1.56e-07 0 1.59e-07 3 1.79e-07 3 
+ 1.82e-07 0 2.08e-07 0 2.11e-07 3 2.31e-07 3 
+ 2.34e-07 0 2.6e-07 0 2.63e-07 3 2.83e-07 3 
+ 2.86e-07 0 3.12e-07 0 3.15e-07 3 3.35e-07 3 
+ 3.38e-07 0 3.64e-07 0 3.67e-07 3 3.87e-07 3 
+ 3.9e-07 0 4.16e-07 0 4.19e-07 3 4.39e-07 3 
+ 4.42e-07 0 5.2e-07 0 5.23e-07 3 5.43e-07 3 
+ 5.46e-07 0 6.24e-07 0 6.27e-07 3 6.47e-07 3 
+ 6.5e-07 0 7.28e-07 0 7.31e-07 3 7.51e-07 3 
+ 7.54e-07 0 8.32e-07 0 8.35e-07 3 8.55e-07 3 
+ 8.58e-07 0 9.36e-07 0 9.39e-07 3 9.59e-07 3 
+ 9.62e-07 0 1.04e-06 0 1.043e-06 3 1.063e-06 3 
+ 1.066e-06 0 1.144e-06 0 1.147e-06 3 1.167e-06 3 
+ 1.17e-06 0 1.248e-06 0 1.251e-06 3 1.271e-06 3 
+ 1.274e-06 0 1.352e-06 0 1.355e-06 3 1.375e-06 3 
+ 1.378e-06 0 1.404e-06 0 1.407e-06 3 1.427e-06 3 
+ 1.43e-06 0 1.456e-06 0 1.459e-06 3 1.479e-06 3 
+ 1.482e-06 0 1.508e-06 0 1.511e-06 3 1.531e-06 3 
+ 1.534e-06 0 1.56e-06 0 1.563e-06 3 1.583e-06 3 
+ 1.586e-06 0 1.612e-06 0 1.615e-06 3 1.635e-06 3 
+ 1.638e-06 0 1.664e-06 0 1.667e-06 3 1.687e-06 3 
+ 1.69e-06 0 1.716e-06 0 1.719e-06 3 1.739e-06 3 
+ 1.742e-06 0 1.82e-06 0 1.823e-06 3 1.843e-06 3 
+ 1.846e-06 0 1.872e-06 0 1.875e-06 3 1.895e-06 3 
+ 1.898e-06 0 1.924e-06 0 1.927e-06 3 1.947e-06 3 
+ 1.95e-06 0 1.976e-06 0 1.979e-06 3 1.999e-06 3 
+ 2.002e-06 0 2.028e-06 0 2.031e-06 3 2.051e-06 3 
+ 2.054e-06 0 2.08e-06 0 2.083e-06 3 2.103e-06 3 
+ 2.106e-06 0 2.132e-06 0 2.135e-06 3 2.155e-06 3 
+ 2.158e-06 0 2.184e-06 0 2.187e-06 3 2.207e-06 3 
+ 2.21e-06 0 2.288e-06 0 2.291e-06 3 2.311e-06 3 
+ 2.314e-06 0 2.34e-06 0 2.343e-06 3 2.363e-06 3 
+ 2.366e-06 0 2.392e-06 0 2.395e-06 3 2.415e-06 3 
+ 2.418e-06 0 2.444e-06 0 2.447e-06 3 2.467e-06 3 
+ 2.47e-06 0 2.496e-06 0 2.499e-06 3 2.519e-06 3 
+ 2.522e-06 0 2.548e-06 0 2.551e-06 3 2.571e-06 3 
+ 2.574e-06 0 2.6e-06 0 2.603e-06 3 2.623e-06 3 
+ 2.626e-06 0 2.652e-06 0 2.655e-06 3 2.675e-06 3 
+ 2.678e-06 0 2.756e-06 0 2.759e-06 3 2.779e-06 3 
+ 2.782e-06 0 2.808e-06 0 2.811e-06 3 2.831e-06 3 
+ 2.834e-06 0 2.86e-06 0 2.863e-06 3 2.883e-06 3 
+ 2.886e-06 0 2.912e-06 0 2.915e-06 3 2.935e-06 3 
+ 2.938e-06 0 2.964e-06 0 2.967e-06 3 2.987e-06 3 
+ 2.99e-06 0 3.016e-06 0 3.019e-06 3 3.039e-06 3 
+ 3.042e-06 0 3.068e-06 0 3.071e-06 3 3.091e-06 3 
+ 3.094e-06 0 3.12e-06 0 3.123e-06 3 3.143e-06 3 
+ 3.146e-06 0 3.224e-06 0 3.227e-06 3 3.247e-06 3 
+ 3.25e-06 0 3.276e-06 0 3.279e-06 3 3.299e-06 3 
+ 3.302e-06 0 3.328e-06 0 3.331e-06 3 3.351e-06 3 
+ 3.354e-06 0 3.38e-06 0 3.383e-06 3 3.403e-06 3 
+ 3.406e-06 0 3.432e-06 0 3.435e-06 3 3.455e-06 3 
+ 3.458e-06 0 3.484e-06 0 3.487e-06 3 3.507e-06 3 
+ 3.51e-06 0 3.536e-06 0 3.539e-06 3 3.559e-06 3 
+ 3.562e-06 0 3.588e-06 0 3.591e-06 3 3.611e-06 3 
+ 3.614e-06 0 3.692e-06 0 3.695e-06 3 3.715e-06 3 
+ 3.718e-06 0 3.744e-06 0 3.747e-06 3 3.767e-06 3 
+ 3.77e-06 0 3.796e-06 0 3.799e-06 3 3.819e-06 3 
+ 3.822e-06 0 3.848e-06 0 3.851e-06 3 3.871e-06 3 
+ 3.874e-06 0 3.9e-06 0 3.903e-06 3 3.923e-06 3 
+ 3.926e-06 0 3.952e-06 0 3.955e-06 3 3.975e-06 3 
+ 3.978e-06 0 4.004e-06 0 4.007e-06 3 4.027e-06 3 
+ 4.03e-06 0 4.056e-06 0 4.059e-06 3 4.079e-06 3 
+ 4.082e-06 0 4.16e-06 0 4.163e-06 3 4.183e-06 3 
+ 4.186e-06 0 4.212e-06 0 4.215e-06 3 4.235e-06 3 
+ 4.238e-06 0 4.264e-06 0 4.267e-06 3 4.287e-06 3 
+ 4.29e-06 0 4.316e-06 0 4.319e-06 3 4.339e-06 3 
+ 4.342e-06 0 4.368e-06 0 4.371e-06 3 4.391e-06 3 
+ 4.394e-06 0 4.42e-06 0 4.423e-06 3 4.443e-06 3 
+ 4.446e-06 0 4.472e-06 0 4.475e-06 3 4.495e-06 3 
+ 4.498e-06 0 4.524e-06 0 4.527e-06 3 4.547e-06 3 
+ 4.55e-06 0 4.628e-06 0 4.631e-06 3 4.651e-06 3 
+ 4.654e-06 0 4.68e-06 0 4.683e-06 3 4.703e-06 3 
+ 4.706e-06 0 4.732e-06 0 4.735e-06 3 4.755e-06 3 
+ 4.758e-06 0 4.784e-06 0 4.787e-06 3 4.807e-06 3 
+ 4.81e-06 0 4.836e-06 0 4.839e-06 3 4.859e-06 3 
+ 4.862e-06 0 4.888e-06 0 4.891e-06 3 4.911e-06 3 
+ 4.914e-06 0 4.94e-06 0 4.943e-06 3 4.963e-06 3 
+ 4.966e-06 0 4.992e-06 0 4.995e-06 3 5.015e-06 3 
+ 5.018e-06 0 6.5e-06 0 )
VDLoadL 299 0 pwl (0 3 5.2e-08 3 5.5e-08 0 7.5e-08 0 
+ 7.8e-08 3 1.04e-07 3 1.07e-07 0 1.27e-07 0 
+ 1.3e-07 3 1.56e-07 3 1.59e-07 0 1.79e-07 0 
+ 1.82e-07 3 2.08e-07 3 2.11e-07 0 2.31e-07 0 
+ 2.34e-07 3 2.6e-07 3 2.63e-07 0 2.83e-07 0 
+ 2.86e-07 3 3.12e-07 3 3.15e-07 0 3.35e-07 0 
+ 3.38e-07 3 3.64e-07 3 3.67e-07 0 3.87e-07 0 
+ 3.9e-07 3 4.16e-07 3 4.19e-07 0 4.39e-07 0 
+ 4.42e-07 3 5.2e-07 3 5.23e-07 0 5.43e-07 0 
+ 5.46e-07 3 6.24e-07 3 6.27e-07 0 6.47e-07 0 
+ 6.5e-07 3 7.28e-07 3 7.31e-07 0 7.51e-07 0 
+ 7.54e-07 3 8.32e-07 3 8.35e-07 0 8.55e-07 0 
+ 8.58e-07 3 9.36e-07 3 9.39e-07 0 9.59e-07 0 
+ 9.62e-07 3 1.04e-06 3 1.043e-06 0 1.063e-06 0 
+ 1.066e-06 3 1.144e-06 3 1.147e-06 0 1.167e-06 0 
+ 1.17e-06 3 1.248e-06 3 1.251e-06 0 1.271e-06 0 
+ 1.274e-06 3 1.352e-06 3 1.355e-06 0 1.375e-06 0 
+ 1.378e-06 3 1.404e-06 3 1.407e-06 0 1.427e-06 0 
+ 1.43e-06 3 1.456e-06 3 1.459e-06 0 1.479e-06 0 
+ 1.482e-06 3 1.508e-06 3 1.511e-06 0 1.531e-06 0 
+ 1.534e-06 3 1.56e-06 3 1.563e-06 0 1.583e-06 0 
+ 1.586e-06 3 1.612e-06 3 1.615e-06 0 1.635e-06 0 
+ 1.638e-06 3 1.664e-06 3 1.667e-06 0 1.687e-06 0 
+ 1.69e-06 3 1.716e-06 3 1.719e-06 0 1.739e-06 0 
+ 1.742e-06 3 1.82e-06 3 1.823e-06 0 1.843e-06 0 
+ 1.846e-06 3 1.872e-06 3 1.875e-06 0 1.895e-06 0 
+ 1.898e-06 3 1.924e-06 3 1.927e-06 0 1.947e-06 0 
+ 1.95e-06 3 1.976e-06 3 1.979e-06 0 1.999e-06 0 
+ 2.002e-06 3 2.028e-06 3 2.031e-06 0 2.051e-06 0 
+ 2.054e-06 3 2.08e-06 3 2.083e-06 0 2.103e-06 0 
+ 2.106e-06 3 2.132e-06 3 2.135e-06 0 2.155e-06 0 
+ 2.158e-06 3 2.184e-06 3 2.187e-06 0 2.207e-06 0 
+ 2.21e-06 3 2.288e-06 3 2.291e-06 0 2.311e-06 0 
+ 2.314e-06 3 2.34e-06 3 2.343e-06 0 2.363e-06 0 
+ 2.366e-06 3 2.392e-06 3 2.395e-06 0 2.415e-06 0 
+ 2.418e-06 3 2.444e-06 3 2.447e-06 0 2.467e-06 0 
+ 2.47e-06 3 2.496e-06 3 2.499e-06 0 2.519e-06 0 
+ 2.522e-06 3 2.548e-06 3 2.551e-06 0 2.571e-06 0 
+ 2.574e-06 3 2.6e-06 3 2.603e-06 0 2.623e-06 0 
+ 2.626e-06 3 2.652e-06 3 2.655e-06 0 2.675e-06 0 
+ 2.678e-06 3 2.756e-06 3 2.759e-06 0 2.779e-06 0 
+ 2.782e-06 3 2.808e-06 3 2.811e-06 0 2.831e-06 0 
+ 2.834e-06 3 2.86e-06 3 2.863e-06 0 2.883e-06 0 
+ 2.886e-06 3 2.912e-06 3 2.915e-06 0 2.935e-06 0 
+ 2.938e-06 3 2.964e-06 3 2.967e-06 0 2.987e-06 0 
+ 2.99e-06 3 3.016e-06 3 3.019e-06 0 3.039e-06 0 
+ 3.042e-06 3 3.068e-06 3 3.071e-06 0 3.091e-06 0 
+ 3.094e-06 3 3.12e-06 3 3.123e-06 0 3.143e-06 0 
+ 3.146e-06 3 3.224e-06 3 3.227e-06 0 3.247e-06 0 
+ 3.25e-06 3 3.276e-06 3 3.279e-06 0 3.299e-06 0 
+ 3.302e-06 3 3.328e-06 3 3.331e-06 0 3.351e-06 0 
+ 3.354e-06 3 3.38e-06 3 3.383e-06 0 3.403e-06 0 
+ 3.406e-06 3 3.432e-06 3 3.435e-06 0 3.455e-06 0 
+ 3.458e-06 3 3.484e-06 3 3.487e-06 0 3.507e-06 0 
+ 3.51e-06 3 3.536e-06 3 3.539e-06 0 3.559e-06 0 
+ 3.562e-06 3 3.588e-06 3 3.591e-06 0 3.611e-06 0 
+ 3.614e-06 3 3.692e-06 3 3.695e-06 0 3.715e-06 0 
+ 3.718e-06 3 3.744e-06 3 3.747e-06 0 3.767e-06 0 
+ 3.77e-06 3 3.796e-06 3 3.799e-06 0 3.819e-06 0 
+ 3.822e-06 3 3.848e-06 3 3.851e-06 0 3.871e-06 0 
+ 3.874e-06 3 3.9e-06 3 3.903e-06 0 3.923e-06 0 
+ 3.926e-06 3 3.952e-06 3 3.955e-06 0 3.975e-06 0 
+ 3.978e-06 3 4.004e-06 3 4.007e-06 0 4.027e-06 0 
+ 4.03e-06 3 4.056e-06 3 4.059e-06 0 4.079e-06 0 
+ 4.082e-06 3 4.16e-06 3 4.163e-06 0 4.183e-06 0 
+ 4.186e-06 3 4.212e-06 3 4.215e-06 0 4.235e-06 0 
+ 4.238e-06 3 4.264e-06 3 4.267e-06 0 4.287e-06 0 
+ 4.29e-06 3 4.316e-06 3 4.319e-06 0 4.339e-06 0 
+ 4.342e-06 3 4.368e-06 3 4.371e-06 0 4.391e-06 0 
+ 4.394e-06 3 4.42e-06 3 4.423e-06 0 4.443e-06 0 
+ 4.446e-06 3 4.472e-06 3 4.475e-06 0 4.495e-06 0 
+ 4.498e-06 3 4.524e-06 3 4.527e-06 0 4.547e-06 0 
+ 4.55e-06 3 4.628e-06 3 4.631e-06 0 4.651e-06 0 
+ 4.654e-06 3 4.68e-06 3 4.683e-06 0 4.703e-06 0 
+ 4.706e-06 3 4.732e-06 3 4.735e-06 0 4.755e-06 0 
+ 4.758e-06 3 4.784e-06 3 4.787e-06 0 4.807e-06 0 
+ 4.81e-06 3 4.836e-06 3 4.839e-06 0 4.859e-06 0 
+ 4.862e-06 3 4.888e-06 3 4.891e-06 0 4.911e-06 0 
+ 4.914e-06 3 4.94e-06 3 4.943e-06 0 4.963e-06 0 
+ 4.966e-06 3 4.992e-06 3 4.995e-06 0 5.015e-06 0 
+ 5.018e-06 3 6.5e-06 3 )
VReadH 297 0 pwl (0 0 1.3e-06 0 1.303e-06 3 1.323e-06 3 
+ 1.326e-06 0 1.768e-06 0 1.771e-06 3 1.791e-06 3 
+ 1.794e-06 0 2.236e-06 0 2.239e-06 3 2.259e-06 3 
+ 2.262e-06 0 2.704e-06 0 2.707e-06 3 2.727e-06 3 
+ 2.73e-06 0 3.172e-06 0 3.175e-06 3 3.195e-06 3 
+ 3.198e-06 0 3.64e-06 0 3.643e-06 3 3.663e-06 3 
+ 3.666e-06 0 4.108e-06 0 4.111e-06 3 4.131e-06 3 
+ 4.134e-06 0 4.576e-06 0 4.579e-06 3 4.599e-06 3 
+ 4.602e-06 0 6.5e-06 0 )
VReadL 300 0 pwl (0 3 1.3e-06 3 1.303e-06 0 1.323e-06 0 
+ 1.326e-06 3 1.768e-06 3 1.771e-06 0 1.791e-06 0 
+ 1.794e-06 3 2.236e-06 3 2.239e-06 0 2.259e-06 0 
+ 2.262e-06 3 2.704e-06 3 2.707e-06 0 2.727e-06 0 
+ 2.73e-06 3 3.172e-06 3 3.175e-06 0 3.195e-06 0 
+ 3.198e-06 3 3.64e-06 3 3.643e-06 0 3.663e-06 0 
+ 3.666e-06 3 4.108e-06 3 4.111e-06 0 4.131e-06 0 
+ 4.134e-06 3 4.576e-06 3 4.579e-06 0 4.599e-06 0 
+ 4.602e-06 3 6.5e-06 3 )
VAShiftIn 340 0 pwl (0 0 3.77e-07 0 3.8e-07 3 4.27e-07 3 
+ 4.3e-07 0 1.26e-06 0 1.263e-06 3 1.31e-06 3 
+ 1.313e-06 0 6.5e-06 0 )
VDShiftIn 344 0 pwl (0 0 3.5e-08 0 3.8e-08 3 1.4e-07 3 
+ 1.43e-07 0 2.47e-07 0 2.5e-07 3 3e-07 3 
+ 3.03e-07 0 6.5e-06 0 )
VVdd 1 0 3.3 
.print TRAN v(285) v(4) v(219) v(17) v(340) v(295) 
+v(344) v(297) v(338) v(342) 
*.options limpts=50000 itl5=50000
.TRAN 1e-09 6.5e-06
.end
