******************************************************************
* For testing -o (SON Bug 911), the key point is that the -r
* command line option takes precedence over -o if both are
* specified on the command line in the .sh file.
******************************************************************

V1 1 0 PWL 0 0 1 1
R1 1 0 1

.TRAN 0 1
.PRINT TRAN V(1)
.OPTIONS OUTPUT INITIAL_INTERVAL=0.2 

.END


