************************************************************************
* Unit test for a Xyce warning message from .IC on a global node in a
* subcircuit, when the translated Xyce netlist is run. 
*
* This "gold" Xyce netlist is not actually run, just the translated
* Xyce netlist.
*
* See SRN Bug 1991
************************************************************************

*Analysis directives: 
.TRAN  0 10ms  
.PRINT TRAN V(N16554) V(N16997)

*RC Decay with IC in subcircuit
V_V3         N16554 0  PULSE(0 1 0 1e-3 1e-3 5e-3 1s)
R_R7         N16554 N16997  1k  
X_X1          N16997 N17112  IC_Subckt
R_R8         0 N17112  10 

.SUBCKT IC_Subckt in out
R1          in  mid 10 
C1          mid out 1u 
.IC         V(mid)=0.5
* setting IC on global node here should cause warning when
* Xyce netlist is run.  This uses $G_TL_VCC, so we can tell
* which netlist (this one, or the translated one) was tested.
.IC         V($G_TL_VCC)=0.0;
.ENDS

.END
