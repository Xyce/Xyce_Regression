* Test DC mode support for MAX, MIN and PP Measures
*
* This bug covers:
*   1) The case of two variables on the .DC line.  (Note:
*      since there is no .STEP statement, the output is treated
*      like one STEP, and the max is computed over all values
*      of vsrc1 and vsrc2.
*
*   2) the use of FROM and TO statements, where the FROM
*      value is always less than TO value.  If there are
*      more than one variable on the .DC line, then the
*      first variable (vsrc1) is used with the FROM-TO
*      qualifiers.
*
*   3) Have one sweep variable (vsrc1) be monotonically decreasing,
*      while the other (vsrc2) is monotonically increasing 
*
* See SON Bug 884 for more details.
**************************************************************

vsrc1   1a 0 1
rload1a 1a 1b 0.1
rload1b 1b 0 1

vsrc2   2a 0 1
rload2a 2a 1b 0.2

.DC vsrc1 5 1 -1 vsrc2 2 5 3

* Note: vsrc1:DCV0 is the syntax for printing the DC value of vsrc1,
* as it is swept. 
.print dc vsrc1:DCV0 vsrc2:DCV0 v(1a) v(2a) v(1b)

* MAX measure
.measure dc maxv1b   max v(1b)
.measure dc maxv1bFT max v(1b) FROM=2 TO=4

*MIN measure
.measure dc minv1b   min v(1b)
.measure dc minv1bFT min v(1b) FROM=2 TO=4

* PP measure
.measure dc ppv1b   pp v(1b)
.measure dc ppv1bFT pp v(1b) FROM=2 TO=4

.end


