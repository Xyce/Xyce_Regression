Test parameer file substitution and response file generation
*
* run this with Xyce -prf <param file> -rsf <respone file> rc_template.cir
*
* Xyce will fill in var "dakota_C1C" with value from param file
* and output .measure responese 

V1  1  0  pulse (1  0  2e-4  1e-9 1e-9  1 1 100)
R1  1  OBJ  dakota_R1R
C1  OBJ 0   dakota_C1C

.measure tran TimeAt2 when v(OBJ)=0.35 MINVAL=0.02

.tran 0 1e-3
.print tran V(OBJ)
.end
