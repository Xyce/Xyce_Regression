level=1 diode circuit
*
* ERK.  1/22/2014.
*
V2 2 0 0.21
D2 2 0 DA lambertw=0

.MODEL DA D  (IS=1.0e-12  RS=0.25  N=1.0)

*.STEP DA:IS 1.0e-12 1.0e-12 1.0e-12
*.STEP DA:RS 0.25 0.25 1.0e-1
*.SENS objfunc={-I(V2)} param=DA:IS,DA:RS
*.options DEVICE DEBUGLEVEL=2 
*.options SENSITIVITY DAKOTAFILE=1  direct=1 adjoint=0  STDOUTPUT=0
*.DC V2 0.0 1.0 0.01 
.rol V2 0.0 1.0 0.01  
.options device voltlim=0
*.OPTIONS TIMEINT RELTOL=1e-8 ABSTOL=1e-12
*.OPTIONS TIMEINT ERROPTION=1 DELMAX=1.0e-4
*.TRAN 1us 100ms NOOP 
.print DC v(2) {-I(V2)}
*.print tran v(2) {-I(V2)}
*.print SENS format=std 

.END

