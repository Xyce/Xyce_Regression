Test circuit for AC output through expressions

v1 a 0 AC 1
R1 a b 1
R2 b 0 2
C1 a b 1u

.ac dec 10 1 1e5
.print ac V(A) V(B) V(A,B) VR(A,B) VI(A,B) VM(A,B) VDB(A,B) VP(A,B)
.end
