* Gold Xyce netlist for testing .DC analysis and printing

*Analysis directives: 
.DC V1 LIST 1 3 5
.PRINT DC FORMAT=PROBE V(1) V(2a) V(2b) I(R1) W(R1) I(R3) W(R3) V(*)

*simple resistor divider
V1 1 0 1
R1 1  2a 1
R2 2a 2b 1
R3 2b 0 3
R4 2b 0 1

.END

