* Test voltage difference operator, after fix
* for SON Bug 718.  This netlist uses GND as a
* synonym for node 0.  This netlist also tests
* SON Bug 1030, which was about using N(1) inside
* of an expression.

.PREPROCESS REPLACEGROUND TRUE
.TRAN 0 1
.OPTIONS OUTPUT INITIAL_INTERVAL=0.2
.PRINT TRAN PRECISION=3 
+ V(1,0) V(1,1) V(1,2) V(1,3) V(1,4)
+ V(2,0) V(2,1) V(2,2) V(2,3) V(2,4)
+ V(GND,3) V(3,1) V(3,2) V(3,3) V(3,4)
+ {V(0,4)} {V(4,1)} {V(4,2)} {V(4,3)} {V(4,4)}
+ V(0) {V(1)}  
+ N(1) {N(1)} N(GND)
V1 1 0 PWL 0 0 1 1
R1 1 2 1
R2 2 3 1
R3 3 4 1
R4 4 0 1

.END
