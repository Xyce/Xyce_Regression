* Test NOISE mode support for the FIND-AT, FIND-WHEN and WHEN measures.
* It was deemed sufficient to mostly just test with the VR and VI operators.
* Expressions are also tested. One current operator (IM) is tested for a
* branch current.
*
* See SON Bug 1301 for more details.
********************************************************************

* RESISTOR DIVIDER
V1  1 0 DC 5.0 AC  1.0
R1  1 2 100K
R2  2 0 100K
*
* AMP AND LP FILTER
EAMP   3 0 2 0 1
CLP1   3 4  2e-4
RLP1a  4 5 50
RLP1b  5 0 50

.NOISE  V(4)  V1  DEC  10 1 100
.STEP RLP1a 50 100 50
.PRINT NOISE VM(4) VR(4) VI(4) VM(5) VR(5) VI(5)

* WHEN
.MEASURE NOISE whenvr4 WHEN vr(4)=0.4
.MEASURE NOISE whenvi4 WHEN vi(4)=0.15

* FIND-WHEN
.MEASURE NOISE whenvr3 FIND VM(5) WHEN vr(4)=0.4
.MEASURE NOISE whenvi3 FIND VM(5) WHEN vi(4)=0.15

* FIND-AT
.MEASURE NOISE at30 FIND vi(4) at 3e1
.MEASURE NOISE at50 FIND {vi(4)+1} at 5e1

* Expressions, with FIND-WHEN measure
.MEASURE NOISE findvm3awhenvm4Exp1 find vm(5) when {vm(4)+0.1}=0.5
.MEASURE NOISE findvm3awhenvm4Exp2 find vm(5) when vm(4)={0.3+0.1}
.MEASURE NOISE findvm3awhenvm4Exp3 find {vm(5)+1} when {vm(4)+0.1}=0.5
.MEASURE NOISE findvm3awhenvm4Exp4 find {vm(5)+1} when vm(4)={0.3+0.1}
.MEASURE NOISE findvr3awhenvm4Exp5 find vr(5) when vr(4)=vi(4)

* Signifies end of test. .sh file looks for a measure named lastMeasure.
* This is needed for compatibility for testing with a verbose build, which
* is often used by the Xyce developers.
.measure noise lastMeasure max vm(4)

.END
