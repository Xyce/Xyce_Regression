* Netlist to test MPDE output in CSV format.
* This version has explicit .print lines for each type of
* MPDE output.  See SON Bug 969 for more details.

*simple LC Tank Oscillator

.mpde 0 1.0e-8
.print mpde FORMAT=CSV {v(1)+2}
.print mpde_ic FORMAT=CSV {v(1)+3}
.print mpde_startup FORMAT=CSV {v(1)+4}
.print tran {v(1)+3}

.param pi = 3.1415926
.param L = {4.869e-7/2/pi}
.param C = {2e-12/2/pi}
.param R = 20k
.param Gn = {-1.1*1/R}
.param satval = {1/R}

.options mpdeint startupperiods=2 ic=4 auton2=true T2=9.8681e-10 saveicdata=1 diff=1 wampde=1 phase=1 phasecoeff=0 oscout="I(L1)"
.options timeint-mpde method=8 erroption=1 delmax=1e-9
.options timeint method=7 newlte=1

r1 1 0 R
c1 1 0 C
l1 1 0 L
B1 1 0 I={satval*tanh(Gn/satval*V(1))}

.ic V(1)=0.58

.end
