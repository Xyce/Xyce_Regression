Power test for resistor
*
iIN  1 0 sin(0 1 4 0 0 ) 
R1   1 2 1K
R2   0 2 100

.options timeint method=gear
.options nonlin-tran rhstol=1.0e-7
.TRAN 0.5U 400ms
.PRINT TRAN v(1) {I(IIN)*v(1)} p(iin) w(iin) p(r1) p(r2) w(r1) w(r2)
.END
