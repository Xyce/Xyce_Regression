*-------------------------------------------------------------------------
* Copyright Notice
*
* Copyright (c) 2000, Sandia Corporation, Albuquerque, NM.
*-------------------------------------------------------------------------
*
*-------------------------------------------------------------------------
* Filename       : $RCSfile$
*
* Purpose        : PDE Diode test circuit , transient.
*
* Special Notes  : This is in the test suite to test out the PDE capability
*                  for the transient case.  It is a very simple voltage
*                  regulator, with one diode, and an input sinewave that
*                  goes for half a period.
*
*                  This is also a partial test of the new doping
*                  specificaiton, and the new electrode specification,
*                  which both depend on the metadata "vector composite".
*
* Creator        : Eric R. Keiter, 9233, Computational Sciences
*
* Creation Date  : 02/17/04
*
* Revision Information:
* ---------------------
*
* Revision Number: $Revision$
*
* Revision Date  : $Date$
*
* Current Owner  : $Author$
*-------------------------------------------------------------------------
R 1 2 1000.0
VP 1 0 PULSE(0 1.5 0.0 1.0e-2 0.0 1.0e+20 1.2e+20)
VF 2 1 SIN(0 0.5 50 1.0e-2)
VT1 4 0 0V
R1 2 3 1k
*------------- Diode PDE device ------------------
.param CERTPARAM=2.5e-4
YPDE Z1DIODE 3 4 PDEDIODE  
+ tecplotlevel=2 
+ l={2*CERTPARAM} nx=11 
* ELECTRODES:
*+ node = {name           =     anode, cathode
*+         bc             = dirichlet, dirichlet
*+         material       =   neutral, neutral
*+         oxideBndryFlag =         0, 0         }
*DOPING REGIONS:
+ region= {name     =    nreg,    preg
+          function =    step,    step
+          type     =   ntype,    ptype
+          nmax     = 1.0e+19,  1.0e+19
+          nmin     = 0.0e+00,    0.0 
+          xloc     =    {CERTPARAM},  2.5e-4
+          flatx    =    -1  ,       1  }
*--------end of  Diode PDE device ----------------
.model PDEDIODE  ZOD  level=1 

.tran 1.0e-3 2.0e-2
.print tran v(1) v(2) v(3) v(4) 
*COMP v(3) RELTOL=0.02
.options nonlin maxstep=100 maxsearchstep=3 
+ searchmethod=2  nox=1 debuglevel=-10
+ auger=false

* Set transient nonlinear solver options to be 
* the same as the DCOP options:
.options nonlin-tran maxstep=100 maxsearchstep=3 
+ searchmethod=2  nox=1 debuglevel=-10
+ abstol=1.0E-12
+ reltol=1.0E-3
+ deltaxtol=1.0
+ smallupdatetol=1.0e-6
+ rhstol=1.0E-6

.options device debuglevel=-10

.END
