% Flattened test of hierarhical libraries

vd d 0 dc 1.8
vg g 0 dc 0
vf f 0 dc 1.5

r1 g d 1k
r2 g f 2k

.dc vg 0 1.8 0.01

.print dc i(vd) i(vf)

.param x = 1
.param x2  = '(x)/3.0'

.end

